
-- ARCHIVO AUTOGENERADO CON generate_weights_package.py

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.perceptron_package.perceptron_input;

package mnist_weights is
    function GetWeights(Dummy: natural)
    return perceptron_input;
end package mnist_weights;

package body mnist_weights is
    function GetWeights(Dummy: natural) return perceptron_input is
        variable pesos_i : perceptron_input(25855 downto 0);
    begin
	pesos_i(0) := b"1111111111111111_1111111111111111_1111011111100111_1110000010111100"; -- -0.03161807452713447
	pesos_i(1) := b"1111111111111111_1111111111111111_1111101100000011_1100010110011100"; -- -0.01947369528305214
	pesos_i(2) := b"1111111111111111_1111111111111111_1110000111011001_0100111001011011"; -- -0.11777792236813982
	pesos_i(3) := b"1111111111111111_1111111111111111_1110000011001110_1110111010100101"; -- -0.12184246523535161
	pesos_i(4) := b"0000000000000000_0000000000000000_0000100001100101_0111010001100100"; -- 0.03279807503565847
	pesos_i(5) := b"1111111111111111_1111111111111111_1111010111111010_0000101110100010"; -- -0.03915335927399165
	pesos_i(6) := b"1111111111111111_1111111111111111_1111000000010110_1110101111110110"; -- -0.06215024223537822
	pesos_i(7) := b"1111111111111111_1111111111111111_1110001100111000_1000011101101110"; -- -0.11241868556472205
	pesos_i(8) := b"1111111111111111_1111111111111111_1110011000110101_0010111111111000"; -- -0.10075092511134867
	pesos_i(9) := b"0000000000000000_0000000000000000_0001010010101001_1111111010101001"; -- 0.08071891417679866
	pesos_i(10) := b"0000000000000000_0000000000000000_0001000111101000_1000111111110111"; -- 0.06995487008955312
	pesos_i(11) := b"1111111111111111_1111111111111111_1110110101000001_0001000111110001"; -- -0.07322585927018169
	pesos_i(12) := b"0000000000000000_0000000000000000_0000110111000111_0111001100111110"; -- 0.053824618031184226
	pesos_i(13) := b"1111111111111111_1111111111111111_1101100111110000_1010001010100010"; -- -0.14867194685785493
	pesos_i(14) := b"0000000000000000_0000000000000000_0000110011011111_1000100100011111"; -- 0.050285882927378824
	pesos_i(15) := b"1111111111111111_1111111111111111_1110100110110111_1010011111100110"; -- -0.08704138398434234
	pesos_i(16) := b"1111111111111111_1111111111111111_1110001001110001_0111111101000011"; -- -0.11545567146168145
	pesos_i(17) := b"0000000000000000_0000000000000000_0010011101100000_0001101011111110"; -- 0.1538102025736196
	pesos_i(18) := b"1111111111111111_1111111111111111_1110110110001100_1110101111100010"; -- -0.07206845981159245
	pesos_i(19) := b"1111111111111111_1111111111111111_1101110011011100_0111110000111100"; -- -0.13726066141080057
	pesos_i(20) := b"1111111111111111_1111111111111111_1101110011010100_0110101001100111"; -- -0.137383794600872
	pesos_i(21) := b"0000000000000000_0000000000000000_0010100100111110_0001001001011101"; -- 0.16110338935531468
	pesos_i(22) := b"0000000000000000_0000000000000000_0000110000101110_0110111010101011"; -- 0.047583500698610746
	pesos_i(23) := b"1111111111111111_1111111111111111_1111101000011001_1110010001010101"; -- -0.02304242058749427
	pesos_i(24) := b"1111111111111111_1111111111111111_1110101010001011_1001001011100011"; -- -0.08380777316003643
	pesos_i(25) := b"1111111111111111_1111111111111111_1111111100110110_0010101011111101"; -- -0.0030797130788295254
	pesos_i(26) := b"1111111111111111_1111111111111111_1101111010100001_1100110110110010"; -- -0.13034357446985304
	pesos_i(27) := b"0000000000000000_0000000000000000_0010000101110010_0001010000001010"; -- 0.13064694626488924
	pesos_i(28) := b"0000000000000000_0000000000000000_0010011110110000_0101100001010111"; -- 0.15503456229516235
	pesos_i(29) := b"0000000000000000_0000000000000000_0010011100100010_0010101011011000"; -- 0.1528651025093835
	pesos_i(30) := b"1111111111111111_1111111111111111_1111011110111001_0000101111011001"; -- -0.03233266778054181
	pesos_i(31) := b"0000000000000000_0000000000000000_0010101101000100_1001100011111101"; -- 0.16901546639199108
	pesos_i(32) := b"1111111111111111_1111111111111111_1111010110010101_1011111110100101"; -- -0.040683767411660327
	pesos_i(33) := b"0000000000000000_0000000000000000_0010000100000010_0111000101011101"; -- 0.12894352461056824
	pesos_i(34) := b"1111111111111111_1111111111111111_1101111010010010_0011101101100101"; -- -0.13058117658970406
	pesos_i(35) := b"1111111111111111_1111111111111111_1101100001001001_1100100001111001"; -- -0.15512415936702767
	pesos_i(36) := b"0000000000000000_0000000000000000_0000000110111010_0000010001111100"; -- 0.006744652132289993
	pesos_i(37) := b"0000000000000000_0000000000000000_0001001101110111_0110001000111101"; -- 0.0760404014305612
	pesos_i(38) := b"0000000000000000_0000000000000000_0001111111010010_1011001101010000"; -- 0.12430878354311159
	pesos_i(39) := b"1111111111111111_1111111111111111_1111000101100100_1000001010111111"; -- -0.057060078073315784
	pesos_i(40) := b"1111111111111111_1111111111111111_1110100111100111_1111111000101000"; -- -0.08630382082424717
	pesos_i(41) := b"1111111111111111_1111111111111111_1111101000001000_1100100011011110"; -- -0.023303457150714302
	pesos_i(42) := b"1111111111111111_1111111111111111_1110101100110000_1011110011101011"; -- -0.08128756766046309
	pesos_i(43) := b"0000000000000000_0000000000000000_0001001100010110_0101010000110111"; -- 0.07455946300757708
	pesos_i(44) := b"0000000000000000_0000000000000000_0010001101110110_0011101110001100"; -- 0.13852283638107207
	pesos_i(45) := b"0000000000000000_0000000000000000_0001111001111000_0111111010010010"; -- 0.11902609897853393
	pesos_i(46) := b"0000000000000000_0000000000000000_0001100011011111_0101000011000010"; -- 0.09715752356480374
	pesos_i(47) := b"1111111111111111_1111111111111111_1110100101100010_1001001001110100"; -- -0.08833965948457989
	pesos_i(48) := b"1111111111111111_1111111111111111_1110101111011100_0110011100111011"; -- -0.07866816332513815
	pesos_i(49) := b"1111111111111111_1111111111111111_1110000100101010_1001011010101110"; -- -0.12044389953798829
	pesos_i(50) := b"1111111111111111_1111111111111111_1111110101110101_1100100111101110"; -- -0.00992143575741833
	pesos_i(51) := b"1111111111111111_1111111111111111_1110101010011111_1111001100001001"; -- -0.08349686647420292
	pesos_i(52) := b"0000000000000000_0000000000000000_0001101010000101_1111001111001101"; -- 0.1036064506383856
	pesos_i(53) := b"0000000000000000_0000000000000000_0010010001001100_1101011011010100"; -- 0.1417974728129746
	pesos_i(54) := b"1111111111111111_1111111111111111_1110011100110000_1010011111100110"; -- -0.09691382052213748
	pesos_i(55) := b"1111111111111111_1111111111111111_1110001100111100_1100011110010111"; -- -0.11235382608639428
	pesos_i(56) := b"1111111111111111_1111111111111111_1111010000010011_1101100100001100"; -- -0.04657214603772061
	pesos_i(57) := b"1111111111111111_1111111111111111_1110011001101100_0001101001011011"; -- -0.0999129799545747
	pesos_i(58) := b"1111111111111111_1111111111111111_1110001110001000_1101010111110110"; -- -0.1111933016060094
	pesos_i(59) := b"0000000000000000_0000000000000000_0010101010011001_0011100011010110"; -- 0.16640048233912832
	pesos_i(60) := b"1111111111111111_1111111111111111_1111111001001000_1001011110011110"; -- -0.006704830114390124
	pesos_i(61) := b"1111111111111111_1111111111111111_1111110110100100_0010100110011111"; -- -0.009213827708677966
	pesos_i(62) := b"0000000000000000_0000000000000000_0000011001110110_0010111110110100"; -- 0.02524088053339395
	pesos_i(63) := b"1111111111111111_1111111111111111_1101100010011010_0111000010111001"; -- -0.15389342779038537
	pesos_i(64) := b"0000000000000000_0000000000000000_0010011110111010_1001011101001110"; -- 0.15519090324651766
	pesos_i(65) := b"1111111111111111_1111111111111111_1101100100110100_1000111011001001"; -- -0.1515417822969979
	pesos_i(66) := b"0000000000000000_0000000000000000_0000111111101010_0110111010011010"; -- 0.06217089907476693
	pesos_i(67) := b"1111111111111111_1111111111111111_1111110011101001_0011101010100101"; -- -0.012066206647882403
	pesos_i(68) := b"1111111111111111_1111111111111111_1111010110010101_1011001000001100"; -- -0.040684578067774285
	pesos_i(69) := b"1111111111111111_1111111111111111_1101010011110011_0000100000011010"; -- -0.16816663147054772
	pesos_i(70) := b"0000000000000000_0000000000000000_0000101010000110_1010111101110111"; -- 0.041117636146111976
	pesos_i(71) := b"1111111111111111_1111111111111111_1101110011110101_0101110000010001"; -- -0.13688110912228257
	pesos_i(72) := b"0000000000000000_0000000000000000_0000101001010010_0110110010101100"; -- 0.040320198117852514
	pesos_i(73) := b"1111111111111111_1111111111111111_1111100010101010_1111000110000001"; -- -0.02864161118524658
	pesos_i(74) := b"0000000000000000_0000000000000000_0010010110001100_0100010011011010"; -- 0.14667158429612237
	pesos_i(75) := b"1111111111111111_1111111111111111_1111010101100000_0100010100100011"; -- -0.041499785302347214
	pesos_i(76) := b"0000000000000000_0000000000000000_0010110010000101_0100000111001000"; -- 0.17390833984951415
	pesos_i(77) := b"0000000000000000_0000000000000000_0000111010011000_1111100011100000"; -- 0.05702166993907242
	pesos_i(78) := b"0000000000000000_0000000000000000_0000011101101011_0011100111111111"; -- 0.02897989728585714
	pesos_i(79) := b"1111111111111111_1111111111111111_1111001110000100_0010110010100101"; -- -0.048764428832682574
	pesos_i(80) := b"1111111111111111_1111111111111111_1110110111100100_1011110111001011"; -- -0.07072843348991041
	pesos_i(81) := b"1111111111111111_1111111111111111_1101110101111000_1011001101111100"; -- -0.1348769971034041
	pesos_i(82) := b"1111111111111111_1111111111111111_1111100111111011_0111001100111100"; -- -0.02350692553589578
	pesos_i(83) := b"1111111111111111_1111111111111111_1110000101000000_0000001011011001"; -- -0.12011701773347103
	pesos_i(84) := b"0000000000000000_0000000000000000_0001111110111111_0000001111111001"; -- 0.12400841552645711
	pesos_i(85) := b"0000000000000000_0000000000000000_0010101001111100_0000100111001100"; -- 0.16595517377933489
	pesos_i(86) := b"0000000000000000_0000000000000000_0000000100110000_0001110111011100"; -- 0.004640451563308637
	pesos_i(87) := b"1111111111111111_1111111111111111_1110100010001001_1111011111010001"; -- -0.09164477494532536
	pesos_i(88) := b"0000000000000000_0000000000000000_0010010100010111_0010000011001101"; -- 0.14488415727968038
	pesos_i(89) := b"0000000000000000_0000000000000000_0010101100010111_0000011001010111"; -- 0.1683200800804979
	pesos_i(90) := b"0000000000000000_0000000000000000_0000010111000110_1010110000011010"; -- 0.022562748191338685
	pesos_i(91) := b"0000000000000000_0000000000000000_0001111000000100_1001010010000010"; -- 0.11725738681044703
	pesos_i(92) := b"0000000000000000_0000000000000000_0001000010111101_0100000100110011"; -- 0.06538779726844132
	pesos_i(93) := b"0000000000000000_0000000000000000_0000100000011011_0101011100001000"; -- 0.031667174694084636
	pesos_i(94) := b"0000000000000000_0000000000000000_0010100001111100_1010111100001101"; -- 0.1581525237418916
	pesos_i(95) := b"0000000000000000_0000000000000000_0000110110000101_0111001100001110"; -- 0.05281752662491576
	pesos_i(96) := b"0000000000000000_0000000000000000_0010010011111011_1110000010111001"; -- 0.1444683506472623
	pesos_i(97) := b"1111111111111111_1111111111111111_1101111001111111_1000000001010010"; -- -0.13086698534584745
	pesos_i(98) := b"0000000000000000_0000000000000000_0000000011100000_0000010001101001"; -- 0.0034182316113617723
	pesos_i(99) := b"1111111111111111_1111111111111111_1110111011101010_1101010111101110"; -- -0.06672919218617751
	pesos_i(100) := b"1111111111111111_1111111111111111_1110111111101101_0101000110111110"; -- -0.06278504474145974
	pesos_i(101) := b"1111111111111111_1111111111111111_1111010100100111_1001110011110011"; -- -0.04236430240028495
	pesos_i(102) := b"0000000000000000_0000000000000000_0010011011000110_0010011110101101"; -- 0.15146110520144546
	pesos_i(103) := b"1111111111111111_1111111111111111_1111101101010000_0001000100011101"; -- -0.018309526841973733
	pesos_i(104) := b"1111111111111111_1111111111111111_1110100011101100_1111100000011001"; -- -0.09013413794888693
	pesos_i(105) := b"1111111111111111_1111111111111111_1111111101011011_1001010111110100"; -- -0.0025087622826053097
	pesos_i(106) := b"0000000000000000_0000000000000000_0010011010000100_1010010001100011"; -- 0.15046145832677915
	pesos_i(107) := b"1111111111111111_1111111111111111_1111011000101010_1001001011011101"; -- -0.03841287714367793
	pesos_i(108) := b"1111111111111111_1111111111111111_1101011111100011_1000011010111011"; -- -0.15668447430522883
	pesos_i(109) := b"0000000000000000_0000000000000000_0010100111101011_0111111010110011"; -- 0.1637496172357607
	pesos_i(110) := b"0000000000000000_0000000000000000_0010011011110100_0011111111011100"; -- 0.15216445083381483
	pesos_i(111) := b"0000000000000000_0000000000000000_0001000000000001_0101110100100000"; -- 0.0625208095208895
	pesos_i(112) := b"0000000000000000_0000000000000000_0010000010110010_0001001001000000"; -- 0.12771715215931154
	pesos_i(113) := b"0000000000000000_0000000000000000_0001110011001000_0001111110111110"; -- 0.11242864968784878
	pesos_i(114) := b"1111111111111111_1111111111111111_1111000101111010_0111100011011011"; -- -0.05672497407237017
	pesos_i(115) := b"0000000000000000_0000000000000000_0010010100110110_1001100100001101"; -- 0.14536434710703258
	pesos_i(116) := b"0000000000000000_0000000000000000_0000101100001000_0111110001100000"; -- 0.043098233586403606
	pesos_i(117) := b"1111111111111111_1111111111111111_1101100000011011_0011111011001111"; -- -0.15583426895873165
	pesos_i(118) := b"1111111111111111_1111111111111111_1110000101101001_0011011111011001"; -- -0.11948824846098795
	pesos_i(119) := b"1111111111111111_1111111111111111_1111111000100110_0010100001001001"; -- -0.007230264747085677
	pesos_i(120) := b"0000000000000000_0000000000000000_0000010101011000_1101011001011110"; -- 0.020886800731319766
	pesos_i(121) := b"1111111111111111_1111111111111111_1111101001001000_1110101000111110"; -- -0.02232490526281942
	pesos_i(122) := b"1111111111111111_1111111111111111_1111001101101011_1010100011000111"; -- -0.0491384997592164
	pesos_i(123) := b"0000000000000000_0000000000000000_0001111111000011_0111011011100111"; -- 0.12407630110278903
	pesos_i(124) := b"1111111111111111_1111111111111111_1111101101111011_0000010010000111"; -- -0.017654148982354498
	pesos_i(125) := b"0000000000000000_0000000000000000_0001010110111101_1011111011010101"; -- 0.08492653562149738
	pesos_i(126) := b"0000000000000000_0000000000000000_0001101111100001_0001001011001111"; -- 0.10890309852375922
	pesos_i(127) := b"0000000000000000_0000000000000000_0001101010101110_1101010001110110"; -- 0.10423019290690229
	pesos_i(128) := b"1111111111111111_1111111111111111_1101011101110011_1110101101000110"; -- -0.15838746583236896
	pesos_i(129) := b"1111111111111111_1111111111111111_1111011110110100_1110101010110101"; -- -0.03239567840474004
	pesos_i(130) := b"0000000000000000_0000000000000000_0000011011101001_0011001011011000"; -- 0.026995828462315154
	pesos_i(131) := b"1111111111111111_1111111111111111_1110010100110001_1011101111011101"; -- -0.10470987172913979
	pesos_i(132) := b"0000000000000000_0000000000000000_0001010110001000_1000101001000010"; -- 0.0841146861116127
	pesos_i(133) := b"0000000000000000_0000000000000000_0001100011111111_1110110101010101"; -- 0.09765513722379732
	pesos_i(134) := b"1111111111111111_1111111111111111_1111101100000101_1000111100111001"; -- -0.019446419417629878
	pesos_i(135) := b"0000000000000000_0000000000000000_0001100101100100_0101101001010100"; -- 0.09918751288142337
	pesos_i(136) := b"0000000000000000_0000000000000000_0000010111000101_0001101010111100"; -- 0.02253882489719633
	pesos_i(137) := b"1111111111111111_1111111111111111_1111000110111000_1111101101001110"; -- -0.05577115392836534
	pesos_i(138) := b"0000000000000000_0000000000000000_0000110110100110_1110000110011101"; -- 0.05332765658880942
	pesos_i(139) := b"1111111111111111_1111111111111111_1110100000111111_0110001000110110"; -- -0.09278284240853368
	pesos_i(140) := b"1111111111111111_1111111111111111_1111010011111101_1011011110000010"; -- -0.043003588529584934
	pesos_i(141) := b"0000000000000000_0000000000000000_0000001110110101_1001010110100101"; -- 0.014489510356614341
	pesos_i(142) := b"1111111111111111_1111111111111111_1110010101010001_0111011100101100"; -- -0.10422568490221053
	pesos_i(143) := b"1111111111111111_1111111111111111_1110101101111010_1110001010000100"; -- -0.08015617636732993
	pesos_i(144) := b"0000000000000000_0000000000000000_0000001001010000_0010101101110101"; -- 0.009035793391107688
	pesos_i(145) := b"1111111111111111_1111111111111111_1101011011100011_0011010111100010"; -- -0.16059554317421706
	pesos_i(146) := b"0000000000000000_0000000000000000_0001010001011100_0110000111111101"; -- 0.0795346491063194
	pesos_i(147) := b"1111111111111111_1111111111111111_1111111100111101_0111011101010001"; -- -0.0029683520069822646
	pesos_i(148) := b"0000000000000000_0000000000000000_0010001010101000_0110000111010001"; -- 0.1353818067607306
	pesos_i(149) := b"0000000000000000_0000000000000000_0000111011011011_0100111011111011"; -- 0.05803388230332562
	pesos_i(150) := b"0000000000000000_0000000000000000_0010011110010001_0010100010100110"; -- 0.15455869736560968
	pesos_i(151) := b"0000000000000000_0000000000000000_0001000001101110_0011000100101000"; -- 0.06418139674111388
	pesos_i(152) := b"1111111111111111_1111111111111111_1101010111110100_0011011001110110"; -- -0.16424235942616722
	pesos_i(153) := b"1111111111111111_1111111111111111_1110101101000111_0110001111101100"; -- -0.08094192019193068
	pesos_i(154) := b"1111111111111111_1111111111111111_1110010001101110_1100010001011001"; -- -0.10768483003587107
	pesos_i(155) := b"1111111111111111_1111111111111111_1110100011001011_0110111101011001"; -- -0.09064582889310192
	pesos_i(156) := b"1111111111111111_1111111111111111_1101111101101010_1001110000100011"; -- -0.12727951193946224
	pesos_i(157) := b"0000000000000000_0000000000000000_0000001000010100_1010100001100100"; -- 0.00812771264788688
	pesos_i(158) := b"1111111111111111_1111111111111111_1101111101000010_0010111101110100"; -- -0.12789634146079912
	pesos_i(159) := b"0000000000000000_0000000000000000_0010000111110100_0101110101001001"; -- 0.13263495477460227
	pesos_i(160) := b"1111111111111111_1111111111111111_1110100011000011_0010001000101001"; -- -0.09077250008746324
	pesos_i(161) := b"1111111111111111_1111111111111111_1101000110101001_0101110000101101"; -- -0.1810095205933277
	pesos_i(162) := b"0000000000000000_0000000000000000_0001100010100001_1000110110100000"; -- 0.09621510644674874
	pesos_i(163) := b"1111111111111111_1111111111111111_1111011011101110_1110010001001011"; -- -0.035417300901119664
	pesos_i(164) := b"1111111111111111_1111111111111111_1111101101111001_0110000100011100"; -- -0.017679148342255854
	pesos_i(165) := b"1111111111111111_1111111111111111_1111100110101011_1101110010100100"; -- -0.024721345976198107
	pesos_i(166) := b"1111111111111111_1111111111111111_1110110000000010_1100110101011101"; -- -0.07808224177096122
	pesos_i(167) := b"1111111111111111_1111111111111111_1110100101110000_0110101110001001"; -- -0.08812835606733095
	pesos_i(168) := b"0000000000000000_0000000000000000_0001010011001111_1010010111110101"; -- 0.0812934610472694
	pesos_i(169) := b"0000000000000000_0000000000000000_0001000010111010_1000001000000101"; -- 0.06534588460482914
	pesos_i(170) := b"1111111111111111_1111111111111111_1110010101110101_1011111000001000"; -- -0.10367214491903091
	pesos_i(171) := b"1111111111111111_1111111111111111_1101010110010101_1010100001100100"; -- -0.16568515364111994
	pesos_i(172) := b"0000000000000000_0000000000000000_0000100000000011_0001001000011110"; -- 0.03129685621226707
	pesos_i(173) := b"0000000000000000_0000000000000000_0000100100001110_0101100011001010"; -- 0.03537516526162151
	pesos_i(174) := b"0000000000000000_0000000000000000_0001011110110011_1110110000111101"; -- 0.09258915420404536
	pesos_i(175) := b"0000000000000000_0000000000000000_0010101000000011_1111000111010000"; -- 0.16412268952321776
	pesos_i(176) := b"1111111111111111_1111111111111111_1111000000100110_1001011000000100"; -- -0.06191122448300908
	pesos_i(177) := b"1111111111111111_1111111111111111_1110101001011111_1101110111100001"; -- -0.08447469013089583
	pesos_i(178) := b"0000000000000000_0000000000000000_0010010100100101_0101111100011111"; -- 0.14510149481718737
	pesos_i(179) := b"0000000000000000_0000000000000000_0010001001010111_0000001010010111"; -- 0.1341401690160611
	pesos_i(180) := b"1111111111111111_1111111111111111_1110100111010000_1001001110011101"; -- -0.08666112338440242
	pesos_i(181) := b"0000000000000000_0000000000000000_0001011111001100_1111100000001101"; -- 0.09297132791198619
	pesos_i(182) := b"1111111111111111_1111111111111111_1111010101010110_1011011111000000"; -- -0.04164554188857661
	pesos_i(183) := b"0000000000000000_0000000000000000_0001011010000100_1100110111101101"; -- 0.08796393426397094
	pesos_i(184) := b"0000000000000000_0000000000000000_0010011101001011_0001101001101110"; -- 0.1534897344117587
	pesos_i(185) := b"1111111111111111_1111111111111111_1111100011100110_0001101010000110"; -- -0.027738897597606026
	pesos_i(186) := b"1111111111111111_1111111111111111_1111111010111001_0000001000001100"; -- -0.004989502026141195
	pesos_i(187) := b"0000000000000000_0000000000000000_0001001000000000_1110111110010011"; -- 0.07032677977775435
	pesos_i(188) := b"1111111111111111_1111111111111111_1111001000011101_1100011100101111"; -- -0.05423312288171147
	pesos_i(189) := b"0000000000000000_0000000000000000_0001000100110001_0001001001000110"; -- 0.06715501977517652
	pesos_i(190) := b"0000000000000000_0000000000000000_0001010000111000_1111101100001000"; -- 0.07899445483540474
	pesos_i(191) := b"1111111111111111_1111111111111111_1110111101000111_1110011010001011"; -- -0.06530913460628344
	pesos_i(192) := b"1111111111111111_1111111111111111_1101110011010011_1000011100011001"; -- -0.13739734306990312
	pesos_i(193) := b"1111111111111111_1111111111111111_1111001001010001_0111001101000001"; -- -0.0534446684720573
	pesos_i(194) := b"0000000000000000_0000000000000000_0001011110110101_0001000101011001"; -- 0.09260662474991492
	pesos_i(195) := b"1111111111111111_1111111111111111_1111010110000011_1000111111110110"; -- -0.04096126796867747
	pesos_i(196) := b"1111111111111111_1111111111111111_1111110100001100_0100001010111010"; -- -0.011531667332216307
	pesos_i(197) := b"1111111111111111_1111111111111111_1101010000010100_0100000001010101"; -- -0.17156598982153295
	pesos_i(198) := b"0000000000000000_0000000000000000_0000100100110000_1001100010011001"; -- 0.03589776732057269
	pesos_i(199) := b"0000000000000000_0000000000000000_0001011001111100_0111011100000111"; -- 0.08783668432710856
	pesos_i(200) := b"0000000000000000_0000000000000000_0010011101100111_1000100111001110"; -- 0.15392361912086602
	pesos_i(201) := b"1111111111111111_1111111111111111_1101100011010000_1001011111001101"; -- -0.15306712380037074
	pesos_i(202) := b"1111111111111111_1111111111111111_1110111001000110_1110010111100001"; -- -0.06923068288344228
	pesos_i(203) := b"0000000000000000_0000000000000000_0001011001110100_0000101110100110"; -- 0.08770821385159641
	pesos_i(204) := b"0000000000000000_0000000000000000_0000010101110000_0100100000010110"; -- 0.02124453091528691
	pesos_i(205) := b"1111111111111111_1111111111111111_1111000110010000_1011011100110001"; -- -0.0563855653791534
	pesos_i(206) := b"1111111111111111_1111111111111111_1101110010001000_0011000100111000"; -- -0.13854687110789277
	pesos_i(207) := b"0000000000000000_0000000000000000_0010110010110011_0111010010111000"; -- 0.17461328028196293
	pesos_i(208) := b"1111111111111111_1111111111111111_1111110100010100_0101001111110110"; -- -0.011408569820678283
	pesos_i(209) := b"1111111111111111_1111111111111111_1110101110111000_1110111011101110"; -- -0.07920939152722957
	pesos_i(210) := b"1111111111111111_1111111111111111_1111000111100000_0010010011110101"; -- -0.05517357846778466
	pesos_i(211) := b"1111111111111111_1111111111111111_1111000000011010_0010000100000010"; -- -0.062101304133883865
	pesos_i(212) := b"1111111111111111_1111111111111111_1111101110001101_1010010101000010"; -- -0.017369910556244823
	pesos_i(213) := b"0000000000000000_0000000000000000_0000111000010001_0111000000101001"; -- 0.05495358471591151
	pesos_i(214) := b"1111111111111111_1111111111111111_1111000111010010_0010010101101000"; -- -0.05538717475750325
	pesos_i(215) := b"1111111111111111_1111111111111111_1110011000100000_1001010000101010"; -- -0.10106538756009088
	pesos_i(216) := b"0000000000000000_0000000000000000_0001111101010000_0010000111001110"; -- 0.12231646793250418
	pesos_i(217) := b"1111111111111111_1111111111111111_1101001001000101_0100010110000011"; -- -0.17863050039792477
	pesos_i(218) := b"0000000000000000_0000000000000000_0010100011110011_1110000101010010"; -- 0.159971315974598
	pesos_i(219) := b"1111111111111111_1111111111111111_1110101000100101_1111001100101101"; -- -0.08535843039130087
	pesos_i(220) := b"0000000000000000_0000000000000000_0000000011011110_0101000110111011"; -- 0.0033923226042471095
	pesos_i(221) := b"0000000000000000_0000000000000000_0000011000111100_0010100010011001"; -- 0.02435544713000558
	pesos_i(222) := b"0000000000000000_0000000000000000_0001000011101101_0010010110000011"; -- 0.06611856895319214
	pesos_i(223) := b"0000000000000000_0000000000000000_0000011101010011_0000100000000000"; -- 0.028610706248465095
	pesos_i(224) := b"0000000000000000_0000000000000000_0010001010110010_0000100001100000"; -- 0.13552906371573162
	pesos_i(225) := b"0000000000000000_0000000000000000_0000100010011101_0001100111001111"; -- 0.03364716815122836
	pesos_i(226) := b"0000000000000000_0000000000000000_0000011111111010_0011100010001110"; -- 0.03116181815900578
	pesos_i(227) := b"1111111111111111_1111111111111111_1101100011000000_1111000001001010"; -- -0.15330599011931093
	pesos_i(228) := b"0000000000000000_0000000000000000_0010011110000001_1101100101100001"; -- 0.15432509051673887
	pesos_i(229) := b"0000000000000000_0000000000000000_0000111000110101_0110100100101111"; -- 0.05550248517205107
	pesos_i(230) := b"1111111111111111_1111111111111111_1111010111000010_1000010011111111"; -- -0.040000617710600685
	pesos_i(231) := b"0000000000000000_0000000000000000_0010000110000110_1011111110001010"; -- 0.1309623442664589
	pesos_i(232) := b"0000000000000000_0000000000000000_0001011101101110_0100000010010000"; -- 0.09152606499540991
	pesos_i(233) := b"0000000000000000_0000000000000000_0000010000000110_1111110110101111"; -- 0.01573167353886719
	pesos_i(234) := b"1111111111111111_1111111111111111_1101101110010101_0010000010100001"; -- -0.14225574567742158
	pesos_i(235) := b"1111111111111111_1111111111111111_1110001111111000_0011001000011111"; -- -0.10949408290820845
	pesos_i(236) := b"0000000000000000_0000000000000000_0010001010011111_1001110111100011"; -- 0.1352480581734796
	pesos_i(237) := b"0000000000000000_0000000000000000_0001111011111100_0010110111010011"; -- 0.12103544624578834
	pesos_i(238) := b"0000000000000000_0000000000000000_0000010100101011_1010011000010011"; -- 0.020197276661974767
	pesos_i(239) := b"1111111111111111_1111111111111111_1111011101011111_0001111001110100"; -- -0.03370484981737307
	pesos_i(240) := b"0000000000000000_0000000000000000_0010011110101101_1000100000000100"; -- 0.15499162761596239
	pesos_i(241) := b"0000000000000000_0000000000000000_0000101110011111_0111110101001111"; -- 0.045402366364238646
	pesos_i(242) := b"1111111111111111_1111111111111111_1111011001000001_0100011111111011"; -- -0.03806638827157381
	pesos_i(243) := b"0000000000000000_0000000000000000_0010110101110101_0110111011011001"; -- 0.17757313541821587
	pesos_i(244) := b"1111111111111111_1111111111111111_1101100101111100_0001001100111000"; -- -0.15045051472407936
	pesos_i(245) := b"0000000000000000_0000000000000000_0000111100000000_0110101011100000"; -- 0.05860012033393054
	pesos_i(246) := b"0000000000000000_0000000000000000_0001000011000111_1111011001001001"; -- 0.06555117867017869
	pesos_i(247) := b"0000000000000000_0000000000000000_0001000111110001_0000010101010010"; -- 0.07008393534534987
	pesos_i(248) := b"0000000000000000_0000000000000000_0001101010010000_1000001101101101"; -- 0.10376759927762305
	pesos_i(249) := b"0000000000000000_0000000000000000_0010000100111110_1000110000001010"; -- 0.12986064194347927
	pesos_i(250) := b"1111111111111111_1111111111111111_1101111000101010_0010100100101101"; -- -0.13216917649190182
	pesos_i(251) := b"0000000000000000_0000000000000000_0010100010000010_0110111100011000"; -- 0.15824026426302557
	pesos_i(252) := b"1111111111111111_1111111111111111_1111011101000011_0011001000001011"; -- -0.03413092836189944
	pesos_i(253) := b"0000000000000000_0000000000000000_0001011001110011_0110111010001110"; -- 0.08769885029857828
	pesos_i(254) := b"0000000000000000_0000000000000000_0000101110110001_1001001110001001"; -- 0.045678349541710205
	pesos_i(255) := b"0000000000000000_0000000000000000_0001111010100101_0010010010011101"; -- 0.11970738246236931
	pesos_i(256) := b"0000000000000000_0000000000000000_0000000010010101_0101000000101001"; -- 0.002278337373153666
	pesos_i(257) := b"0000000000000000_0000000000000000_0001001100101111_1011100000000111"; -- 0.07494688200380349
	pesos_i(258) := b"1111111111111111_1111111111111111_1110110111100110_1101101000100100"; -- -0.07069622620669734
	pesos_i(259) := b"0000000000000000_0000000000000000_0000011011111111_0111000111011000"; -- 0.027335276747618778
	pesos_i(260) := b"0000000000000000_0000000000000000_0010000110010001_0001001010010011"; -- 0.1311198814638493
	pesos_i(261) := b"1111111111111111_1111111111111111_1110100111110001_1100010100011001"; -- -0.08615463398642852
	pesos_i(262) := b"0000000000000000_0000000000000000_0000100100101101_0111111001101111"; -- 0.035850431474785956
	pesos_i(263) := b"0000000000000000_0000000000000000_0000011000000111_0011000010010111"; -- 0.02354720763930745
	pesos_i(264) := b"1111111111111111_1111111111111111_1110011011111100_0111101010110101"; -- -0.09770997113613636
	pesos_i(265) := b"0000000000000000_0000000000000000_0000111110100110_1101110001001011"; -- 0.061139839443428955
	pesos_i(266) := b"1111111111111111_1111111111111111_1111100110000011_0011101110010101"; -- -0.02534129716049488
	pesos_i(267) := b"1111111111111111_1111111111111111_1111011000001101_1101001110011010"; -- -0.038851523333126255
	pesos_i(268) := b"0000000000000000_0000000000000000_0001010010011001_0010010011111101"; -- 0.08046179950217798
	pesos_i(269) := b"0000000000000000_0000000000000000_0000111000111111_0101110000011110"; -- 0.055654294287861526
	pesos_i(270) := b"1111111111111111_1111111111111111_1101011001001111_1010100001101000"; -- -0.1628470179147042
	pesos_i(271) := b"1111111111111111_1111111111111111_1110011110010011_0011100110111110"; -- -0.09540976630569473
	pesos_i(272) := b"0000000000000000_0000000000000000_0010100110000010_1110101001111101"; -- 0.16215386909158955
	pesos_i(273) := b"0000000000000000_0000000000000000_0000010100010111_1010101101100110"; -- 0.0198924182711254
	pesos_i(274) := b"0000000000000000_0000000000000000_0000001001111010_0110111110101111"; -- 0.009680729172073306
	pesos_i(275) := b"1111111111111111_1111111111111111_1111111101101000_1011101110110000"; -- -0.002308148860144503
	pesos_i(276) := b"0000000000000000_0000000000000000_0010010101011110_0010010111001001"; -- 0.14596782842034878
	pesos_i(277) := b"0000000000000000_0000000000000000_0001000000000110_1101011001011011"; -- 0.06260432937611655
	pesos_i(278) := b"0000000000000000_0000000000000000_0010011001001101_1110000011100001"; -- 0.14962583050155356
	pesos_i(279) := b"1111111111111111_1111111111111111_1100111111101101_1010110000010100"; -- -0.18777966022160256
	pesos_i(280) := b"0000000000000000_0000000000000000_0000101000001010_0010101001000010"; -- 0.03921760658768966
	pesos_i(281) := b"1111111111111111_1111111111111111_1111101000001000_1101001001110100"; -- -0.023302885590882057
	pesos_i(282) := b"0000000000000000_0000000000000000_0000110000111110_0111101001101110"; -- 0.047828342376348164
	pesos_i(283) := b"1111111111111111_1111111111111111_1110110010000011_1110101100111110"; -- -0.07611207710792402
	pesos_i(284) := b"1111111111111111_1111111111111111_1110101000001110_0001010001000110"; -- -0.08572266846472301
	pesos_i(285) := b"0000000000000000_0000000000000000_0000100010101101_0110000110110101"; -- 0.03389559427381334
	pesos_i(286) := b"1111111111111111_1111111111111111_1111110100010000_1001011001100110"; -- -0.01146564483627677
	pesos_i(287) := b"0000000000000000_0000000000000000_0001101111110011_0001000111110001"; -- 0.10917770517039779
	pesos_i(288) := b"1111111111111111_1111111111111111_1110110010101001_1110100101110001"; -- -0.07553235055880705
	pesos_i(289) := b"1111111111111111_1111111111111111_1101001011001101_0111111111010010"; -- -0.17655182951276518
	pesos_i(290) := b"1111111111111111_1111111111111111_1111100011100011_1001010110100001"; -- -0.027777336280727514
	pesos_i(291) := b"0000000000000000_0000000000000000_0001101001010110_1101001101100010"; -- 0.10288735517897983
	pesos_i(292) := b"0000000000000000_0000000000000000_0000110010001010_1010011111100100"; -- 0.048990719980346376
	pesos_i(293) := b"0000000000000000_0000000000000000_0001011100011011_0110111101010100"; -- 0.09026237286165137
	pesos_i(294) := b"1111111111111111_1111111111111111_1101001000011000_0000111101011000"; -- -0.17932037451847366
	pesos_i(295) := b"1111111111111111_1111111111111111_1110100100101101_0011000001111001"; -- -0.08915421538356086
	pesos_i(296) := b"0000000000000000_0000000000000000_0010000111011101_1000000111110000"; -- 0.13228618715182686
	pesos_i(297) := b"1111111111111111_1111111111111111_1110010000111010_1000000111110110"; -- -0.10848224391637255
	pesos_i(298) := b"0000000000000000_0000000000000000_0000010001110010_1010011001000111"; -- 0.01737441276388578
	pesos_i(299) := b"1111111111111111_1111111111111111_1101100010110010_1000001010110100"; -- -0.1535261450570129
	pesos_i(300) := b"1111111111111111_1111111111111111_1110101000001100_1010010010001000"; -- -0.08574458781781957
	pesos_i(301) := b"1111111111111111_1111111111111111_1111000010000100_1001000000010111"; -- -0.06047725144041826
	pesos_i(302) := b"1111111111111111_1111111111111111_1111010111011100_0010101001110011"; -- -0.03960928614644421
	pesos_i(303) := b"1111111111111111_1111111111111111_1110110101110001_1100001001110001"; -- -0.07248291730686882
	pesos_i(304) := b"0000000000000000_0000000000000000_0000000010111010_0010011100111000"; -- 0.002840472465131555
	pesos_i(305) := b"0000000000000000_0000000000000000_0001110101101110_1111001000100010"; -- 0.11497414900917349
	pesos_i(306) := b"1111111111111111_1111111111111111_1111111001001100_0111100000011011"; -- -0.006645673233416066
	pesos_i(307) := b"1111111111111111_1111111111111111_1111110111110110_0010111011100000"; -- -0.007962293911088934
	pesos_i(308) := b"0000000000000000_0000000000000000_0000011111010001_1011100011100001"; -- 0.030543856594827307
	pesos_i(309) := b"1111111111111111_1111111111111111_1111011111110100_0100011110000111"; -- -0.03142884201769076
	pesos_i(310) := b"1111111111111111_1111111111111111_1110001000010011_0010100111101001"; -- -0.11689508507862442
	pesos_i(311) := b"1111111111111111_1111111111111111_1100111110110111_1101001111001000"; -- -0.1886012684542979
	pesos_i(312) := b"1111111111111111_1111111111111111_1101111101100100_1100111000001000"; -- -0.12736809057697748
	pesos_i(313) := b"0000000000000000_0000000000000000_0010000000010010_0110110001110100"; -- 0.12528112253415075
	pesos_i(314) := b"0000000000000000_0000000000000000_0001011011111101_0111100000010010"; -- 0.08980513037566427
	pesos_i(315) := b"1111111111111111_1111111111111111_1111100001010001_0001001101110100"; -- -0.030012878704691652
	pesos_i(316) := b"0000000000000000_0000000000000000_0010101010101101_0111101111100111"; -- 0.16670965561891193
	pesos_i(317) := b"0000000000000000_0000000000000000_0001000100000000_0000000001011010"; -- 0.06640627093407876
	pesos_i(318) := b"1111111111111111_1111111111111111_1111011100110010_1110101111100000"; -- -0.03437925131752839
	pesos_i(319) := b"1111111111111111_1111111111111111_1101110000011101_1010101111111001"; -- -0.1401722446370988
	pesos_i(320) := b"0000000000000000_0000000000000000_0000001101101000_1101101010100010"; -- 0.013318695692692506
	pesos_i(321) := b"0000000000000000_0000000000000000_0000010010110010_0111100100100011"; -- 0.018348284751329613
	pesos_i(322) := b"1111111111111111_1111111111111111_1101111010001111_1110010011111100"; -- -0.1306168446510942
	pesos_i(323) := b"0000000000000000_0000000000000000_0010011001111011_0010101110100100"; -- 0.15031693214253136
	pesos_i(324) := b"0000000000000000_0000000000000000_0000000101101010_0110100010101110"; -- 0.005529921053628277
	pesos_i(325) := b"0000000000000000_0000000000000000_0000000110010100_0111110100010110"; -- 0.006172006520847229
	pesos_i(326) := b"0000000000000000_0000000000000000_0000001010001001_0101000010100011"; -- 0.009907760493372724
	pesos_i(327) := b"0000000000000000_0000000000000000_0000100001001000_1101101101001100"; -- 0.03236170400634885
	pesos_i(328) := b"1111111111111111_1111111111111111_1111101011001101_1100011101000011"; -- -0.020297571356121046
	pesos_i(329) := b"1111111111111111_1111111111111111_1111011100001100_1101101100110000"; -- -0.034960079966835866
	pesos_i(330) := b"1111111111111111_1111111111111111_1111101111111110_0100110100011000"; -- -0.015650922424965418
	pesos_i(331) := b"0000000000000000_0000000000000000_0010000001011110_1111101011110011"; -- 0.12644928386338009
	pesos_i(332) := b"0000000000000000_0000000000000000_0000101010111010_1101001101101001"; -- 0.04191323584579137
	pesos_i(333) := b"0000000000000000_0000000000000000_0000101110011111_1100000101110100"; -- 0.04540642812997995
	pesos_i(334) := b"0000000000000000_0000000000000000_0000011100001110_1011101101101110"; -- 0.027568544775501892
	pesos_i(335) := b"1111111111111111_1111111111111111_1110001011010110_0111011101101000"; -- -0.11391500208973046
	pesos_i(336) := b"0000000000000000_0000000000000000_0000111111101010_0100111011110110"; -- 0.062169013019626324
	pesos_i(337) := b"0000000000000000_0000000000000000_0000001110010100_1110100110010001"; -- 0.013990972529227274
	pesos_i(338) := b"0000000000000000_0000000000000000_0000110101111011_0110100110110001"; -- 0.05266438084187584
	pesos_i(339) := b"1111111111111111_1111111111111111_1110101111010111_1111101100010110"; -- -0.07873564441363581
	pesos_i(340) := b"1111111111111111_1111111111111111_1101101100100101_0110100111111100"; -- -0.143960357714001
	pesos_i(341) := b"1111111111111111_1111111111111111_1110101001011000_0110101101111000"; -- -0.08458832096499368
	pesos_i(342) := b"0000000000000000_0000000000000000_0001000000000010_1011000110111111"; -- 0.06254111198085298
	pesos_i(343) := b"1111111111111111_1111111111111111_1101111010000011_1001100011100100"; -- -0.13080448554834845
	pesos_i(344) := b"1111111111111111_1111111111111111_1100100001101110_1101000000010011"; -- -0.21705913107492936
	pesos_i(345) := b"1111111111111111_1111111111111111_1111100101011001_0010001001111011"; -- -0.025983662480647474
	pesos_i(346) := b"0000000000000000_0000000000000000_0001000110100010_0011101101110111"; -- 0.06888171812643276
	pesos_i(347) := b"0000000000000000_0000000000000000_0000100010011010_0011010110000110"; -- 0.03360304364921644
	pesos_i(348) := b"0000000000000000_0000000000000000_0001001001111110_0000110101000001"; -- 0.07223589733106756
	pesos_i(349) := b"1111111111111111_1111111111111111_1111111111011100_1111111101110101"; -- -0.0005340898821312816
	pesos_i(350) := b"0000000000000000_0000000000000000_0000001101110100_1000110010100111"; -- 0.013497153028020084
	pesos_i(351) := b"0000000000000000_0000000000000000_0001100001011010_0100100110100001"; -- 0.09512767954182114
	pesos_i(352) := b"1111111111111111_1111111111111111_1110000111001000_0000000101010010"; -- -0.11804191345681825
	pesos_i(353) := b"0000000000000000_0000000000000000_0001111001010011_0000011001100101"; -- 0.11845436074934154
	pesos_i(354) := b"1111111111111111_1111111111111111_1101000100110001_0100101101011001"; -- -0.1828415783179143
	pesos_i(355) := b"1111111111111111_1111111111111111_1111000110000001_0101011010001010"; -- -0.05662020813235459
	pesos_i(356) := b"1111111111111111_1111111111111111_1110000001000011_1110100110000101"; -- -0.123963742272798
	pesos_i(357) := b"0000000000000000_0000000000000000_0001100000111001_1110100111011101"; -- 0.09463369033696759
	pesos_i(358) := b"1111111111111111_1111111111111111_1111101101110001_0001111111100110"; -- -0.017805105489237406
	pesos_i(359) := b"1111111111111111_1111111111111111_1111001100001110_0101100010010101"; -- -0.050562346940084685
	pesos_i(360) := b"1111111111111111_1111111111111111_1110111000001001_1111111010010100"; -- -0.07015999691143052
	pesos_i(361) := b"0000000000000000_0000000000000000_0001010001011000_0101011111100100"; -- 0.07947301204928169
	pesos_i(362) := b"1111111111111111_1111111111111111_1110001101111011_1100111000101110"; -- -0.11139212970688742
	pesos_i(363) := b"1111111111111111_1111111111111111_1101011100000001_1000000111100010"; -- -0.16013324967292342
	pesos_i(364) := b"1111111111111111_1111111111111111_1110110011100001_1100011000000110"; -- -0.07467996935240206
	pesos_i(365) := b"1111111111111111_1111111111111111_1110010001000111_0100000011000000"; -- -0.10828776647781718
	pesos_i(366) := b"0000000000000000_0000000000000000_0000000111001000_1000101100111010"; -- 0.0069663062973987985
	pesos_i(367) := b"1111111111111111_1111111111111111_1111110111101100_1011101000100000"; -- -0.008106581927993467
	pesos_i(368) := b"1111111111111111_1111111111111111_1111100011101110_0010100111000111"; -- -0.027615918020007207
	pesos_i(369) := b"0000000000000000_0000000000000000_0010110000101110_1000001101001010"; -- 0.1725847296554488
	pesos_i(370) := b"0000000000000000_0000000000000000_0010101011000001_1000111010000110"; -- 0.16701594131389574
	pesos_i(371) := b"0000000000000000_0000000000000000_0000110001100100_0011000100011011"; -- 0.04840380586342835
	pesos_i(372) := b"1111111111111111_1111111111111111_1110100101111100_0010011111010110"; -- -0.08794928585175649
	pesos_i(373) := b"1111111111111111_1111111111111111_1111001111110010_1111010000001000"; -- -0.04707407772231334
	pesos_i(374) := b"0000000000000000_0000000000000000_0001000010101100_1100001010111010"; -- 0.06513611839741702
	pesos_i(375) := b"0000000000000000_0000000000000000_0001100110111101_0000111111011001"; -- 0.10054110567830656
	pesos_i(376) := b"1111111111111111_1111111111111111_1110101001001110_1000101011000101"; -- -0.08473904311533784
	pesos_i(377) := b"1111111111111111_1111111111111111_1110010001000111_1010001011101110"; -- -0.10828191449519213
	pesos_i(378) := b"1111111111111111_1111111111111111_1110100101001001_1010101101100100"; -- -0.0887196427620318
	pesos_i(379) := b"1111111111111111_1111111111111111_1111010001001000_1110010111110000"; -- -0.04576266193529348
	pesos_i(380) := b"0000000000000000_0000000000000000_0001010111100100_1110010111111011"; -- 0.08552396191026229
	pesos_i(381) := b"0000000000000000_0000000000000000_0000111111110001_1110100011111101"; -- 0.0622850052944261
	pesos_i(382) := b"1111111111111111_1111111111111111_1110011000101010_0001111110011101"; -- -0.10091974655548533
	pesos_i(383) := b"1111111111111111_1111111111111111_1110110001001010_0001011100101110"; -- -0.07699446806079613
	pesos_i(384) := b"0000000000000000_0000000000000000_0000001100111110_0101110111001101"; -- 0.01267038591312264
	pesos_i(385) := b"0000000000000000_0000000000000000_0010000110010111_1011111000010010"; -- 0.13122165620740997
	pesos_i(386) := b"1111111111111111_1111111111111111_1110110101110110_1110101000110000"; -- -0.07240425431828539
	pesos_i(387) := b"0000000000000000_0000000000000000_0010100100101100_0000011111010101"; -- 0.16082810365971278
	pesos_i(388) := b"0000000000000000_0000000000000000_0000101110011101_0110100111011001"; -- 0.04537068878431376
	pesos_i(389) := b"1111111111111111_1111111111111111_1110101111000100_1010011001011101"; -- -0.07903061135436863
	pesos_i(390) := b"0000000000000000_0000000000000000_0010011010000010_0011101110100010"; -- 0.15042469692361843
	pesos_i(391) := b"1111111111111111_1111111111111111_1111000111111101_0110111001000111"; -- -0.05472670343241091
	pesos_i(392) := b"0000000000000000_0000000000000000_0000010010100101_0011110101100011"; -- 0.018146359103483677
	pesos_i(393) := b"0000000000000000_0000000000000000_0001110101110111_0111101001010000"; -- 0.11510433624543094
	pesos_i(394) := b"1111111111111111_1111111111111111_1101100000000011_1000100010110110"; -- -0.156196075048623
	pesos_i(395) := b"0000000000000000_0000000000000000_0010100010110110_0011101010111110"; -- 0.15903060099392913
	pesos_i(396) := b"0000000000000000_0000000000000000_0001010001000000_0000010010010110"; -- 0.07910183584908718
	pesos_i(397) := b"1111111111111111_1111111111111111_1101110001100000_1100011101100000"; -- -0.13914827262908117
	pesos_i(398) := b"1111111111111111_1111111111111111_1101111000100111_1000011010001011"; -- -0.13220938779149638
	pesos_i(399) := b"0000000000000000_0000000000000000_0010000011101100_1111110100110100"; -- 0.12861616619255772
	pesos_i(400) := b"1111111111111111_1111111111111111_1111101100111000_0101110100011111"; -- -0.018671207311157678
	pesos_i(401) := b"0000000000000000_0000000000000000_0000100001101000_0100001101001010"; -- 0.0328409248673109
	pesos_i(402) := b"1111111111111111_1111111111111111_1111100011111001_1001010011010000"; -- -0.027441691701444483
	pesos_i(403) := b"0000000000000000_0000000000000000_0010101001101110_1100110000001101"; -- 0.16575312915274887
	pesos_i(404) := b"0000000000000000_0000000000000000_0010001100100111_0110011001110011"; -- 0.13731994932045122
	pesos_i(405) := b"0000000000000000_0000000000000000_0001101101000001_0100011010010100"; -- 0.10646477810581183
	pesos_i(406) := b"1111111111111111_1111111111111111_1101100100101011_0001001010110101"; -- -0.15168650700537567
	pesos_i(407) := b"0000000000000000_0000000000000000_0000110110001011_1111100110001000"; -- 0.0529170947862537
	pesos_i(408) := b"1111111111111111_1111111111111111_1110100110100111_0111111011101000"; -- -0.08728796796021414
	pesos_i(409) := b"0000000000000000_0000000000000000_0000101110110111_0001111101110000"; -- 0.04576298213211745
	pesos_i(410) := b"0000000000000000_0000000000000000_0001010111100001_1100001110000011"; -- 0.08547613102627218
	pesos_i(411) := b"1111111111111111_1111111111111111_1101011111101001_1111000100000010"; -- -0.15658658690437252
	pesos_i(412) := b"1111111111111111_1111111111111111_1101100111011111_0001110010011110"; -- -0.1489393343656949
	pesos_i(413) := b"1111111111111111_1111111111111111_1110000100111011_1110000110101101"; -- -0.12018003022711304
	pesos_i(414) := b"1111111111111111_1111111111111111_1110011000110101_1111101001010111"; -- -0.10073886266434155
	pesos_i(415) := b"0000000000000000_0000000000000000_0010110010010000_1011011101000000"; -- 0.1740831881131836
	pesos_i(416) := b"0000000000000000_0000000000000000_0000100011010111_1011010000110001"; -- 0.03454137988011083
	pesos_i(417) := b"1111111111111111_1111111111111111_1111000101110100_1010100010000011"; -- -0.056813686464887506
	pesos_i(418) := b"0000000000000000_0000000000000000_0010100000111100_1011000100101000"; -- 0.1571760866168729
	pesos_i(419) := b"0000000000000000_0000000000000000_0001100110001100_0000010111001010"; -- 0.09979282541069469
	pesos_i(420) := b"1111111111111111_1111111111111111_1110010110001010_0100111111010100"; -- -0.10335827891612952
	pesos_i(421) := b"0000000000000000_0000000000000000_0001010110111111_1110001101110110"; -- 0.08495923637268968
	pesos_i(422) := b"0000000000000000_0000000000000000_0010011010111101_0000010010111100"; -- 0.15132169337723578
	pesos_i(423) := b"0000000000000000_0000000000000000_0001011011101001_0111110011101110"; -- 0.08950024432738687
	pesos_i(424) := b"1111111111111111_1111111111111111_1101100010111100_0001100011011110"; -- -0.15337986544368515
	pesos_i(425) := b"0000000000000000_0000000000000000_0000100101000100_0101010011001000"; -- 0.036198901036993456
	pesos_i(426) := b"1111111111111111_1111111111111111_1110101011011111_0010111110100000"; -- -0.08253195137657823
	pesos_i(427) := b"1111111111111111_1111111111111111_1110011101110101_1100100010010011"; -- -0.09585901644708528
	pesos_i(428) := b"1111111111111111_1111111111111111_1111111000011110_1101111010011000"; -- -0.0073414688068240445
	pesos_i(429) := b"1111111111111111_1111111111111111_1111111001100000_1111010111000011"; -- -0.006333007662983911
	pesos_i(430) := b"1111111111111111_1111111111111111_1111010101111100_0000010110000010"; -- -0.04107633184970902
	pesos_i(431) := b"0000000000000000_0000000000000000_0001000110001101_1100110101100010"; -- 0.0685699810295428
	pesos_i(432) := b"1111111111111111_1111111111111111_1110111011001011_0111000110011011"; -- -0.06720819440690433
	pesos_i(433) := b"1111111111111111_1111111111111111_1111100001010101_0110000100011001"; -- -0.029947215405014223
	pesos_i(434) := b"1111111111111111_1111111111111111_1111101111001001_0000011000010110"; -- -0.016463870645285587
	pesos_i(435) := b"0000000000000000_0000000000000000_0000110011000100_0111011111101010"; -- 0.049872870077835245
	pesos_i(436) := b"1111111111111111_1111111111111111_1101101001111110_0001011101100011"; -- -0.146513498613748
	pesos_i(437) := b"0000000000000000_0000000000000000_0000101011101111_1111011110110011"; -- 0.04272411453886019
	pesos_i(438) := b"1111111111111111_1111111111111111_1110011000000100_0101010111000110"; -- -0.10149635239394086
	pesos_i(439) := b"1111111111111111_1111111111111111_1110111011001010_0000010100000010"; -- -0.06722992618127474
	pesos_i(440) := b"0000000000000000_0000000000000000_0000011010110000_0010101101011001"; -- 0.026125630623397844
	pesos_i(441) := b"0000000000000000_0000000000000000_0000010110011100_1001111010111010"; -- 0.02192108199348413
	pesos_i(442) := b"1111111111111111_1111111111111111_1110110100100110_0001010010011000"; -- -0.0736376885646495
	pesos_i(443) := b"0000000000000000_0000000000000000_0001111001000101_1010010011110111"; -- 0.11825018907543443
	pesos_i(444) := b"1111111111111111_1111111111111111_1101001101100101_0001010010010111"; -- -0.17423888497296597
	pesos_i(445) := b"1111111111111111_1111111111111111_1111001100100100_0101001111001001"; -- -0.05022693972354388
	pesos_i(446) := b"1111111111111111_1111111111111111_1111110001110011_1001010001000000"; -- -0.01386140276433208
	pesos_i(447) := b"1111111111111111_1111111111111111_1110111101111001_0100100000000110"; -- -0.06455564355525148
	pesos_i(448) := b"1111111111111111_1111111111111111_1111110000010011_0011010010011100"; -- -0.01533194733677326
	pesos_i(449) := b"1111111111111111_1111111111111111_1110110010110110_1110101111110111"; -- -0.07533383568386882
	pesos_i(450) := b"1111111111111111_1111111111111111_1101101101010101_0101110011001110"; -- -0.14322872122390717
	pesos_i(451) := b"0000000000000000_0000000000000000_0000010101000110_1101100010111110"; -- 0.020612284190549782
	pesos_i(452) := b"0000000000000000_0000000000000000_0000100001111100_1001010001111010"; -- 0.03315093984647777
	pesos_i(453) := b"0000000000000000_0000000000000000_0010000110101010_1010000001011011"; -- 0.13150980216050778
	pesos_i(454) := b"1111111111111111_1111111111111111_1110011100101001_1100111010110011"; -- -0.09701831943489204
	pesos_i(455) := b"0000000000000000_0000000000000000_0010111011001101_1000000010101000"; -- 0.18282322027187392
	pesos_i(456) := b"1111111111111111_1111111111111111_1111011101101111_1111110101101001"; -- -0.03344742000092908
	pesos_i(457) := b"1111111111111111_1111111111111111_1111110010010111_0101101010101101"; -- -0.01331551824031108
	pesos_i(458) := b"0000000000000000_0000000000000000_0010010010000010_0101101000100001"; -- 0.1426140145695108
	pesos_i(459) := b"1111111111111111_1111111111111111_1101111011110101_0001101001100011"; -- -0.12907252398872107
	pesos_i(460) := b"0000000000000000_0000000000000000_0000110011111011_0000001010101001"; -- 0.05070511460926
	pesos_i(461) := b"0000000000000000_0000000000000000_0000000100111111_0111011001000101"; -- 0.004874603237548726
	pesos_i(462) := b"1111111111111111_1111111111111111_1111010000110000_0111000101101011"; -- -0.046135817939145396
	pesos_i(463) := b"0000000000000000_0000000000000000_0011000001111001_0110111000111101"; -- 0.18935288413707088
	pesos_i(464) := b"0000000000000000_0000000000000000_0000111000111101_0110101011011000"; -- 0.05562465456995347
	pesos_i(465) := b"1111111111111111_1111111111111111_1101111000110111_1111100011101100"; -- -0.13195842962949333
	pesos_i(466) := b"0000000000000000_0000000000000000_0010100001111001_1110110010110000"; -- 0.15811042109361104
	pesos_i(467) := b"0000000000000000_0000000000000000_0000000011011001_0110001000010000"; -- 0.003317002156014653
	pesos_i(468) := b"0000000000000000_0000000000000000_0010100010110111_0011000100000111"; -- 0.15904528075807214
	pesos_i(469) := b"1111111111111111_1111111111111111_1111010000010010_0111001100000101"; -- -0.04659348621230288
	pesos_i(470) := b"1111111111111111_1111111111111111_1101100110111011_1111101011010000"; -- -0.14947540685514707
	pesos_i(471) := b"1111111111111111_1111111111111111_1111010000101011_0111111111101100"; -- -0.0462112474469473
	pesos_i(472) := b"1111111111111111_1111111111111111_1110011111000100_1101000000110000"; -- -0.0946531183851616
	pesos_i(473) := b"1111111111111111_1111111111111111_1110110111101110_0011000100101101"; -- -0.07058422709553137
	pesos_i(474) := b"1111111111111111_1111111111111111_1111000100110001_1111010010110100"; -- -0.057831483857320475
	pesos_i(475) := b"0000000000000000_0000000000000000_0010101000111111_0110111011011101"; -- 0.1650304117737058
	pesos_i(476) := b"0000000000000000_0000000000000000_0000101000100001_1111011010111001"; -- 0.03958074586820405
	pesos_i(477) := b"0000000000000000_0000000000000000_0001001001111101_1101101100001101"; -- 0.07223290517168025
	pesos_i(478) := b"1111111111111111_1111111111111111_1110000101110111_0110111011000110"; -- -0.1192713514016224
	pesos_i(479) := b"0000000000000000_0000000000000000_0000001101011011_0010101110011111"; -- 0.013109899929091201
	pesos_i(480) := b"1111111111111111_1111111111111111_1111101101001010_1101000101100100"; -- -0.018389618863705187
	pesos_i(481) := b"0000000000000000_0000000000000000_0001001001011011_0010100001101000"; -- 0.07170345830326186
	pesos_i(482) := b"1111111111111111_1111111111111111_1101010110011010_0110101100101010"; -- -0.1656125089946691
	pesos_i(483) := b"1111111111111111_1111111111111111_1101011000010110_0011011100011000"; -- -0.16372352283612066
	pesos_i(484) := b"0000000000000000_0000000000000000_0000011011111001_0001001011111101"; -- 0.02723807031287583
	pesos_i(485) := b"0000000000000000_0000000000000000_0001110100001001_0011001100011110"; -- 0.11342162595075476
	pesos_i(486) := b"1111111111111111_1111111111111111_1101011110010100_1010001011101111"; -- -0.15788823765633492
	pesos_i(487) := b"1111111111111111_1111111111111111_1101011000010011_0010001000110101"; -- -0.16377054411563924
	pesos_i(488) := b"0000000000000000_0000000000000000_0000101011100011_1000101010100001"; -- 0.04253450797350533
	pesos_i(489) := b"0000000000000000_0000000000000000_0000110111001010_0111000001010101"; -- 0.053870220882675825
	pesos_i(490) := b"0000000000000000_0000000000000000_0000000001101100_1110001110001010"; -- 0.001661511670496053
	pesos_i(491) := b"1111111111111111_1111111111111111_1110000100101110_1010100011000011"; -- -0.1203817866813029
	pesos_i(492) := b"1111111111111111_1111111111111111_1110110010111000_0101011010001110"; -- -0.07531222372222846
	pesos_i(493) := b"0000000000000000_0000000000000000_0001100001011100_1010000001000001"; -- 0.095163360367006
	pesos_i(494) := b"0000000000000000_0000000000000000_0000010101111110_1001101110000101"; -- 0.02146312699829045
	pesos_i(495) := b"0000000000000000_0000000000000000_0001111110100001_1001010110110011"; -- 0.12355933784023215
	pesos_i(496) := b"1111111111111111_1111111111111111_1101110111111010_1101010001101111"; -- -0.132891390798526
	pesos_i(497) := b"1111111111111111_1111111111111111_1110000010110100_0011110100100111"; -- -0.12224977291323824
	pesos_i(498) := b"1111111111111111_1111111111111111_1101101001001110_1100000101111011"; -- -0.1472357821514689
	pesos_i(499) := b"0000000000000000_0000000000000000_0001010110010010_1000000011101010"; -- 0.08426671714617524
	pesos_i(500) := b"1111111111111111_1111111111111111_1101100101111001_1010111111100111"; -- -0.15048695196146133
	pesos_i(501) := b"1111111111111111_1111111111111111_1110100000000110_0011110010101001"; -- -0.09365483160440766
	pesos_i(502) := b"0000000000000000_0000000000000000_0010000011110111_1110001101111000"; -- 0.12878247910432644
	pesos_i(503) := b"1111111111111111_1111111111111111_1110011111111111_0010101011100101"; -- -0.09376270203718139
	pesos_i(504) := b"0000000000000000_0000000000000000_0010001001110101_1101110001000101"; -- 0.1346109075063381
	pesos_i(505) := b"1111111111111111_1111111111111111_1110110101011100_0101011111000110"; -- -0.07280970964551217
	pesos_i(506) := b"1111111111111111_1111111111111111_1110111101010110_1110001111001010"; -- -0.06508041678643696
	pesos_i(507) := b"1111111111111111_1111111111111111_1111110001001011_0111011011111010"; -- -0.014473499353162046
	pesos_i(508) := b"1111111111111111_1111111111111111_1101100100010100_0010001010010001"; -- -0.1520365139865774
	pesos_i(509) := b"1111111111111111_1111111111111111_1111000000110011_1100001011001111"; -- -0.061710190358504134
	pesos_i(510) := b"1111111111111111_1111111111111111_1101100101001000_0011010110000110"; -- -0.1512419268286145
	pesos_i(511) := b"1111111111111111_1111111111111111_1111011010000111_0100010110001000"; -- -0.03699841909315402
	pesos_i(512) := b"0000000000000000_0000000000000000_0000000001010111_0001100100101010"; -- 0.0013290144374279167
	pesos_i(513) := b"1111111111111111_1111111111111111_1111010100001101_0111100100001001"; -- -0.042763171388989316
	pesos_i(514) := b"1111111111111111_1111111111111111_1110110010010011_1010101100111000"; -- -0.07587175252424407
	pesos_i(515) := b"1111111111111111_1111111111111111_1110111110000010_0100011101011100"; -- -0.06441835396030934
	pesos_i(516) := b"0000000000000000_0000000000000000_0010101111010110_0111001111001110"; -- 0.17124103324298492
	pesos_i(517) := b"1111111111111111_1111111111111111_1110100111011101_0101000011110101"; -- -0.08646673221716226
	pesos_i(518) := b"0000000000000000_0000000000000000_0000010010001111_1010011011011110"; -- 0.017816952803078826
	pesos_i(519) := b"0000000000000000_0000000000000000_0010000110101011_1000010000111110"; -- 0.13152338520349358
	pesos_i(520) := b"1111111111111111_1111111111111111_1111110111110010_1000001000100100"; -- -0.008018365965286024
	pesos_i(521) := b"1111111111111111_1111111111111111_1111100100110111_1011110101001001"; -- -0.02649323438595049
	pesos_i(522) := b"1111111111111111_1111111111111111_1110111111100000_0011111000100010"; -- -0.06298457795789515
	pesos_i(523) := b"1111111111111111_1111111111111111_1110000000011000_0111000010000100"; -- -0.12462708259253737
	pesos_i(524) := b"0000000000000000_0000000000000000_0001000000111111_0111100101010001"; -- 0.06346853483735126
	pesos_i(525) := b"1111111111111111_1111111111111111_1111101001101110_1100001010000011"; -- -0.02174743940495029
	pesos_i(526) := b"1111111111111111_1111111111111111_1111000100000110_0101110100111010"; -- -0.05849664053196309
	pesos_i(527) := b"1111111111111111_1111111111111111_1101110110101011_1010000010110101"; -- -0.13409991818247474
	pesos_i(528) := b"1111111111111111_1111111111111111_1111111101111100_0101110110111011"; -- -0.002008573437284389
	pesos_i(529) := b"0000000000000000_0000000000000000_0001001010110001_1110110000011111"; -- 0.0730273796689701
	pesos_i(530) := b"1111111111111111_1111111111111111_1101111000110000_0000000111010000"; -- -0.13207997003484961
	pesos_i(531) := b"0000000000000000_0000000000000000_0000011010001001_0001010101101001"; -- 0.02552923025929379
	pesos_i(532) := b"1111111111111111_1111111111111111_1101101000101100_1011111101110011"; -- -0.1477547020847112
	pesos_i(533) := b"0000000000000000_0000000000000000_0010011010110111_0100110011000110"; -- 0.1512344344247598
	pesos_i(534) := b"0000000000000000_0000000000000000_0010011000001010_0011100001010000"; -- 0.1485934444576774
	pesos_i(535) := b"0000000000000000_0000000000000000_0001000001010100_0001110001011110"; -- 0.06378342905885094
	pesos_i(536) := b"1111111111111111_1111111111111111_1110100111001011_1111101110100110"; -- -0.08673121632425862
	pesos_i(537) := b"0000000000000000_0000000000000000_0000101001101011_1011101000111110"; -- 0.040706291316836375
	pesos_i(538) := b"1111111111111111_1111111111111111_1110111010111011_0010111100111000"; -- -0.06745629187221723
	pesos_i(539) := b"1111111111111111_1111111111111111_1111110001110011_0111110000010101"; -- -0.013862843505927838
	pesos_i(540) := b"1111111111111111_1111111111111111_1110000000110101_1000110010000000"; -- -0.1241829098406435
	pesos_i(541) := b"1111111111111111_1111111111111111_1111010010111010_1110001101100111"; -- -0.04402331090227748
	pesos_i(542) := b"0000000000000000_0000000000000000_0010100110011011_1101011101010001"; -- 0.16253419625678614
	pesos_i(543) := b"1111111111111111_1111111111111111_1111011110111010_1011111110110101"; -- -0.03230668861794206
	pesos_i(544) := b"1111111111111111_1111111111111111_1111111101110101_0000011000110100"; -- -0.002120601959403695
	pesos_i(545) := b"0000000000000000_0000000000000000_0000010001001000_1011111111011111"; -- 0.01673506923245809
	pesos_i(546) := b"1111111111111111_1111111111111111_1111111100111000_1010100110000100"; -- -0.0030416537892086733
	pesos_i(547) := b"1111111111111111_1111111111111111_1111101101100111_0100001111100011"; -- -0.017955548289636337
	pesos_i(548) := b"0000000000000000_0000000000000000_0010010010101110_0111010110000011"; -- 0.14328703363566345
	pesos_i(549) := b"0000000000000000_0000000000000000_0001010110000111_1101000001011111"; -- 0.08410360643226465
	pesos_i(550) := b"0000000000000000_0000000000000000_0001111100101100_0100001011000111"; -- 0.12176911703452688
	pesos_i(551) := b"0000000000000000_0000000000000000_0001000111111101_1000111101110001"; -- 0.0702752734990913
	pesos_i(552) := b"1111111111111111_1111111111111111_1111001001101110_1111001010011000"; -- -0.05299457359047541
	pesos_i(553) := b"0000000000000000_0000000000000000_0001011001011101_1101001111110101"; -- 0.08736920099335131
	pesos_i(554) := b"1111111111111111_1111111111111111_1101111100010011_0010111011010111"; -- -0.1286135411854639
	pesos_i(555) := b"1111111111111111_1111111111111111_1111000000000001_0111000100001011"; -- -0.062478003391997924
	pesos_i(556) := b"1111111111111111_1111111111111111_1111100101000000_1011111100110101"; -- -0.02635579067868956
	pesos_i(557) := b"0000000000000000_0000000000000000_0000110101010011_1001000000111111"; -- 0.052056327249324755
	pesos_i(558) := b"1111111111111111_1111111111111111_1110001100101010_0010010110101100"; -- -0.11263813549885032
	pesos_i(559) := b"1111111111111111_1111111111111111_1111011101011011_0101000100101111"; -- -0.03376286133690925
	pesos_i(560) := b"1111111111111111_1111111111111111_1101010110000010_1000101000011110"; -- -0.16597687488036414
	pesos_i(561) := b"0000000000000000_0000000000000000_0000000111100010_1010010111010010"; -- 0.007364620025200559
	pesos_i(562) := b"0000000000000000_0000000000000000_0001110001000111_1000100011001001"; -- 0.11046652699942044
	pesos_i(563) := b"1111111111111111_1111111111111111_1110001000100010_0000001011000110"; -- -0.11666853592366255
	pesos_i(564) := b"1111111111111111_1111111111111111_1111100111011110_1001110000110110"; -- -0.02394698803871375
	pesos_i(565) := b"1111111111111111_1111111111111111_1111001000010001_0001001010101000"; -- -0.05442698857521127
	pesos_i(566) := b"1111111111111111_1111111111111111_1111110111111101_1100111010010100"; -- -0.007845963388397957
	pesos_i(567) := b"1111111111111111_1111111111111111_1110010010100110_0000011010000111"; -- -0.10684165199152586
	pesos_i(568) := b"1111111111111111_1111111111111111_1101010101101110_0011001100100110"; -- -0.16628723441346
	pesos_i(569) := b"0000000000000000_0000000000000000_0000001100001000_0010001000110101"; -- 0.0118428592315597
	pesos_i(570) := b"1111111111111111_1111111111111111_1110111110000000_0110111011000000"; -- -0.06444652385106316
	pesos_i(571) := b"1111111111111111_1111111111111111_1111101111000110_0001110001011001"; -- -0.016508320172470003
	pesos_i(572) := b"1111111111111111_1111111111111111_1110011110000101_0010010010110111"; -- -0.09562464262810048
	pesos_i(573) := b"0000000000000000_0000000000000000_0001100001011011_1110011011011000"; -- 0.09515230923690285
	pesos_i(574) := b"1111111111111111_1111111111111111_1110010010110100_1000011001111111"; -- -0.1066204013710376
	pesos_i(575) := b"0000000000000000_0000000000000000_0000101100001001_0001111001001010"; -- 0.04310788442796491
	pesos_i(576) := b"1111111111111111_1111111111111111_1111011001010101_1101001111110001"; -- -0.03775287033654967
	pesos_i(577) := b"1111111111111111_1111111111111111_1101100000100111_0011101101000011"; -- -0.1556513749234236
	pesos_i(578) := b"0000000000000000_0000000000000000_0000010001110001_1011011111101100"; -- 0.017360205839113196
	pesos_i(579) := b"1111111111111111_1111111111111111_1101011000000110_1111010111001100"; -- -0.1639562965925202
	pesos_i(580) := b"0000000000000000_0000000000000000_0001101000010100_1000011110001011"; -- 0.10187575473360869
	pesos_i(581) := b"0000000000000000_0000000000000000_0001110110110101_1011001110100011"; -- 0.11605379794059088
	pesos_i(582) := b"0000000000000000_0000000000000000_0000100000000011_0111011111100011"; -- 0.03130292205750122
	pesos_i(583) := b"1111111111111111_1111111111111111_1101001000001101_0010000110110001"; -- -0.17948712760633886
	pesos_i(584) := b"0000000000000000_0000000000000000_0010101110101010_1101001101111010"; -- 0.1705753491628184
	pesos_i(585) := b"0000000000000000_0000000000000000_0010010110011000_1001011011010111"; -- 0.14685957662846028
	pesos_i(586) := b"1111111111111111_1111111111111111_1111000110101100_1010010010100111"; -- -0.055959424277333
	pesos_i(587) := b"0000000000000000_0000000000000000_0000110110111111_1110101101000101"; -- 0.053709701791982804
	pesos_i(588) := b"1111111111111111_1111111111111111_1111111001010100_1011111101110110"; -- -0.006519349777997984
	pesos_i(589) := b"0000000000000000_0000000000000000_0001000001001011_0011110001010110"; -- 0.06364800540619119
	pesos_i(590) := b"0000000000000000_0000000000000000_0001101100110100_1000001001110100"; -- 0.1062699827309407
	pesos_i(591) := b"0000000000000000_0000000000000000_0010011100111010_0110110011001110"; -- 0.15323524500933794
	pesos_i(592) := b"1111111111111111_1111111111111111_1101110101010001_1010111000000001"; -- -0.1354724166562596
	pesos_i(593) := b"0000000000000000_0000000000000000_0001000110010100_0100001111111111"; -- 0.06866860366377359
	pesos_i(594) := b"0000000000000000_0000000000000000_0010001011011000_1101011000011010"; -- 0.13612115978578457
	pesos_i(595) := b"1111111111111111_1111111111111111_1110011010101110_1011110010101110"; -- -0.09889622460124779
	pesos_i(596) := b"0000000000000000_0000000000000000_0001001011101001_1100001100001111"; -- 0.07387942416520815
	pesos_i(597) := b"0000000000000000_0000000000000000_0000000111101101_0001110001000010"; -- 0.007524267316898777
	pesos_i(598) := b"0000000000000000_0000000000000000_0010001000101000_0000010001000000"; -- 0.13342310491625864
	pesos_i(599) := b"0000000000000000_0000000000000000_0000010000010000_1111001110001010"; -- 0.015883656789655663
	pesos_i(600) := b"1111111111111111_1111111111111111_1111011001000001_1000010110100100"; -- -0.03806271305945191
	pesos_i(601) := b"1111111111111111_1111111111111111_1101001011100111_1101011110111110"; -- -0.1761498603995838
	pesos_i(602) := b"0000000000000000_0000000000000000_0001100111000011_0000011100011100"; -- 0.10063213758848301
	pesos_i(603) := b"1111111111111111_1111111111111111_1111110011011011_0010000001100101"; -- -0.012281394215930141
	pesos_i(604) := b"0000000000000000_0000000000000000_0000001010001010_1101100010010001"; -- 0.009931121336491173
	pesos_i(605) := b"0000000000000000_0000000000000000_0001000011101101_1111101101001001"; -- 0.06613131070602965
	pesos_i(606) := b"0000000000000000_0000000000000000_0001010111000000_1011100010010101"; -- 0.08497193950443362
	pesos_i(607) := b"0000000000000000_0000000000000000_0001010110010011_0101110101111000"; -- 0.08427986323927986
	pesos_i(608) := b"1111111111111111_1111111111111111_1110100010010010_1111000111010011"; -- -0.09150780290760546
	pesos_i(609) := b"0000000000000000_0000000000000000_0001110111011111_0001100110010011"; -- 0.11668548433804532
	pesos_i(610) := b"0000000000000000_0000000000000000_0000101000100111_1001110101010001"; -- 0.039666969446875845
	pesos_i(611) := b"1111111111111111_1111111111111111_1110100110000111_1111001100101010"; -- -0.08776931974826833
	pesos_i(612) := b"0000000000000000_0000000000000000_0001000101100000_0000111110100101"; -- 0.06787202614316251
	pesos_i(613) := b"0000000000000000_0000000000000000_0000101000010001_1001100010000111"; -- 0.03933099074718706
	pesos_i(614) := b"1111111111111111_1111111111111111_1111100010110100_0001100111010011"; -- -0.028501878774738493
	pesos_i(615) := b"1111111111111111_1111111111111111_1101001100010110_1111000100111011"; -- -0.17543117809849576
	pesos_i(616) := b"1111111111111111_1111111111111111_1111001100111100_0111011111000001"; -- -0.049858584751122065
	pesos_i(617) := b"1111111111111111_1111111111111111_1101001101011001_0000100111110110"; -- -0.17442262416728013
	pesos_i(618) := b"1111111111111111_1111111111111111_1111111101100111_0100101010001010"; -- -0.00233015182587026
	pesos_i(619) := b"0000000000000000_0000000000000000_0001010101111001_0110101100010001"; -- 0.08388394512490488
	pesos_i(620) := b"1111111111111111_1111111111111111_1101100111010000_1100011100001010"; -- -0.14915805826027542
	pesos_i(621) := b"0000000000000000_0000000000000000_0000100011011001_0000101001110110"; -- 0.03456178084736198
	pesos_i(622) := b"1111111111111111_1111111111111111_1110011101010000_1110110111001001"; -- -0.09642137383307403
	pesos_i(623) := b"0000000000000000_0000000000000000_0010000010101100_0001110011111011"; -- 0.1276262390985352
	pesos_i(624) := b"1111111111111111_1111111111111111_1101100010110100_1100001100001111"; -- -0.15349179152769415
	pesos_i(625) := b"0000000000000000_0000000000000000_0001011111101110_0000100010111010"; -- 0.09347586190192606
	pesos_i(626) := b"1111111111111111_1111111111111111_1111001100011000_1010111000111100"; -- -0.05040465389581916
	pesos_i(627) := b"0000000000000000_0000000000000000_0001010000000101_0101001000111001"; -- 0.07820619474670903
	pesos_i(628) := b"0000000000000000_0000000000000000_0001000001110110_1111010110000100"; -- 0.06431517088043665
	pesos_i(629) := b"1111111111111111_1111111111111111_1101101000000011_0101000001010111"; -- -0.14838693491749158
	pesos_i(630) := b"1111111111111111_1111111111111111_1111100001111001_1001011011100011"; -- -0.02939469299482397
	pesos_i(631) := b"1111111111111111_1111111111111111_1110110110111111_0000010101011111"; -- -0.07130400115474445
	pesos_i(632) := b"0000000000000000_0000000000000000_0001010110110001_1010101110011001"; -- 0.08474228357066313
	pesos_i(633) := b"1111111111111111_1111111111111111_1111000001111000_0011101100111110"; -- -0.06066541409070134
	pesos_i(634) := b"0000000000000000_0000000000000000_0001000010111001_1010011011100001"; -- 0.06533282283662055
	pesos_i(635) := b"0000000000000000_0000000000000000_0001011001101111_0001111001111001"; -- 0.08763304180180712
	pesos_i(636) := b"0000000000000000_0000000000000000_0010100100100001_0001001010100001"; -- 0.1606609004156315
	pesos_i(637) := b"1111111111111111_1111111111111111_1110001100011001_0111001010000111"; -- -0.11289295388655776
	pesos_i(638) := b"0000000000000000_0000000000000000_0000000001110110_1001110110000110"; -- 0.0018099263258727742
	pesos_i(639) := b"0000000000000000_0000000000000000_0000110111001111_1001101001010100"; -- 0.053949017926418284
	pesos_i(640) := b"0000000000000000_0000000000000000_0001011010010110_1110100000101110"; -- 0.08824015739403054
	pesos_i(641) := b"0000000000000000_0000000000000000_0000010011100010_0011101111001100"; -- 0.019077050532061744
	pesos_i(642) := b"1111111111111111_1111111111111111_1101110001000001_1101110011010110"; -- -0.1396200158930832
	pesos_i(643) := b"0000000000000000_0000000000000000_0001110010101011_1000100100111111"; -- 0.11199243333726844
	pesos_i(644) := b"1111111111111111_1111111111111111_1111011111100011_1111011101110101"; -- -0.03167775527664038
	pesos_i(645) := b"0000000000000000_0000000000000000_0000100010011100_1000010000100001"; -- 0.03363824655656167
	pesos_i(646) := b"0000000000000000_0000000000000000_0000000100101010_0101111100010111"; -- 0.004552786855949614
	pesos_i(647) := b"0000000000000000_0000000000000000_0001001001011011_1100100001010000"; -- 0.07171298928842226
	pesos_i(648) := b"0000000000000000_0000000000000000_0000000001010000_0100011011010100"; -- 0.0012249248673728904
	pesos_i(649) := b"1111111111111111_1111111111111111_1101001010001100_1011000010100110"; -- -0.17754074043478102
	pesos_i(650) := b"1111111111111111_1111111111111111_1111000010011001_0010111101100011"; -- -0.06016258088891046
	pesos_i(651) := b"0000000000000000_0000000000000000_0010010011110001_1011111000110101"; -- 0.14431370537461788
	pesos_i(652) := b"1111111111111111_1111111111111111_1110101010101101_0000111111001101"; -- -0.08329678772507333
	pesos_i(653) := b"0000000000000000_0000000000000000_0010001000000101_1000101111100000"; -- 0.13289713110849832
	pesos_i(654) := b"1111111111111111_1111111111111111_1110110110100010_0111100011100110"; -- -0.07173962004649183
	pesos_i(655) := b"1111111111111111_1111111111111111_1101000010110111_0101011111110101"; -- -0.18470239904289049
	pesos_i(656) := b"0000000000000000_0000000000000000_0001101011000000_1001010010110110"; -- 0.10450105135655804
	pesos_i(657) := b"0000000000000000_0000000000000000_0000000101101001_0011101001010100"; -- 0.005511899491295283
	pesos_i(658) := b"1111111111111111_1111111111111111_1111100010100001_1011111111001011"; -- -0.02878190312722175
	pesos_i(659) := b"1111111111111111_1111111111111111_1110101010000110_1101010011110011"; -- -0.08388012954366404
	pesos_i(660) := b"1111111111111111_1111111111111111_1111100101111101_0001000110001111"; -- -0.025435354865724763
	pesos_i(661) := b"1111111111111111_1111111111111111_1111000111010011_1111110011100100"; -- -0.055359072078673806
	pesos_i(662) := b"0000000000000000_0000000000000000_0000000101101111_1010111000111001"; -- 0.005610359981518082
	pesos_i(663) := b"1111111111111111_1111111111111111_1111110000110111_0001001100101001"; -- -0.014784624561879471
	pesos_i(664) := b"0000000000000000_0000000000000000_0000111000000100_1001000100011011"; -- 0.05475718407655232
	pesos_i(665) := b"0000000000000000_0000000000000000_0000101010010001_1111111110010101"; -- 0.041290258296140206
	pesos_i(666) := b"1111111111111111_1111111111111111_1110011111101101_1100000101000100"; -- -0.09402839736364377
	pesos_i(667) := b"0000000000000000_0000000000000000_0001001011111011_1011111010001111"; -- 0.07415381427970177
	pesos_i(668) := b"1111111111111111_1111111111111111_1110100110011110_0111110110100101"; -- -0.08742537228104925
	pesos_i(669) := b"0000000000000000_0000000000000000_0001101110000001_1110010110101010"; -- 0.10745082286904252
	pesos_i(670) := b"0000000000000000_0000000000000000_0000001101101010_1010011010011001"; -- 0.013346111587319482
	pesos_i(671) := b"0000000000000000_0000000000000000_0000111100010001_1100101101100110"; -- 0.058865272929847307
	pesos_i(672) := b"1111111111111111_1111111111111111_1101110100100100_0011111001011111"; -- -0.13616571602512711
	pesos_i(673) := b"1111111111111111_1111111111111111_1110111100001111_0101011001110100"; -- -0.06617221504164002
	pesos_i(674) := b"0000000000000000_0000000000000000_0000010110001110_0011010000000010"; -- 0.021701097869629007
	pesos_i(675) := b"0000000000000000_0000000000000000_0000000000010111_1111100011111111"; -- 0.00036579350526725165
	pesos_i(676) := b"1111111111111111_1111111111111111_1110100000110100_1110110100010001"; -- -0.09294241272820408
	pesos_i(677) := b"1111111111111111_1111111111111111_1111110101101100_0101111101100010"; -- -0.010065115542706893
	pesos_i(678) := b"0000000000000000_0000000000000000_0001100011101001_1000001000011100"; -- 0.09731305304140818
	pesos_i(679) := b"0000000000000000_0000000000000000_0010100101010111_0100000001001010"; -- 0.16148759667644383
	pesos_i(680) := b"0000000000000000_0000000000000000_0010010111010001_1111001111110111"; -- 0.14773487826168832
	pesos_i(681) := b"0000000000000000_0000000000000000_0010100101100001_1011101101010111"; -- 0.16164751880962738
	pesos_i(682) := b"0000000000000000_0000000000000000_0001011001100010_1000111100101000"; -- 0.08744139402296933
	pesos_i(683) := b"1111111111111111_1111111111111111_1101001100010000_1111110010010001"; -- -0.17552205523345837
	pesos_i(684) := b"0000000000000000_0000000000000000_0001110111101011_1101101011001110"; -- 0.11688010711053684
	pesos_i(685) := b"0000000000000000_0000000000000000_0010100001010111_0010110101111010"; -- 0.1575802253786452
	pesos_i(686) := b"0000000000000000_0000000000000000_0001001000000011_0010110101001011"; -- 0.07036097612285032
	pesos_i(687) := b"1111111111111111_1111111111111111_1111011110010110_0001100011010001"; -- -0.03286595255082978
	pesos_i(688) := b"1111111111111111_1111111111111111_1110100111111010_0111001101001001"; -- -0.08602218115714079
	pesos_i(689) := b"0000000000000000_0000000000000000_0010111000010001_0111001000110001"; -- 0.1799537058454888
	pesos_i(690) := b"1111111111111111_1111111111111111_1101110111001101_1001010101111101"; -- -0.13358178796101294
	pesos_i(691) := b"1111111111111111_1111111111111111_1111011011011101_0001010001110110"; -- -0.03568908808043661
	pesos_i(692) := b"0000000000000000_0000000000000000_0010011011000110_0001100111111101"; -- 0.1514602892934048
	pesos_i(693) := b"0000000000000000_0000000000000000_0001000101100111_1011000100101111"; -- 0.06798846621101973
	pesos_i(694) := b"0000000000000000_0000000000000000_0001001110000100_0111010100100111"; -- 0.07623989290573803
	pesos_i(695) := b"0000000000000000_0000000000000000_0010100001010010_0000101001000101"; -- 0.1575018329074574
	pesos_i(696) := b"1111111111111111_1111111111111111_1101101010110011_0010110001100001"; -- -0.14570353160486801
	pesos_i(697) := b"1111111111111111_1111111111111111_1100110110101011_0010110110010100"; -- -0.19660678049803448
	pesos_i(698) := b"0000000000000000_0000000000000000_0001111110111001_1010111001010000"; -- 0.12392701577561205
	pesos_i(699) := b"1111111111111111_1111111111111111_1101010101011001_1000100110100011"; -- -0.1666025140444962
	pesos_i(700) := b"1111111111111111_1111111111111111_1110101111010111_1111000010110110"; -- -0.07873626283475374
	pesos_i(701) := b"1111111111111111_1111111111111111_1111110011111001_1010110110001000"; -- -0.011815218301188198
	pesos_i(702) := b"1111111111111111_1111111111111111_1110011100010010_0110011111110111"; -- -0.09737539497893369
	pesos_i(703) := b"1111111111111111_1111111111111111_1111001000001001_1010111001010111"; -- -0.05453977949685018
	pesos_i(704) := b"1111111111111111_1111111111111111_1101010010111110_1100101111110110"; -- -0.16896367297292353
	pesos_i(705) := b"0000000000000000_0000000000000000_0001101101010011_0001110011011111"; -- 0.10673695042078116
	pesos_i(706) := b"1111111111111111_1111111111111111_1110001101010111_1110000001010101"; -- -0.11194036420749337
	pesos_i(707) := b"1111111111111111_1111111111111111_1111110110011011_0111000011010101"; -- -0.00934691236608223
	pesos_i(708) := b"1111111111111111_1111111111111111_1111011111010010_0001010011000011"; -- -0.03195066677217223
	pesos_i(709) := b"0000000000000000_0000000000000000_0000100111011000_0101110000001010"; -- 0.03845763436057793
	pesos_i(710) := b"0000000000000000_0000000000000000_0001001110101001_0000001101101001"; -- 0.07679768852792963
	pesos_i(711) := b"0000000000000000_0000000000000000_0001111010001100_0100101011110010"; -- 0.11932819766289479
	pesos_i(712) := b"1111111111111111_1111111111111111_1101101000101010_1110111000111011"; -- -0.14778243120492376
	pesos_i(713) := b"1111111111111111_1111111111111111_1110001111011001_1111011000100001"; -- -0.10995542232952782
	pesos_i(714) := b"1111111111111111_1111111111111111_1101101110100010_1000010000101111"; -- -0.1420514473389469
	pesos_i(715) := b"1111111111111111_1111111111111111_1111100010001010_0010011011011001"; -- -0.029141971541423693
	pesos_i(716) := b"1111111111111111_1111111111111111_1111011001011000_1111011100101000"; -- -0.03770499499643162
	pesos_i(717) := b"1111111111111111_1111111111111111_1110000100101000_1101110110110010"; -- -0.1204701844371957
	pesos_i(718) := b"0000000000000000_0000000000000000_0010010101111100_0111001110000111"; -- 0.1464302258304404
	pesos_i(719) := b"0000000000000000_0000000000000000_0001000101111010_1110010110001001"; -- 0.0682815037241553
	pesos_i(720) := b"0000000000000000_0000000000000000_0001111111101011_1011101101001111"; -- 0.12469072986772786
	pesos_i(721) := b"0000000000000000_0000000000000000_0000000010110110_1101101110101001"; -- 0.0027901924828218623
	pesos_i(722) := b"0000000000000000_0000000000000000_0000111100110001_0111110001011011"; -- 0.05934884286156734
	pesos_i(723) := b"1111111111111111_1111111111111111_1101010001000000_1100000010100111"; -- -0.17088695457095548
	pesos_i(724) := b"0000000000000000_0000000000000000_0000110010101101_0010010110001000"; -- 0.04951700762876007
	pesos_i(725) := b"0000000000000000_0000000000000000_0001011010100100_0001111001010000"; -- 0.08844174822252306
	pesos_i(726) := b"0000000000000000_0000000000000000_0010001000110110_1111111111001001"; -- 0.1336517207081711
	pesos_i(727) := b"0000000000000000_0000000000000000_0010000011001111_0111001111001011"; -- 0.12816547109598334
	pesos_i(728) := b"1111111111111111_1111111111111111_1111100101111111_1011110000001101"; -- -0.025394675102071957
	pesos_i(729) := b"1111111111111111_1111111111111111_1101110111100000_1001101000111100"; -- -0.13329158811250222
	pesos_i(730) := b"0000000000000000_0000000000000000_0010011111001011_1101011100000100"; -- 0.15545410018047495
	pesos_i(731) := b"1111111111111111_1111111111111111_1111001011011110_0111101111101000"; -- -0.05129266344070909
	pesos_i(732) := b"0000000000000000_0000000000000000_0010010111001111_1110010110010011"; -- 0.14770350298284177
	pesos_i(733) := b"0000000000000000_0000000000000000_0000000011011101_0000000001011110"; -- 0.003372214341333454
	pesos_i(734) := b"1111111111111111_1111111111111111_1111001101000001_1101000000101110"; -- -0.04977702027626591
	pesos_i(735) := b"0000000000000000_0000000000000000_0000110111110100_0010011001111011"; -- 0.05450668824862842
	pesos_i(736) := b"1111111111111111_1111111111111111_1101100111100101_0010000000000010"; -- -0.1488475794060196
	pesos_i(737) := b"1111111111111111_1111111111111111_1110000010110101_0100010010001111"; -- -0.12223407274617638
	pesos_i(738) := b"1111111111111111_1111111111111111_1101100110110001_1000101101111111"; -- -0.14963462971190558
	pesos_i(739) := b"1111111111111111_1111111111111111_1111100001001000_1110001011000011"; -- -0.03013785105300284
	pesos_i(740) := b"1111111111111111_1111111111111111_1110010101110000_0111001011010000"; -- -0.10375292221580915
	pesos_i(741) := b"1111111111111111_1111111111111111_1101101001000000_0110101111100100"; -- -0.1474545067440846
	pesos_i(742) := b"1111111111111111_1111111111111111_1101010000100000_0000101110110001"; -- -0.17138602193471036
	pesos_i(743) := b"1111111111111111_1111111111111111_1110001001100111_0111011100110101"; -- -0.11560873934920513
	pesos_i(744) := b"1111111111111111_1111111111111111_1111001010111110_0001110110100010"; -- -0.05178656372923439
	pesos_i(745) := b"0000000000000000_0000000000000000_0010010001101110_1001100100100111"; -- 0.14231259539972077
	pesos_i(746) := b"0000000000000000_0000000000000000_0000110001100101_0001111001110110"; -- 0.04841795332878018
	pesos_i(747) := b"0000000000000000_0000000000000000_0010000011000000_0001011000101010"; -- 0.1279310085879287
	pesos_i(748) := b"0000000000000000_0000000000000000_0000110001101101_1101001011010011"; -- 0.04855077412336125
	pesos_i(749) := b"1111111111111111_1111111111111111_1111111110101000_1100100101111010"; -- -0.0013307644584613473
	pesos_i(750) := b"0000000000000000_0000000000000000_0010001100000110_0111001100001100"; -- 0.13681716005238914
	pesos_i(751) := b"0000000000000000_0000000000000000_0010011001011101_0001000011101001"; -- 0.14985757522137105
	pesos_i(752) := b"1111111111111111_1111111111111111_1111010010010111_0111100101010001"; -- -0.0445636917510705
	pesos_i(753) := b"1111111111111111_1111111111111111_1101001001011001_1001100111001101"; -- -0.17832030049792483
	pesos_i(754) := b"0000000000000000_0000000000000000_0000011010111000_1111101010010100"; -- 0.026260052910086065
	pesos_i(755) := b"0000000000000000_0000000000000000_0001000111100110_0100110101111001"; -- 0.06992038928178243
	pesos_i(756) := b"1111111111111111_1111111111111111_1110000001101111_1001101100000111"; -- -0.12329703398947679
	pesos_i(757) := b"1111111111111111_1111111111111111_1111110011101000_1010111011011001"; -- -0.012074539300097605
	pesos_i(758) := b"0000000000000000_0000000000000000_0010100010000110_0001100110111010"; -- 0.15829621121047616
	pesos_i(759) := b"0000000000000000_0000000000000000_0000110011001101_0111100101101001"; -- 0.05001028848285987
	pesos_i(760) := b"1111111111111111_1111111111111111_1110101111100110_1011010110100001"; -- -0.07851090250136859
	pesos_i(761) := b"1111111111111111_1111111111111111_1101101100001000_1100100111110001"; -- -0.14439714293474815
	pesos_i(762) := b"0000000000000000_0000000000000000_0001000111001110_0010010000111010"; -- 0.0695517199157254
	pesos_i(763) := b"0000000000000000_0000000000000000_0000010001110101_0001010100010101"; -- 0.017411534862264735
	pesos_i(764) := b"0000000000000000_0000000000000000_0010100110110010_1101010011101101"; -- 0.1628850058626223
	pesos_i(765) := b"0000000000000000_0000000000000000_0001001001000101_0011011010000000"; -- 0.07136860500002953
	pesos_i(766) := b"0000000000000000_0000000000000000_0001011001101001_1011100110001101"; -- 0.08755073256932848
	pesos_i(767) := b"1111111111111111_1111111111111111_1101110111100111_1111101010011011"; -- -0.13317903258349675
	pesos_i(768) := b"0000000000000000_0000000000000000_0001111110101000_1010011110100110"; -- 0.12366721915108278
	pesos_i(769) := b"1111111111111111_1111111111111111_1111111011100010_0111001101110001"; -- -0.004357132746424896
	pesos_i(770) := b"1111111111111111_1111111111111111_1111110101000111_0011100100110110"; -- -0.010631965976244256
	pesos_i(771) := b"1111111111111111_1111111111111111_1110111011001010_0011001101100110"; -- -0.06722716110913199
	pesos_i(772) := b"1111111111111111_1111111111111111_1111101101101001_1010101011001111"; -- -0.017918896157120733
	pesos_i(773) := b"1111111111111111_1111111111111111_1111010000100100_1101101101101100"; -- -0.04631260494959249
	pesos_i(774) := b"0000000000000000_0000000000000000_0001000101000100_1000111011010010"; -- 0.06745236046086295
	pesos_i(775) := b"0000000000000000_0000000000000000_0000110100011000_0100101000000101"; -- 0.05115187277438035
	pesos_i(776) := b"1111111111111111_1111111111111111_1110000110010010_1110010111010000"; -- -0.11885226898918272
	pesos_i(777) := b"0000000000000000_0000000000000000_0010011001110001_0011100001111100"; -- 0.15016510990831522
	pesos_i(778) := b"1111111111111111_1111111111111111_1101110101111111_0110001000010010"; -- -0.13477503826000622
	pesos_i(779) := b"0000000000000000_0000000000000000_0010001011010000_1011011001011001"; -- 0.13599719679231267
	pesos_i(780) := b"1111111111111111_1111111111111111_1110010110100111_1101110101011011"; -- -0.10290733837427517
	pesos_i(781) := b"1111111111111111_1111111111111111_1110110110111101_1101010111110001"; -- -0.07132208696506037
	pesos_i(782) := b"1111111111111111_1111111111111111_1111110111001011_1000010110111111"; -- -0.008613244045393311
	pesos_i(783) := b"1111111111111111_1111111111111111_1110000111111101_0111100001001011"; -- -0.11722610643356678
	pesos_i(784) := b"0000000000000000_0000000000000000_0001001001001110_1100100011110110"; -- 0.07151466374792312
	pesos_i(785) := b"0000000000000000_0000000000000000_0000111111000000_1110110000100111"; -- 0.06153751321953872
	pesos_i(786) := b"1111111111111111_1111111111111111_1111100111010110_1100111000000110"; -- -0.024066089098849476
	pesos_i(787) := b"0000000000000000_0000000000000000_0001000110001101_0001001011000111"; -- 0.06855885848540014
	pesos_i(788) := b"0000000000000000_0000000000000000_0001001111011100_1100001000010010"; -- 0.07758725101481041
	pesos_i(789) := b"1111111111111111_1111111111111111_1101111110110100_0101010101000100"; -- -0.1261545858168314
	pesos_i(790) := b"0000000000000000_0000000000000000_0001100011010011_1001101100001010"; -- 0.09697884545574342
	pesos_i(791) := b"1111111111111111_1111111111111111_1110000000010010_0101011110101010"; -- -0.12472011652973249
	pesos_i(792) := b"1111111111111111_1111111111111111_1111011010010010_1010001101001010"; -- -0.03682498410122764
	pesos_i(793) := b"0000000000000000_0000000000000000_0010010101000000_1111011001100010"; -- 0.14552249805683407
	pesos_i(794) := b"0000000000000000_0000000000000000_0000111011111111_0101110111000001"; -- 0.05858407936911923
	pesos_i(795) := b"0000000000000000_0000000000000000_0001110100011110_0111011011111110"; -- 0.11374610614558163
	pesos_i(796) := b"1111111111111111_1111111111111111_1111111101001010_0110000101001000"; -- -0.0027713013108452474
	pesos_i(797) := b"0000000000000000_0000000000000000_0000110101101001_1001110010100111"; -- 0.05239276004381879
	pesos_i(798) := b"0000000000000000_0000000000000000_0001010101001010_0110100101011111"; -- 0.08316668089345508
	pesos_i(799) := b"1111111111111111_1111111111111111_1111010011001111_0011101111000010"; -- -0.04371286877465136
	pesos_i(800) := b"1111111111111111_1111111111111111_1111101100011011_0101010111010010"; -- -0.019114147292084382
	pesos_i(801) := b"0000000000000000_0000000000000000_0000001110101101_0011000000010011"; -- 0.014361385917294479
	pesos_i(802) := b"0000000000000000_0000000000000000_0000100010101000_1000010111011011"; -- 0.03382145498658313
	pesos_i(803) := b"0000000000000000_0000000000000000_0010011011000111_1100000100110100"; -- 0.15148551479384298
	pesos_i(804) := b"1111111111111111_1111111111111111_1101010000111000_1011011101010110"; -- -0.1710095801931925
	pesos_i(805) := b"0000000000000000_0000000000000000_0001111011011001_1010000011010111"; -- 0.12050824405530217
	pesos_i(806) := b"0000000000000000_0000000000000000_0001101000000111_0100000110111011"; -- 0.10167322944215644
	pesos_i(807) := b"1111111111111111_1111111111111111_1110010000111111_0101110111101100"; -- -0.10840809813470195
	pesos_i(808) := b"1111111111111111_1111111111111111_1110100110111100_1001110001100100"; -- -0.08696577604989092
	pesos_i(809) := b"0000000000000000_0000000000000000_0000000100100111_0010000000110100"; -- 0.004503262310566006
	pesos_i(810) := b"1111111111111111_1111111111111111_1111000110100111_0111000101111110"; -- -0.056038767530678595
	pesos_i(811) := b"0000000000000000_0000000000000000_0001111110101101_1011010011110000"; -- 0.12374430516946586
	pesos_i(812) := b"1111111111111111_1111111111111111_1101001111110000_1110010110001110"; -- -0.17210545813215666
	pesos_i(813) := b"1111111111111111_1111111111111111_1101101011111010_0111101010101101"; -- -0.14461549072003194
	pesos_i(814) := b"1111111111111111_1111111111111111_1110001010011101_1001011110101011"; -- -0.11478283004650847
	pesos_i(815) := b"0000000000000000_0000000000000000_0000111100101010_0000110111011001"; -- 0.059235444597905695
	pesos_i(816) := b"0000000000000000_0000000000000000_0001010010011011_0110100111001000"; -- 0.0804964174607877
	pesos_i(817) := b"1111111111111111_1111111111111111_1111100000100001_1010100010111011"; -- -0.03073640284414772
	pesos_i(818) := b"1111111111111111_1111111111111111_1101110101101011_1111110001100110"; -- -0.13507101536099902
	pesos_i(819) := b"0000000000000000_0000000000000000_0010110001111101_0111010100001010"; -- 0.17378932472160735
	pesos_i(820) := b"0000000000000000_0000000000000000_0000011001100100_1011010001110000"; -- 0.02497413389352191
	pesos_i(821) := b"1111111111111111_1111111111111111_1110110111011010_0110011110101010"; -- -0.07088615502064029
	pesos_i(822) := b"1111111111111111_1111111111111111_1101100110100101_1100101100001010"; -- -0.1498139477186992
	pesos_i(823) := b"0000000000000000_0000000000000000_0000111011001111_1100100010100000"; -- 0.05785802759925492
	pesos_i(824) := b"0000000000000000_0000000000000000_0000110100011111_0010100101001111"; -- 0.05125673458330807
	pesos_i(825) := b"0000000000000000_0000000000000000_0000110101010100_0000001001011001"; -- 0.052063128175626756
	pesos_i(826) := b"1111111111111111_1111111111111111_1111100011100110_0101010100111001"; -- -0.027735398744463912
	pesos_i(827) := b"1111111111111111_1111111111111111_1111011000001100_0001101000100001"; -- -0.038877837148296464
	pesos_i(828) := b"1111111111111111_1111111111111111_1101110100110111_0000000011110000"; -- -0.1358794608111569
	pesos_i(829) := b"0000000000000000_0000000000000000_0001100011011011_1000101110010010"; -- 0.09709999373451395
	pesos_i(830) := b"1111111111111111_1111111111111111_1111000001000011_1001001101010010"; -- -0.06146888021770889
	pesos_i(831) := b"1111111111111111_1111111111111111_1101011111110110_0100010001001111"; -- -0.15639851638875096
	pesos_i(832) := b"1111111111111111_1111111111111111_1110111111000010_0101101011000100"; -- -0.06344063482587034
	pesos_i(833) := b"0000000000000000_0000000000000000_0000001000001000_1001100011010110"; -- 0.007943680050830354
	pesos_i(834) := b"1111111111111111_1111111111111111_1111000011010101_1011001011011100"; -- -0.059239216989002565
	pesos_i(835) := b"1111111111111111_1111111111111111_1111100111110101_1010011010001001"; -- -0.0235954203979614
	pesos_i(836) := b"0000000000000000_0000000000000000_0000101000011101_0001100101000000"; -- 0.03950650991198381
	pesos_i(837) := b"0000000000000000_0000000000000000_0001011010010101_1011100011110001"; -- 0.08822208301981757
	pesos_i(838) := b"0000000000000000_0000000000000000_0000110100010110_0000111010010111"; -- 0.05111781295796908
	pesos_i(839) := b"0000000000000000_0000000000000000_0001010000111100_0110011000010000"; -- 0.07904661085782963
	pesos_i(840) := b"1111111111111111_1111111111111111_1110110011110101_1100010111111010"; -- -0.07437479645948329
	pesos_i(841) := b"0000000000000000_0000000000000000_0001010100100000_0111110010010101"; -- 0.08252695687619047
	pesos_i(842) := b"0000000000000000_0000000000000000_0000000001001000_0110000011011111"; -- 0.0011044068530546396
	pesos_i(843) := b"0000000000000000_0000000000000000_0000101111000111_1000011100011000"; -- 0.04601330125414807
	pesos_i(844) := b"0000000000000000_0000000000000000_0000000111011001_1110111010001011"; -- 0.007231625447656433
	pesos_i(845) := b"1111111111111111_1111111111111111_1111000101010011_1100111101111111"; -- -0.05731490286712338
	pesos_i(846) := b"1111111111111111_1111111111111111_1101010101001001_1111000111000100"; -- -0.16684044806300882
	pesos_i(847) := b"0000000000000000_0000000000000000_0001100111110101_1000011110101001"; -- 0.10140273935640397
	pesos_i(848) := b"0000000000000000_0000000000000000_0010011010111000_1110010010000011"; -- 0.15125873760905253
	pesos_i(849) := b"0000000000000000_0000000000000000_0001110110111101_1011110111011000"; -- 0.11617647670881379
	pesos_i(850) := b"1111111111111111_1111111111111111_1110110101111010_1110110110001000"; -- -0.07234301973268403
	pesos_i(851) := b"0000000000000000_0000000000000000_0000011100100101_1111000000001011"; -- 0.02792263289323387
	pesos_i(852) := b"1111111111111111_1111111111111111_1101111001001110_0111010100111010"; -- -0.1316153273128208
	pesos_i(853) := b"0000000000000000_0000000000000000_0010101111110110_0111011111100100"; -- 0.17172955811248045
	pesos_i(854) := b"0000000000000000_0000000000000000_0010011110010110_1100101101110100"; -- 0.15464469512791318
	pesos_i(855) := b"1111111111111111_1111111111111111_1111101110011110_0000100111000001"; -- -0.017119779843974815
	pesos_i(856) := b"1111111111111111_1111111111111111_1111101000001100_0101011010010001"; -- -0.023249234799289146
	pesos_i(857) := b"0000000000000000_0000000000000000_0001000000111101_1011110011111101"; -- 0.06344205070712047
	pesos_i(858) := b"1111111111111111_1111111111111111_1101110011010000_0010110111100111"; -- -0.1374484358432456
	pesos_i(859) := b"1111111111111111_1111111111111111_1110110000100101_1001010100011000"; -- -0.07755153807348278
	pesos_i(860) := b"0000000000000000_0000000000000000_0001100100001111_1110001000000100"; -- 0.09789860333696228
	pesos_i(861) := b"1111111111111111_1111111111111111_1101100101011101_0010101100000101"; -- -0.150922118483189
	pesos_i(862) := b"0000000000000000_0000000000000000_0010000011111000_1001000110001001"; -- 0.12879285436326046
	pesos_i(863) := b"1111111111111111_1111111111111111_1101010100111001_0101101111110001"; -- -0.167093518983213
	pesos_i(864) := b"0000000000000000_0000000000000000_0001100010000001_1100010101011010"; -- 0.09573014682643752
	pesos_i(865) := b"1111111111111111_1111111111111111_1110000111101010_0001010110111100"; -- -0.11752189786021153
	pesos_i(866) := b"1111111111111111_1111111111111111_1101011001011100_0100010100000010"; -- -0.1626545781457472
	pesos_i(867) := b"1111111111111111_1111111111111111_1101110100010110_0100100011111010"; -- -0.13637870679600303
	pesos_i(868) := b"1111111111111111_1111111111111111_1101101011100000_1100000001011110"; -- -0.14500806525013873
	pesos_i(869) := b"1111111111111111_1111111111111111_1111000101000011_0011011010111001"; -- -0.0575681494963201
	pesos_i(870) := b"0000000000000000_0000000000000000_0000001111111000_1100011100010001"; -- 0.015514794929305813
	pesos_i(871) := b"0000000000000000_0000000000000000_0001100010010111_0110110011111110"; -- 0.09606057368974844
	pesos_i(872) := b"1111111111111111_1111111111111111_1110011110000010_0000001010101101"; -- -0.09567244798627057
	pesos_i(873) := b"1111111111111111_1111111111111111_1110011101111110_0100111100111010"; -- -0.0957289202964078
	pesos_i(874) := b"1111111111111111_1111111111111111_1111101111000001_0100010010001010"; -- -0.016582218483500166
	pesos_i(875) := b"1111111111111111_1111111111111111_1101100111101101_0001101001110000"; -- -0.1487258411355398
	pesos_i(876) := b"0000000000000000_0000000000000000_0010100001010000_0111110111111101"; -- 0.15747821261120148
	pesos_i(877) := b"1111111111111111_1111111111111111_1111001000000011_0010100000100101"; -- -0.05463933091081873
	pesos_i(878) := b"1111111111111111_1111111111111111_1111011000001100_1101101010001100"; -- -0.038866368170657715
	pesos_i(879) := b"1111111111111111_1111111111111111_1101010101010011_1100100101100000"; -- -0.16669026754454852
	pesos_i(880) := b"0000000000000000_0000000000000000_0010101111111110_0000001000000001"; -- 0.17184460182796815
	pesos_i(881) := b"1111111111111111_1111111111111111_1110001011100111_0000001001010001"; -- -0.11366258157698335
	pesos_i(882) := b"1111111111111111_1111111111111111_1111001111110010_0100010110011010"; -- -0.04708447445928824
	pesos_i(883) := b"0000000000000000_0000000000000000_0000101100011111_1001100100011001"; -- 0.043450897812600524
	pesos_i(884) := b"1111111111111111_1111111111111111_1101111100001000_0101011100111110"; -- -0.12877897954173478
	pesos_i(885) := b"0000000000000000_0000000000000000_0001111000011010_1000101001100100"; -- 0.11759247714866204
	pesos_i(886) := b"1111111111111111_1111111111111111_1111111011110100_0001110010000100"; -- -0.004087655775818721
	pesos_i(887) := b"0000000000000000_0000000000000000_0001110111100111_0000001001010000"; -- 0.11680616800211596
	pesos_i(888) := b"1111111111111111_1111111111111111_1101001111101111_1100001110000111"; -- -0.1721227451622295
	pesos_i(889) := b"0000000000000000_0000000000000000_0000010101001001_0110010000100001"; -- 0.020651109779786014
	pesos_i(890) := b"0000000000000000_0000000000000000_0001010000011101_1110101001010111"; -- 0.07858147260301382
	pesos_i(891) := b"0000000000000000_0000000000000000_0000000111011010_1101111110111010"; -- 0.007246001271448968
	pesos_i(892) := b"0000000000000000_0000000000000000_0010100111100000_1100011101101001"; -- 0.16358610456743772
	pesos_i(893) := b"0000000000000000_0000000000000000_0000011010100001_0001011011011100"; -- 0.025895527672539834
	pesos_i(894) := b"1111111111111111_1111111111111111_1101111010000110_0101101100010010"; -- -0.13076239414947252
	pesos_i(895) := b"1111111111111111_1111111111111111_1111111110101111_0100110110110111"; -- -0.0012313298432161971
	pesos_i(896) := b"0000000000000000_0000000000000000_0010101110110101_1000110010100111"; -- 0.17073897433169474
	pesos_i(897) := b"0000000000000000_0000000000000000_0010000110110000_1001101001011100"; -- 0.13160099752033952
	pesos_i(898) := b"0000000000000000_0000000000000000_0000110101001111_1111111100001110"; -- 0.05200189680183818
	pesos_i(899) := b"1111111111111111_1111111111111111_1110101010001111_1000000110011110"; -- -0.08374776731858345
	pesos_i(900) := b"1111111111111111_1111111111111111_1101001001001001_1111100110000110"; -- -0.17855873561094135
	pesos_i(901) := b"1111111111111111_1111111111111111_1111011001010011_0110100111111011"; -- -0.03778970358226091
	pesos_i(902) := b"1111111111111111_1111111111111111_1111100000110001_0100000101011111"; -- -0.03049842292378512
	pesos_i(903) := b"0000000000000000_0000000000000000_0000011100110001_1010001100101010"; -- 0.028101156039147496
	pesos_i(904) := b"0000000000000000_0000000000000000_0000101110111100_0101100000010001"; -- 0.045842651625184826
	pesos_i(905) := b"1111111111111111_1111111111111111_1111000100110110_0000100110010100"; -- -0.05776920455408073
	pesos_i(906) := b"1111111111111111_1111111111111111_1111001011100111_0011101000011001"; -- -0.051159256873167726
	pesos_i(907) := b"1111111111111111_1111111111111111_1110001010110111_0011011100111010"; -- -0.11439184972896503
	pesos_i(908) := b"1111111111111111_1111111111111111_1110001000001100_0111111101000001"; -- -0.11699680958009948
	pesos_i(909) := b"0000000000000000_0000000000000000_0001010101010111_1110001111011011"; -- 0.08337234598110002
	pesos_i(910) := b"1111111111111111_1111111111111111_1110101011110101_1010011111011111"; -- -0.0821890908846683
	pesos_i(911) := b"0000000000000000_0000000000000000_0001110001001010_0010001100000100"; -- 0.11050623740063563
	pesos_i(912) := b"0000000000000000_0000000000000000_0010010101111001_1100111101101001"; -- 0.14638992604729753
	pesos_i(913) := b"1111111111111111_1111111111111111_1111001010001100_0011110010001000"; -- -0.052547661671679444
	pesos_i(914) := b"0000000000000000_0000000000000000_0001101011110111_1110011110011010"; -- 0.10534522533935639
	pesos_i(915) := b"1111111111111111_1111111111111111_1110011110010010_0100110000001100"; -- -0.09542393407803625
	pesos_i(916) := b"0000000000000000_0000000000000000_0000110001111001_0111110111100001"; -- 0.04872881634915506
	pesos_i(917) := b"1111111111111111_1111111111111111_1110011000100001_0011011111011001"; -- -0.10105563121128963
	pesos_i(918) := b"0000000000000000_0000000000000000_0001111011110101_1001010101000000"; -- 0.1209347992010761
	pesos_i(919) := b"1111111111111111_1111111111111111_1101110010011111_0011110000101001"; -- -0.13819526660210796
	pesos_i(920) := b"1111111111111111_1111111111111111_1110100010110101_0010001111100001"; -- -0.09098602070969443
	pesos_i(921) := b"1111111111111111_1111111111111111_1101100011010000_1011111100101011"; -- -0.15306477742724428
	pesos_i(922) := b"1111111111111111_1111111111111111_1111010011001110_0001000110000000"; -- -0.04373064629283415
	pesos_i(923) := b"0000000000000000_0000000000000000_0000110111011111_1101010110101010"; -- 0.05419669536150581
	pesos_i(924) := b"0000000000000000_0000000000000000_0010010010011011_1110101101000110"; -- 0.14300413573730397
	pesos_i(925) := b"0000000000000000_0000000000000000_0000000011010110_1111011000101000"; -- 0.003280052944684043
	pesos_i(926) := b"0000000000000000_0000000000000000_0001011001011111_1000110100111001"; -- 0.08739550245943863
	pesos_i(927) := b"1111111111111111_1111111111111111_1110111011100001_0101111111111110"; -- -0.06687355083218247
	pesos_i(928) := b"0000000000000000_0000000000000000_0010011001100110_1110111011011001"; -- 0.15000813283808853
	pesos_i(929) := b"1111111111111111_1111111111111111_1111010110000110_1001101111101100"; -- -0.04091477863857343
	pesos_i(930) := b"0000000000000000_0000000000000000_0001110101111010_0110100000100111"; -- 0.11514903030817668
	pesos_i(931) := b"1111111111111111_1111111111111111_1101000110101011_0000000101001010"; -- -0.1809844203089488
	pesos_i(932) := b"0000000000000000_0000000000000000_0000101001000111_1010001110011001"; -- 0.04015562522444885
	pesos_i(933) := b"0000000000000000_0000000000000000_0001101101011111_1011000011101011"; -- 0.10692888009902053
	pesos_i(934) := b"0000000000000000_0000000000000000_0000100100010111_0010011110011100"; -- 0.03550956296807226
	pesos_i(935) := b"1111111111111111_1111111111111111_1110000100100010_0011101101110101"; -- -0.12057140719901431
	pesos_i(936) := b"1111111111111111_1111111111111111_1111110100011010_1110110000011010"; -- -0.01130794862778467
	pesos_i(937) := b"0000000000000000_0000000000000000_0000101110001110_1110101111110010"; -- 0.0451495614873866
	pesos_i(938) := b"1111111111111111_1111111111111111_1101100001011010_1010101010110011"; -- -0.15486653447355864
	pesos_i(939) := b"0000000000000000_0000000000000000_0000100111100010_0111100101010001"; -- 0.03861196728055762
	pesos_i(940) := b"0000000000000000_0000000000000000_0000101111101010_0110001011011001"; -- 0.04654519837166531
	pesos_i(941) := b"0000000000000000_0000000000000000_0010011001000011_1101001011101110"; -- 0.14947241121446986
	pesos_i(942) := b"0000000000000000_0000000000000000_0010010000000110_0111110100110111"; -- 0.1407240161202302
	pesos_i(943) := b"1111111111111111_1111111111111111_1101001111110110_1010001010110000"; -- -0.17201789088692646
	pesos_i(944) := b"1111111111111111_1111111111111111_1111000100110111_1001101001000100"; -- -0.057745321764647375
	pesos_i(945) := b"1111111111111111_1111111111111111_1101010001001010_1001011001001101"; -- -0.17073689090647298
	pesos_i(946) := b"0000000000000000_0000000000000000_0001100100101011_0001000110100110"; -- 0.0983134298650192
	pesos_i(947) := b"0000000000000000_0000000000000000_0010100011000000_1001111011111000"; -- 0.15918916278478967
	pesos_i(948) := b"0000000000000000_0000000000000000_0001000111011111_0000001110111001"; -- 0.06980918187832305
	pesos_i(949) := b"0000000000000000_0000000000000000_0000011011101110_0000010011100100"; -- 0.027069383240578716
	pesos_i(950) := b"0000000000000000_0000000000000000_0001111000011110_0110011010101100"; -- 0.11765138346105981
	pesos_i(951) := b"0000000000000000_0000000000000000_0010000101000111_0001110001110101"; -- 0.12999132028975657
	pesos_i(952) := b"0000000000000000_0000000000000000_0001011111101001_0100000011000011"; -- 0.09340290792742786
	pesos_i(953) := b"0000000000000000_0000000000000000_0001100011110101_1101101100111100"; -- 0.09750147070829636
	pesos_i(954) := b"0000000000000000_0000000000000000_0001000110100101_0010110100100000"; -- 0.06892663975813187
	pesos_i(955) := b"1111111111111111_1111111111111111_1111001100010111_1001110000010000"; -- -0.05042099580333223
	pesos_i(956) := b"0000000000000000_0000000000000000_0001110000111010_0100111001111000"; -- 0.11026468678776773
	pesos_i(957) := b"0000000000000000_0000000000000000_0010100111111000_0111110000000011"; -- 0.16394782127023338
	pesos_i(958) := b"0000000000000000_0000000000000000_0001110010000010_0100000110110010"; -- 0.11136255823744279
	pesos_i(959) := b"0000000000000000_0000000000000000_0000001101011011_0011011010100100"; -- 0.013110556684168781
	pesos_i(960) := b"0000000000000000_0000000000000000_0001000111111000_0111101000100100"; -- 0.07019770974888073
	pesos_i(961) := b"0000000000000000_0000000000000000_0000101101001011_0110011111010011"; -- 0.04411934766166213
	pesos_i(962) := b"0000000000000000_0000000000000000_0000010101001101_1011100001010000"; -- 0.020717162570812145
	pesos_i(963) := b"0000000000000000_0000000000000000_0001011101001111_1010111011010110"; -- 0.09105961546145004
	pesos_i(964) := b"0000000000000000_0000000000000000_0001000101110110_1011011101100111"; -- 0.06821771869365159
	pesos_i(965) := b"1111111111111111_1111111111111111_1111110111111010_0010001000010000"; -- -0.007902022507136291
	pesos_i(966) := b"0000000000000000_0000000000000000_0000010100001011_0101000011011100"; -- 0.019703916270843364
	pesos_i(967) := b"0000000000000000_0000000000000000_0010011000011110_1010001111101111"; -- 0.14890503495547225
	pesos_i(968) := b"0000000000000000_0000000000000000_0000110100010000_1101111000010001"; -- 0.051038626754335965
	pesos_i(969) := b"1111111111111111_1111111111111111_1101111000111000_0111001100100001"; -- -0.13195114558458548
	pesos_i(970) := b"0000000000000000_0000000000000000_0001001110110000_1111000101100010"; -- 0.07691868449962873
	pesos_i(971) := b"0000000000000000_0000000000000000_0000001110010101_0010101000110101"; -- 0.013994825400417271
	pesos_i(972) := b"1111111111111111_1111111111111111_1111101111100011_1010000000111010"; -- -0.016057954548344397
	pesos_i(973) := b"0000000000000000_0000000000000000_0000100010000110_0010010010000011"; -- 0.03329685404059239
	pesos_i(974) := b"1111111111111111_1111111111111111_1110000000101001_1101111000010100"; -- -0.12436115280573827
	pesos_i(975) := b"0000000000000000_0000000000000000_0000000111010111_1010000010000001"; -- 0.0071964564141046095
	pesos_i(976) := b"0000000000000000_0000000000000000_0000010011000111_1111000110001001"; -- 0.01867589559148311
	pesos_i(977) := b"1111111111111111_1111111111111111_1111100111011011_0110001011000011"; -- -0.023996188532650155
	pesos_i(978) := b"1111111111111111_1111111111111111_1101110001011011_0110011010110100"; -- -0.13923032862792614
	pesos_i(979) := b"1111111111111111_1111111111111111_1110000010111100_0110000001101101"; -- -0.12212560025523436
	pesos_i(980) := b"0000000000000000_0000000000000000_0010011001110111_0101010011110011"; -- 0.1502583593502044
	pesos_i(981) := b"1111111111111111_1111111111111111_1110000100101010_0001100111100011"; -- -0.12045133793170394
	pesos_i(982) := b"0000000000000000_0000000000000000_0001010011000110_1100100001110110"; -- 0.08115818871634617
	pesos_i(983) := b"1111111111111111_1111111111111111_1111011000111001_1000111111000110"; -- -0.03818417951339282
	pesos_i(984) := b"0000000000000000_0000000000000000_0001000000011010_1001100111111110"; -- 0.06290590725932983
	pesos_i(985) := b"0000000000000000_0000000000000000_0010011100110010_0101110111101010"; -- 0.1531122872200887
	pesos_i(986) := b"0000000000000000_0000000000000000_0000100011001010_1111100010100011"; -- 0.03434709528007327
	pesos_i(987) := b"0000000000000000_0000000000000000_0000011010011111_0001010101101000"; -- 0.02586492336208613
	pesos_i(988) := b"0000000000000000_0000000000000000_0001111001011010_0010010010100101"; -- 0.11856297531622313
	pesos_i(989) := b"1111111111111111_1111111111111111_1111111101100010_1101001101111101"; -- -0.002398282961991609
	pesos_i(990) := b"1111111111111111_1111111111111111_1110000001000111_0100001111111100"; -- -0.1239125737975966
	pesos_i(991) := b"1111111111111111_1111111111111111_1101100100100011_1000000110011011"; -- -0.15180196736220275
	pesos_i(992) := b"0000000000000000_0000000000000000_0000110000001010_0110010011011101"; -- 0.04703359971010365
	pesos_i(993) := b"1111111111111111_1111111111111111_1110111101001110_0111101101101111"; -- -0.06520870728439884
	pesos_i(994) := b"0000000000000000_0000000000000000_0001110111110101_0101000110110101"; -- 0.11702452354775619
	pesos_i(995) := b"1111111111111111_1111111111111111_1110001011100111_0010010010110000"; -- -0.11366053296014592
	pesos_i(996) := b"0000000000000000_0000000000000000_0001001100011110_1111001001011110"; -- 0.07469095983919247
	pesos_i(997) := b"1111111111111111_1111111111111111_1111000000111001_0111010001101111"; -- -0.06162330895310244
	pesos_i(998) := b"1111111111111111_1111111111111111_1110100100111100_0111110111111101"; -- -0.08892071328556261
	pesos_i(999) := b"0000000000000000_0000000000000000_0010010000001010_0000001000111000"; -- 0.1407777201269175
	pesos_i(1000) := b"1111111111111111_1111111111111111_1110000000001111_0100010110100010"; -- -0.12476696781377863
	pesos_i(1001) := b"0000000000000000_0000000000000000_0001100011010010_1100101111001110"; -- 0.09696649351774628
	pesos_i(1002) := b"1111111111111111_1111111111111111_1110111110010111_0101000110011101"; -- -0.06409730827124133
	pesos_i(1003) := b"0000000000000000_0000000000000000_0010000101000111_1010110000010100"; -- 0.1299998805774685
	pesos_i(1004) := b"0000000000000000_0000000000000000_0001000100101011_0100101000101011"; -- 0.0670667986730814
	pesos_i(1005) := b"1111111111111111_1111111111111111_1111100001010011_1011101100000010"; -- -0.029972374008333722
	pesos_i(1006) := b"1111111111111111_1111111111111111_1101010101100000_1101001101000100"; -- -0.16649131394462202
	pesos_i(1007) := b"1111111111111111_1111111111111111_1101011001110111_1001110111110010"; -- -0.1622372897864117
	pesos_i(1008) := b"0000000000000000_0000000000000000_0000001101100010_0110110111110010"; -- 0.013220664687207756
	pesos_i(1009) := b"1111111111111111_1111111111111111_1111110101010100_0110111100000001"; -- -0.010430395458739672
	pesos_i(1010) := b"0000000000000000_0000000000000000_0000111011101110_0101001010010111"; -- 0.05832401442157792
	pesos_i(1011) := b"1111111111111111_1111111111111111_1110010101010011_0010000011101111"; -- -0.1042003075331717
	pesos_i(1012) := b"0000000000000000_0000000000000000_0000100001010110_1011011110110110"; -- 0.03257320589143734
	pesos_i(1013) := b"0000000000000000_0000000000000000_0000100100111000_1000001100101000"; -- 0.036018559696013905
	pesos_i(1014) := b"1111111111111111_1111111111111111_1101010101111100_1000101011011011"; -- -0.1660683837289574
	pesos_i(1015) := b"0000000000000000_0000000000000000_0010011011100110_1011010010001111"; -- 0.1519577835496657
	pesos_i(1016) := b"1111111111111111_1111111111111111_1101011101100100_1010000100011010"; -- -0.1586207687533583
	pesos_i(1017) := b"1111111111111111_1111111111111111_1111100100010011_1001100010111000"; -- -0.027044730239610848
	pesos_i(1018) := b"0000000000000000_0000000000000000_0010001001100010_0000011110011100"; -- 0.1343083148441811
	pesos_i(1019) := b"1111111111111111_1111111111111111_1111001111000101_1011011011101000"; -- -0.047764366405149195
	pesos_i(1020) := b"0000000000000000_0000000000000000_0010000000110000_0100101011001101"; -- 0.1257368802925497
	pesos_i(1021) := b"1111111111111111_1111111111111111_1101110011010100_0000111011111001"; -- -0.13738924418938445
	pesos_i(1022) := b"0000000000000000_0000000000000000_0000110000010111_1110110101011000"; -- 0.047240099026694356
	pesos_i(1023) := b"1111111111111111_1111111111111111_1110010110000000_0001000101000101"; -- -0.10351459564546166
	pesos_i(1024) := b"1111111111111111_1111111111111111_1111100001111011_0001101000001111"; -- -0.029371615626410358
	pesos_i(1025) := b"0000000000000000_0000000000000000_0010001111100010_0110110001010000"; -- 0.14017369218703396
	pesos_i(1026) := b"0000000000000000_0000000000000000_0000111110101000_1111111110000000"; -- 0.061172455626024975
	pesos_i(1027) := b"0000000000000000_0000000000000000_0001001000011001_0111110000110110"; -- 0.07070137320531802
	pesos_i(1028) := b"0000000000000000_0000000000000000_0000111100111101_1011100000101000"; -- 0.059535512774792604
	pesos_i(1029) := b"0000000000000000_0000000000000000_0010000110110000_1011111011101010"; -- 0.13160317619609696
	pesos_i(1030) := b"0000000000000000_0000000000000000_0010010011011110_1000101000100101"; -- 0.14402068532749307
	pesos_i(1031) := b"1111111111111111_1111111111111111_1101100011001010_1101111000110000"; -- -0.1531544812405344
	pesos_i(1032) := b"0000000000000000_0000000000000000_0010010100101000_1000010000101101"; -- 0.14514947994958374
	pesos_i(1033) := b"1111111111111111_1111111111111111_1101101110000001_0010011110001110"; -- -0.1425605086809183
	pesos_i(1034) := b"0000000000000000_0000000000000000_0001011100111010_1010110010101111"; -- 0.09073905248910058
	pesos_i(1035) := b"1111111111111111_1111111111111111_1101110010100001_1111110001000101"; -- -0.13815329845629756
	pesos_i(1036) := b"0000000000000000_0000000000000000_0001101011100011_1100001011011000"; -- 0.10503785865434691
	pesos_i(1037) := b"1111111111111111_1111111111111111_1111010000101010_0000011001101001"; -- -0.04623374869740005
	pesos_i(1038) := b"1111111111111111_1111111111111111_1110010000010110_0000110110001111"; -- -0.10903849848006371
	pesos_i(1039) := b"0000000000000000_0000000000000000_0001011101101011_0100010101001000"; -- 0.09148056987243915
	pesos_i(1040) := b"1111111111111111_1111111111111111_1101101110110110_1010101101101000"; -- -0.1417439336770398
	pesos_i(1041) := b"0000000000000000_0000000000000000_0000111101000011_1010001001010101"; -- 0.059625764709500054
	pesos_i(1042) := b"0000000000000000_0000000000000000_0000000001101100_1000110100001000"; -- 0.001656355241862361
	pesos_i(1043) := b"1111111111111111_1111111111111111_1110001011000100_0110010000011110"; -- -0.11419080985080851
	pesos_i(1044) := b"0000000000000000_0000000000000000_0000110001101001_0101011110001110"; -- 0.04848239147688567
	pesos_i(1045) := b"1111111111111111_1111111111111111_1111110100000000_1110100010011011"; -- -0.011704885723392837
	pesos_i(1046) := b"0000000000000000_0000000000000000_0001101100110100_1101010111100001"; -- 0.1062749551301437
	pesos_i(1047) := b"0000000000000000_0000000000000000_0000101011111010_0011110100001110"; -- 0.042880836314044476
	pesos_i(1048) := b"1111111111111111_1111111111111111_1111010101100001_1110010000001000"; -- -0.041475055680299557
	pesos_i(1049) := b"1111111111111111_1111111111111111_1101100000110010_1111110111110101"; -- -0.15547192346445596
	pesos_i(1050) := b"0000000000000000_0000000000000000_0001111010100000_1101000110100011"; -- 0.11964140154400138
	pesos_i(1051) := b"0000000000000000_0000000000000000_0001111110110011_1111111000111010"; -- 0.12384022642931496
	pesos_i(1052) := b"0000000000000000_0000000000000000_0001011111010101_1011111110110110"; -- 0.09310529892611435
	pesos_i(1053) := b"1111111111111111_1111111111111111_1101111001000110_0110110000000111"; -- -0.1317379459085808
	pesos_i(1054) := b"1111111111111111_1111111111111111_1110000011010111_0011000010101110"; -- -0.12171645875110396
	pesos_i(1055) := b"0000000000000000_0000000000000000_0001011011100110_1101011110000100"; -- 0.08945986721582447
	pesos_i(1056) := b"0000000000000000_0000000000000000_0000101010000011_1111110100101000"; -- 0.04107649072379463
	pesos_i(1057) := b"1111111111111111_1111111111111111_1110000000011111_0111000101011110"; -- -0.12452022030891345
	pesos_i(1058) := b"1111111111111111_1111111111111111_1101100100111010_0001111000000110"; -- -0.15145695079635196
	pesos_i(1059) := b"1111111111111111_1111111111111111_1110110000110111_1100011111011100"; -- -0.0772738541541417
	pesos_i(1060) := b"0000000000000000_0000000000000000_0001010100100110_0000010101110101"; -- 0.08261140936048167
	pesos_i(1061) := b"1111111111111111_1111111111111111_1110110000011100_1000100011110000"; -- -0.07768959171256615
	pesos_i(1062) := b"1111111111111111_1111111111111111_1110000001100110_1111111100110110"; -- -0.12342839174414251
	pesos_i(1063) := b"1111111111111111_1111111111111111_1111010111110011_1101111110100010"; -- -0.03924753475223866
	pesos_i(1064) := b"1111111111111111_1111111111111111_1101011111010100_1101011001011100"; -- -0.15690860995661499
	pesos_i(1065) := b"0000000000000000_0000000000000000_0010000111001011_0010110010111111"; -- 0.1320064512770979
	pesos_i(1066) := b"0000000000000000_0000000000000000_0001000000011010_1001001010010010"; -- 0.06290546470669559
	pesos_i(1067) := b"1111111111111111_1111111111111111_1110100011010011_1100001001010100"; -- -0.09051881272047253
	pesos_i(1068) := b"0000000000000000_0000000000000000_0001100010011100_1100111011001100"; -- 0.09614269726048849
	pesos_i(1069) := b"0000000000000000_0000000000000000_0000011000110111_1111100111011000"; -- 0.0242916253212646
	pesos_i(1070) := b"0000000000000000_0000000000000000_0010001011101001_0100011000110011"; -- 0.13637198207881257
	pesos_i(1071) := b"1111111111111111_1111111111111111_1110011000100110_1001011100100011"; -- -0.10097365766726703
	pesos_i(1072) := b"0000000000000000_0000000000000000_0010001100111100_1011111100110110"; -- 0.13764567444968076
	pesos_i(1073) := b"0000000000000000_0000000000000000_0001100111111100_0001111001000101"; -- 0.10150326911793069
	pesos_i(1074) := b"0000000000000000_0000000000000000_0001101010001111_1000111000101110"; -- 0.10375298146113439
	pesos_i(1075) := b"0000000000000000_0000000000000000_0000000000101110_1011101000100111"; -- 0.0007129998783904695
	pesos_i(1076) := b"0000000000000000_0000000000000000_0000100010000100_0000111101110011"; -- 0.0332650810863608
	pesos_i(1077) := b"1111111111111111_1111111111111111_1110001111001010_0011101101101100"; -- -0.11019543274549973
	pesos_i(1078) := b"0000000000000000_0000000000000000_0000010000010101_1101010001011000"; -- 0.01595809129182092
	pesos_i(1079) := b"0000000000000000_0000000000000000_0000011110100011_1100011001111111"; -- 0.029842763929716434
	pesos_i(1080) := b"1111111111111111_1111111111111111_1101101001101011_1101010000011010"; -- -0.1467921674368406
	pesos_i(1081) := b"1111111111111111_1111111111111111_1110011001100100_0011010001010001"; -- -0.10003350288931986
	pesos_i(1082) := b"1111111111111111_1111111111111111_1111101000011101_0101011011011100"; -- -0.02298981796201989
	pesos_i(1083) := b"0000000000000000_0000000000000000_0001100111111010_1010110100100101"; -- 0.10148126748623226
	pesos_i(1084) := b"0000000000000000_0000000000000000_0001101011000011_1001000100101100"; -- 0.10454661679182674
	pesos_i(1085) := b"0000000000000000_0000000000000000_0001011001100100_0000011011000110"; -- 0.08746378263288276
	pesos_i(1086) := b"0000000000000000_0000000000000000_0010001100111111_0001110010100010"; -- 0.13768176028969073
	pesos_i(1087) := b"0000000000000000_0000000000000000_0011001000011111_0000010011000010"; -- 0.19578580596167938
	pesos_i(1088) := b"1111111111111111_1111111111111111_1111000000010111_0111101110010111"; -- -0.062141681303501145
	pesos_i(1089) := b"0000000000000000_0000000000000000_0010011011011110_1100111111111010"; -- 0.1518373476402046
	pesos_i(1090) := b"0000000000000000_0000000000000000_0001100000000011_1101101110111010"; -- 0.09380887301061541
	pesos_i(1091) := b"1111111111111111_1111111111111111_1111000110110111_0011000001001101"; -- -0.05579851268291205
	pesos_i(1092) := b"1111111111111111_1111111111111111_1101111101100010_1000000110101111"; -- -0.12740315893032314
	pesos_i(1093) := b"0000000000000000_0000000000000000_0001010100011010_0011101110110001"; -- 0.08243153647482088
	pesos_i(1094) := b"0000000000000000_0000000000000000_0010110011101111_1001111000000011"; -- 0.17553126888886778
	pesos_i(1095) := b"1111111111111111_1111111111111111_1101100011000000_0000001101010101"; -- -0.15332011394312026
	pesos_i(1096) := b"0000000000000000_0000000000000000_0001000010010101_1110001100000011"; -- 0.0647870904606332
	pesos_i(1097) := b"0000000000000000_0000000000000000_0000100101000000_1110110101100001"; -- 0.03614696149822145
	pesos_i(1098) := b"0000000000000000_0000000000000000_0001101010010100_1011110101101111"; -- 0.1038320917882333
	pesos_i(1099) := b"0000000000000000_0000000000000000_0001000111011000_1011110101111110"; -- 0.06971344301231185
	pesos_i(1100) := b"0000000000000000_0000000000000000_0000100010000111_0110010001001001"; -- 0.033315913988632526
	pesos_i(1101) := b"0000000000000000_0000000000000000_0001011101110000_0000011011011110"; -- 0.09155314368494728
	pesos_i(1102) := b"0000000000000000_0000000000000000_0000000011100111_1001101001001001"; -- 0.003533976301165074
	pesos_i(1103) := b"1111111111111111_1111111111111111_1110001101100110_1111111101000000"; -- -0.1117096394601885
	pesos_i(1104) := b"1111111111111111_1111111111111111_1101011001101001_0101000100011000"; -- -0.16245549352907301
	pesos_i(1105) := b"0000000000000000_0000000000000000_0000001000001010_0101110111001101"; -- 0.007970678812188277
	pesos_i(1106) := b"0000000000000000_0000000000000000_0010011000011100_0000110010110111"; -- 0.14886550389172967
	pesos_i(1107) := b"1111111111111111_1111111111111111_1111010001010111_1010000100101000"; -- -0.045537879805916566
	pesos_i(1108) := b"0000000000000000_0000000000000000_0000101001101111_0001001111000101"; -- 0.0407574038913465
	pesos_i(1109) := b"0000000000000000_0000000000000000_0001011001110111_1110001101000111"; -- 0.08776684268341342
	pesos_i(1110) := b"1111111111111111_1111111111111111_1101101010111010_0001001100101000"; -- -0.14559822347038875
	pesos_i(1111) := b"0000000000000000_0000000000000000_0000100100000111_0101111010100100"; -- 0.03526870253841933
	pesos_i(1112) := b"1111111111111111_1111111111111111_1110101100101010_1101101101001111"; -- -0.0813773089408512
	pesos_i(1113) := b"1111111111111111_1111111111111111_1111101100101000_0100010100001011"; -- -0.018916783193475884
	pesos_i(1114) := b"0000000000000000_0000000000000000_0001000111000000_1001011011101101"; -- 0.06934493326921343
	pesos_i(1115) := b"1111111111111111_1111111111111111_1110000110010011_1001000001010101"; -- -0.11884210514799401
	pesos_i(1116) := b"1111111111111111_1111111111111111_1111111110110110_0111000010100110"; -- -0.0011224360054096197
	pesos_i(1117) := b"0000000000000000_0000000000000000_0000110100011010_1111011001010010"; -- 0.0511926604489079
	pesos_i(1118) := b"0000000000000000_0000000000000000_0010110100110100_1100001101000011"; -- 0.17658634553559108
	pesos_i(1119) := b"1111111111111111_1111111111111111_1111000001010001_0010000111010011"; -- -0.061262021903824085
	pesos_i(1120) := b"1111111111111111_1111111111111111_1110100000100101_1101100011010101"; -- -0.0931725005940282
	pesos_i(1121) := b"1111111111111111_1111111111111111_1101111001110011_0010010110101000"; -- -0.13105549484903997
	pesos_i(1122) := b"1111111111111111_1111111111111111_1111011100011011_1100010100000001"; -- -0.03473252038576531
	pesos_i(1123) := b"1111111111111111_1111111111111111_1111100000001111_0001100111000111"; -- -0.031019581662910845
	pesos_i(1124) := b"0000000000000000_0000000000000000_0000101101110110_1100110100111011"; -- 0.04478151974901622
	pesos_i(1125) := b"0000000000000000_0000000000000000_0001101101101100_0111001100110000"; -- 0.10712356491491445
	pesos_i(1126) := b"1111111111111111_1111111111111111_1111110010011010_0101001100111000"; -- -0.013270186359987338
	pesos_i(1127) := b"1111111111111111_1111111111111111_1101110000010111_1010001001111000"; -- -0.14026436399576522
	pesos_i(1128) := b"1111111111111111_1111111111111111_1110101010101000_0000010101001101"; -- -0.08337370748851744
	pesos_i(1129) := b"1111111111111111_1111111111111111_1111000110111000_0101100010001111"; -- -0.05578085440627674
	pesos_i(1130) := b"0000000000000000_0000000000000000_0000101101010110_0110100000001010"; -- 0.04428720703979871
	pesos_i(1131) := b"0000000000000000_0000000000000000_0010001110010001_0000001101010100"; -- 0.13893147283988627
	pesos_i(1132) := b"0000000000000000_0000000000000000_0001001100111111_1010000100101111"; -- 0.07518966097050211
	pesos_i(1133) := b"1111111111111111_1111111111111111_1111100100111100_1111001001101001"; -- -0.026413773814103644
	pesos_i(1134) := b"1111111111111111_1111111111111111_1101101101011111_1101101111000000"; -- -0.1430685669209774
	pesos_i(1135) := b"1111111111111111_1111111111111111_1110001011011000_0101111010001111"; -- -0.11388596552251337
	pesos_i(1136) := b"0000000000000000_0000000000000000_0001111110101110_1011101111110001"; -- 0.12375998142201602
	pesos_i(1137) := b"1111111111111111_1111111111111111_1111100101001000_0011101000010000"; -- -0.026241656297896113
	pesos_i(1138) := b"1111111111111111_1111111111111111_1101110000111001_0010100011110101"; -- -0.13975280790301667
	pesos_i(1139) := b"0000000000000000_0000000000000000_0001010111011010_1010101100001111"; -- 0.08536786201029656
	pesos_i(1140) := b"1111111111111111_1111111111111111_1111111111010001_0100101000000101"; -- -0.0007127512810992773
	pesos_i(1141) := b"1111111111111111_1111111111111111_1111110001001111_0011111101100000"; -- -0.014415778145021586
	pesos_i(1142) := b"1111111111111111_1111111111111111_1111110000101101_0101000100011001"; -- -0.014933520695321036
	pesos_i(1143) := b"0000000000000000_0000000000000000_0001000110111101_0101000000100000"; -- 0.06929493702103105
	pesos_i(1144) := b"0000000000000000_0000000000000000_0001111000001110_0110101110001011"; -- 0.11740753315287031
	pesos_i(1145) := b"1111111111111111_1111111111111111_1111000100011110_1011001111100001"; -- -0.0581252646125757
	pesos_i(1146) := b"0000000000000000_0000000000000000_0001100010111111_0011111111100001"; -- 0.09666823620750238
	pesos_i(1147) := b"1111111111111111_1111111111111111_1111000001101011_0010011001010010"; -- -0.06086502549881775
	pesos_i(1148) := b"1111111111111111_1111111111111111_1101011001100010_0000011101000101"; -- -0.16256670535804824
	pesos_i(1149) := b"1111111111111111_1111111111111111_1111111000101011_1101111111001110"; -- -0.007143032183832135
	pesos_i(1150) := b"1111111111111111_1111111111111111_1101111001000100_0100011011011101"; -- -0.13177067858064115
	pesos_i(1151) := b"1111111111111111_1111111111111111_1101101010000010_0001011001000111"; -- -0.1464525296973559
	pesos_i(1152) := b"0000000000000000_0000000000000000_0000000010011001_0011001010000111"; -- 0.002337606291235278
	pesos_i(1153) := b"1111111111111111_1111111111111111_1111111110101110_0010111101001001"; -- -0.0012484022681855513
	pesos_i(1154) := b"1111111111111111_1111111111111111_1110111110001010_0101101110110010"; -- -0.06429507168371348
	pesos_i(1155) := b"1111111111111111_1111111111111111_1101101001010111_0100001111010011"; -- -0.14710594268337482
	pesos_i(1156) := b"0000000000000000_0000000000000000_0001101110100001_0001111101010100"; -- 0.10792728241858524
	pesos_i(1157) := b"1111111111111111_1111111111111111_1110011101001010_1101001001111011"; -- -0.09651455410679612
	pesos_i(1158) := b"0000000000000000_0000000000000000_0000101010110010_0110010110011111"; -- 0.04178462144996392
	pesos_i(1159) := b"0000000000000000_0000000000000000_0000010110011111_0110100010000111"; -- 0.021963627715750316
	pesos_i(1160) := b"0000000000000000_0000000000000000_0001100110011111_1001101101100101"; -- 0.10009165973545638
	pesos_i(1161) := b"0000000000000000_0000000000000000_0000010010100000_0000111000110000"; -- 0.01806725183412221
	pesos_i(1162) := b"0000000000000000_0000000000000000_0000001011100011_1001110110000011"; -- 0.011285633537608782
	pesos_i(1163) := b"1111111111111111_1111111111111111_1111011001101011_0101000001101011"; -- -0.03742501622662745
	pesos_i(1164) := b"1111111111111111_1111111111111111_1110110111101111_0101111001100001"; -- -0.07056627394340169
	pesos_i(1165) := b"0000000000000000_0000000000000000_0001101111001111_1001101101100111"; -- 0.10863658192679479
	pesos_i(1166) := b"1111111111111111_1111111111111111_1101011011001001_0001011110001010"; -- -0.16099408031034487
	pesos_i(1167) := b"0000000000000000_0000000000000000_0001000110100101_1100000011011100"; -- 0.06893544541104417
	pesos_i(1168) := b"1111111111111111_1111111111111111_1111101000000000_1101000101010110"; -- -0.02342502267306884
	pesos_i(1169) := b"0000000000000000_0000000000000000_0001001101011100_1111110111101100"; -- 0.07563769357471141
	pesos_i(1170) := b"1111111111111111_1111111111111111_1111110011010010_0000001100001000"; -- -0.012420473568435394
	pesos_i(1171) := b"1111111111111111_1111111111111111_1111011010000101_0100110000110011"; -- -0.037028539306852445
	pesos_i(1172) := b"1111111111111111_1111111111111111_1111011000111011_1110000001001110"; -- -0.03814886175514512
	pesos_i(1173) := b"1111111111111111_1111111111111111_1101111100011000_1010111111100001"; -- -0.12852955581256797
	pesos_i(1174) := b"0000000000000000_0000000000000000_0000011110100111_0111100111101101"; -- 0.029899235060162194
	pesos_i(1175) := b"1111111111111111_1111111111111111_1111101010101101_0010110011011110"; -- -0.020795055254373782
	pesos_i(1176) := b"0000000000000000_0000000000000000_0001100100101011_0101000010010100"; -- 0.0983171808381428
	pesos_i(1177) := b"1111111111111111_1111111111111111_1101001000111001_1101010010101010"; -- -0.17880507327090908
	pesos_i(1178) := b"0000000000000000_0000000000000000_0001011100001100_0011101100000010"; -- 0.090030372642189
	pesos_i(1179) := b"1111111111111111_1111111111111111_1110001011110100_1100010111010010"; -- -0.11345256442257862
	pesos_i(1180) := b"1111111111111111_1111111111111111_1111011110010101_1011110010111110"; -- -0.032871440413394515
	pesos_i(1181) := b"1111111111111111_1111111111111111_1101111111011111_0010101000010110"; -- -0.125501031512598
	pesos_i(1182) := b"1111111111111111_1111111111111111_1111110100111000_1011001111110010"; -- -0.010853532321409579
	pesos_i(1183) := b"1111111111111111_1111111111111111_1101001111110101_1100100100010011"; -- -0.17203086162961373
	pesos_i(1184) := b"1111111111111111_1111111111111111_1101101001000001_0011101000000010"; -- -0.14744222118930397
	pesos_i(1185) := b"1111111111111111_1111111111111111_1110110000001010_0001110101111010"; -- -0.07797065521849962
	pesos_i(1186) := b"1111111111111111_1111111111111111_1101110101100100_1001110011111011"; -- -0.1351835142237894
	pesos_i(1187) := b"1111111111111111_1111111111111111_1111001001110001_1101100110100001"; -- -0.0529502851087421
	pesos_i(1188) := b"1111111111111111_1111111111111111_1110010100100110_0101000111001001"; -- -0.1048840413234074
	pesos_i(1189) := b"0000000000000000_0000000000000000_0001101111111001_1111111100011101"; -- 0.1092833945289607
	pesos_i(1190) := b"0000000000000000_0000000000000000_0001110000010001_1110001010000011"; -- 0.10964790052822307
	pesos_i(1191) := b"1111111111111111_1111111111111111_1111100001110111_1000100100011011"; -- -0.0294260320166585
	pesos_i(1192) := b"0000000000000000_0000000000000000_0001011110111000_0011100000001111"; -- 0.09265470862506978
	pesos_i(1193) := b"1111111111111111_1111111111111111_1111001011111000_0011001110010001"; -- -0.05090024673742306
	pesos_i(1194) := b"1111111111111111_1111111111111111_1110110111111001_0011111001001110"; -- -0.07041559797038667
	pesos_i(1195) := b"0000000000000000_0000000000000000_0001110101000101_0100001101110000"; -- 0.11433812600059691
	pesos_i(1196) := b"1111111111111111_1111111111111111_1110110111101011_0010110001010110"; -- -0.0706302919705694
	pesos_i(1197) := b"0000000000000000_0000000000000000_0010000010110000_1011100000101110"; -- 0.12769652484858343
	pesos_i(1198) := b"0000000000000000_0000000000000000_0001101111011000_1011100011100000"; -- 0.108775667914741
	pesos_i(1199) := b"1111111111111111_1111111111111111_1111101100100111_1010011000001110"; -- -0.018926259504240466
	pesos_i(1200) := b"1111111111111111_1111111111111111_1111100101010101_1010111001011010"; -- -0.026036360775222256
	pesos_i(1201) := b"0000000000000000_0000000000000000_0001111000001111_1111100000000011"; -- 0.1174311645692227
	pesos_i(1202) := b"1111111111111111_1111111111111111_1111011100011010_1110100110101111"; -- -0.03474559281429697
	pesos_i(1203) := b"0000000000000000_0000000000000000_0010100000000001_1110000100010100"; -- 0.15627867442538088
	pesos_i(1204) := b"1111111111111111_1111111111111111_1110010111111101_0000010110111011"; -- -0.10160793471692914
	pesos_i(1205) := b"0000000000000000_0000000000000000_0000010001001111_1100000100100011"; -- 0.016841956101475
	pesos_i(1206) := b"0000000000000000_0000000000000000_0000100001110000_1110101011011101"; -- 0.03297298334873026
	pesos_i(1207) := b"0000000000000000_0000000000000000_0000001000011101_0100101101101110"; -- 0.008259500952870653
	pesos_i(1208) := b"0000000000000000_0000000000000000_0000011101000110_0111111100100001"; -- 0.0284194426449996
	pesos_i(1209) := b"0000000000000000_0000000000000000_0001100001011010_1101000011101101"; -- 0.09513574386549578
	pesos_i(1210) := b"1111111111111111_1111111111111111_1110011101011110_1100000011100111"; -- -0.09621042594463389
	pesos_i(1211) := b"0000000000000000_0000000000000000_0010000000011001_1001101101110100"; -- 0.12539073539989848
	pesos_i(1212) := b"1111111111111111_1111111111111111_1111100111111011_1001010110001010"; -- -0.02350488064172348
	pesos_i(1213) := b"1111111111111111_1111111111111111_1111110101001000_1110111110011000"; -- -0.0106058363871168
	pesos_i(1214) := b"0000000000000000_0000000000000000_0000011000100100_1000011001001111"; -- 0.023994821795371015
	pesos_i(1215) := b"0000000000000000_0000000000000000_0010000111111100_1010101110000101"; -- 0.13276168826488907
	pesos_i(1216) := b"0000000000000000_0000000000000000_0010011011011100_0101101110111011"; -- 0.15179990112927946
	pesos_i(1217) := b"1111111111111111_1111111111111111_1111111100011011_1100000100110101"; -- -0.003482746655846362
	pesos_i(1218) := b"1111111111111111_1111111111111111_1111000100011000_1001010010000110"; -- -0.05821868628806524
	pesos_i(1219) := b"0000000000000000_0000000000000000_0000001101101010_0100111011100000"; -- 0.013340883040759598
	pesos_i(1220) := b"0000000000000000_0000000000000000_0000101111101101_0111001011001000"; -- 0.04659192449964596
	pesos_i(1221) := b"1111111111111111_1111111111111111_1101111111001001_0100111100000101"; -- -0.1258345234059421
	pesos_i(1222) := b"0000000000000000_0000000000000000_0001100001100100_1100110110111111"; -- 0.09528814226152477
	pesos_i(1223) := b"1111111111111111_1111111111111111_1111101001000011_1001001000110100"; -- -0.02240644666105325
	pesos_i(1224) := b"0000000000000000_0000000000000000_0011000100000001_1111111100010101"; -- 0.1914367127609186
	pesos_i(1225) := b"1111111111111111_1111111111111111_1111001111100000_0101111110011111"; -- -0.04735758177273395
	pesos_i(1226) := b"0000000000000000_0000000000000000_0001010111110011_1110100101101111"; -- 0.08575304956226039
	pesos_i(1227) := b"0000000000000000_0000000000000000_0001101101100100_1000000011011101"; -- 0.10700230983122339
	pesos_i(1228) := b"1111111111111111_1111111111111111_1110100100010011_0110010111010011"; -- -0.08954776371804739
	pesos_i(1229) := b"0000000000000000_0000000000000000_0001010010000010_1001100000011111"; -- 0.08011770977182944
	pesos_i(1230) := b"0000000000000000_0000000000000000_0001001111001011_0010111001000000"; -- 0.07731904088580577
	pesos_i(1231) := b"1111111111111111_1111111111111111_1111011100111101_0010011110100110"; -- -0.03422310070233853
	pesos_i(1232) := b"0000000000000000_0000000000000000_0000110011000101_1010001110111100"; -- 0.049890740838643505
	pesos_i(1233) := b"0000000000000000_0000000000000000_0000100110000100_1011001000101011"; -- 0.03718102975201969
	pesos_i(1234) := b"1111111111111111_1111111111111111_1101110110011001_1000011111001011"; -- -0.13437606142699438
	pesos_i(1235) := b"0000000000000000_0000000000000000_0001101111101100_0000001000000111"; -- 0.10906994508647856
	pesos_i(1236) := b"0000000000000000_0000000000000000_0010011011011111_1001000110011001"; -- 0.1518488883053215
	pesos_i(1237) := b"0000000000000000_0000000000000000_0000110010011110_1100110001111000"; -- 0.049298075869819075
	pesos_i(1238) := b"1111111111111111_1111111111111111_1111100001110100_1111000000000011"; -- -0.029465674709684808
	pesos_i(1239) := b"1111111111111111_1111111111111111_1110111001101001_1011000001111101"; -- -0.06869980772240818
	pesos_i(1240) := b"1111111111111111_1111111111111111_1111101101011001_0011101000111110"; -- -0.018169746245811004
	pesos_i(1241) := b"0000000000000000_0000000000000000_0001101100110011_1001100101111100"; -- 0.10625609651407723
	pesos_i(1242) := b"1111111111111111_1111111111111111_1110100101001010_0000001101000000"; -- -0.08871440592105213
	pesos_i(1243) := b"0000000000000000_0000000000000000_0010011110111110_1010011000010000"; -- 0.15525281812137737
	pesos_i(1244) := b"1111111111111111_1111111111111111_1111010100001110_0011001100000000"; -- -0.04275208701566593
	pesos_i(1245) := b"1111111111111111_1111111111111111_1111110001101110_0111011010110010"; -- -0.013939458436019125
	pesos_i(1246) := b"0000000000000000_0000000000000000_0001101000001110_1110000010001110"; -- 0.10178950760883991
	pesos_i(1247) := b"1111111111111111_1111111111111111_1110011000110010_0100110000000001"; -- -0.10079503034417492
	pesos_i(1248) := b"0000000000000000_0000000000000000_0001110010111001_0001011000110000"; -- 0.11219919849951057
	pesos_i(1249) := b"1111111111111111_1111111111111111_1110000100010011_1101110000000101"; -- -0.12079071892710082
	pesos_i(1250) := b"0000000000000000_0000000000000000_0010001101000101_0110010101101110"; -- 0.1377776522209121
	pesos_i(1251) := b"1111111111111111_1111111111111111_1111101000011010_1100100010100101"; -- -0.023028812208200515
	pesos_i(1252) := b"1111111111111111_1111111111111111_1111111101011111_0000110100010010"; -- -0.0024558859857456467
	pesos_i(1253) := b"0000000000000000_0000000000000000_0010001000010110_1001000100101111"; -- 0.13315684687259471
	pesos_i(1254) := b"1111111111111111_1111111111111111_1111010001101101_1000101110010110"; -- -0.04520347201525157
	pesos_i(1255) := b"0000000000000000_0000000000000000_0001001111010001_0111010000100110"; -- 0.07741475988826538
	pesos_i(1256) := b"0000000000000000_0000000000000000_0001010101001010_1111011011101000"; -- 0.08317511721125073
	pesos_i(1257) := b"0000000000000000_0000000000000000_0001100100110001_1011111000000011"; -- 0.09841525614942846
	pesos_i(1258) := b"1111111111111111_1111111111111111_1110111011000011_1011110101010001"; -- -0.06732575190912576
	pesos_i(1259) := b"0000000000000000_0000000000000000_0000100010101001_1111111110000010"; -- 0.03384396490834079
	pesos_i(1260) := b"0000000000000000_0000000000000000_0010011110110101_1011101001011010"; -- 0.1551166982414183
	pesos_i(1261) := b"1111111111111111_1111111111111111_1110111101111011_0001001000001001"; -- -0.0645283439174801
	pesos_i(1262) := b"0000000000000000_0000000000000000_0000100110101111_1110010101101010"; -- 0.037840212323099906
	pesos_i(1263) := b"1111111111111111_1111111111111111_1101110100011010_0010110010010100"; -- -0.13631936451358395
	pesos_i(1264) := b"1111111111111111_1111111111111111_1111110110110000_1011110100010001"; -- -0.009021933779509494
	pesos_i(1265) := b"1111111111111111_1111111111111111_1101101001010011_1011000101001100"; -- -0.14716045275534897
	pesos_i(1266) := b"1111111111111111_1111111111111111_1111000000001010_0100000011011010"; -- -0.062343546608620314
	pesos_i(1267) := b"1111111111111111_1111111111111111_1111000110010110_1000111010010001"; -- -0.05629643392429125
	pesos_i(1268) := b"0000000000000000_0000000000000000_0000011111101110_0001010000111110"; -- 0.030976548289499025
	pesos_i(1269) := b"0000000000000000_0000000000000000_0010000111000001_1100101100111111"; -- 0.1318633106804483
	pesos_i(1270) := b"0000000000000000_0000000000000000_0000100100001100_1111011100011110"; -- 0.035354084823807926
	pesos_i(1271) := b"1111111111111111_1111111111111111_1110110011010001_0011011000110110"; -- -0.07493268177281764
	pesos_i(1272) := b"0000000000000000_0000000000000000_0001111110010101_0000111101100000"; -- 0.123368225878742
	pesos_i(1273) := b"1111111111111111_1111111111111111_1101100001100000_1000000011001000"; -- -0.15477748026527466
	pesos_i(1274) := b"1111111111111111_1111111111111111_1101011111001001_1111110000100111"; -- -0.15707420390868845
	pesos_i(1275) := b"1111111111111111_1111111111111111_1110010010101101_1100110110100000"; -- -0.10672297323920263
	pesos_i(1276) := b"0000000000000000_0000000000000000_0010010101101010_1111010000100100"; -- 0.1461632334682011
	pesos_i(1277) := b"1111111111111111_1111111111111111_1111011011100010_0110101010100001"; -- -0.035607658204118764
	pesos_i(1278) := b"1111111111111111_1111111111111111_1111100001010100_1011111111000100"; -- -0.02995683168250412
	pesos_i(1279) := b"0000000000000000_0000000000000000_0001011000101111_1001000101001100"; -- 0.08666332356568919
	pesos_i(1280) := b"0000000000000000_0000000000000000_0000101011110010_1010111010010000"; -- 0.04276553159520349
	pesos_i(1281) := b"1111111111111111_1111111111111111_1111101100001001_0111011000011111"; -- -0.01938688039620407
	pesos_i(1282) := b"0000000000000000_0000000000000000_0000011001111010_0001100000100100"; -- 0.02530051119086736
	pesos_i(1283) := b"0000000000000000_0000000000000000_0001101111000101_1010000000001100"; -- 0.10848427093820602
	pesos_i(1284) := b"0000000000000000_0000000000000000_0001010111011001_1100010101110100"; -- 0.08535417635514109
	pesos_i(1285) := b"0000000000000000_0000000000000000_0000000101010000_0010010100110110"; -- 0.005129171115688733
	pesos_i(1286) := b"0000000000000000_0000000000000000_0001110111001111_1000111011001010"; -- 0.11644833026971015
	pesos_i(1287) := b"1111111111111111_1111111111111111_1101111011110101_0101001100100101"; -- -0.1290691409787865
	pesos_i(1288) := b"1111111111111111_1111111111111111_1111101111010011_1011111001001010"; -- -0.016300303398960492
	pesos_i(1289) := b"1111111111111111_1111111111111111_1101001110110001_0001011011110010"; -- -0.17307907667180744
	pesos_i(1290) := b"0000000000000000_0000000000000000_0000111001000100_0110011100011000"; -- 0.05573124247044859
	pesos_i(1291) := b"0000000000000000_0000000000000000_0010000010110101_1000100100010111"; -- 0.12777001199818228
	pesos_i(1292) := b"1111111111111111_1111111111111111_1101111101010100_0010111010010010"; -- -0.12762173588072945
	pesos_i(1293) := b"0000000000000000_0000000000000000_0001101110011100_1001110111111010"; -- 0.10785853718883537
	pesos_i(1294) := b"1111111111111111_1111111111111111_1111111110010011_1101011010000010"; -- -0.001650422304258596
	pesos_i(1295) := b"0000000000000000_0000000000000000_0010001011011010_1101010101011000"; -- 0.13615163219257878
	pesos_i(1296) := b"1111111111111111_1111111111111111_1101100110101110_1110100011001101"; -- -0.14967484459757321
	pesos_i(1297) := b"0000000000000000_0000000000000000_0000010011101110_1010001100111011"; -- 0.019266321106987203
	pesos_i(1298) := b"1111111111111111_1111111111111111_1101011110010000_1000001010011111"; -- -0.15795119871832328
	pesos_i(1299) := b"1111111111111111_1111111111111111_1101010110100000_0010100011111100"; -- -0.16552490085534596
	pesos_i(1300) := b"0000000000000000_0000000000000000_0010000110101010_1001101000000000"; -- 0.13150942323356501
	pesos_i(1301) := b"0000000000000000_0000000000000000_0010100011101100_1011001010000101"; -- 0.15986171473154762
	pesos_i(1302) := b"0000000000000000_0000000000000000_0001000000100000_1010010111111110"; -- 0.06299817522297732
	pesos_i(1303) := b"0000000000000000_0000000000000000_0001100111111011_0011101001111100"; -- 0.10148969207520638
	pesos_i(1304) := b"0000000000000000_0000000000000000_0000100101100000_1100110001001011"; -- 0.036633270604428024
	pesos_i(1305) := b"0000000000000000_0000000000000000_0000101011101001_1111111110001011"; -- 0.04263302947573486
	pesos_i(1306) := b"0000000000000000_0000000000000000_0001111011101101_0100001000110111"; -- 0.12080777973859788
	pesos_i(1307) := b"1111111111111111_1111111111111111_1101110000010100_0100010101010001"; -- -0.14031569254959636
	pesos_i(1308) := b"0000000000000000_0000000000000000_0010000101010000_0111010011100111"; -- 0.13013392102909663
	pesos_i(1309) := b"1111111111111111_1111111111111111_1101111011010110_0110001010011000"; -- -0.12954124256878652
	pesos_i(1310) := b"0000000000000000_0000000000000000_0010100110111111_1011100111001101"; -- 0.1630817532110542
	pesos_i(1311) := b"0000000000000000_0000000000000000_0000100001110011_0010101110100100"; -- 0.033007361892992026
	pesos_i(1312) := b"0000000000000000_0000000000000000_0010000011110001_0101000110100111"; -- 0.12868223496721462
	pesos_i(1313) := b"0000000000000000_0000000000000000_0000100001110111_0110110001100010"; -- 0.03307225592497272
	pesos_i(1314) := b"0000000000000000_0000000000000000_0000001111100000_0001001001001100"; -- 0.01513780936811522
	pesos_i(1315) := b"1111111111111111_1111111111111111_1111101011111000_1101010001110011"; -- -0.019640657293828176
	pesos_i(1316) := b"1111111111111111_1111111111111111_1111100000100111_1101011011001001"; -- -0.03064210507587653
	pesos_i(1317) := b"0000000000000000_0000000000000000_0001010001011101_1110100100011001"; -- 0.07955796102287715
	pesos_i(1318) := b"1111111111111111_1111111111111111_1111001100000001_0011111010010011"; -- -0.05076226158507875
	pesos_i(1319) := b"0000000000000000_0000000000000000_0001010100110110_1011010101110011"; -- 0.08286603983580107
	pesos_i(1320) := b"1111111111111111_1111111111111111_1101100001111001_1011001110001100"; -- -0.1543929847484598
	pesos_i(1321) := b"1111111111111111_1111111111111111_1111110111101001_1011101111111000"; -- -0.008152248225090418
	pesos_i(1322) := b"0000000000000000_0000000000000000_0001100110101001_1110011010010010"; -- 0.10024872835881014
	pesos_i(1323) := b"0000000000000000_0000000000000000_0000001011011000_1011111010011001"; -- 0.01111975898536505
	pesos_i(1324) := b"1111111111111111_1111111111111111_1110100111100111_0101001111101100"; -- -0.0863139675356131
	pesos_i(1325) := b"1111111111111111_1111111111111111_1111010000101001_0111010000101100"; -- -0.04624246516241446
	pesos_i(1326) := b"0000000000000000_0000000000000000_0010001101001111_1001000100100100"; -- 0.13793284531823757
	pesos_i(1327) := b"0000000000000000_0000000000000000_0001111100111101_0111001001011100"; -- 0.122031352558409
	pesos_i(1328) := b"1111111111111111_1111111111111111_1111110000001111_1100101011010100"; -- -0.015384028682761869
	pesos_i(1329) := b"1111111111111111_1111111111111111_1110111101100101_1001100001110001"; -- -0.06485602619204102
	pesos_i(1330) := b"0000000000000000_0000000000000000_0010100011010111_1001001100111010"; -- 0.1595394151242215
	pesos_i(1331) := b"1111111111111111_1111111111111111_1101100000000010_1010000010000001"; -- -0.15620991553856706
	pesos_i(1332) := b"1111111111111111_1111111111111111_1111110111110100_0000001110011101"; -- -0.0079953901395753
	pesos_i(1333) := b"0000000000000000_0000000000000000_0000010110100011_0111111001101000"; -- 0.022025966988561886
	pesos_i(1334) := b"1111111111111111_1111111111111111_1101011100111100_0000001110010000"; -- -0.15924051022625796
	pesos_i(1335) := b"0000000000000000_0000000000000000_0001110000011111_1111001000011100"; -- 0.1098624532522395
	pesos_i(1336) := b"1111111111111111_1111111111111111_1101010101001101_1101000110111110"; -- -0.1667813215247173
	pesos_i(1337) := b"1111111111111111_1111111111111111_1110010111111101_1111011110000101"; -- -0.10159352293875362
	pesos_i(1338) := b"1111111111111111_1111111111111111_1110010110000110_0101001101001101"; -- -0.10341910721826779
	pesos_i(1339) := b"1111111111111111_1111111111111111_1101011011111010_1111111011001100"; -- -0.16023261567707173
	pesos_i(1340) := b"0000000000000000_0000000000000000_0010000110010111_0110000010110000"; -- 0.13121609008728014
	pesos_i(1341) := b"1111111111111111_1111111111111111_1101011011100010_0001100010100110"; -- -0.16061254453472404
	pesos_i(1342) := b"1111111111111111_1111111111111111_1110111101001000_1110001111101110"; -- -0.06529403154036373
	pesos_i(1343) := b"0000000000000000_0000000000000000_0000000011000111_0011001010111111"; -- 0.003039523709191594
	pesos_i(1344) := b"1111111111111111_1111111111111111_1101111110011100_1110000101110101"; -- -0.12651244054235602
	pesos_i(1345) := b"1111111111111111_1111111111111111_1101101011011001_0000000000001111"; -- -0.14512633932571636
	pesos_i(1346) := b"0000000000000000_0000000000000000_0000110111100000_0100011000110010"; -- 0.05420340265978549
	pesos_i(1347) := b"1111111111111111_1111111111111111_1111100101011101_0100111110111000"; -- -0.025919931111506377
	pesos_i(1348) := b"1111111111111111_1111111111111111_1101110001101000_1100100110101111"; -- -0.13902606468108378
	pesos_i(1349) := b"0000000000000000_0000000000000000_0000000100001010_0100011111010111"; -- 0.0040631199246186425
	pesos_i(1350) := b"1111111111111111_1111111111111111_1111101001011111_0101111110101101"; -- -0.02198221232761423
	pesos_i(1351) := b"1111111111111111_1111111111111111_1110100111110101_0000001110011001"; -- -0.08610513235456653
	pesos_i(1352) := b"0000000000000000_0000000000000000_0010000001001110_0110001100011000"; -- 0.12619609201840892
	pesos_i(1353) := b"0000000000000000_0000000000000000_0000011101111110_0100001010011101"; -- 0.029270327953271547
	pesos_i(1354) := b"1111111111111111_1111111111111111_1101101101001100_0111000111011110"; -- -0.1433647950419243
	pesos_i(1355) := b"1111111111111111_1111111111111111_1111101010010010_1011001010111000"; -- -0.021199064412575432
	pesos_i(1356) := b"0000000000000000_0000000000000000_0000101110000000_1110000110110010"; -- 0.04493532742636473
	pesos_i(1357) := b"1111111111111111_1111111111111111_1110011001011001_1111011101111101"; -- -0.10018971640204155
	pesos_i(1358) := b"1111111111111111_1111111111111111_1101101011010100_1110101111100101"; -- -0.14518857634988988
	pesos_i(1359) := b"1111111111111111_1111111111111111_1100110100101101_0000010110101111"; -- -0.19853176573204492
	pesos_i(1360) := b"1111111111111111_1111111111111111_1110110000111011_0110111011111101"; -- -0.07721811593802522
	pesos_i(1361) := b"0000000000000000_0000000000000000_0010001110101111_0011011010001100"; -- 0.1393922893598111
	pesos_i(1362) := b"0000000000000000_0000000000000000_0000100111100001_1010011011101101"; -- 0.038599427136880984
	pesos_i(1363) := b"0000000000000000_0000000000000000_0010011111101001_1100011001110010"; -- 0.15591087618148874
	pesos_i(1364) := b"1111111111111111_1111111111111111_1111000000011100_1001011011110111"; -- -0.06206375574285512
	pesos_i(1365) := b"0000000000000000_0000000000000000_0001111010101110_0001100111001110"; -- 0.11984406745618574
	pesos_i(1366) := b"0000000000000000_0000000000000000_0000010111101111_1111100001110111"; -- 0.023192910198639692
	pesos_i(1367) := b"0000000000000000_0000000000000000_0001000010110001_0011100000101101"; -- 0.06520415410853125
	pesos_i(1368) := b"1111111111111111_1111111111111111_1111111011000111_0110011001010111"; -- -0.00476990113350311
	pesos_i(1369) := b"1111111111111111_1111111111111111_1110011111110001_1000010010110100"; -- -0.09397097209632463
	pesos_i(1370) := b"0000000000000000_0000000000000000_0000100001111011_1100100101100000"; -- 0.03313883404651477
	pesos_i(1371) := b"0000000000000000_0000000000000000_0010100111010101_1001101001010100"; -- 0.16341557065138315
	pesos_i(1372) := b"0000000000000000_0000000000000000_0010000001101001_0110000100101110"; -- 0.12660796524889512
	pesos_i(1373) := b"0000000000000000_0000000000000000_0000110110111001_1110110011010100"; -- 0.05361824197551446
	pesos_i(1374) := b"0000000000000000_0000000000000000_0010101101010011_0010010001010100"; -- 0.16923739492849355
	pesos_i(1375) := b"0000000000000000_0000000000000000_0000001010101100_1101110111110111"; -- 0.010450241814872419
	pesos_i(1376) := b"1111111111111111_1111111111111111_1101101101110110_0001011001000101"; -- -0.14272938558957052
	pesos_i(1377) := b"1111111111111111_1111111111111111_1111001110110000_0110100010111111"; -- -0.04808945973197331
	pesos_i(1378) := b"1111111111111111_1111111111111111_1110101011100001_0110101010110010"; -- -0.08249791285618134
	pesos_i(1379) := b"1111111111111111_1111111111111111_1110111110110111_1110100011010110"; -- -0.06360001345108039
	pesos_i(1380) := b"0000000000000000_0000000000000000_0010000010001000_1101000111000111"; -- 0.12708769890872404
	pesos_i(1381) := b"0000000000000000_0000000000000000_0001000010111100_0001010100000001"; -- 0.06536990423471094
	pesos_i(1382) := b"1111111111111111_1111111111111111_1110100010110010_0000010010101011"; -- -0.09103365740980116
	pesos_i(1383) := b"0000000000000000_0000000000000000_0000111100100011_1101111001100110"; -- 0.05914106358107599
	pesos_i(1384) := b"1111111111111111_1111111111111111_1101001100111100_1000001100011100"; -- -0.1748579079534582
	pesos_i(1385) := b"1111111111111111_1111111111111111_1111001010010001_1001111101001111"; -- -0.05246548012753523
	pesos_i(1386) := b"0000000000000000_0000000000000000_0001101010101001_0111110001011101"; -- 0.10414864792663685
	pesos_i(1387) := b"0000000000000000_0000000000000000_0010011001011111_0111010100011011"; -- 0.14989406497657315
	pesos_i(1388) := b"0000000000000000_0000000000000000_0010001100110100_0000110000010000"; -- 0.13751292598628106
	pesos_i(1389) := b"0000000000000000_0000000000000000_0001110001010000_1001001001001010"; -- 0.1106044226451222
	pesos_i(1390) := b"0000000000000000_0000000000000000_0010011011011101_1101011110101100"; -- 0.15182254731313724
	pesos_i(1391) := b"1111111111111111_1111111111111111_1101111101011110_1000001111000110"; -- -0.12746406944806116
	pesos_i(1392) := b"1111111111111111_1111111111111111_1110100110100111_0010111100000011"; -- -0.08729273000615706
	pesos_i(1393) := b"1111111111111111_1111111111111111_1111000111110010_1110110011110100"; -- -0.05488699958877671
	pesos_i(1394) := b"1111111111111111_1111111111111111_1101111011010010_1101001110010000"; -- -0.1295955442673766
	pesos_i(1395) := b"0000000000000000_0000000000000000_0010101101010000_1011100010011101"; -- 0.16920045698354272
	pesos_i(1396) := b"0000000000000000_0000000000000000_0010001110101000_0011011011101101"; -- 0.13928550041942656
	pesos_i(1397) := b"0000000000000000_0000000000000000_0000100110011101_0101100010000110"; -- 0.03755715623984721
	pesos_i(1398) := b"1111111111111111_1111111111111111_1111111001010100_1110100101000101"; -- -0.006516857884123608
	pesos_i(1399) := b"0000000000000000_0000000000000000_0001010010000010_1011111111010111"; -- 0.08012007720859987
	pesos_i(1400) := b"1111111111111111_1111111111111111_1111010110010000_1101111101100101"; -- -0.040758168910632275
	pesos_i(1401) := b"1111111111111111_1111111111111111_1111100111011111_1000000010000011"; -- -0.023933380147273493
	pesos_i(1402) := b"0000000000000000_0000000000000000_0000100110000110_1101001011110011"; -- 0.03721350139391898
	pesos_i(1403) := b"0000000000000000_0000000000000000_0000110000000010_0000010011010001"; -- 0.04690580454344309
	pesos_i(1404) := b"0000000000000000_0000000000000000_0000001111100101_0000011101100111"; -- 0.015213453829348073
	pesos_i(1405) := b"1111111111111111_1111111111111111_1110010100010011_0010000010100110"; -- -0.10517688699095049
	pesos_i(1406) := b"0000000000000000_0000000000000000_0001011000110000_1110001001111110"; -- 0.08668342178437871
	pesos_i(1407) := b"0000000000000000_0000000000000000_0001011011100010_1111111000001000"; -- 0.08940112773612881
	pesos_i(1408) := b"1111111111111111_1111111111111111_1111110010011001_1100010011101000"; -- -0.013278668862101356
	pesos_i(1409) := b"1111111111111111_1111111111111111_1111101111111000_1101101110011111"; -- -0.01573397976718499
	pesos_i(1410) := b"0000000000000000_0000000000000000_0010101100111100_1001111100101000"; -- 0.1688937637185877
	pesos_i(1411) := b"1111111111111111_1111111111111111_1101010010010001_0010000111010000"; -- -0.1696604601287605
	pesos_i(1412) := b"1111111111111111_1111111111111111_1110100011100010_1100011111001000"; -- -0.09028960572446644
	pesos_i(1413) := b"1111111111111111_1111111111111111_1110110111001101_1100000110101001"; -- -0.07107915518194273
	pesos_i(1414) := b"1111111111111111_1111111111111111_1101110110001000_0011001000001110"; -- -0.1346405710835612
	pesos_i(1415) := b"0000000000000000_0000000000000000_0001110001111001_1011010101111010"; -- 0.11123213025014736
	pesos_i(1416) := b"0000000000000000_0000000000000000_0001101001011001_0110001110111011"; -- 0.10292647666951618
	pesos_i(1417) := b"0000000000000000_0000000000000000_0001100111010011_1110001010000011"; -- 0.10088935567064004
	pesos_i(1418) := b"1111111111111111_1111111111111111_1110000110010001_0100100001111001"; -- -0.11887690595406261
	pesos_i(1419) := b"1111111111111111_1111111111111111_1111001011111111_1001001111010010"; -- -0.05078769796006155
	pesos_i(1420) := b"1111111111111111_1111111111111111_1111110011011110_0001100000011001"; -- -0.012236112504219994
	pesos_i(1421) := b"1111111111111111_1111111111111111_1101011110100011_1111101111010111"; -- -0.15765405652080303
	pesos_i(1422) := b"0000000000000000_0000000000000000_0000111101001001_0101010001000010"; -- 0.05971266376399204
	pesos_i(1423) := b"1111111111111111_1111111111111111_1101110111111000_1110011101011100"; -- -0.13292078021014284
	pesos_i(1424) := b"1111111111111111_1111111111111111_1101101111011011_0001111001001000"; -- -0.14118777028599544
	pesos_i(1425) := b"1111111111111111_1111111111111111_1110101101010001_0000111111100011"; -- -0.08079434107796146
	pesos_i(1426) := b"0000000000000000_0000000000000000_0010010111110000_0000110011110101"; -- 0.14819413166440615
	pesos_i(1427) := b"1111111111111111_1111111111111111_1110001110100001_1101100000011010"; -- -0.11081170422466279
	pesos_i(1428) := b"1111111111111111_1111111111111111_1111010100111100_1010010100111100"; -- -0.04204337391483849
	pesos_i(1429) := b"0000000000000000_0000000000000000_0001010001000000_0011100010101110"; -- 0.0791049408046827
	pesos_i(1430) := b"1111111111111111_1111111111111111_1111011010001100_0010101001001110"; -- -0.03692374805540363
	pesos_i(1431) := b"1111111111111111_1111111111111111_1110010100100110_1001100001000001"; -- -0.10487984092669289
	pesos_i(1432) := b"1111111111111111_1111111111111111_1101101010011000_0100111100010111"; -- -0.14611344983634847
	pesos_i(1433) := b"0000000000000000_0000000000000000_0001000101011011_0111101010000111"; -- 0.06780210292788551
	pesos_i(1434) := b"1111111111111111_1111111111111111_1110111001010010_0111011101001010"; -- -0.06905416901845901
	pesos_i(1435) := b"0000000000000000_0000000000000000_0000110000010101_1111010111010011"; -- 0.04721008672514851
	pesos_i(1436) := b"0000000000000000_0000000000000000_0010110000110111_1101010100111100"; -- 0.17272694325256105
	pesos_i(1437) := b"1111111111111111_1111111111111111_1101101011110111_1000011010111011"; -- -0.1446605485813584
	pesos_i(1438) := b"0000000000000000_0000000000000000_0010000111010011_1010100110000011"; -- 0.13213595807816175
	pesos_i(1439) := b"0000000000000000_0000000000000000_0000111000000011_1110111111011001"; -- 0.054747572380922344
	pesos_i(1440) := b"0000000000000000_0000000000000000_0001110110100101_0100101110110101"; -- 0.11580346266417416
	pesos_i(1441) := b"1111111111111111_1111111111111111_1111001100001110_1100110011000011"; -- -0.05055542211734372
	pesos_i(1442) := b"0000000000000000_0000000000000000_0001100010101101_1000000111110011"; -- 0.09639751599752817
	pesos_i(1443) := b"1111111111111111_1111111111111111_1101101000001010_1100011111011101"; -- -0.14827299934023624
	pesos_i(1444) := b"0000000000000000_0000000000000000_0010010001110010_0011110010100010"; -- 0.14236811585372422
	pesos_i(1445) := b"0000000000000000_0000000000000000_0000100110010000_1010101011110101"; -- 0.03736370537346079
	pesos_i(1446) := b"0000000000000000_0000000000000000_0000111111011001_0110000001101110"; -- 0.06191065491784439
	pesos_i(1447) := b"1111111111111111_1111111111111111_1101011111011011_0000101110110111"; -- -0.1568138770485229
	pesos_i(1448) := b"0000000000000000_0000000000000000_0001111001101001_1010011001111101"; -- 0.11879959633738671
	pesos_i(1449) := b"0000000000000000_0000000000000000_0010110011000011_0110010101011010"; -- 0.17485650497126082
	pesos_i(1450) := b"0000000000000000_0000000000000000_0000111110000110_0010010001100000"; -- 0.06064059589045318
	pesos_i(1451) := b"0000000000000000_0000000000000000_0010100010100011_0011011100010000"; -- 0.158740464689045
	pesos_i(1452) := b"0000000000000000_0000000000000000_0001000111101011_0010011000001110"; -- 0.06999433361438268
	pesos_i(1453) := b"0000000000000000_0000000000000000_0000101110110101_0101101101100010"; -- 0.04573603771667624
	pesos_i(1454) := b"0000000000000000_0000000000000000_0000101010110010_1001000111100101"; -- 0.0417872605573172
	pesos_i(1455) := b"0000000000000000_0000000000000000_0001101001111001_1111110001101000"; -- 0.10342385800253419
	pesos_i(1456) := b"1111111111111111_1111111111111111_1110001111010101_1000011110111000"; -- -0.1100230383587985
	pesos_i(1457) := b"0000000000000000_0000000000000000_0010000110011111_0111100101001101"; -- 0.13133962762100404
	pesos_i(1458) := b"0000000000000000_0000000000000000_0001110100011101_1101011011011110"; -- 0.11373656185135209
	pesos_i(1459) := b"1111111111111111_1111111111111111_1111001100001100_1000101010000111"; -- -0.05058988772443047
	pesos_i(1460) := b"0000000000000000_0000000000000000_0000001001101101_0111000101000000"; -- 0.009482458297754065
	pesos_i(1461) := b"1111111111111111_1111111111111111_1101100101101000_0110101000111100"; -- -0.15075050398587733
	pesos_i(1462) := b"1111111111111111_1111111111111111_1111001001110000_1011000010101100"; -- -0.05296798520231169
	pesos_i(1463) := b"1111111111111111_1111111111111111_1110000101011100_1001001110110100"; -- -0.11968113770344639
	pesos_i(1464) := b"1111111111111111_1111111111111111_1101101101111100_1011110010001000"; -- -0.14262792290802662
	pesos_i(1465) := b"0000000000000000_0000000000000000_0010011010111001_0111100111101000"; -- 0.15126764224580613
	pesos_i(1466) := b"0000000000000000_0000000000000000_0000011100110111_1001111000101000"; -- 0.028192410206378367
	pesos_i(1467) := b"1111111111111111_1111111111111111_1111111101111001_1110100001000011"; -- -0.0020460926212142174
	pesos_i(1468) := b"0000000000000000_0000000000000000_0000001001000000_1001001100110000"; -- 0.00879783550006186
	pesos_i(1469) := b"0000000000000000_0000000000000000_0000111100001001_1101010110011100"; -- 0.05874381113552146
	pesos_i(1470) := b"1111111111111111_1111111111111111_1111001101100000_1000010000110100"; -- -0.049308526407119246
	pesos_i(1471) := b"0000000000000000_0000000000000000_0001111011111000_1101101111001111"; -- 0.12098478141568982
	pesos_i(1472) := b"0000000000000000_0000000000000000_0001001100001101_0010101111101101"; -- 0.07441973253595566
	pesos_i(1473) := b"1111111111111111_1111111111111111_1111100101100101_0100001011011001"; -- -0.025798627958875563
	pesos_i(1474) := b"1111111111111111_1111111111111111_1101100000010000_1100010100111000"; -- -0.15599410418208484
	pesos_i(1475) := b"0000000000000000_0000000000000000_0001110111110000_0000111000000101"; -- 0.11694419507916474
	pesos_i(1476) := b"0000000000000000_0000000000000000_0001100001010000_0101110011101011"; -- 0.09497624151371147
	pesos_i(1477) := b"0000000000000000_0000000000000000_0000110100101110_0001111110000011"; -- 0.05148503263658059
	pesos_i(1478) := b"1111111111111111_1111111111111111_1110101110000100_0010001011111111"; -- -0.08001500382120623
	pesos_i(1479) := b"0000000000000000_0000000000000000_0001110000001110_0111101110101100"; -- 0.10959599454704713
	pesos_i(1480) := b"0000000000000000_0000000000000000_0000001001011001_1001001100001110"; -- 0.009179297353057512
	pesos_i(1481) := b"1111111111111111_1111111111111111_1110010000100001_0111101110011100"; -- -0.10886409216337593
	pesos_i(1482) := b"0000000000000000_0000000000000000_0001111000011101_1011000000000110"; -- 0.11764049667224935
	pesos_i(1483) := b"0000000000000000_0000000000000000_0001010111000011_1110110001110000"; -- 0.08502080661421133
	pesos_i(1484) := b"0000000000000000_0000000000000000_0001000101001111_0101011011101111"; -- 0.0676168758799843
	pesos_i(1485) := b"1111111111111111_1111111111111111_1111110000001101_1100101111110111"; -- -0.015414478544384654
	pesos_i(1486) := b"1111111111111111_1111111111111111_1111011000001111_1000110110111010"; -- -0.03882517055386468
	pesos_i(1487) := b"1111111111111111_1111111111111111_1111010101110010_1100101111010111"; -- -0.041217098327316695
	pesos_i(1488) := b"0000000000000000_0000000000000000_0010001010011000_0110001000111101"; -- 0.13513769128647227
	pesos_i(1489) := b"0000000000000000_0000000000000000_0001001011010100_1011111001101111"; -- 0.07355871403066844
	pesos_i(1490) := b"0000000000000000_0000000000000000_0000000011100010_0011100111000101"; -- 0.003451929616748911
	pesos_i(1491) := b"0000000000000000_0000000000000000_0001000111010000_0101100011001000"; -- 0.06958536999819209
	pesos_i(1492) := b"0000000000000000_0000000000000000_0001101011111101_0101100100011100"; -- 0.10542828496563426
	pesos_i(1493) := b"0000000000000000_0000000000000000_0010001010100110_0011111110101000"; -- 0.13534925312414234
	pesos_i(1494) := b"1111111111111111_1111111111111111_1110011111100000_0010111101111101"; -- -0.0942354508299196
	pesos_i(1495) := b"1111111111111111_1111111111111111_1110110101101101_0110000010110011"; -- -0.07254977825247401
	pesos_i(1496) := b"0000000000000000_0000000000000000_0010001100101110_0001000100101100"; -- 0.13742167775747346
	pesos_i(1497) := b"0000000000000000_0000000000000000_0010000011001000_1011110101100001"; -- 0.12806304568522994
	pesos_i(1498) := b"1111111111111111_1111111111111111_1101101110011011_0101110100010110"; -- -0.1421605892954243
	pesos_i(1499) := b"0000000000000000_0000000000000000_0010011001010011_0010000001100011"; -- 0.14970590986401788
	pesos_i(1500) := b"1111111111111111_1111111111111111_1110011010001110_1101101101110111"; -- -0.09938267075355905
	pesos_i(1501) := b"1111111111111111_1111111111111111_1110011011011100_1111010000011010"; -- -0.09819101680223177
	pesos_i(1502) := b"1111111111111111_1111111111111111_1111001000101010_1010001000101110"; -- -0.05403696413907124
	pesos_i(1503) := b"1111111111111111_1111111111111111_1110010110100010_0000000010101110"; -- -0.10299678559819266
	pesos_i(1504) := b"1111111111111111_1111111111111111_1101110011100100_0111011111001101"; -- -0.1371388553482898
	pesos_i(1505) := b"1111111111111111_1111111111111111_1101110100011110_1101110111011100"; -- -0.13624776246315656
	pesos_i(1506) := b"0000000000000000_0000000000000000_0001100101100100_0100101111101101"; -- 0.0991866544069247
	pesos_i(1507) := b"0000000000000000_0000000000000000_0010100101110000_0001001111101010"; -- 0.1618664214335292
	pesos_i(1508) := b"0000000000000000_0000000000000000_0001111001011010_0101011101111001"; -- 0.11856600472860077
	pesos_i(1509) := b"0000000000000000_0000000000000000_0001110101101011_1110001110101011"; -- 0.11492751051210386
	pesos_i(1510) := b"1111111111111111_1111111111111111_1110001110100110_0111010000001011"; -- -0.11074137424017433
	pesos_i(1511) := b"0000000000000000_0000000000000000_0000111111111001_0001101101110010"; -- 0.06239482424044315
	pesos_i(1512) := b"1111111111111111_1111111111111111_1111110101010001_1010110000111111"; -- -0.010472521309740968
	pesos_i(1513) := b"0000000000000000_0000000000000000_0000100101010111_1111100010000010"; -- 0.036498576953487794
	pesos_i(1514) := b"1111111111111111_1111111111111111_1110001110001000_1110101101101001"; -- -0.11119202323590589
	pesos_i(1515) := b"1111111111111111_1111111111111111_1101100100101101_1001101101011001"; -- -0.1516478451002289
	pesos_i(1516) := b"0000000000000000_0000000000000000_0001000000111111_1111010001000100"; -- 0.06347586302369615
	pesos_i(1517) := b"1111111111111111_1111111111111111_1101111101000100_0010100011111001"; -- -0.12786621027579462
	pesos_i(1518) := b"1111111111111111_1111111111111111_1110101011001001_1110111110000111"; -- -0.08285620637961842
	pesos_i(1519) := b"0000000000000000_0000000000000000_0000110111110100_1011110000110010"; -- 0.05451561174380962
	pesos_i(1520) := b"0000000000000000_0000000000000000_0010001111111011_0110111110011000"; -- 0.1405553575623215
	pesos_i(1521) := b"0000000000000000_0000000000000000_0000011100001111_1100101010000111"; -- 0.027584703324793763
	pesos_i(1522) := b"0000000000000000_0000000000000000_0010100000001111_0111100111000000"; -- 0.156486138766912
	pesos_i(1523) := b"0000000000000000_0000000000000000_0001011111110101_0001101001011001"; -- 0.09358372367532522
	pesos_i(1524) := b"0000000000000000_0000000000000000_0001101100100100_1010011001110011"; -- 0.10602798758140433
	pesos_i(1525) := b"1111111111111111_1111111111111111_1111100001111011_1101110101001011"; -- -0.02935997894010956
	pesos_i(1526) := b"0000000000000000_0000000000000000_0001111011111111_0000011100100001"; -- 0.12107891615746898
	pesos_i(1527) := b"0000000000000000_0000000000000000_0000011101011110_1101011111101010"; -- 0.028790945631174077
	pesos_i(1528) := b"1111111111111111_1111111111111111_1110110000001001_1010111000110011"; -- -0.07797728779619574
	pesos_i(1529) := b"0000000000000000_0000000000000000_0000101001001001_1001111111001110"; -- 0.040185916787461196
	pesos_i(1530) := b"1111111111111111_1111111111111111_1111110111111010_0111010010001110"; -- -0.007897105576707497
	pesos_i(1531) := b"0000000000000000_0000000000000000_0000101011001101_0110011010101110"; -- 0.04219667185280419
	pesos_i(1532) := b"1111111111111111_1111111111111111_1101110001011000_1010100101100000"; -- -0.13927213097206048
	pesos_i(1533) := b"1111111111111111_1111111111111111_1110010111100111_1100111010010111"; -- -0.10193165611859425
	pesos_i(1534) := b"1111111111111111_1111111111111111_1110110100101110_1010001011111111"; -- -0.07350713046353763
	pesos_i(1535) := b"0000000000000000_0000000000000000_0000010110000110_1000010001010101"; -- 0.021583815325923274
	pesos_i(1536) := b"0000000000000000_0000000000000000_0001001010001010_0010111011110001"; -- 0.07242101086843017
	pesos_i(1537) := b"1111111111111111_1111111111111111_1101000001010111_1110111100011110"; -- -0.18615823293427064
	pesos_i(1538) := b"1111111111111111_1111111111111111_1111001000001101_1001011110110001"; -- -0.05448009432882497
	pesos_i(1539) := b"1111111111111111_1111111111111111_1110101011111101_0100101110111111"; -- -0.08207251149910073
	pesos_i(1540) := b"0000000000000000_0000000000000000_0000110010011000_1000010000011111"; -- 0.049202211030093014
	pesos_i(1541) := b"0000000000000000_0000000000000000_0000011010111100_1110101101101101"; -- 0.026320184872515747
	pesos_i(1542) := b"1111111111111111_1111111111111111_1111000110010001_1100101110000001"; -- -0.056369095694087164
	pesos_i(1543) := b"1111111111111111_1111111111111111_1111001110110010_1100000100000000"; -- -0.04805368185775476
	pesos_i(1544) := b"1111111111111111_1111111111111111_1110101111111110_1010100100001011"; -- -0.07814544172620369
	pesos_i(1545) := b"1111111111111111_1111111111111111_1111111011001110_1000010110100101"; -- -0.004661223687441292
	pesos_i(1546) := b"0000000000000000_0000000000000000_0001110101000001_0111001110101011"; -- 0.11427996567288064
	pesos_i(1547) := b"1111111111111111_1111111111111111_1111010001100111_1101001110101101"; -- -0.04529072783678372
	pesos_i(1548) := b"0000000000000000_0000000000000000_0001111011011001_0110111101010110"; -- 0.12050529327281653
	pesos_i(1549) := b"1111111111111111_1111111111111111_1111011000101100_1100001011010111"; -- -0.038379500032615456
	pesos_i(1550) := b"1111111111111111_1111111111111111_1111001101001010_0010100110010001"; -- -0.04964962208533988
	pesos_i(1551) := b"1111111111111111_1111111111111111_1101101001001011_0000100001101111"; -- -0.14729258816141166
	pesos_i(1552) := b"0000000000000000_0000000000000000_0010010111111110_0100111011101010"; -- 0.1484116859573766
	pesos_i(1553) := b"0000000000000000_0000000000000000_0001100000111011_1001101000001100"; -- 0.0946594503813804
	pesos_i(1554) := b"0000000000000000_0000000000000000_0001011111110000_0010110011111101"; -- 0.09350854090866338
	pesos_i(1555) := b"1111111111111111_1111111111111111_1101110011110110_0000000011100101"; -- -0.1368712845938695
	pesos_i(1556) := b"0000000000000000_0000000000000000_0010001101111000_0100000011101110"; -- 0.13855367469847976
	pesos_i(1557) := b"1111111111111111_1111111111111111_1110000001101001_0100110011010001"; -- -0.12339324852928989
	pesos_i(1558) := b"1111111111111111_1111111111111111_1110011001101011_0111011000111001"; -- -0.0999227630375
	pesos_i(1559) := b"1111111111111111_1111111111111111_1111110101101010_1110000111010110"; -- -0.010087857463353852
	pesos_i(1560) := b"0000000000000000_0000000000000000_0010110010100101_1010001010001001"; -- 0.17440238792958937
	pesos_i(1561) := b"1111111111111111_1111111111111111_1110011011111110_0101110000011110"; -- -0.09768127689915708
	pesos_i(1562) := b"0000000000000000_0000000000000000_0001111010101000_1100110100100010"; -- 0.11976320341938296
	pesos_i(1563) := b"0000000000000000_0000000000000000_0010010100101100_1001100100001101"; -- 0.14521175923604768
	pesos_i(1564) := b"1111111111111111_1111111111111111_1111110011101100_1010011110010011"; -- -0.012013937677343016
	pesos_i(1565) := b"0000000000000000_0000000000000000_0010101101000010_0000100001011001"; -- 0.16897632765169393
	pesos_i(1566) := b"0000000000000000_0000000000000000_0001000000100111_1001100111010101"; -- 0.06310426198965498
	pesos_i(1567) := b"0000000000000000_0000000000000000_0001010011001000_1001101011110011"; -- 0.08118599339311414
	pesos_i(1568) := b"1111111111111111_1111111111111111_1110100001101001_0101111100110100"; -- -0.0921421525437715
	pesos_i(1569) := b"0000000000000000_0000000000000000_0001001010111010_0010001010111101"; -- 0.0731527052395837
	pesos_i(1570) := b"1111111111111111_1111111111111111_1110011000100101_0100000101101010"; -- -0.10099402586940837
	pesos_i(1571) := b"1111111111111111_1111111111111111_1111110010001001_1010001110011101"; -- -0.013524793883072001
	pesos_i(1572) := b"0000000000000000_0000000000000000_0010010101010010_0000111110001010"; -- 0.14578339700348228
	pesos_i(1573) := b"0000000000000000_0000000000000000_0001101111001101_0011111011010000"; -- 0.10860054570717927
	pesos_i(1574) := b"1111111111111111_1111111111111111_1101111101000110_1011000000011101"; -- -0.12782763768310035
	pesos_i(1575) := b"0000000000000000_0000000000000000_0001110101111011_1000100110111110"; -- 0.11516629104034723
	pesos_i(1576) := b"0000000000000000_0000000000000000_0001111111011000_1101100010010111"; -- 0.12440255830462102
	pesos_i(1577) := b"1111111111111111_1111111111111111_1110111101001111_0110100010111010"; -- -0.06519456336846631
	pesos_i(1578) := b"1111111111111111_1111111111111111_1101011000000001_0111100100010001"; -- -0.16404002510402696
	pesos_i(1579) := b"1111111111111111_1111111111111111_1101101101001111_1010010110100101"; -- -0.14331593244634977
	pesos_i(1580) := b"0000000000000000_0000000000000000_0000101011010001_0111110011010001"; -- 0.042259026534208224
	pesos_i(1581) := b"1111111111111111_1111111111111111_1101000100101101_0000111110101111"; -- -0.1829061696347009
	pesos_i(1582) := b"1111111111111111_1111111111111111_1101011100001010_1010100101110010"; -- -0.15999356226793737
	pesos_i(1583) := b"0000000000000000_0000000000000000_0010111001100000_1011011001000001"; -- 0.1811632070126796
	pesos_i(1584) := b"0000000000000000_0000000000000000_0010011101011111_0111000000000100"; -- 0.15380001161149878
	pesos_i(1585) := b"0000000000000000_0000000000000000_0000100011101101_1001010001011000"; -- 0.03487517487970226
	pesos_i(1586) := b"0000000000000000_0000000000000000_0001110010100011_0110010011001110"; -- 0.111868190970999
	pesos_i(1587) := b"1111111111111111_1111111111111111_1111100101000111_0011100011111110"; -- -0.026256978915797136
	pesos_i(1588) := b"1111111111111111_1111111111111111_1111000011101010_1101001111111001"; -- -0.0589168087744835
	pesos_i(1589) := b"1111111111111111_1111111111111111_1111111100111001_1011011110010111"; -- -0.003025556277480208
	pesos_i(1590) := b"0000000000000000_0000000000000000_0001010100100101_0100001010111110"; -- 0.08259980324522095
	pesos_i(1591) := b"0000000000000000_0000000000000000_0010111011010011_1110011010111011"; -- 0.18292085711260664
	pesos_i(1592) := b"0000000000000000_0000000000000000_0001111010100101_0010110001001001"; -- 0.11970783971480473
	pesos_i(1593) := b"0000000000000000_0000000000000000_0001100110101001_0010110101110111"; -- 0.10023769533250597
	pesos_i(1594) := b"0000000000000000_0000000000000000_0010001011101011_0111101010011110"; -- 0.13640562391927913
	pesos_i(1595) := b"0000000000000000_0000000000000000_0010100000010001_1000010001001000"; -- 0.15651728409901156
	pesos_i(1596) := b"1111111111111111_1111111111111111_1110011010100111_1000010000000001"; -- -0.09900641428655838
	pesos_i(1597) := b"1111111111111111_1111111111111111_1110100011100101_0011111110111111"; -- -0.09025193782503402
	pesos_i(1598) := b"1111111111111111_1111111111111111_1110000110100111_1000001101110010"; -- -0.11853769753300611
	pesos_i(1599) := b"1111111111111111_1111111111111111_1111011001101110_1101100010100001"; -- -0.03737112117899798
	pesos_i(1600) := b"1111111111111111_1111111111111111_1110000111010101_1001011100101100"; -- -0.11783461749366261
	pesos_i(1601) := b"0000000000000000_0000000000000000_0001000111011100_1000101101100100"; -- 0.06977149185673014
	pesos_i(1602) := b"0000000000000000_0000000000000000_0010001110011100_1101001111111111"; -- 0.13911175707394233
	pesos_i(1603) := b"1111111111111111_1111111111111111_1111010000101110_1111001011000011"; -- -0.04615862596451571
	pesos_i(1604) := b"0000000000000000_0000000000000000_0000110000101010_1010101001100010"; -- 0.047526024780223546
	pesos_i(1605) := b"0000000000000000_0000000000000000_0010000000011001_0001101110101010"; -- 0.12538311864532012
	pesos_i(1606) := b"1111111111111111_1111111111111111_1110111111000000_1001001000100111"; -- -0.06346785110083203
	pesos_i(1607) := b"1111111111111111_1111111111111111_1110001101010110_0110101001101011"; -- -0.11196265114164303
	pesos_i(1608) := b"0000000000000000_0000000000000000_0001111101110010_1011110001110100"; -- 0.12284448464915818
	pesos_i(1609) := b"0000000000000000_0000000000000000_0010101101001010_1000110110010101"; -- 0.16910633945087133
	pesos_i(1610) := b"1111111111111111_1111111111111111_1101011010110011_1010001111001111"; -- -0.16132141307001535
	pesos_i(1611) := b"1111111111111111_1111111111111111_1111111111101100_1011010101100010"; -- -0.00029436458121298326
	pesos_i(1612) := b"0000000000000000_0000000000000000_0010101001100010_0111011000000010"; -- 0.1655648951924642
	pesos_i(1613) := b"1111111111111111_1111111111111111_1101101101101111_1011001011101001"; -- -0.14282686051184482
	pesos_i(1614) := b"1111111111111111_1111111111111111_1101011010000001_1100011101010111"; -- -0.1620822345632368
	pesos_i(1615) := b"1111111111111111_1111111111111111_1111000010100101_1000110110001100"; -- -0.05997386306915585
	pesos_i(1616) := b"1111111111111111_1111111111111111_1110111000111011_1001101101001101"; -- -0.06940297485704491
	pesos_i(1617) := b"1111111111111111_1111111111111111_1101100101000111_0110111010010100"; -- -0.15125378511166063
	pesos_i(1618) := b"1111111111111111_1111111111111111_1111101101011100_0100110110110101"; -- -0.018122809686085567
	pesos_i(1619) := b"1111111111111111_1111111111111111_1111010010111000_1111110111111010"; -- -0.044052244737564646
	pesos_i(1620) := b"0000000000000000_0000000000000000_0001001110010101_0011100100010100"; -- 0.07649571159108653
	pesos_i(1621) := b"0000000000000000_0000000000000000_0001001100001010_0110011011110000"; -- 0.0743774734654623
	pesos_i(1622) := b"0000000000000000_0000000000000000_0001100100011110_1110011001110101"; -- 0.09812775002488817
	pesos_i(1623) := b"0000000000000000_0000000000000000_0000001100101111_0101000110101111"; -- 0.012440781750575326
	pesos_i(1624) := b"1111111111111111_1111111111111111_1101000101001110_1001101001110001"; -- -0.18239435910522767
	pesos_i(1625) := b"1111111111111111_1111111111111111_1101100101100100_1010100010010110"; -- -0.15080782266826473
	pesos_i(1626) := b"0000000000000000_0000000000000000_0001000000000110_1010100001100111"; -- 0.06260159037080251
	pesos_i(1627) := b"1111111111111111_1111111111111111_1110101100000110_0011101000011111"; -- -0.08193623299300233
	pesos_i(1628) := b"0000000000000000_0000000000000000_0001001111010111_0010010010011000"; -- 0.0775015707181565
	pesos_i(1629) := b"0000000000000000_0000000000000000_0010001100000110_0110110111111011"; -- 0.1368168581636795
	pesos_i(1630) := b"0000000000000000_0000000000000000_0001101010101011_1011111100010001"; -- 0.10418314146162916
	pesos_i(1631) := b"1111111111111111_1111111111111111_1101011101110110_0000011110110010"; -- -0.15835525427164257
	pesos_i(1632) := b"1111111111111111_1111111111111111_1111010001111110_0010101001010001"; -- -0.04494987037941697
	pesos_i(1633) := b"0000000000000000_0000000000000000_0000101001101001_1010111011001100"; -- 0.04067509156454189
	pesos_i(1634) := b"0000000000000000_0000000000000000_0010100011111000_0000101110100010"; -- 0.16003487314578102
	pesos_i(1635) := b"0000000000000000_0000000000000000_0001100011011011_1100010101111010"; -- 0.09710344522081768
	pesos_i(1636) := b"0000000000000000_0000000000000000_0001011111001010_0110100010001000"; -- 0.09293225595060478
	pesos_i(1637) := b"0000000000000000_0000000000000000_0001001000111110_1000010011001000"; -- 0.07126645933339879
	pesos_i(1638) := b"1111111111111111_1111111111111111_1111000110010001_1110010010110010"; -- -0.056367594208592116
	pesos_i(1639) := b"1111111111111111_1111111111111111_1110101110100011_0101111101011111"; -- -0.07953838280999884
	pesos_i(1640) := b"0000000000000000_0000000000000000_0010011001101011_0110101001000110"; -- 0.15007652475577085
	pesos_i(1641) := b"1111111111111111_1111111111111111_1110000110101011_0110000001001001"; -- -0.11847875807816005
	pesos_i(1642) := b"1111111111111111_1111111111111111_1111010111010111_1110011000110011"; -- -0.03967438951913745
	pesos_i(1643) := b"1111111111111111_1111111111111111_1111101001101100_1101010110111101"; -- -0.02177681100756982
	pesos_i(1644) := b"1111111111111111_1111111111111111_1111010101011101_1110101010000101"; -- -0.04153570408409577
	pesos_i(1645) := b"1111111111111111_1111111111111111_1111101100101111_1001100111011010"; -- -0.01880491656900183
	pesos_i(1646) := b"1111111111111111_1111111111111111_1101110001101010_1101001100001111"; -- -0.13899498831957208
	pesos_i(1647) := b"0000000000000000_0000000000000000_0000000101101001_1011011011101110"; -- 0.005519326309785933
	pesos_i(1648) := b"1111111111111111_1111111111111111_1111101110010100_0100111100111011"; -- -0.017268226808916542
	pesos_i(1649) := b"0000000000000000_0000000000000000_0001001001110100_0110010001011010"; -- 0.0720885010000439
	pesos_i(1650) := b"0000000000000000_0000000000000000_0001010010101111_1010101010101001"; -- 0.08080546025607255
	pesos_i(1651) := b"1111111111111111_1111111111111111_1101111101000011_0000010111101001"; -- -0.12788355876090512
	pesos_i(1652) := b"0000000000000000_0000000000000000_0010001111001101_0100011000001111"; -- 0.13985097753435793
	pesos_i(1653) := b"1111111111111111_1111111111111111_1111101011001101_1001010011100111"; -- -0.020300572978915528
	pesos_i(1654) := b"1111111111111111_1111111111111111_1101110111011000_1101110011000101"; -- -0.1334096925843481
	pesos_i(1655) := b"0000000000000000_0000000000000000_0000000101010100_0110001001000110"; -- 0.005193845823801729
	pesos_i(1656) := b"1111111111111111_1111111111111111_1110111011101110_1111010001000010"; -- -0.06666634923362731
	pesos_i(1657) := b"0000000000000000_0000000000000000_0001111011011111_0100010101001100"; -- 0.12059434034219793
	pesos_i(1658) := b"0000000000000000_0000000000000000_0010001011111100_0100111111110100"; -- 0.13666248051747515
	pesos_i(1659) := b"0000000000000000_0000000000000000_0001001010001110_1001011100010100"; -- 0.07248825300567227
	pesos_i(1660) := b"1111111111111111_1111111111111111_1111101111001011_1001100110010110"; -- -0.016424561479831547
	pesos_i(1661) := b"0000000000000000_0000000000000000_0000001010000001_0000101111110001"; -- 0.009781595442857333
	pesos_i(1662) := b"0000000000000000_0000000000000000_0010010000000000_0001000111111111"; -- 0.14062607264034713
	pesos_i(1663) := b"1111111111111111_1111111111111111_1111111110100110_0111011111010010"; -- -0.0013661492271885053
	pesos_i(1664) := b"1111111111111111_1111111111111111_1110000010100100_0000010101110011"; -- -0.122497233773259
	pesos_i(1665) := b"0000000000000000_0000000000000000_0001011000100101_1001110110100110"; -- 0.08651147178853008
	pesos_i(1666) := b"0000000000000000_0000000000000000_0001001100111011_1111101101100000"; -- 0.0751340017786345
	pesos_i(1667) := b"0000000000000000_0000000000000000_0000001101100011_1011000001000001"; -- 0.013239875659387548
	pesos_i(1668) := b"1111111111111111_1111111111111111_1110110001110110_1010101101000111"; -- -0.07631425387373018
	pesos_i(1669) := b"0000000000000000_0000000000000000_0010011011111101_1011101010111000"; -- 0.15230910298832026
	pesos_i(1670) := b"1111111111111111_1111111111111111_1110010111011100_0101001000110100"; -- -0.10210691668618345
	pesos_i(1671) := b"0000000000000000_0000000000000000_0000111110010001_1000100000010011"; -- 0.06081438505476355
	pesos_i(1672) := b"1111111111111111_1111111111111111_1101101010010110_0110010101011110"; -- -0.14614263960953777
	pesos_i(1673) := b"0000000000000000_0000000000000000_0000111010011010_1111101010101011"; -- 0.057052294450006834
	pesos_i(1674) := b"1111111111111111_1111111111111111_1101111010101000_1000011111101100"; -- -0.13024092195316753
	pesos_i(1675) := b"0000000000000000_0000000000000000_0010011011111000_0101010111100101"; -- 0.15222679935916228
	pesos_i(1676) := b"1111111111111111_1111111111111111_1101011101011100_0000111011011000"; -- -0.15875155674247246
	pesos_i(1677) := b"1111111111111111_1111111111111111_1111110101110010_0010110101110111"; -- -0.009976538205408269
	pesos_i(1678) := b"1111111111111111_1111111111111111_1111100000110010_1100100001011010"; -- -0.030475118586755424
	pesos_i(1679) := b"1111111111111111_1111111111111111_1111100010100101_1110111110110110"; -- -0.028718012015135578
	pesos_i(1680) := b"0000000000000000_0000000000000000_0010100111100010_0101001100110011"; -- 0.16360969550364426
	pesos_i(1681) := b"1111111111111111_1111111111111111_1101110010000101_0001101100000010"; -- -0.13859397126916925
	pesos_i(1682) := b"0000000000000000_0000000000000000_0010000100010111_0101111111001111"; -- 0.12926291275915416
	pesos_i(1683) := b"1111111111111111_1111111111111111_1111001110111100_0000001001111100"; -- -0.04791244946644244
	pesos_i(1684) := b"0000000000000000_0000000000000000_0000010001110001_0011100111110011"; -- 0.01735269711155372
	pesos_i(1685) := b"1111111111111111_1111111111111111_1101010011100001_0001100001110001"; -- -0.16844031572489973
	pesos_i(1686) := b"0000000000000000_0000000000000000_0001000110011101_0111110111011101"; -- 0.06880938180413204
	pesos_i(1687) := b"1111111111111111_1111111111111111_1100111001001101_0100010001101011"; -- -0.19413349514748343
	pesos_i(1688) := b"1111111111111111_1111111111111111_1101111010010100_1011000100100111"; -- -0.13054364015120679
	pesos_i(1689) := b"0000000000000000_0000000000000000_0000010100000101_0000101110110011"; -- 0.019608241158234372
	pesos_i(1690) := b"1111111111111111_1111111111111111_1111000011001100_1101100000100100"; -- -0.05937432393017713
	pesos_i(1691) := b"1111111111111111_1111111111111111_1110100101000111_1010100000110110"; -- -0.08875034978092226
	pesos_i(1692) := b"0000000000000000_0000000000000000_0000110101100111_0011010111111110"; -- 0.05235612354420385
	pesos_i(1693) := b"1111111111111111_1111111111111111_1110001001001110_0011100100100000"; -- -0.11599390958417267
	pesos_i(1694) := b"1111111111111111_1111111111111111_1110001001001010_1011010101101110"; -- -0.11604753562648328
	pesos_i(1695) := b"1111111111111111_1111111111111111_1111011101010011_0101010010110001"; -- -0.033884722585367205
	pesos_i(1696) := b"1111111111111111_1111111111111111_1101011001001011_0110001100000101"; -- -0.16291218870892316
	pesos_i(1697) := b"0000000000000000_0000000000000000_0000101100011111_1100101101110110"; -- 0.04345389972018923
	pesos_i(1698) := b"1111111111111111_1111111111111111_1111100100101001_0101111010111101"; -- -0.026712492844401747
	pesos_i(1699) := b"1111111111111111_1111111111111111_1110011001011111_0010100011011001"; -- -0.10011048021276733
	pesos_i(1700) := b"0000000000000000_0000000000000000_0010101110111100_1010110010110001"; -- 0.17084769550333187
	pesos_i(1701) := b"0000000000000000_0000000000000000_0000100101010101_1000111100111100"; -- 0.03646178450797864
	pesos_i(1702) := b"0000000000000000_0000000000000000_0000110000100111_1000001100100011"; -- 0.04747790915195806
	pesos_i(1703) := b"1111111111111111_1111111111111111_1111001111000101_1001111001001111"; -- -0.04776583254224803
	pesos_i(1704) := b"1111111111111111_1111111111111111_1110101101101100_0111101011111100"; -- -0.08037597028182111
	pesos_i(1705) := b"0000000000000000_0000000000000000_0001011011101001_1101101100001001"; -- 0.08950585331629737
	pesos_i(1706) := b"0000000000000000_0000000000000000_0001101001110110_0110110001001111"; -- 0.10336949286876392
	pesos_i(1707) := b"0000000000000000_0000000000000000_0000101011101010_0100011010000000"; -- 0.04263725870978892
	pesos_i(1708) := b"1111111111111111_1111111111111111_1111010011110110_1001110000001101"; -- -0.04311203653549442
	pesos_i(1709) := b"1111111111111111_1111111111111111_1110111010000111_0101010010110000"; -- -0.06824751578431343
	pesos_i(1710) := b"1111111111111111_1111111111111111_1110010011011111_0000001110100110"; -- -0.10597207254762298
	pesos_i(1711) := b"1111111111111111_1111111111111111_1111100110110111_0011000001000001"; -- -0.024548515486286414
	pesos_i(1712) := b"0000000000000000_0000000000000000_0000001111101111_0011100011000100"; -- 0.015368984103385358
	pesos_i(1713) := b"0000000000000000_0000000000000000_0001001110000111_0111010111001001"; -- 0.07628570711618393
	pesos_i(1714) := b"1111111111111111_1111111111111111_1111000010000100_0101010001100101"; -- -0.06048080956709835
	pesos_i(1715) := b"0000000000000000_0000000000000000_0000101110011110_1100100110001000"; -- 0.045391650766388125
	pesos_i(1716) := b"0000000000000000_0000000000000000_0000011100011101_0110011001000010"; -- 0.027792349836650472
	pesos_i(1717) := b"1111111111111111_1111111111111111_1110101101011110_0010000100100111"; -- -0.08059494778622878
	pesos_i(1718) := b"1111111111111111_1111111111111111_1111110011100010_0101011000011010"; -- -0.012171381586737893
	pesos_i(1719) := b"0000000000000000_0000000000000000_0000100000011011_0111111011010111"; -- 0.03166954762233951
	pesos_i(1720) := b"0000000000000000_0000000000000000_0000111000001101_1111101101010100"; -- 0.05490084468158957
	pesos_i(1721) := b"1111111111111111_1111111111111111_1110111100011000_1011001000110011"; -- -0.06602941758624375
	pesos_i(1722) := b"1111111111111111_1111111111111111_1110111101000010_0100000010001010"; -- -0.06539532319975083
	pesos_i(1723) := b"1111111111111111_1111111111111111_1111000010101100_1011101001011011"; -- -0.05986438073234359
	pesos_i(1724) := b"1111111111111111_1111111111111111_1110000011001010_1111001111110010"; -- -0.1219031842503005
	pesos_i(1725) := b"0000000000000000_0000000000000000_0001101011011001_0111010010010101"; -- 0.10488060599968406
	pesos_i(1726) := b"0000000000000000_0000000000000000_0010100101111110_1100011110010110"; -- 0.16209075357895067
	pesos_i(1727) := b"1111111111111111_1111111111111111_1111000101010110_1000110000010010"; -- -0.05727314522607506
	pesos_i(1728) := b"1111111111111111_1111111111111111_1111011000100111_1111000101101111"; -- -0.03845301661284323
	pesos_i(1729) := b"1111111111111111_1111111111111111_1101011100110110_0011111111101011"; -- -0.1593284656256263
	pesos_i(1730) := b"1111111111111111_1111111111111111_1101110101001110_1010001111010010"; -- -0.1355188000758308
	pesos_i(1731) := b"0000000000000000_0000000000000000_0001110100000011_1010101000101111"; -- 0.11333717007353517
	pesos_i(1732) := b"1111111111111111_1111111111111111_1111010010000001_1011011001110100"; -- -0.04489574116779477
	pesos_i(1733) := b"0000000000000000_0000000000000000_0010110000011011_1010111111011011"; -- 0.17229746916311714
	pesos_i(1734) := b"0000000000000000_0000000000000000_0001111110011011_1100110100110111"; -- 0.1234710940713675
	pesos_i(1735) := b"0000000000000000_0000000000000000_0000110110101111_0001010001100111"; -- 0.05345275427279884
	pesos_i(1736) := b"0000000000000000_0000000000000000_0001011010010010_0011011000110000"; -- 0.08816851300651578
	pesos_i(1737) := b"1111111111111111_1111111111111111_1101010011110101_1110101011000110"; -- -0.16812260311299998
	pesos_i(1738) := b"1111111111111111_1111111111111111_1111011010011001_0101111011100100"; -- -0.03672224944742039
	pesos_i(1739) := b"1111111111111111_1111111111111111_1111110011101011_0000010010010010"; -- -0.012038912057633843
	pesos_i(1740) := b"1111111111111111_1111111111111111_1110010111001000_1111011100011111"; -- -0.10240226267821327
	pesos_i(1741) := b"0000000000000000_0000000000000000_0010100101110110_1110010110100010"; -- 0.16197047419562854
	pesos_i(1742) := b"0000000000000000_0000000000000000_0001011001001010_0110101010100010"; -- 0.0870730061469591
	pesos_i(1743) := b"0000000000000000_0000000000000000_0001101010110101_0000110111010000"; -- 0.10432516414759743
	pesos_i(1744) := b"1111111111111111_1111111111111111_1111010101011000_0110000100101010"; -- -0.04162018522555008
	pesos_i(1745) := b"1111111111111111_1111111111111111_1111100100111111_1100110110010111"; -- -0.026370192116421866
	pesos_i(1746) := b"0000000000000000_0000000000000000_0000111110100001_1100111111001001"; -- 0.06106280000717198
	pesos_i(1747) := b"1111111111111111_1111111111111111_1111001001011010_0001111111100100"; -- -0.05331230814613898
	pesos_i(1748) := b"0000000000000000_0000000000000000_0010000001100101_0111000000010011"; -- 0.12654781793751385
	pesos_i(1749) := b"1111111111111111_1111111111111111_1101100100110100_1110011100011110"; -- -0.1515365172085427
	pesos_i(1750) := b"0000000000000000_0000000000000000_0000111101111000_1110000100110010"; -- 0.0604382273159712
	pesos_i(1751) := b"0000000000000000_0000000000000000_0000101111001101_0001001001011111"; -- 0.046097896716454353
	pesos_i(1752) := b"1111111111111111_1111111111111111_1111001011100111_0111000000101011"; -- -0.051156034099918465
	pesos_i(1753) := b"1111111111111111_1111111111111111_1110101111110011_1001111000010010"; -- -0.07831394252674984
	pesos_i(1754) := b"1111111111111111_1111111111111111_1101011000100101_0110101000100100"; -- -0.16349159834058172
	pesos_i(1755) := b"0000000000000000_0000000000000000_0000011001011001_1110001111111001"; -- 0.024809120459511946
	pesos_i(1756) := b"0000000000000000_0000000000000000_0010000111110011_1001110111101100"; -- 0.1326235486777246
	pesos_i(1757) := b"0000000000000000_0000000000000000_0001111100001101_1001010110100101"; -- 0.12130103366063097
	pesos_i(1758) := b"1111111111111111_1111111111111111_1111010001111001_1010011010111111"; -- -0.045018747792254586
	pesos_i(1759) := b"0000000000000000_0000000000000000_0010000110011011_1000110101100010"; -- 0.13127978934532133
	pesos_i(1760) := b"1111111111111111_1111111111111111_1110011110001100_1101000111111010"; -- -0.09550750388797836
	pesos_i(1761) := b"0000000000000000_0000000000000000_0001110011000101_1011011010000001"; -- 0.1123918594842255
	pesos_i(1762) := b"1111111111111111_1111111111111111_1101110101110000_1001110010110001"; -- -0.13500042610885793
	pesos_i(1763) := b"0000000000000000_0000000000000000_0000010010111001_0100000001011110"; -- 0.018451712597916333
	pesos_i(1764) := b"0000000000000000_0000000000000000_0010000111010111_0001111110101000"; -- 0.1321887765563023
	pesos_i(1765) := b"1111111111111111_1111111111111111_1110011100001101_0101010001011101"; -- -0.09745285723470995
	pesos_i(1766) := b"0000000000000000_0000000000000000_0000111000100100_1100101010000110"; -- 0.05524888771111467
	pesos_i(1767) := b"1111111111111111_1111111111111111_1111101100111000_1111000000001010"; -- -0.018662450407631148
	pesos_i(1768) := b"1111111111111111_1111111111111111_1101111110100101_0100100010010010"; -- -0.12638422429838198
	pesos_i(1769) := b"1111111111111111_1111111111111111_1110010000100101_1111011001001100"; -- -0.10879574430371376
	pesos_i(1770) := b"1111111111111111_1111111111111111_1111010110000111_0010100000110011"; -- -0.04090641751498286
	pesos_i(1771) := b"0000000000000000_0000000000000000_0000011110111101_1000011111011111"; -- 0.03023575959925087
	pesos_i(1772) := b"1111111111111111_1111111111111111_1110000001101100_0010110000100001"; -- -0.12334942050056123
	pesos_i(1773) := b"0000000000000000_0000000000000000_0000010010100110_1001010000111000"; -- 0.018166793613920734
	pesos_i(1774) := b"0000000000000000_0000000000000000_0000000011110110_1001011010001100"; -- 0.0037626353157841613
	pesos_i(1775) := b"1111111111111111_1111111111111111_1101110100110111_0011000011111101"; -- -0.1358765965583113
	pesos_i(1776) := b"0000000000000000_0000000000000000_0010100010100001_1011001011000000"; -- 0.15871731925290158
	pesos_i(1777) := b"1111111111111111_1111111111111111_1101100100011001_1001000101101000"; -- -0.15195361330994867
	pesos_i(1778) := b"0000000000000000_0000000000000000_0000100100011000_0111100111011001"; -- 0.035529723548524385
	pesos_i(1779) := b"0000000000000000_0000000000000000_0010010000010101_1110000001001111"; -- 0.14095880431426588
	pesos_i(1780) := b"1111111111111111_1111111111111111_1101010011000101_0011000010111000"; -- -0.16886611468830187
	pesos_i(1781) := b"1111111111111111_1111111111111111_1111010110111101_0111000001011001"; -- -0.040078142477419455
	pesos_i(1782) := b"1111111111111111_1111111111111111_1111100000010000_0101101001001111"; -- -0.031000476678396865
	pesos_i(1783) := b"1111111111111111_1111111111111111_1111010100010011_1010000011101110"; -- -0.04266924088583227
	pesos_i(1784) := b"0000000000000000_0000000000000000_0000101010001100_1011111111100111"; -- 0.041210168649053525
	pesos_i(1785) := b"1111111111111111_1111111111111111_1101100000010000_0010101100001011"; -- -0.15600329372667626
	pesos_i(1786) := b"1111111111111111_1111111111111111_1101101000111110_0001101000100000"; -- -0.14748989794568867
	pesos_i(1787) := b"0000000000000000_0000000000000000_0010000000110110_1101010001100010"; -- 0.1258366336592297
	pesos_i(1788) := b"1111111111111111_1111111111111111_1111111100000101_0001100100001111"; -- -0.003828462415301818
	pesos_i(1789) := b"0000000000000000_0000000000000000_0000011010010101_0101000010100010"; -- 0.025715865763377817
	pesos_i(1790) := b"0000000000000000_0000000000000000_0001001110011111_0010000101101101"; -- 0.07664688985657614
	pesos_i(1791) := b"0000000000000000_0000000000000000_0000010011101011_1110101010110011"; -- 0.019224804598258004
	pesos_i(1792) := b"0000000000000000_0000000000000000_0010000111001001_0111111001010010"; -- 0.13198079586838893
	pesos_i(1793) := b"1111111111111111_1111111111111111_1101001111100010_1110100101001010"; -- -0.1723188586704799
	pesos_i(1794) := b"1111111111111111_1111111111111111_1111000011110111_1010110110011001"; -- -0.0587207318377147
	pesos_i(1795) := b"0000000000000000_0000000000000000_0001000101011011_1010101000001000"; -- 0.06780493444588742
	pesos_i(1796) := b"1111111111111111_1111111111111111_1101111001101010_0001001111011110"; -- -0.13119388410074398
	pesos_i(1797) := b"1111111111111111_1111111111111111_1111101111101100_0110100010111110"; -- -0.015923932601687146
	pesos_i(1798) := b"0000000000000000_0000000000000000_0010001001011000_1111011001010100"; -- 0.13416995565659845
	pesos_i(1799) := b"0000000000000000_0000000000000000_0001111000011111_1100110100010101"; -- 0.11767274620009865
	pesos_i(1800) := b"1111111111111111_1111111111111111_1111011101110011_1101111101000000"; -- -0.03338818249570981
	pesos_i(1801) := b"1111111111111111_1111111111111111_1101011010011001_1011101110111001"; -- -0.16171671604433832
	pesos_i(1802) := b"0000000000000000_0000000000000000_0000011101110101_0100010010100110"; -- 0.02913312008329773
	pesos_i(1803) := b"0000000000000000_0000000000000000_0010101010110111_1011110010000100"; -- 0.16686609482763168
	pesos_i(1804) := b"1111111111111111_1111111111111111_1110100100111001_0011001100111111"; -- -0.08897094445600502
	pesos_i(1805) := b"0000000000000000_0000000000000000_0010101101001010_0111101001001011"; -- 0.1691051896273272
	pesos_i(1806) := b"0000000000000000_0000000000000000_0000001010000011_1001110101111100"; -- 0.009820788202911641
	pesos_i(1807) := b"1111111111111111_1111111111111111_1100111010110111_1111000011001101"; -- -0.1925057887898869
	pesos_i(1808) := b"1111111111111111_1111111111111111_1111000010010110_0101011000111000"; -- -0.06020604259451859
	pesos_i(1809) := b"1111111111111111_1111111111111111_1110111011001111_1010100101100110"; -- -0.06714383377147304
	pesos_i(1810) := b"0000000000000000_0000000000000000_0001011001000101_1100001001111110"; -- 0.08700194904791758
	pesos_i(1811) := b"0000000000000000_0000000000000000_0001101001011110_1011011100000011"; -- 0.10300773455901709
	pesos_i(1812) := b"0000000000000000_0000000000000000_0000101000101001_1100111111011010"; -- 0.039700499174571635
	pesos_i(1813) := b"0000000000000000_0000000000000000_0001111100100011_1011101101001110"; -- 0.12163897178972698
	pesos_i(1814) := b"0000000000000000_0000000000000000_0001100011100001_0101000101010000"; -- 0.09718807421213115
	pesos_i(1815) := b"1111111111111111_1111111111111111_1101111111101000_0100001011101111"; -- -0.12536222130813082
	pesos_i(1816) := b"0000000000000000_0000000000000000_0001111010100001_1101000110111111"; -- 0.1196566668171128
	pesos_i(1817) := b"0000000000000000_0000000000000000_0010000010110100_0000010100101011"; -- 0.12774689014179366
	pesos_i(1818) := b"1111111111111111_1111111111111111_1111010100111011_0011010001110100"; -- -0.04206535508587636
	pesos_i(1819) := b"1111111111111111_1111111111111111_1111101111100110_1001100000101111"; -- -0.016012657719384572
	pesos_i(1820) := b"0000000000000000_0000000000000000_0001100000101110_1110101100111010"; -- 0.09446592499151243
	pesos_i(1821) := b"0000000000000000_0000000000000000_0000100001111010_0111000111111111"; -- 0.03311836684803099
	pesos_i(1822) := b"1111111111111111_1111111111111111_1101011010000100_0111010001000001"; -- -0.16204141063678823
	pesos_i(1823) := b"0000000000000000_0000000000000000_0001101010010000_0000100010000111"; -- 0.10376027386071404
	pesos_i(1824) := b"1111111111111111_1111111111111111_1110011110111101_0100011000010001"; -- -0.09476816265617055
	pesos_i(1825) := b"0000000000000000_0000000000000000_0000010000000000_0001000000110100"; -- 0.01562596587044637
	pesos_i(1826) := b"0000000000000000_0000000000000000_0000000001111011_0111001110011110"; -- 0.0018837223665772614
	pesos_i(1827) := b"0000000000000000_0000000000000000_0000001000000110_0110101001011110"; -- 0.007910392742396985
	pesos_i(1828) := b"1111111111111111_1111111111111111_1101100101101001_0101001000001100"; -- -0.1507366868305642
	pesos_i(1829) := b"1111111111111111_1111111111111111_1110011101110100_0100110111100101"; -- -0.09588158756727669
	pesos_i(1830) := b"1111111111111111_1111111111111111_1101110111100111_1111011101001010"; -- -0.1331792301318111
	pesos_i(1831) := b"1111111111111111_1111111111111111_1101011011001011_0010110101010011"; -- -0.16096226434238015
	pesos_i(1832) := b"0000000000000000_0000000000000000_0001010110111111_1000001100000001"; -- 0.08495348712463299
	pesos_i(1833) := b"1111111111111111_1111111111111111_1101110110010100_1110001010011111"; -- -0.13444694150812841
	pesos_i(1834) := b"1111111111111111_1111111111111111_1111111110000100_1111000101001010"; -- -0.0018777079177558942
	pesos_i(1835) := b"0000000000000000_0000000000000000_0000010010000000_1011111011101110"; -- 0.017589505386794945
	pesos_i(1836) := b"0000000000000000_0000000000000000_0001010101110001_0111100001100011"; -- 0.08376266888485796
	pesos_i(1837) := b"1111111111111111_1111111111111111_1110111001000000_1101111010010000"; -- -0.06932267174191926
	pesos_i(1838) := b"1111111111111111_1111111111111111_1110100000011010_1000000011011101"; -- -0.093345590598226
	pesos_i(1839) := b"0000000000000000_0000000000000000_0000011010010011_0011110101000001"; -- 0.025684193085950005
	pesos_i(1840) := b"1111111111111111_1111111111111111_1101011101000101_0110110111001100"; -- -0.15909684915307198
	pesos_i(1841) := b"0000000000000000_0000000000000000_0001001001111000_0001000111100010"; -- 0.07214462059819689
	pesos_i(1842) := b"0000000000000000_0000000000000000_0001001111010101_1111110001010000"; -- 0.07748391116804505
	pesos_i(1843) := b"0000000000000000_0000000000000000_0010010111000011_0010100101010110"; -- 0.14750917758238014
	pesos_i(1844) := b"1111111111111111_1111111111111111_1111101001100011_0011101100010000"; -- -0.021923359427500105
	pesos_i(1845) := b"0000000000000000_0000000000000000_0001100111100010_1001110011001000"; -- 0.10111408116455944
	pesos_i(1846) := b"1111111111111111_1111111111111111_1111101100011010_0001000000101101"; -- -0.019133557345113687
	pesos_i(1847) := b"0000000000000000_0000000000000000_0001110101111000_0000011111100111"; -- 0.11511277577092394
	pesos_i(1848) := b"1111111111111111_1111111111111111_1110101100111001_1110101101000111"; -- -0.08114747545236695
	pesos_i(1849) := b"1111111111111111_1111111111111111_1111110110111111_1110101000000111"; -- -0.008790372276924717
	pesos_i(1850) := b"1111111111111111_1111111111111111_1101100111111000_1101101000000100"; -- -0.148546575475651
	pesos_i(1851) := b"1111111111111111_1111111111111111_1101110000100110_1101110000010101"; -- -0.14003204815189385
	pesos_i(1852) := b"1111111111111111_1111111111111111_1111110100110111_1101111111010111"; -- -0.010866174757844741
	pesos_i(1853) := b"0000000000000000_0000000000000000_0000010011001011_0011000101011010"; -- 0.018725475847672826
	pesos_i(1854) := b"0000000000000000_0000000000000000_0000011100100110_0111101111101001"; -- 0.027930969571676605
	pesos_i(1855) := b"0000000000000000_0000000000000000_0010000101011100_0111001010000110"; -- 0.13031688475080883
	pesos_i(1856) := b"0000000000000000_0000000000000000_0010000010110111_0101110100111111"; -- 0.12779791626613632
	pesos_i(1857) := b"1111111111111111_1111111111111111_1101011000111110_1011101100111111"; -- -0.16310529439657676
	pesos_i(1858) := b"1111111111111111_1111111111111111_1111000001111110_1110011001010001"; -- -0.060563664644403714
	pesos_i(1859) := b"0000000000000000_0000000000000000_0000111110000110_1111100101011001"; -- 0.06065329010372004
	pesos_i(1860) := b"0000000000000000_0000000000000000_0001100111001001_0110011011100000"; -- 0.10072939846203788
	pesos_i(1861) := b"0000000000000000_0000000000000000_0010000111000001_1110111101010111"; -- 0.1318654620006511
	pesos_i(1862) := b"1111111111111111_1111111111111111_1110000100001011_0110100101111110"; -- -0.12091961557833697
	pesos_i(1863) := b"1111111111111111_1111111111111111_1101101011001111_1000010010010001"; -- -0.1452710289931798
	pesos_i(1864) := b"1111111111111111_1111111111111111_1110110000000000_1011010111011001"; -- -0.07811416105391421
	pesos_i(1865) := b"0000000000000000_0000000000000000_0001100011010010_1001111000010101"; -- 0.09696376824046417
	pesos_i(1866) := b"1111111111111111_1111111111111111_1111111100111001_0111010010000111"; -- -0.003029553355061769
	pesos_i(1867) := b"1111111111111111_1111111111111111_1111000111000010_1011110010000100"; -- -0.05562230852232404
	pesos_i(1868) := b"1111111111111111_1111111111111111_1110010011110001_1111010011001110"; -- -0.10568304045056634
	pesos_i(1869) := b"1111111111111111_1111111111111111_1111110101000001_1101011001011111"; -- -0.010714151281509496
	pesos_i(1870) := b"0000000000000000_0000000000000000_0000001110100111_0010010000110111"; -- 0.014269126253154789
	pesos_i(1871) := b"1111111111111111_1111111111111111_1111101100011101_0110110111001100"; -- -0.01908220060890086
	pesos_i(1872) := b"0000000000000000_0000000000000000_0010101101100101_0000110000011110"; -- 0.16951060998284387
	pesos_i(1873) := b"1111111111111111_1111111111111111_1101011110000010_1110000010101111"; -- -0.15815921529573296
	pesos_i(1874) := b"1111111111111111_1111111111111111_1110101011001110_1101111101010010"; -- -0.08278087863657863
	pesos_i(1875) := b"1111111111111111_1111111111111111_1110011110101011_1010100011000011"; -- -0.095036938196234
	pesos_i(1876) := b"1111111111111111_1111111111111111_1110011101011101_0100110111111010"; -- -0.09623253485517387
	pesos_i(1877) := b"0000000000000000_0000000000000000_0010011101111000_1111111100011111"; -- 0.15419001119887388
	pesos_i(1878) := b"1111111111111111_1111111111111111_1110110011010011_0000100010011001"; -- -0.0749048831548542
	pesos_i(1879) := b"0000000000000000_0000000000000000_0001101110001100_1110100000011111"; -- 0.10761881592090725
	pesos_i(1880) := b"1111111111111111_1111111111111111_1111110010110000_1100001100100000"; -- -0.012927822809858271
	pesos_i(1881) := b"0000000000000000_0000000000000000_0001000101101101_0111000001000010"; -- 0.06807614907806729
	pesos_i(1882) := b"0000000000000000_0000000000000000_0001101111011001_1001010111000100"; -- 0.10878883386142436
	pesos_i(1883) := b"1111111111111111_1111111111111111_1110011111010011_1101101101001010"; -- -0.09442357491772427
	pesos_i(1884) := b"1111111111111111_1111111111111111_1111111100000101_1110001011000101"; -- -0.003816439643316971
	pesos_i(1885) := b"0000000000000000_0000000000000000_0010001011110100_1110010000110100"; -- 0.13654924638601124
	pesos_i(1886) := b"1111111111111111_1111111111111111_1101111101100101_1100010000010000"; -- -0.1273534261135107
	pesos_i(1887) := b"0000000000000000_0000000000000000_0001010100011010_1011011101111011"; -- 0.08243891482340646
	pesos_i(1888) := b"1111111111111111_1111111111111111_1101011011001000_0101110100000101"; -- -0.1610051978553582
	pesos_i(1889) := b"1111111111111111_1111111111111111_1110100111010101_1010100101011000"; -- -0.0865835343440649
	pesos_i(1890) := b"1111111111111111_1111111111111111_1101111000101001_1011000010010010"; -- -0.132176365270151
	pesos_i(1891) := b"1111111111111111_1111111111111111_1111101010101101_0111110100011011"; -- -0.020790272567405614
	pesos_i(1892) := b"0000000000000000_0000000000000000_0010011000001000_0110100001000101"; -- 0.14856578528341527
	pesos_i(1893) := b"1111111111111111_1111111111111111_1110110101010110_0010001111100101"; -- -0.07290435454812372
	pesos_i(1894) := b"1111111111111111_1111111111111111_1110100000111010_0010100001101011"; -- -0.09286258107508383
	pesos_i(1895) := b"0000000000000000_0000000000000000_0000001101100100_1101111101010000"; -- 0.013257939263954271
	pesos_i(1896) := b"1111111111111111_1111111111111111_1101111110001000_1100100101110110"; -- -0.12681904667505864
	pesos_i(1897) := b"1111111111111111_1111111111111111_1111001010011100_0101010011100011"; -- -0.05230206919781484
	pesos_i(1898) := b"1111111111111111_1111111111111111_1111111000001110_1100010110100011"; -- -0.007587096854381203
	pesos_i(1899) := b"1111111111111111_1111111111111111_1110000001011101_0100111100100000"; -- -0.1235762163333854
	pesos_i(1900) := b"0000000000000000_0000000000000000_0001001110111100_1000010101010001"; -- 0.07709534857855437
	pesos_i(1901) := b"1111111111111111_1111111111111111_1101100000100011_1101100111101010"; -- -0.1557029536544849
	pesos_i(1902) := b"1111111111111111_1111111111111111_1111000010110010_1111110011011000"; -- -0.0597688648696477
	pesos_i(1903) := b"1111111111111111_1111111111111111_1111000101011011_0011010100101001"; -- -0.05720203163597732
	pesos_i(1904) := b"0000000000000000_0000000000000000_0000110010100111_0010100100011101"; -- 0.049425668216166035
	pesos_i(1905) := b"1111111111111111_1111111111111111_1110111111110110_1110110110111010"; -- -0.06263841830214763
	pesos_i(1906) := b"1111111111111111_1111111111111111_1110010110010011_1011010000011000"; -- -0.103214973474151
	pesos_i(1907) := b"1111111111111111_1111111111111111_1110001110010110_1010111110111011"; -- -0.11098195739486454
	pesos_i(1908) := b"0000000000000000_0000000000000000_0001110110100000_0111001101100010"; -- 0.11572953368790156
	pesos_i(1909) := b"0000000000000000_0000000000000000_0000010111000100_1010100110001111"; -- 0.0225320792091502
	pesos_i(1910) := b"0000000000000000_0000000000000000_0010011100111110_1011100010011011"; -- 0.153300798357582
	pesos_i(1911) := b"1111111111111111_1111111111111111_1110101010110010_1011001100100010"; -- -0.08321075840569216
	pesos_i(1912) := b"1111111111111111_1111111111111111_1110111000010101_1000011110010101"; -- -0.06998398420390302
	pesos_i(1913) := b"0000000000000000_0000000000000000_0001110011011111_1000110111000101"; -- 0.11278616002442139
	pesos_i(1914) := b"1111111111111111_1111111111111111_1101111110011001_1110011001001000"; -- -0.12655792940834526
	pesos_i(1915) := b"0000000000000000_0000000000000000_0010100010101101_0000000101101011"; -- 0.15888985513153478
	pesos_i(1916) := b"0000000000000000_0000000000000000_0001100100010101_0111110010111111"; -- 0.09798411995562245
	pesos_i(1917) := b"1111111111111111_1111111111111111_1101011100001111_0101010110100110"; -- -0.15992226316608812
	pesos_i(1918) := b"0000000000000000_0000000000000000_0010110110101001_0011101100001110"; -- 0.17836350518139776
	pesos_i(1919) := b"0000000000000000_0000000000000000_0010101111100010_0000110010011111"; -- 0.17141798867115005
	pesos_i(1920) := b"1111111111111111_1111111111111111_1101011100111011_1100010100000100"; -- -0.15924423849754002
	pesos_i(1921) := b"0000000000000000_0000000000000000_0000000011100100_1101011010001001"; -- 0.0034917911879460486
	pesos_i(1922) := b"1111111111111111_1111111111111111_1110100100100001_1111110011001011"; -- -0.08932514236223744
	pesos_i(1923) := b"1111111111111111_1111111111111111_1111000001001101_0011100001101101"; -- -0.06132171010835932
	pesos_i(1924) := b"1111111111111111_1111111111111111_1111010010011101_0011100111100000"; -- -0.04447592044619911
	pesos_i(1925) := b"1111111111111111_1111111111111111_1101110010110101_0110111000111010"; -- -0.13785658925419841
	pesos_i(1926) := b"0000000000000000_0000000000000000_0010000011011111_1010000010000001"; -- 0.12841227672613306
	pesos_i(1927) := b"1111111111111111_1111111111111111_1111000100110001_1101000001111101"; -- -0.05783364253763638
	pesos_i(1928) := b"1111111111111111_1111111111111111_1110011010011000_0001010110010111"; -- -0.09924187709950791
	pesos_i(1929) := b"1111111111111111_1111111111111111_1111111101011101_1101110001011001"; -- -0.0024740489855051033
	pesos_i(1930) := b"1111111111111111_1111111111111111_1110110110100010_0000010011111111"; -- -0.07174652830415885
	pesos_i(1931) := b"1111111111111111_1111111111111111_1110000000010101_0011111111100011"; -- -0.12467575752513758
	pesos_i(1932) := b"0000000000000000_0000000000000000_0001010000000110_1010000011011011"; -- 0.07822614041982702
	pesos_i(1933) := b"0000000000000000_0000000000000000_0001101001001110_1101010001000011"; -- 0.10276533724216531
	pesos_i(1934) := b"0000000000000000_0000000000000000_0001100000100110_1100010111001100"; -- 0.09434162371039712
	pesos_i(1935) := b"1111111111111111_1111111111111111_1110111110000100_0100110100011001"; -- -0.0643874943652874
	pesos_i(1936) := b"0000000000000000_0000000000000000_0001010001010111_0001110100010011"; -- 0.07945424761017847
	pesos_i(1937) := b"0000000000000000_0000000000000000_0010110000100110_1001010001011000"; -- 0.17246367594713977
	pesos_i(1938) := b"1111111111111111_1111111111111111_1111100000010000_0110001101111000"; -- -0.030999930488518748
	pesos_i(1939) := b"0000000000000000_0000000000000000_0001011100001110_0010110001000110"; -- 0.09006001186923947
	pesos_i(1940) := b"1111111111111111_1111111111111111_1101111111100110_0100111110011000"; -- -0.1253919843306623
	pesos_i(1941) := b"0000000000000000_0000000000000000_0000100101111011_1000011110100101"; -- 0.0370411660444991
	pesos_i(1942) := b"1111111111111111_1111111111111111_1111111000100111_0111011001100100"; -- -0.007210350585071143
	pesos_i(1943) := b"1111111111111111_1111111111111111_1111000110100010_1010110001111010"; -- -0.05611154583615654
	pesos_i(1944) := b"0000000000000000_0000000000000000_0010010110010101_1111110100011010"; -- 0.14681989558599917
	pesos_i(1945) := b"1111111111111111_1111111111111111_1110110110001101_0111101110100011"; -- -0.07205989149085493
	pesos_i(1946) := b"1111111111111111_1111111111111111_1101101000001010_0101100001000101"; -- -0.14827965092954828
	pesos_i(1947) := b"0000000000000000_0000000000000000_0010011000100000_1100101110110010"; -- 0.14893792245645354
	pesos_i(1948) := b"1111111111111111_1111111111111111_1111011110101111_0010110000101011"; -- -0.03248332919076236
	pesos_i(1949) := b"1111111111111111_1111111111111111_1110100110100110_1011110000011011"; -- -0.08729957911968644
	pesos_i(1950) := b"0000000000000000_0000000000000000_0000111011110000_1110101001011000"; -- 0.05836357733825527
	pesos_i(1951) := b"1111111111111111_1111111111111111_1110000101100111_1011101101000011"; -- -0.11951093298122888
	pesos_i(1952) := b"1111111111111111_1111111111111111_1101101001101100_1000001110111001"; -- -0.14678169953661735
	pesos_i(1953) := b"0000000000000000_0000000000000000_0010110111011100_0111111001001110"; -- 0.17914571191301917
	pesos_i(1954) := b"1111111111111111_1111111111111111_1111111010010010_1011101101101010"; -- -0.005573546127854735
	pesos_i(1955) := b"1111111111111111_1111111111111111_1111101110001100_1111111101000011"; -- -0.0173798046413774
	pesos_i(1956) := b"1111111111111111_1111111111111111_1110011001011000_1100101111001110"; -- -0.10020757878827509
	pesos_i(1957) := b"1111111111111111_1111111111111111_1110010000110101_0101010001110101"; -- -0.10856125016442485
	pesos_i(1958) := b"1111111111111111_1111111111111111_1111110100111110_0111111001111011"; -- -0.010765166162464772
	pesos_i(1959) := b"0000000000000000_0000000000000000_0000000100111100_0001100000001101"; -- 0.004823210803887229
	pesos_i(1960) := b"0000000000000000_0000000000000000_0000001100010110_1010000000000111"; -- 0.012063981708459265
	pesos_i(1961) := b"1111111111111111_1111111111111111_1101011011011110_1011001010001001"; -- -0.16066440725482303
	pesos_i(1962) := b"0000000000000000_0000000000000000_0000110001001001_1100110001001001"; -- 0.0480010680434443
	pesos_i(1963) := b"1111111111111111_1111111111111111_1110011001010110_0011000101010011"; -- -0.10024730413619386
	pesos_i(1964) := b"1111111111111111_1111111111111111_1110101011001001_1001000101111101"; -- -0.08286181169209741
	pesos_i(1965) := b"1111111111111111_1111111111111111_1101010001000010_0001111001110011"; -- -0.17086610509910985
	pesos_i(1966) := b"1111111111111111_1111111111111111_1101010010101010_1010101000111010"; -- -0.16927085957547633
	pesos_i(1967) := b"0000000000000000_0000000000000000_0001111100100000_1111111101101101"; -- 0.12159725580315017
	pesos_i(1968) := b"1111111111111111_1111111111111111_1110110001010110_1111100010011011"; -- -0.0767979261965812
	pesos_i(1969) := b"1111111111111111_1111111111111111_1110101001111001_1011100100101111"; -- -0.08408014873856957
	pesos_i(1970) := b"0000000000000000_0000000000000000_0000000100111111_0001000001101001"; -- 0.004868531930395089
	pesos_i(1971) := b"0000000000000000_0000000000000000_0000111001011101_1000010111110110"; -- 0.05611455213156265
	pesos_i(1972) := b"0000000000000000_0000000000000000_0000111001111100_1111010100001100"; -- 0.05659419582872207
	pesos_i(1973) := b"1111111111111111_1111111111111111_1101110100011011_0111000000010110"; -- -0.1363000817481632
	pesos_i(1974) := b"1111111111111111_1111111111111111_1110001001010011_0001100000011111"; -- -0.11591958268742476
	pesos_i(1975) := b"1111111111111111_1111111111111111_1110011010011000_0001011001011001"; -- -0.09924183213642498
	pesos_i(1976) := b"0000000000000000_0000000000000000_0010011011010100_0001011000010010"; -- 0.15167367882025032
	pesos_i(1977) := b"0000000000000000_0000000000000000_0000101001100000_1101101111001100"; -- 0.040540444627557466
	pesos_i(1978) := b"0000000000000000_0000000000000000_0001111111100001_0111110010100111"; -- 0.12453440733814485
	pesos_i(1979) := b"1111111111111111_1111111111111111_1111000111100110_0011111011101000"; -- -0.05508047892759786
	pesos_i(1980) := b"0000000000000000_0000000000000000_0001010011110011_0000001011101001"; -- 0.08183305915301424
	pesos_i(1981) := b"1111111111111111_1111111111111111_1111111010110111_0100101000110100"; -- -0.005015718829405172
	pesos_i(1982) := b"0000000000000000_0000000000000000_0010000000101111_0000001001101101"; -- 0.12571730774264214
	pesos_i(1983) := b"1111111111111111_1111111111111111_1111101011011110_0110001111001101"; -- -0.020044100219744083
	pesos_i(1984) := b"1111111111111111_1111111111111111_1101111110101010_1001100001110101"; -- -0.1263031687336466
	pesos_i(1985) := b"0000000000000000_0000000000000000_0001100110100100_1001101101010101"; -- 0.1001679499661726
	pesos_i(1986) := b"0000000000000000_0000000000000000_0000011001010100_1111010101110011"; -- 0.02473386823859587
	pesos_i(1987) := b"1111111111111111_1111111111111111_1111100100001011_0100010001000010"; -- -0.027171834925375858
	pesos_i(1988) := b"1111111111111111_1111111111111111_1111111100011000_1110100000001100"; -- -0.003526208084061375
	pesos_i(1989) := b"0000000000000000_0000000000000000_0000011110100111_1000010110101111"; -- 0.02989993583290889
	pesos_i(1990) := b"1111111111111111_1111111111111111_1111101110110111_1100110000100100"; -- -0.016726723893280133
	pesos_i(1991) := b"1111111111111111_1111111111111111_1111000110010001_0111000010111101"; -- -0.05637450587105356
	pesos_i(1992) := b"0000000000000000_0000000000000000_0001001100100000_1000100000000011"; -- 0.07471513811719194
	pesos_i(1993) := b"0000000000000000_0000000000000000_0010010001100100_1000101111011010"; -- 0.14215921476616722
	pesos_i(1994) := b"1111111111111111_1111111111111111_1110100010101011_1110110111000001"; -- -0.09112657584700477
	pesos_i(1995) := b"1111111111111111_1111111111111111_1110000101001010_0100000010011011"; -- -0.11996074885217814
	pesos_i(1996) := b"0000000000000000_0000000000000000_0010100110010001_0010111010000001"; -- 0.16237154621223432
	pesos_i(1997) := b"0000000000000000_0000000000000000_0000001111010011_1101010010011000"; -- 0.014951025957454284
	pesos_i(1998) := b"0000000000000000_0000000000000000_0010001111101000_0011001101110000"; -- 0.14026185488128748
	pesos_i(1999) := b"1111111111111111_1111111111111111_1101100010110010_1100000101010010"; -- -0.15352241275296039
	pesos_i(2000) := b"1111111111111111_1111111111111111_1111110110101001_0101101011100100"; -- -0.009134597251897025
	pesos_i(2001) := b"1111111111111111_1111111111111111_1110000101111010_0001010010100001"; -- -0.11923094819844259
	pesos_i(2002) := b"0000000000000000_0000000000000000_0010011001001101_0010111101010000"; -- 0.1496152467531761
	pesos_i(2003) := b"1111111111111111_1111111111111111_1110000001000100_1110001101001010"; -- -0.12394885477981424
	pesos_i(2004) := b"0000000000000000_0000000000000000_0001100111110000_1111011110000111"; -- 0.10133311318010392
	pesos_i(2005) := b"1111111111111111_1111111111111111_1111100011110001_1100011111000101"; -- -0.02756072462387605
	pesos_i(2006) := b"0000000000000000_0000000000000000_0001000001110101_1110011110011111"; -- 0.06429908390627018
	pesos_i(2007) := b"1111111111111111_1111111111111111_1110100010111100_0011111010011100"; -- -0.09087761594395913
	pesos_i(2008) := b"0000000000000000_0000000000000000_0001000001101110_0001101001011111"; -- 0.0641800386552224
	pesos_i(2009) := b"0000000000000000_0000000000000000_0000100011101000_1111010010111010"; -- 0.034804625943248374
	pesos_i(2010) := b"1111111111111111_1111111111111111_1111100101010101_0010100101001011"; -- -0.026044291560822986
	pesos_i(2011) := b"0000000000000000_0000000000000000_0000001001100101_0110101111011001"; -- 0.009360065862227002
	pesos_i(2012) := b"0000000000000000_0000000000000000_0001100001001111_1000011100011111"; -- 0.09496349824613241
	pesos_i(2013) := b"1111111111111111_1111111111111111_1111000101110101_1000000011111101"; -- -0.05680078335407003
	pesos_i(2014) := b"1111111111111111_1111111111111111_1110111111101101_1100000001011000"; -- -0.06277845239431554
	pesos_i(2015) := b"0000000000000000_0000000000000000_0000101010100001_0010000010100101"; -- 0.04152111077820875
	pesos_i(2016) := b"0000000000000000_0000000000000000_0001110111101101_1100111100001011"; -- 0.11690992362496924
	pesos_i(2017) := b"0000000000000000_0000000000000000_0010001101101100_1110010001100110"; -- 0.13838031294238662
	pesos_i(2018) := b"0000000000000000_0000000000000000_0000111010010101_1101100000101000"; -- 0.05697394351988721
	pesos_i(2019) := b"0000000000000000_0000000000000000_0001010011110110_0101000100110110"; -- 0.08188350259699985
	pesos_i(2020) := b"0000000000000000_0000000000000000_0010000100010001_1011110011000000"; -- 0.12917689971846774
	pesos_i(2021) := b"0000000000000000_0000000000000000_0001011010111111_1010001110000100"; -- 0.08886167508082464
	pesos_i(2022) := b"0000000000000000_0000000000000000_0000000110110100_0111011110010100"; -- 0.006659959554493342
	pesos_i(2023) := b"0000000000000000_0000000000000000_0010010100011100_0001111110101111"; -- 0.14496038462502667
	pesos_i(2024) := b"0000000000000000_0000000000000000_0001001011110000_0111100011101001"; -- 0.0739818162191008
	pesos_i(2025) := b"0000000000000000_0000000000000000_0001011010011001_0100110101000110"; -- 0.08827670060631372
	pesos_i(2026) := b"0000000000000000_0000000000000000_0010101100000010_0000000011000101"; -- 0.16799931348578823
	pesos_i(2027) := b"0000000000000000_0000000000000000_0000111011011110_0111011000010111"; -- 0.0580819898009194
	pesos_i(2028) := b"1111111111111111_1111111111111111_1111101110110101_1001010010011101"; -- -0.016760551042810094
	pesos_i(2029) := b"1111111111111111_1111111111111111_1110111000110100_1111010010011010"; -- -0.0695044636442258
	pesos_i(2030) := b"0000000000000000_0000000000000000_0010100110011111_1000101101111000"; -- 0.1625907105435185
	pesos_i(2031) := b"0000000000000000_0000000000000000_0001001000100000_1100011011001110"; -- 0.07081263100829467
	pesos_i(2032) := b"0000000000000000_0000000000000000_0010101000001110_0101000110011001"; -- 0.16428098673040611
	pesos_i(2033) := b"1111111111111111_1111111111111111_1110000110110011_1010100011000011"; -- -0.11835236787834673
	pesos_i(2034) := b"1111111111111111_1111111111111111_1111000011001011_1000011100000110"; -- -0.0593944178414288
	pesos_i(2035) := b"1111111111111111_1111111111111111_1110101100010101_1001010100010001"; -- -0.08170193040390286
	pesos_i(2036) := b"1111111111111111_1111111111111111_1101110111110111_1100000000010001"; -- -0.13293838106002992
	pesos_i(2037) := b"1111111111111111_1111111111111111_1110101000000100_1000100001011101"; -- -0.08586833687899427
	pesos_i(2038) := b"0000000000000000_0000000000000000_0010011000010100_0100010100011000"; -- 0.14874679418581316
	pesos_i(2039) := b"1111111111111111_1111111111111111_1110110011010010_1000111111010110"; -- -0.07491208094365474
	pesos_i(2040) := b"1111111111111111_1111111111111111_1111000011111001_1000110110010111"; -- -0.05869212221854035
	pesos_i(2041) := b"0000000000000000_0000000000000000_0010100000011101_0000110111001011"; -- 0.15669332694103574
	pesos_i(2042) := b"0000000000000000_0000000000000000_0000010111101001_1111011100001010"; -- 0.02310127248992077
	pesos_i(2043) := b"0000000000000000_0000000000000000_0001100101100100_0011001011110010"; -- 0.0991851654727871
	pesos_i(2044) := b"0000000000000000_0000000000000000_0001000000101110_0111010101011111"; -- 0.06320890027457063
	pesos_i(2045) := b"0000000000000000_0000000000000000_0000010011100111_1111010010011000"; -- 0.019164359117108835
	pesos_i(2046) := b"1111111111111111_1111111111111111_1101100001000001_0100111001110111"; -- -0.15525350179374287
	pesos_i(2047) := b"0000000000000000_0000000000000000_0010011010001001_0011001011111001"; -- 0.15053099236835452
	pesos_i(2048) := b"1111111111111111_1111111111111111_1111011111000001_1100101100110101"; -- -0.032199191543766575
	pesos_i(2049) := b"1111111111111111_1111111111111111_1111010011110101_1010100110111011"; -- -0.04312648003690634
	pesos_i(2050) := b"0000000000000000_0000000000000000_0010010101101000_1010110101101110"; -- 0.14612850124709748
	pesos_i(2051) := b"1111111111111111_1111111111111111_1110101101110010_0100010011110011"; -- -0.08028763838491094
	pesos_i(2052) := b"0000000000000000_0000000000000000_0001101100001101_0011010001000101"; -- 0.10567022969319177
	pesos_i(2053) := b"1111111111111111_1111111111111111_1110110110100101_1011000110001000"; -- -0.0716904682038297
	pesos_i(2054) := b"0000000000000000_0000000000000000_0001011100010011_0011100000001000"; -- 0.09013700681446653
	pesos_i(2055) := b"0000000000000000_0000000000000000_0010000100000010_1010000110101001"; -- 0.12894640337976015
	pesos_i(2056) := b"1111111111111111_1111111111111111_1110101010011101_0011111011100000"; -- -0.0835381223922424
	pesos_i(2057) := b"1111111111111111_1111111111111111_1101111011101011_1011000010000010"; -- -0.12921616377815698
	pesos_i(2058) := b"1111111111111111_1111111111111111_1110101000100100_0111000000100101"; -- -0.08538149918162177
	pesos_i(2059) := b"0000000000000000_0000000000000000_0000011010110100_0000001110110011"; -- 0.026184302478221465
	pesos_i(2060) := b"1111111111111111_1111111111111111_1110001110110111_1011101001111000"; -- -0.11047777722593911
	pesos_i(2061) := b"0000000000000000_0000000000000000_0001110001011100_1111010101100100"; -- 0.11079343496030715
	pesos_i(2062) := b"1111111111111111_1111111111111111_1111011100000100_0010000010101001"; -- -0.035093268077501495
	pesos_i(2063) := b"1111111111111111_1111111111111111_1110011010111000_0010011000011001"; -- -0.09875261205068521
	pesos_i(2064) := b"1111111111111111_1111111111111111_1111101101100011_0101111001000111"; -- -0.018015010449247054
	pesos_i(2065) := b"0000000000000000_0000000000000000_0001100011000101_1110111101010111"; -- 0.0967702472131273
	pesos_i(2066) := b"1111111111111111_1111111111111111_1101101101001010_1000110011011001"; -- -0.14339370440665503
	pesos_i(2067) := b"1111111111111111_1111111111111111_1110110110101010_1110111010110001"; -- -0.0716105287033571
	pesos_i(2068) := b"0000000000000000_0000000000000000_0000001010111001_0101010101111111"; -- 0.010640471979559552
	pesos_i(2069) := b"1111111111111111_1111111111111111_1101010101011011_1001001111110011"; -- -0.1665713818213221
	pesos_i(2070) := b"1111111111111111_1111111111111111_1111100011100001_0001000000101101"; -- -0.027815808372241933
	pesos_i(2071) := b"0000000000000000_0000000000000000_0001011100100110_0110110110100010"; -- 0.09043011856507088
	pesos_i(2072) := b"0000000000000000_0000000000000000_0010001110000010_0101101101111100"; -- 0.138707845384404
	pesos_i(2073) := b"1111111111111111_1111111111111111_1110011110110110_1100011001101011"; -- -0.09486732379132712
	pesos_i(2074) := b"0000000000000000_0000000000000000_0001010110110101_0110101110001000"; -- 0.08479950029230941
	pesos_i(2075) := b"1111111111111111_1111111111111111_1110011110101111_1000001111000101"; -- -0.09497810787719278
	pesos_i(2076) := b"1111111111111111_1111111111111111_1101001001000010_1011001111011001"; -- -0.17866970009236616
	pesos_i(2077) := b"1111111111111111_1111111111111111_1111001100100110_1011000010110011"; -- -0.05019088399134547
	pesos_i(2078) := b"1111111111111111_1111111111111111_1110100100010011_1001100001011011"; -- -0.08954475186393761
	pesos_i(2079) := b"0000000000000000_0000000000000000_0010001111010111_1010011111100101"; -- 0.14000939702803397
	pesos_i(2080) := b"1111111111111111_1111111111111111_1110001110000001_0001011110000110"; -- -0.11131146412955445
	pesos_i(2081) := b"1111111111111111_1111111111111111_1110001011010111_0111111101001110"; -- -0.11389927231165355
	pesos_i(2082) := b"1111111111111111_1111111111111111_1101110010100010_1111100110010001"; -- -0.13813820093424897
	pesos_i(2083) := b"1111111111111111_1111111111111111_1101110010010010_0110011010101000"; -- -0.1383910979197388
	pesos_i(2084) := b"0000000000000000_0000000000000000_0001110110000101_1101001110101100"; -- 0.11532328555292373
	pesos_i(2085) := b"0000000000000000_0000000000000000_0010001000000001_1111110000111001"; -- 0.1328427925045326
	pesos_i(2086) := b"1111111111111111_1111111111111111_1110001111010111_0111001000001010"; -- -0.10999381298470876
	pesos_i(2087) := b"1111111111111111_1111111111111111_1101010101100100_0100110100111011"; -- -0.16643826780937637
	pesos_i(2088) := b"0000000000000000_0000000000000000_0001000001001001_0001110100001011"; -- 0.06361562263180814
	pesos_i(2089) := b"1111111111111111_1111111111111111_1110101111111110_0001001111010000"; -- -0.07815433673579276
	pesos_i(2090) := b"0000000000000000_0000000000000000_0010011101010111_0101110011000101"; -- 0.15367679416157573
	pesos_i(2091) := b"1111111111111111_1111111111111111_1101011111100100_0000111000111010"; -- -0.15667639804300226
	pesos_i(2092) := b"1111111111111111_1111111111111111_1110000010001000_0000110010110110"; -- -0.12292404710501907
	pesos_i(2093) := b"1111111111111111_1111111111111111_1101010011111100_1110001110011100"; -- -0.16801621867697833
	pesos_i(2094) := b"1111111111111111_1111111111111111_1101011011101010_1110000101111111"; -- -0.16047850274856923
	pesos_i(2095) := b"0000000000000000_0000000000000000_0000111111001101_1000001010100000"; -- 0.061729587571395225
	pesos_i(2096) := b"1111111111111111_1111111111111111_1101100010100010_0111110101011111"; -- -0.15377060337118245
	pesos_i(2097) := b"0000000000000000_0000000000000000_0001000100110010_1010000111000000"; -- 0.06717883048614581
	pesos_i(2098) := b"1111111111111111_1111111111111111_1111100100101011_1000100010011010"; -- -0.02667947997343454
	pesos_i(2099) := b"0000000000000000_0000000000000000_0000100100011000_0000001100010110"; -- 0.03552264481022545
	pesos_i(2100) := b"1111111111111111_1111111111111111_1111010110111011_1011100111001010"; -- -0.04010428257212204
	pesos_i(2101) := b"0000000000000000_0000000000000000_0000000111000111_1001110110101111"; -- 0.0069521477111676045
	pesos_i(2102) := b"0000000000000000_0000000000000000_0001000011000000_1111010010111001"; -- 0.06544427412652018
	pesos_i(2103) := b"1111111111111111_1111111111111111_1110101100001010_1011101001100011"; -- -0.08186755259156121
	pesos_i(2104) := b"1111111111111111_1111111111111111_1110001101110011_0001011001011001"; -- -0.11152515721028346
	pesos_i(2105) := b"0000000000000000_0000000000000000_0001100110001101_0111100111110010"; -- 0.09981500769813575
	pesos_i(2106) := b"1111111111111111_1111111111111111_1111010010111011_1111111100110000"; -- -0.04400639597970645
	pesos_i(2107) := b"1111111111111111_1111111111111111_1110010110000011_0100110001101000"; -- -0.10346529445758143
	pesos_i(2108) := b"0000000000000000_0000000000000000_0000000110011100_1101011001101111"; -- 0.0062994022842088595
	pesos_i(2109) := b"0000000000000000_0000000000000000_0010010010001000_1111000111000000"; -- 0.1427146048150235
	pesos_i(2110) := b"1111111111111111_1111111111111111_1110011110110100_0101101011011100"; -- -0.09490425226207155
	pesos_i(2111) := b"1111111111111111_1111111111111111_1110011111011100_0111101111111010"; -- -0.0942919268883255
	pesos_i(2112) := b"0000000000000000_0000000000000000_0000111001011010_1001100010001111"; -- 0.05606988422849796
	pesos_i(2113) := b"1111111111111111_1111111111111111_1111111010001100_0000011001010111"; -- -0.0056758915369613215
	pesos_i(2114) := b"0000000000000000_0000000000000000_0000110001100010_0011000111100010"; -- 0.04837333446465047
	pesos_i(2115) := b"1111111111111111_1111111111111111_1110001110110111_0001001011011011"; -- -0.11048776771081183
	pesos_i(2116) := b"0000000000000000_0000000000000000_0000111010111000_1101111111010000"; -- 0.05750845741690934
	pesos_i(2117) := b"0000000000000000_0000000000000000_0001110110011011_1111010100011100"; -- 0.1156609720290887
	pesos_i(2118) := b"1111111111111111_1111111111111111_1101111100111100_1001001010100011"; -- -0.12798198231805802
	pesos_i(2119) := b"0000000000000000_0000000000000000_0001110001010100_1110111001111001"; -- 0.11067095243413409
	pesos_i(2120) := b"0000000000000000_0000000000000000_0000001110010010_1101010100111101"; -- 0.013959243125668767
	pesos_i(2121) := b"0000000000000000_0000000000000000_0000100111101100_0111011000000110"; -- 0.0387643589809331
	pesos_i(2122) := b"0000000000000000_0000000000000000_0000111010010111_1010011101101000"; -- 0.0570015554414578
	pesos_i(2123) := b"0000000000000000_0000000000000000_0000000101000010_0101100100010100"; -- 0.004918639471172719
	pesos_i(2124) := b"0000000000000000_0000000000000000_0001100110111111_1001100100111111"; -- 0.1005798128446777
	pesos_i(2125) := b"1111111111111111_1111111111111111_1101111000100110_1011110010001010"; -- -0.13222142825240793
	pesos_i(2126) := b"1111111111111111_1111111111111111_1110000011111110_1100110010111010"; -- -0.1211120649094268
	pesos_i(2127) := b"1111111111111111_1111111111111111_1101110100010011_0100001010001110"; -- -0.13642486612376323
	pesos_i(2128) := b"0000000000000000_0000000000000000_0000100101011000_0111111010100001"; -- 0.0365065711911392
	pesos_i(2129) := b"0000000000000000_0000000000000000_0010011111011110_0101111001110010"; -- 0.15573683058817603
	pesos_i(2130) := b"1111111111111111_1111111111111111_1110110111011010_0001111001100001"; -- -0.07089052325348688
	pesos_i(2131) := b"1111111111111111_1111111111111111_1110001010001110_0010000111000100"; -- -0.11501873946217124
	pesos_i(2132) := b"1111111111111111_1111111111111111_1111100111010100_0000110010111100"; -- -0.024108127798331675
	pesos_i(2133) := b"0000000000000000_0000000000000000_0001101100000100_1001011000100100"; -- 0.10553873429382853
	pesos_i(2134) := b"0000000000000000_0000000000000000_0001000110011101_0000010011000011"; -- 0.06880216362707738
	pesos_i(2135) := b"0000000000000000_0000000000000000_0001000111111100_1101110000011001"; -- 0.07026458370356838
	pesos_i(2136) := b"0000000000000000_0000000000000000_0001000001000010_1111010100101111"; -- 0.06352169416342782
	pesos_i(2137) := b"0000000000000000_0000000000000000_0000101001001101_0111000101001001"; -- 0.040244179016521664
	pesos_i(2138) := b"0000000000000000_0000000000000000_0000111111101001_1010011001010011"; -- 0.06215896161255617
	pesos_i(2139) := b"0000000000000000_0000000000000000_0010000000010111_0011011010101100"; -- 0.12535421074142009
	pesos_i(2140) := b"1111111111111111_1111111111111111_1111001011000100_0101000010011011"; -- -0.051691972980716344
	pesos_i(2141) := b"1111111111111111_1111111111111111_1101011010000101_0111011100011111"; -- -0.1620259809672244
	pesos_i(2142) := b"0000000000000000_0000000000000000_0001010000010010_0111001010011101"; -- 0.07840648970155581
	pesos_i(2143) := b"1111111111111111_1111111111111111_1101111100100001_0111000010001101"; -- -0.1283960013872941
	pesos_i(2144) := b"1111111111111111_1111111111111111_1111010100111101_0001101000010111"; -- -0.04203640881449974
	pesos_i(2145) := b"0000000000000000_0000000000000000_0000101011110100_0110100010110001"; -- 0.04279188463516184
	pesos_i(2146) := b"0000000000000000_0000000000000000_0000011010000110_1101100010101010"; -- 0.025495091970181606
	pesos_i(2147) := b"0000000000000000_0000000000000000_0000001100000110_0110101111000000"; -- 0.011816725140549014
	pesos_i(2148) := b"0000000000000000_0000000000000000_0000011111101010_1110000001101111"; -- 0.030927683820082714
	pesos_i(2149) := b"1111111111111111_1111111111111111_1110010101101010_0101011100011011"; -- -0.10384612653735124
	pesos_i(2150) := b"0000000000000000_0000000000000000_0010011010100010_0011100101111110"; -- 0.1509128507419302
	pesos_i(2151) := b"0000000000000000_0000000000000000_0001110010001100_0101110000100011"; -- 0.11151672219330463
	pesos_i(2152) := b"0000000000000000_0000000000000000_0001101001110011_0001100100111001"; -- 0.10331876413401184
	pesos_i(2153) := b"1111111111111111_1111111111111111_1101011010010101_0101100000011110"; -- -0.16178368813069288
	pesos_i(2154) := b"1111111111111111_1111111111111111_1110101001011001_1000010101000011"; -- -0.08457152484280947
	pesos_i(2155) := b"1111111111111111_1111111111111111_1101010010110001_0100010110100001"; -- -0.16917004422506784
	pesos_i(2156) := b"1111111111111111_1111111111111111_1111101110011101_1010110010001011"; -- -0.01712533575734937
	pesos_i(2157) := b"1111111111111111_1111111111111111_1111011110010010_1101101010111001"; -- -0.03291542982242496
	pesos_i(2158) := b"1111111111111111_1111111111111111_1111110000111101_0011100000101101"; -- -0.01469086563559354
	pesos_i(2159) := b"0000000000000000_0000000000000000_0010001101010111_1100000100100100"; -- 0.13805777670996286
	pesos_i(2160) := b"0000000000000000_0000000000000000_0000011000010001_0111111001001000"; -- 0.023704426347010088
	pesos_i(2161) := b"1111111111111111_1111111111111111_1111110010001001_0101010011111011"; -- -0.013529480589955067
	pesos_i(2162) := b"1111111111111111_1111111111111111_1101100001001100_1011011111010101"; -- -0.15507937471170755
	pesos_i(2163) := b"0000000000000000_0000000000000000_0000110111010000_1010011010100101"; -- 0.05396501096457277
	pesos_i(2164) := b"0000000000000000_0000000000000000_0001001001101101_0100000110010001"; -- 0.07197961609804783
	pesos_i(2165) := b"0000000000000000_0000000000000000_0000000110010111_1000000100001011"; -- 0.006218018742130979
	pesos_i(2166) := b"0000000000000000_0000000000000000_0000001100010000_0000110001110010"; -- 0.011963632405684337
	pesos_i(2167) := b"1111111111111111_1111111111111111_1111011101101011_0010110101100010"; -- -0.03352085445051778
	pesos_i(2168) := b"1111111111111111_1111111111111111_1110111000011011_1111010001110111"; -- -0.0698859413707213
	pesos_i(2169) := b"1111111111111111_1111111111111111_1110101011110000_1010101110000100"; -- -0.08226516752757596
	pesos_i(2170) := b"1111111111111111_1111111111111111_1101111110111111_0111110110100111"; -- -0.12598433180357113
	pesos_i(2171) := b"0000000000000000_0000000000000000_0001011111011111_0011111011010100"; -- 0.09325020480370579
	pesos_i(2172) := b"1111111111111111_1111111111111111_1111000000000101_0000010111011111"; -- -0.06242335608065897
	pesos_i(2173) := b"1111111111111111_1111111111111111_1111101110111011_1011010100010011"; -- -0.016667063570489953
	pesos_i(2174) := b"1111111111111111_1111111111111111_1101101111001000_1010001001011100"; -- -0.14146981480941254
	pesos_i(2175) := b"0000000000000000_0000000000000000_0000010001100000_0010100011110110"; -- 0.01709228513207814
	pesos_i(2176) := b"0000000000000000_0000000000000000_0000011100111000_1011101010111111"; -- 0.02820937314506325
	pesos_i(2177) := b"0000000000000000_0000000000000000_0000000110101000_1111101001010110"; -- 0.006484647702866262
	pesos_i(2178) := b"0000000000000000_0000000000000000_0001110001000100_1101000001111000"; -- 0.11042502337129928
	pesos_i(2179) := b"1111111111111111_1111111111111111_1101001101110000_1111010010111010"; -- -0.17405767868360134
	pesos_i(2180) := b"0000000000000000_0000000000000000_0010000111001001_0110110010110011"; -- 0.13197974554603636
	pesos_i(2181) := b"1111111111111111_1111111111111111_1111101000010001_1001101000111011"; -- -0.02316890764811847
	pesos_i(2182) := b"0000000000000000_0000000000000000_0001010010100101_0000010011001010"; -- 0.08064298567226723
	pesos_i(2183) := b"0000000000000000_0000000000000000_0000001011001100_0110111100110010"; -- 0.010931920795274355
	pesos_i(2184) := b"1111111111111111_1111111111111111_1111100101100110_0100111111010000"; -- -0.02578259643043994
	pesos_i(2185) := b"0000000000000000_0000000000000000_0001000110100110_1101011010000011"; -- 0.0689519949687386
	pesos_i(2186) := b"0000000000000000_0000000000000000_0000010011010001_0101001000101001"; -- 0.01881898399770544
	pesos_i(2187) := b"1111111111111111_1111111111111111_1110110000000110_1110011111001000"; -- -0.078019631955478
	pesos_i(2188) := b"0000000000000000_0000000000000000_0010011110101011_0110001101110001"; -- 0.15495893004416034
	pesos_i(2189) := b"1111111111111111_1111111111111111_1110011001011110_1010111001111110"; -- -0.10011777335300019
	pesos_i(2190) := b"1111111111111111_1111111111111111_1101001110000000_0101000100000010"; -- -0.17382329656568138
	pesos_i(2191) := b"1111111111111111_1111111111111111_1110101110111001_0101100100011010"; -- -0.07920306312779171
	pesos_i(2192) := b"1111111111111111_1111111111111111_1101110110101000_0110000010010111"; -- -0.13414951629216754
	pesos_i(2193) := b"0000000000000000_0000000000000000_0010011100000000_1111010111000110"; -- 0.1523583992865417
	pesos_i(2194) := b"0000000000000000_0000000000000000_0010000100010000_1010100001100110"; -- 0.12916042791711244
	pesos_i(2195) := b"1111111111111111_1111111111111111_1110110100101001_1000101100111010"; -- -0.07358484120890782
	pesos_i(2196) := b"1111111111111111_1111111111111111_1110001001001010_1000100100100111"; -- -0.1160501745803638
	pesos_i(2197) := b"1111111111111111_1111111111111111_1111000110010100_1001001010000001"; -- -0.05632671681924167
	pesos_i(2198) := b"1111111111111111_1111111111111111_1101010011010101_0110011010010110"; -- -0.1686187632834901
	pesos_i(2199) := b"1111111111111111_1111111111111111_1101010010000101_0110000100000100"; -- -0.16983979835741017
	pesos_i(2200) := b"1111111111111111_1111111111111111_1111110100110001_0010101100100001"; -- -0.0109684987655323
	pesos_i(2201) := b"1111111111111111_1111111111111111_1110011111011101_1000001011100000"; -- -0.09427625677107351
	pesos_i(2202) := b"0000000000000000_0000000000000000_0000001100110011_1101000011111001"; -- 0.012509403979743027
	pesos_i(2203) := b"0000000000000000_0000000000000000_0001111101100011_1001001101011101"; -- 0.12261315370891919
	pesos_i(2204) := b"1111111111111111_1111111111111111_1111110111110000_0111110100001010"; -- -0.008049187737851292
	pesos_i(2205) := b"1111111111111111_1111111111111111_1110010111110011_1011001101111100"; -- -0.10175016614887697
	pesos_i(2206) := b"1111111111111111_1111111111111111_1111110001000100_1100010011000011"; -- -0.014575674325553423
	pesos_i(2207) := b"1111111111111111_1111111111111111_1111100010010011_0011101111111011"; -- -0.029003382915478687
	pesos_i(2208) := b"0000000000000000_0000000000000000_0001111011001011_0000001011100001"; -- 0.1202852057179313
	pesos_i(2209) := b"1111111111111111_1111111111111111_1110001011111011_1001111011111101"; -- -0.11334806744285308
	pesos_i(2210) := b"0000000000000000_0000000000000000_0010001001110010_0000001111110011"; -- 0.1345522373311681
	pesos_i(2211) := b"1111111111111111_1111111111111111_1111001010100001_1100111101100110"; -- -0.05221847302536079
	pesos_i(2212) := b"1111111111111111_1111111111111111_1111101101011110_0011010000101111"; -- -0.01809381352376588
	pesos_i(2213) := b"1111111111111111_1111111111111111_1101011000100000_1100111001011101"; -- -0.16356191849824014
	pesos_i(2214) := b"0000000000000000_0000000000000000_0010001111000110_0010111100011000"; -- 0.1397427971998995
	pesos_i(2215) := b"1111111111111111_1111111111111111_1110101001111101_1110101010110011"; -- -0.08401616228015937
	pesos_i(2216) := b"0000000000000000_0000000000000000_0000111011100110_0111110011000101"; -- 0.05820445830543644
	pesos_i(2217) := b"0000000000000000_0000000000000000_0000110001111110_1101110001100010"; -- 0.048810743266735526
	pesos_i(2218) := b"0000000000000000_0000000000000000_0000010100011100_1101100000101011"; -- 0.01997138061304856
	pesos_i(2219) := b"1111111111111111_1111111111111111_1110010000100010_1010010101101100"; -- -0.1088463412269929
	pesos_i(2220) := b"0000000000000000_0000000000000000_0001000001010100_1001000010011011"; -- 0.06379035734122142
	pesos_i(2221) := b"1111111111111111_1111111111111111_1110000110000011_1101010010111010"; -- -0.11908216923756984
	pesos_i(2222) := b"1111111111111111_1111111111111111_1101011110001001_1101111000101000"; -- -0.1580525543585787
	pesos_i(2223) := b"0000000000000000_0000000000000000_0010111110101111_1001001100111010"; -- 0.18627281356348688
	pesos_i(2224) := b"1111111111111111_1111111111111111_1110010110011111_0011000111011011"; -- -0.10303963100798276
	pesos_i(2225) := b"0000000000000000_0000000000000000_0001110011111010_0100011111100010"; -- 0.11319398171789861
	pesos_i(2226) := b"0000000000000000_0000000000000000_0010000000100100_0010010001111000"; -- 0.12555149002605193
	pesos_i(2227) := b"0000000000000000_0000000000000000_0000000110100001_0011100001110100"; -- 0.006366280023613575
	pesos_i(2228) := b"0000000000000000_0000000000000000_0001000000101001_1011010011110010"; -- 0.06313639558657666
	pesos_i(2229) := b"1111111111111111_1111111111111111_1111100011100111_1111111010100000"; -- -0.027710042921422998
	pesos_i(2230) := b"1111111111111111_1111111111111111_1111110100000010_0111010001101001"; -- -0.011681293887531582
	pesos_i(2231) := b"1111111111111111_1111111111111111_1111110000101011_0111000011110010"; -- -0.014962139963829106
	pesos_i(2232) := b"0000000000000000_0000000000000000_0001010010000011_0001011011010100"; -- 0.08012526212672258
	pesos_i(2233) := b"0000000000000000_0000000000000000_0001101011101001_0010010010000110"; -- 0.10511997490179817
	pesos_i(2234) := b"0000000000000000_0000000000000000_0001001110010111_1101000100010000"; -- 0.07653528818549538
	pesos_i(2235) := b"1111111111111111_1111111111111111_1111001010010111_0100110001100110"; -- -0.052378869113676695
	pesos_i(2236) := b"1111111111111111_1111111111111111_1111111100100001_0001000001010111"; -- -0.003401736012040355
	pesos_i(2237) := b"0000000000000000_0000000000000000_0001100101100100_1111100101000110"; -- 0.09919698677526798
	pesos_i(2238) := b"1111111111111111_1111111111111111_1111101001110011_0000000000001000"; -- -0.021682737463760024
	pesos_i(2239) := b"1111111111111111_1111111111111111_1110111010010000_0101111001100001"; -- -0.06810960885662809
	pesos_i(2240) := b"0000000000000000_0000000000000000_0001011001111101_1010111000001110"; -- 0.08785522307441088
	pesos_i(2241) := b"1111111111111111_1111111111111111_1111001010010001_1001010100100111"; -- -0.05246608545277347
	pesos_i(2242) := b"0000000000000000_0000000000000000_0010001111001010_1010100110100001"; -- 0.13981113616906918
	pesos_i(2243) := b"1111111111111111_1111111111111111_1101010011101101_1100001111001110"; -- -0.16824699602801382
	pesos_i(2244) := b"1111111111111111_1111111111111111_1101101011000101_0001010101001101"; -- -0.14543024899699178
	pesos_i(2245) := b"0000000000000000_0000000000000000_0000111101001111_0010000100100011"; -- 0.05980116935698333
	pesos_i(2246) := b"1111111111111111_1111111111111111_1111010011000100_0100110001101110"; -- -0.04387972180749586
	pesos_i(2247) := b"1111111111111111_1111111111111111_1111000011010111_1101010000010100"; -- -0.05920671958013853
	pesos_i(2248) := b"1111111111111111_1111111111111111_1110111101010000_1010100010100101"; -- -0.06517549493834524
	pesos_i(2249) := b"1111111111111111_1111111111111111_1110110011101010_1100110111101110"; -- -0.0745421688915941
	pesos_i(2250) := b"0000000000000000_0000000000000000_0010001000100011_0011111111110001"; -- 0.1333503687222834
	pesos_i(2251) := b"0000000000000000_0000000000000000_0010011011101011_1010010100111111"; -- 0.152033164918037
	pesos_i(2252) := b"1111111111111111_1111111111111111_1111100111100010_1111110111001011"; -- -0.02388013645668677
	pesos_i(2253) := b"0000000000000000_0000000000000000_0010100010010001_1101010011100000"; -- 0.15847521268996723
	pesos_i(2254) := b"0000000000000000_0000000000000000_0010000000110011_0010000000100110"; -- 0.12578011441130243
	pesos_i(2255) := b"1111111111111111_1111111111111111_1111101011110000_1111110111101001"; -- -0.019760256296296817
	pesos_i(2256) := b"1111111111111111_1111111111111111_1101111010101000_0110100001001101"; -- -0.13024280651860987
	pesos_i(2257) := b"1111111111111111_1111111111111111_1111001010111110_0001100010001111"; -- -0.05178686632344646
	pesos_i(2258) := b"1111111111111111_1111111111111111_1111011111001110_1000001000011000"; -- -0.03200518517442286
	pesos_i(2259) := b"1111111111111111_1111111111111111_1111110000100100_0101010010111000"; -- -0.015070633887710908
	pesos_i(2260) := b"0000000000000000_0000000000000000_0000001100011100_1110111001100101"; -- 0.01216020557848851
	pesos_i(2261) := b"1111111111111111_1111111111111111_1110110111100010_0011100101000100"; -- -0.07076685030779997
	pesos_i(2262) := b"1111111111111111_1111111111111111_1101011011111010_1010110010111010"; -- -0.16023750741888926
	pesos_i(2263) := b"0000000000000000_0000000000000000_0001100001011010_1111001000101101"; -- 0.0951377258769185
	pesos_i(2264) := b"1111111111111111_1111111111111111_1100000100001010_0111001100111111"; -- -0.24593429285314666
	pesos_i(2265) := b"0000000000000000_0000000000000000_0010001000101101_1000010101010000"; -- 0.13350709158622853
	pesos_i(2266) := b"0000000000000000_0000000000000000_0010011110111111_0101111100110000"; -- 0.15526385223424993
	pesos_i(2267) := b"0000000000000000_0000000000000000_0000101111000111_1100011111101100"; -- 0.04601716534955983
	pesos_i(2268) := b"0000000000000000_0000000000000000_0001100011000010_0011010011010010"; -- 0.09671335345591289
	pesos_i(2269) := b"1111111111111111_1111111111111111_1110101000010010_1010010010010100"; -- -0.0856530320964168
	pesos_i(2270) := b"0000000000000000_0000000000000000_0000000101011000_1100011010010010"; -- 0.005260859168152561
	pesos_i(2271) := b"0000000000000000_0000000000000000_0000100001100010_0110011000111001"; -- 0.032751454307100164
	pesos_i(2272) := b"0000000000000000_0000000000000000_0000001000111011_0010101011011110"; -- 0.0087153236920266
	pesos_i(2273) := b"0000000000000000_0000000000000000_0000011110010011_1010011101001111"; -- 0.029596764444227843
	pesos_i(2274) := b"1111111111111111_1111111111111111_1110110011000010_0001001001110011"; -- -0.07516369534969555
	pesos_i(2275) := b"1111111111111111_1111111111111111_1101100010000001_1110100111011100"; -- -0.15426767700157645
	pesos_i(2276) := b"0000000000000000_0000000000000000_0000011101101111_0001100100010110"; -- 0.029038970839566455
	pesos_i(2277) := b"1111111111111111_1111111111111111_1110101111101001_1010000001100100"; -- -0.0784663922203484
	pesos_i(2278) := b"0000000000000000_0000000000000000_0000100000101100_1111001100010100"; -- 0.031935875281141994
	pesos_i(2279) := b"1111111111111111_1111111111111111_1111001100101101_1010011011101101"; -- -0.050084654895995645
	pesos_i(2280) := b"1111111111111111_1111111111111111_1101111000000001_0011111100100110"; -- -0.1327934772544681
	pesos_i(2281) := b"0000000000000000_0000000000000000_0010000011010011_1111001101011011"; -- 0.12823410961125578
	pesos_i(2282) := b"1111111111111111_1111111111111111_1110111110011010_0010011000010100"; -- -0.06405412679676101
	pesos_i(2283) := b"0000000000000000_0000000000000000_0001000000010110_1101100001100001"; -- 0.06284859054794016
	pesos_i(2284) := b"0000000000000000_0000000000000000_0001001011111101_0110000001111111"; -- 0.07417872535885046
	pesos_i(2285) := b"1111111111111111_1111111111111111_1101110000101110_0101101000010110"; -- -0.13991772616067685
	pesos_i(2286) := b"0000000000000000_0000000000000000_0000111010111010_0110100001011011"; -- 0.05753185490852829
	pesos_i(2287) := b"0000000000000000_0000000000000000_0001111101100001_0011011101100101"; -- 0.12257715427218506
	pesos_i(2288) := b"1111111111111111_1111111111111111_1101010110100111_0001010010001001"; -- -0.16541930828768395
	pesos_i(2289) := b"1111111111111111_1111111111111111_1110110001000100_0000110000100110"; -- -0.07708667827280563
	pesos_i(2290) := b"1111111111111111_1111111111111111_1110001101111100_0100011111111000"; -- -0.11138487058536921
	pesos_i(2291) := b"1111111111111111_1111111111111111_1110001010110100_1001100001111000"; -- -0.11443183008550438
	pesos_i(2292) := b"0000000000000000_0000000000000000_0010110110011001_0000110011111110"; -- 0.17811661902190423
	pesos_i(2293) := b"1111111111111111_1111111111111111_1110101110011010_1000111011100101"; -- -0.0796728792610314
	pesos_i(2294) := b"0000000000000000_0000000000000000_0010100100010001_0010000010000011"; -- 0.16041758734995673
	pesos_i(2295) := b"1111111111111111_1111111111111111_1101010110011111_0001011100001010"; -- -0.16554122939185284
	pesos_i(2296) := b"1111111111111111_1111111111111111_1101110110001110_1000000000000111"; -- -0.1345443710238088
	pesos_i(2297) := b"0000000000000000_0000000000000000_0000101100101111_0010011001010110"; -- 0.04368819799716053
	pesos_i(2298) := b"1111111111111111_1111111111111111_1110101110001010_1000100111111001"; -- -0.0799173131928565
	pesos_i(2299) := b"1111111111111111_1111111111111111_1110000111101000_0110101010111011"; -- -0.11754734942120064
	pesos_i(2300) := b"0000000000000000_0000000000000000_0001101001111001_1101011110100101"; -- 0.10342166690829449
	pesos_i(2301) := b"0000000000000000_0000000000000000_0010110011111001_1101110100100110"; -- 0.17568761997799928
	pesos_i(2302) := b"1111111111111111_1111111111111111_1101011111010100_0011100111010000"; -- -0.15691794089934435
	pesos_i(2303) := b"1111111111111111_1111111111111111_1110001011111100_1011000110010110"; -- -0.11333170031517042
	pesos_i(2304) := b"0000000000000000_0000000000000000_0000111110001000_0110110110101100"; -- 0.06067548216133087
	pesos_i(2305) := b"1111111111111111_1111111111111111_1111001101010111_1100101101100011"; -- -0.04944161254167028
	pesos_i(2306) := b"1111111111111111_1111111111111111_1110110101110100_1111010101111111"; -- -0.07243409783997551
	pesos_i(2307) := b"0000000000000000_0000000000000000_0010010001100110_1000011111000011"; -- 0.14218948840227957
	pesos_i(2308) := b"0000000000000000_0000000000000000_0000101000110110_1111000110110111"; -- 0.03990088183862427
	pesos_i(2309) := b"1111111111111111_1111111111111111_1111010000011111_1101011100000100"; -- -0.04638916158992602
	pesos_i(2310) := b"1111111111111111_1111111111111111_1101111011000100_1010110100101011"; -- -0.12981145568141883
	pesos_i(2311) := b"1111111111111111_1111111111111111_1110001000100100_1011111100010001"; -- -0.11662679518196943
	pesos_i(2312) := b"0000000000000000_0000000000000000_0001001101100110_0111100101010000"; -- 0.07578237718680537
	pesos_i(2313) := b"1111111111111111_1111111111111111_1111000111000101_0011011000110010"; -- -0.055584538254260005
	pesos_i(2314) := b"0000000000000000_0000000000000000_0010100010101101_0010011110111000"; -- 0.15889213795769733
	pesos_i(2315) := b"0000000000000000_0000000000000000_0010000011110110_1111100000111011"; -- 0.12876845786741364
	pesos_i(2316) := b"0000000000000000_0000000000000000_0001010110111101_0001001110100001"; -- 0.08491633113595908
	pesos_i(2317) := b"1111111111111111_1111111111111111_1110101110100010_1001011111011101"; -- -0.07955027439980049
	pesos_i(2318) := b"0000000000000000_0000000000000000_0000000010010001_0000111000010010"; -- 0.0022133630626505643
	pesos_i(2319) := b"0000000000000000_0000000000000000_0001100001001110_0100011000001001"; -- 0.09494435993208301
	pesos_i(2320) := b"0000000000000000_0000000000000000_0010110010001101_0100100011011110"; -- 0.17403083244253584
	pesos_i(2321) := b"0000000000000000_0000000000000000_0000011001100000_0100010100110101"; -- 0.024906468864451827
	pesos_i(2322) := b"0000000000000000_0000000000000000_0010010110101110_1001010111001111"; -- 0.1471952086045183
	pesos_i(2323) := b"1111111111111111_1111111111111111_1110001000000011_1101110011001100"; -- -0.11712856301259841
	pesos_i(2324) := b"1111111111111111_1111111111111111_1110100101001010_0011011101100010"; -- -0.08871129864062936
	pesos_i(2325) := b"0000000000000000_0000000000000000_0001100111110100_1010000110001001"; -- 0.10138902284555143
	pesos_i(2326) := b"1111111111111111_1111111111111111_1110010000100000_0100011011001010"; -- -0.10888249939273852
	pesos_i(2327) := b"1111111111111111_1111111111111111_1110001100110010_1000010010000111"; -- -0.11251041126031111
	pesos_i(2328) := b"0000000000000000_0000000000000000_0000001100111110_0101011110000001"; -- 0.012670010496416773
	pesos_i(2329) := b"1111111111111111_1111111111111111_1111000000110001_1111010001010000"; -- -0.06173775718058938
	pesos_i(2330) := b"1111111111111111_1111111111111111_1110001111111011_0011111011001101"; -- -0.1094475506144894
	pesos_i(2331) := b"0000000000000000_0000000000000000_0010010010101000_0110100101101100"; -- 0.14319476024975616
	pesos_i(2332) := b"1111111111111111_1111111111111111_1101011000110011_0010110000111100"; -- -0.16328166506750252
	pesos_i(2333) := b"0000000000000000_0000000000000000_0001111000010001_0000010110001100"; -- 0.1174472300216126
	pesos_i(2334) := b"1111111111111111_1111111111111111_1101001000011100_1101011011011010"; -- -0.17924744766108663
	pesos_i(2335) := b"0000000000000000_0000000000000000_0000100000100101_0001011000111100"; -- 0.03181590044682778
	pesos_i(2336) := b"1111111111111111_1111111111111111_1101110010110011_0101110100010110"; -- -0.13788812836268857
	pesos_i(2337) := b"0000000000000000_0000000000000000_0000100010010111_1000010111101110"; -- 0.03356205989163547
	pesos_i(2338) := b"1111111111111111_1111111111111111_1110011010110010_0100100111011100"; -- -0.09884203307439698
	pesos_i(2339) := b"1111111111111111_1111111111111111_1110101101010100_0110111011100010"; -- -0.08074290252381165
	pesos_i(2340) := b"1111111111111111_1111111111111111_1110001101010110_1010010110101001"; -- -0.11195911999763451
	pesos_i(2341) := b"0000000000000000_0000000000000000_0010011010100010_0101100010111110"; -- 0.15091471317231825
	pesos_i(2342) := b"1111111111111111_1111111111111111_1111011101110000_0011010010001100"; -- -0.03344413348859503
	pesos_i(2343) := b"0000000000000000_0000000000000000_0000010011100001_1111000001001100"; -- 0.01907255037561048
	pesos_i(2344) := b"1111111111111111_1111111111111111_1101110110110010_1101010100101110"; -- -0.13398997908305565
	pesos_i(2345) := b"1111111111111111_1111111111111111_1110100010100100_1100111101011110"; -- -0.09123519855319334
	pesos_i(2346) := b"0000000000000000_0000000000000000_0010110000001011_0111011001111110"; -- 0.172049909329411
	pesos_i(2347) := b"0000000000000000_0000000000000000_0010110011001000_1100100101111001"; -- 0.17493876661519908
	pesos_i(2348) := b"0000000000000000_0000000000000000_0001110000001000_0010101100110111"; -- 0.1094996461797361
	pesos_i(2349) := b"0000000000000000_0000000000000000_0000000011001010_1111011101101110"; -- 0.0030970233186701735
	pesos_i(2350) := b"0000000000000000_0000000000000000_0000010110001100_0100101110100101"; -- 0.02167198917072547
	pesos_i(2351) := b"1111111111111111_1111111111111111_1101001110100011_0100010000011111"; -- -0.1732900070944065
	pesos_i(2352) := b"1111111111111111_1111111111111111_1110010000001011_0111001010110001"; -- -0.10920031720188457
	pesos_i(2353) := b"0000000000000000_0000000000000000_0000001000010011_0000011011001101"; -- 0.008102822237533452
	pesos_i(2354) := b"0000000000000000_0000000000000000_0000001001000110_1011001101111110"; -- 0.008891313848095944
	pesos_i(2355) := b"1111111111111111_1111111111111111_1110010000101000_0000111011010011"; -- -0.10876376480698634
	pesos_i(2356) := b"0000000000000000_0000000000000000_0001100110011010_1010010010111100"; -- 0.10001592256536437
	pesos_i(2357) := b"0000000000000000_0000000000000000_0001010011111101_0010101011100110"; -- 0.08198803053135646
	pesos_i(2358) := b"0000000000000000_0000000000000000_0000010001101110_1111001101011111"; -- 0.017317972765662437
	pesos_i(2359) := b"1111111111111111_1111111111111111_1100101010110100_0110110100001011"; -- -0.2081844185244986
	pesos_i(2360) := b"0000000000000000_0000000000000000_0001101110011010_0010001010111011"; -- 0.1078206735099552
	pesos_i(2361) := b"1111111111111111_1111111111111111_1110101001100001_0010001001110001"; -- -0.08445534451980931
	pesos_i(2362) := b"1111111111111111_1111111111111111_1101111010001100_0000110010000111"; -- -0.13067552291347018
	pesos_i(2363) := b"0000000000000000_0000000000000000_0000101111000000_1001100011011011"; -- 0.045907548333818174
	pesos_i(2364) := b"0000000000000000_0000000000000000_0001001011110101_0110000001001001"; -- 0.07405664227671901
	pesos_i(2365) := b"0000000000000000_0000000000000000_0000111100000101_1111111100001010"; -- 0.05868524552706235
	pesos_i(2366) := b"1111111111111111_1111111111111111_1101111100000101_0100010100100100"; -- -0.1288258349216705
	pesos_i(2367) := b"0000000000000000_0000000000000000_0000000110110101_0100101101001011"; -- 0.0066725787267818085
	pesos_i(2368) := b"0000000000000000_0000000000000000_0001001100110001_0011011010011010"; -- 0.07496968519498645
	pesos_i(2369) := b"0000000000000000_0000000000000000_0001101001001000_0001000000110111"; -- 0.10266209929980524
	pesos_i(2370) := b"0000000000000000_0000000000000000_0000100001001110_1110101001111101"; -- 0.03245416204783854
	pesos_i(2371) := b"1111111111111111_1111111111111111_1111111100111111_1000100010101010"; -- -0.0029368003928921626
	pesos_i(2372) := b"0000000000000000_0000000000000000_0000001110011100_0010111011001100"; -- 0.014101910480961533
	pesos_i(2373) := b"1111111111111111_1111111111111111_1110111010111110_0101100111111111"; -- -0.06740796583750246
	pesos_i(2374) := b"1111111111111111_1111111111111111_1110011110001000_1011110010100000"; -- -0.09556981187040284
	pesos_i(2375) := b"1111111111111111_1111111111111111_1111000101011100_0001010010011101"; -- -0.05718871264675025
	pesos_i(2376) := b"0000000000000000_0000000000000000_0000010010000010_0010111011101000"; -- 0.017611438369142012
	pesos_i(2377) := b"1111111111111111_1111111111111111_1111111000000111_1001010010111100"; -- -0.007696823162230615
	pesos_i(2378) := b"0000000000000000_0000000000000000_0000010100111000_1111111111100010"; -- 0.02040099405457495
	pesos_i(2379) := b"1111111111111111_1111111111111111_1110101000000001_1100100000111001"; -- -0.08591030709772303
	pesos_i(2380) := b"0000000000000000_0000000000000000_0001000001001110_0100101001011111"; -- 0.06369461837266317
	pesos_i(2381) := b"1111111111111111_1111111111111111_1101001011111010_0000011100001000"; -- -0.17587238361356333
	pesos_i(2382) := b"1111111111111111_1111111111111111_1110000111111011_0110110101001000"; -- -0.11725728030913962
	pesos_i(2383) := b"0000000000000000_0000000000000000_0010001101100001_0111010001001011"; -- 0.13820578420574003
	pesos_i(2384) := b"1111111111111111_1111111111111111_1110001110100001_1011001100011101"; -- -0.1108139090916235
	pesos_i(2385) := b"1111111111111111_1111111111111111_1111101001011111_0101110001100010"; -- -0.02198240865473843
	pesos_i(2386) := b"0000000000000000_0000000000000000_0001001101110001_1000000001000100"; -- 0.07595063833148133
	pesos_i(2387) := b"0000000000000000_0000000000000000_0000001011001000_0101010100101010"; -- 0.01086933388122179
	pesos_i(2388) := b"1111111111111111_1111111111111111_1110010101001111_0010001011111001"; -- -0.10426122118054094
	pesos_i(2389) := b"0000000000000000_0000000000000000_0001110111001001_1010111101010110"; -- 0.1163587174760789
	pesos_i(2390) := b"1111111111111111_1111111111111111_1110001011011010_0010101011001010"; -- -0.1138585336513723
	pesos_i(2391) := b"1111111111111111_1111111111111111_1110111010100000_1111111000010110"; -- -0.0678559491573891
	pesos_i(2392) := b"0000000000000000_0000000000000000_0001101000000100_1011011101111011"; -- 0.10163447147557815
	pesos_i(2393) := b"1111111111111111_1111111111111111_1101101000011000_0010101001100011"; -- -0.14806876261564506
	pesos_i(2394) := b"0000000000000000_0000000000000000_0010000011101111_1101110000101111"; -- 0.1286599746390536
	pesos_i(2395) := b"1111111111111111_1111111111111111_1111111000011010_1001010001010101"; -- -0.007406930099222592
	pesos_i(2396) := b"1111111111111111_1111111111111111_1101011101101001_1000011110111011"; -- -0.15854598697481906
	pesos_i(2397) := b"0000000000000000_0000000000000000_0010010111110011_0000101000011100"; -- 0.14823973836718773
	pesos_i(2398) := b"0000000000000000_0000000000000000_0000010010111100_1011001101011011"; -- 0.01850434277651038
	pesos_i(2399) := b"0000000000000000_0000000000000000_0000011001000110_0010010110011001"; -- 0.024507856297112163
	pesos_i(2400) := b"1111111111111111_1111111111111111_1111111110111001_1110001101011011"; -- -0.0010698225789212423
	pesos_i(2401) := b"1111111111111111_1111111111111111_1111110100110101_1111011101101010"; -- -0.010895287143803894
	pesos_i(2402) := b"0000000000000000_0000000000000000_0010100101001100_0101001101100001"; -- 0.16132088785167994
	pesos_i(2403) := b"0000000000000000_0000000000000000_0000100101100001_1110100111111111"; -- 0.03665029971378182
	pesos_i(2404) := b"1111111111111111_1111111111111111_1111111101010100_0111010100011110"; -- -0.0026175309236684385
	pesos_i(2405) := b"1111111111111111_1111111111111111_1110000000000100_1001100000000001"; -- -0.12492990465108891
	pesos_i(2406) := b"1111111111111111_1111111111111111_1111010110111101_0001001001100110"; -- -0.04008374227138509
	pesos_i(2407) := b"0000000000000000_0000000000000000_0000111100001000_0001111110000000"; -- 0.05871769796454701
	pesos_i(2408) := b"1111111111111111_1111111111111111_1111101010001111_0011000111101001"; -- -0.021252518296431794
	pesos_i(2409) := b"1111111111111111_1111111111111111_1110101001000000_1101010011010101"; -- -0.08494825176091567
	pesos_i(2410) := b"1111111111111111_1111111111111111_1101111011011011_0100001101000101"; -- -0.12946681559991438
	pesos_i(2411) := b"1111111111111111_1111111111111111_1111111000010110_1100110101011100"; -- -0.007464566171070058
	pesos_i(2412) := b"0000000000000000_0000000000000000_0000000100010001_1100011011100101"; -- 0.004177504466209688
	pesos_i(2413) := b"0000000000000000_0000000000000000_0000000111000110_1101001110000100"; -- 0.006940097562968186
	pesos_i(2414) := b"0000000000000000_0000000000000000_0010010010000001_0101110100100010"; -- 0.14259893483031585
	pesos_i(2415) := b"1111111111111111_1111111111111111_1111001011001111_1011010001001011"; -- -0.051518184442096555
	pesos_i(2416) := b"0000000000000000_0000000000000000_0000010110110010_1010101010100111"; -- 0.022257486109841712
	pesos_i(2417) := b"0000000000000000_0000000000000000_0010100001110010_1011101101010011"; -- 0.15800066726362572
	pesos_i(2418) := b"0000000000000000_0000000000000000_0000100100111001_0011100010101110"; -- 0.03602937945407792
	pesos_i(2419) := b"1111111111111111_1111111111111111_1111101110000000_0011000000010101"; -- -0.01757525916209993
	pesos_i(2420) := b"1111111111111111_1111111111111111_1110110100110000_0101010111010010"; -- -0.07348121288743843
	pesos_i(2421) := b"0000000000000000_0000000000000000_0010110101001010_1001110010101100"; -- 0.17691973879960374
	pesos_i(2422) := b"1111111111111111_1111111111111111_1110111011011010_0100111110010010"; -- -0.06698134113672025
	pesos_i(2423) := b"0000000000000000_0000000000000000_0010011100101100_0111100001001000"; -- 0.15302230596631605
	pesos_i(2424) := b"0000000000000000_0000000000000000_0001000101011110_0100000001101011"; -- 0.0678444158379051
	pesos_i(2425) := b"1111111111111111_1111111111111111_1111100111101100_1000111100101101"; -- -0.023734141892587348
	pesos_i(2426) := b"1111111111111111_1111111111111111_1110110000000011_1011010010001101"; -- -0.07806846199967463
	pesos_i(2427) := b"0000000000000000_0000000000000000_0000000011100011_1000100110000011"; -- 0.0034719413760932872
	pesos_i(2428) := b"1111111111111111_1111111111111111_1110100111001100_1111100101000000"; -- -0.08671610051257742
	pesos_i(2429) := b"0000000000000000_0000000000000000_0000010110111000_1110101110100100"; -- 0.02235291247445567
	pesos_i(2430) := b"1111111111111111_1111111111111111_1111101101000011_0110101110010111"; -- -0.01850249830392092
	pesos_i(2431) := b"1111111111111111_1111111111111111_1101100111010110_0011100100001110"; -- -0.14907496851662222
	pesos_i(2432) := b"0000000000000000_0000000000000000_0010100000000001_1001001011010000"; -- 0.15627400945669348
	pesos_i(2433) := b"0000000000000000_0000000000000000_0000110011101011_0001000110001100"; -- 0.050461861332326025
	pesos_i(2434) := b"0000000000000000_0000000000000000_0010000011100000_0100100101011011"; -- 0.12842234104203504
	pesos_i(2435) := b"1111111111111111_1111111111111111_1111110000111011_0100101000111100"; -- -0.01472030673373539
	pesos_i(2436) := b"0000000000000000_0000000000000000_0000011000111000_0100101011001000"; -- 0.024296449410352028
	pesos_i(2437) := b"1111111111111111_1111111111111111_1111100101100100_1001011011011101"; -- -0.025808879048641088
	pesos_i(2438) := b"1111111111111111_1111111111111111_1110001001000010_1010111110001111"; -- -0.11616995575742987
	pesos_i(2439) := b"0000000000000000_0000000000000000_0001101001000000_1100100100011010"; -- 0.10255104919416799
	pesos_i(2440) := b"0000000000000000_0000000000000000_0001010101000101_0111100111110110"; -- 0.08309137587807806
	pesos_i(2441) := b"1111111111111111_1111111111111111_1110000000111111_1010001111001000"; -- -0.12402893418111686
	pesos_i(2442) := b"1111111111111111_1111111111111111_1110011111110110_0000011110011001"; -- -0.09390213509589074
	pesos_i(2443) := b"0000000000000000_0000000000000000_0001100001010001_1011101111100101"; -- 0.09499716128234569
	pesos_i(2444) := b"1111111111111111_1111111111111111_1111000100010100_1010001011010001"; -- -0.058278869684652755
	pesos_i(2445) := b"0000000000000000_0000000000000000_0001101101001110_1000010000010110"; -- 0.1066668084906415
	pesos_i(2446) := b"0000000000000000_0000000000000000_0000111100110000_1110011100000010"; -- 0.05933994112131204
	pesos_i(2447) := b"0000000000000000_0000000000000000_0010001111011100_1100001111110010"; -- 0.14008736294389365
	pesos_i(2448) := b"0000000000000000_0000000000000000_0010001110101010_1010010101100111"; -- 0.13932260287530548
	pesos_i(2449) := b"0000000000000000_0000000000000000_0010101011001000_0110110011100101"; -- 0.1671207484398395
	pesos_i(2450) := b"1111111111111111_1111111111111111_1111101110111001_0111011111010001"; -- -0.0167012323304781
	pesos_i(2451) := b"1111111111111111_1111111111111111_1111101110010001_0110000011101101"; -- -0.017312948288739038
	pesos_i(2452) := b"1111111111111111_1111111111111111_1111001011000111_1010111100100101"; -- -0.05164056163058105
	pesos_i(2453) := b"0000000000000000_0000000000000000_0001000101101011_0101101110100110"; -- 0.06804440306319087
	pesos_i(2454) := b"0000000000000000_0000000000000000_0001011110001000_0010100001101010"; -- 0.09192135415908896
	pesos_i(2455) := b"0000000000000000_0000000000000000_0000100111100101_0000010101101011"; -- 0.0386508357202365
	pesos_i(2456) := b"0000000000000000_0000000000000000_0000111101100100_0110011011001110"; -- 0.06012575665879193
	pesos_i(2457) := b"0000000000000000_0000000000000000_0001010011101110_1100111010000111"; -- 0.08176890170473132
	pesos_i(2458) := b"0000000000000000_0000000000000000_0001010100110101_0011111101011111"; -- 0.08284374292187557
	pesos_i(2459) := b"0000000000000000_0000000000000000_0001010000111001_1111011100010111"; -- 0.07900947869933798
	pesos_i(2460) := b"1111111111111111_1111111111111111_1101010011011000_1110110001111100"; -- -0.16856500589224221
	pesos_i(2461) := b"0000000000000000_0000000000000000_0000001101111010_0011011011111010"; -- 0.013583599149065382
	pesos_i(2462) := b"1111111111111111_1111111111111111_1111101001101101_1100100110100111"; -- -0.02176227263809161
	pesos_i(2463) := b"1111111111111111_1111111111111111_1101010011010001_0011101001000110"; -- -0.16868243964392957
	pesos_i(2464) := b"0000000000000000_0000000000000000_0001110000110010_0110100010100010"; -- 0.11014417613324054
	pesos_i(2465) := b"1111111111111111_1111111111111111_1110101111111101_0110111011011110"; -- -0.07816416817160789
	pesos_i(2466) := b"0000000000000000_0000000000000000_0001110110011101_1110001111010101"; -- 0.11569045962946883
	pesos_i(2467) := b"1111111111111111_1111111111111111_1101110011000101_0000101100010010"; -- -0.137618358765779
	pesos_i(2468) := b"0000000000000000_0000000000000000_0000100110011101_0001011001100101"; -- 0.03755321472944009
	pesos_i(2469) := b"0000000000000000_0000000000000000_0001101111111100_1101101100001101"; -- 0.10932702122654295
	pesos_i(2470) := b"1111111111111111_1111111111111111_1111111101000111_1010001011110011"; -- -0.0028131634363117914
	pesos_i(2471) := b"1111111111111111_1111111111111111_1111100100100101_1100110001001111"; -- -0.026766997171456003
	pesos_i(2472) := b"1111111111111111_1111111111111111_1111011001110010_0010001100000110"; -- -0.03732091049499642
	pesos_i(2473) := b"0000000000000000_0000000000000000_0010010000101100_1110000110101001"; -- 0.14130983702366448
	pesos_i(2474) := b"1111111111111111_1111111111111111_1110101001010100_1110011111001001"; -- -0.08464194613379748
	pesos_i(2475) := b"1111111111111111_1111111111111111_1110100000111001_0100111001111111"; -- -0.09287557032665107
	pesos_i(2476) := b"0000000000000000_0000000000000000_0000100010101010_0011110000011111"; -- 0.03384757753474129
	pesos_i(2477) := b"0000000000000000_0000000000000000_0000111111001101_1011000011111111"; -- 0.06173235162762071
	pesos_i(2478) := b"1111111111111111_1111111111111111_1110010110001010_0111101001011101"; -- -0.10335574378519116
	pesos_i(2479) := b"0000000000000000_0000000000000000_0010000001111100_1011111101110000"; -- 0.12690350029740555
	pesos_i(2480) := b"0000000000000000_0000000000000000_0001111001111011_0010100101011101"; -- 0.11906679655513483
	pesos_i(2481) := b"0000000000000000_0000000000000000_0010011001100101_0100101001101001"; -- 0.1499830730010825
	pesos_i(2482) := b"1111111111111111_1111111111111111_1110111110101110_0111000001001001"; -- -0.06374452789041996
	pesos_i(2483) := b"0000000000000000_0000000000000000_0010100101010110_1011100011111010"; -- 0.16147953138355725
	pesos_i(2484) := b"0000000000000000_0000000000000000_0001011100101101_0101111001010110"; -- 0.09053601828442433
	pesos_i(2485) := b"0000000000000000_0000000000000000_0001011100101110_0000001100010100"; -- 0.09054583786779045
	pesos_i(2486) := b"0000000000000000_0000000000000000_0000011110110110_1001100010010111"; -- 0.030129944728371758
	pesos_i(2487) := b"0000000000000000_0000000000000000_0000010111001010_1010001010011000"; -- 0.022623216746480188
	pesos_i(2488) := b"0000000000000000_0000000000000000_0001001001110001_1101001010001000"; -- 0.07204929189401252
	pesos_i(2489) := b"0000000000000000_0000000000000000_0000010101101010_1000010110001101"; -- 0.021156641863028448
	pesos_i(2490) := b"0000000000000000_0000000000000000_0010010010110011_0010110000111100"; -- 0.14335895979669208
	pesos_i(2491) := b"1111111111111111_1111111111111111_1101110001101111_0010011111010010"; -- -0.13892890095228258
	pesos_i(2492) := b"1111111111111111_1111111111111111_1111001110110001_0010000110110110"; -- -0.04807843510135212
	pesos_i(2493) := b"1111111111111111_1111111111111111_1101001000110101_1101000010001100"; -- -0.17886635380521798
	pesos_i(2494) := b"0000000000000000_0000000000000000_0000010010010110_0000011101100111"; -- 0.01791425955249251
	pesos_i(2495) := b"0000000000000000_0000000000000000_0010001110000011_0110000111101001"; -- 0.13872348730373152
	pesos_i(2496) := b"1111111111111111_1111111111111111_1111010010001010_1011000110111010"; -- -0.04475869380361652
	pesos_i(2497) := b"0000000000000000_0000000000000000_0010010100011110_1011101100101101"; -- 0.14500017016393976
	pesos_i(2498) := b"1111111111111111_1111111111111111_1101101011111011_0100011010011000"; -- -0.14460333620268132
	pesos_i(2499) := b"0000000000000000_0000000000000000_0000100101000011_0110011011010000"; -- 0.03618471691425336
	pesos_i(2500) := b"1111111111111111_1111111111111111_1101110100000100_1110111010110101"; -- -0.13664348678909308
	pesos_i(2501) := b"1111111111111111_1111111111111111_1110001011010110_1111100001000111"; -- -0.11390732068168304
	pesos_i(2502) := b"1111111111111111_1111111111111111_1111110100010101_1110000010100001"; -- -0.011384926453230268
	pesos_i(2503) := b"1111111111111111_1111111111111111_1110011101110010_1101000111000001"; -- -0.09590424568749507
	pesos_i(2504) := b"1111111111111111_1111111111111111_1110101110001110_0111011101101101"; -- -0.07985738357260662
	pesos_i(2505) := b"0000000000000000_0000000000000000_0001101010010110_0010111000110111"; -- 0.10385407293985471
	pesos_i(2506) := b"1111111111111111_1111111111111111_1110000001101011_0000100010101001"; -- -0.1233667933076979
	pesos_i(2507) := b"1111111111111111_1111111111111111_1111010100111110_0011101010111111"; -- -0.04201920354622978
	pesos_i(2508) := b"1111111111111111_1111111111111111_1101101101001111_1010101111011011"; -- -0.14331556233731568
	pesos_i(2509) := b"1111111111111111_1111111111111111_1101111101100110_1011001001111111"; -- -0.12733921442293397
	pesos_i(2510) := b"1111111111111111_1111111111111111_1101100001010000_0101110110001010"; -- -0.15502372151254917
	pesos_i(2511) := b"0000000000000000_0000000000000000_0000000001001110_1000000101111111"; -- 0.001197904137951533
	pesos_i(2512) := b"1111111111111111_1111111111111111_1110110110001010_1111101001110111"; -- -0.07209810816659042
	pesos_i(2513) := b"1111111111111111_1111111111111111_1111010110110110_1011101110001000"; -- -0.04018047256675855
	pesos_i(2514) := b"1111111111111111_1111111111111111_1111011101011000_1000001110010101"; -- -0.03380563374816839
	pesos_i(2515) := b"1111111111111111_1111111111111111_1111000010001110_0111000111001001"; -- -0.060326469824871505
	pesos_i(2516) := b"0000000000000000_0000000000000000_0000110110110011_1000001011010010"; -- 0.05352037078576799
	pesos_i(2517) := b"1111111111111111_1111111111111111_1111000001000101_1010111110101000"; -- -0.061436673537694324
	pesos_i(2518) := b"0000000000000000_0000000000000000_0010011011010111_0000011011101111"; -- 0.15171855287966307
	pesos_i(2519) := b"1111111111111111_1111111111111111_1110001011110010_0011101111100111"; -- -0.11349130269043278
	pesos_i(2520) := b"0000000000000000_0000000000000000_0000010010101001_0000000111011000"; -- 0.01820384519778867
	pesos_i(2521) := b"0000000000000000_0000000000000000_0000101000111101_1101010011111011"; -- 0.04000598064598276
	pesos_i(2522) := b"0000000000000000_0000000000000000_0010001001000011_1000100011010000"; -- 0.13384299343446013
	pesos_i(2523) := b"0000000000000000_0000000000000000_0010111110010011_1111110000010110"; -- 0.18585181744144408
	pesos_i(2524) := b"0000000000000000_0000000000000000_0000001010011011_1110110001000111"; -- 0.010191695599196115
	pesos_i(2525) := b"0000000000000000_0000000000000000_0000001101010001_1101100101010110"; -- 0.012967666116758168
	pesos_i(2526) := b"0000000000000000_0000000000000000_0000000101100001_1011000010000110"; -- 0.005396874107690628
	pesos_i(2527) := b"0000000000000000_0000000000000000_0000010001000100_0100001100111011"; -- 0.016666605020399128
	pesos_i(2528) := b"0000000000000000_0000000000000000_0000100001100011_1001011101010010"; -- 0.03276963943272718
	pesos_i(2529) := b"1111111111111111_1111111111111111_1101011001000010_1001001101011110"; -- -0.1630466362079914
	pesos_i(2530) := b"1111111111111111_1111111111111111_1110111111100101_1011100000111001"; -- -0.06290100675977776
	pesos_i(2531) := b"1111111111111111_1111111111111111_1111100101101100_1011011110110111"; -- -0.025684850416534795
	pesos_i(2532) := b"0000000000000000_0000000000000000_0000011000010000_1110000010111100"; -- 0.023695035869283038
	pesos_i(2533) := b"1111111111111111_1111111111111111_1111100001011001_1011010111111110"; -- -0.029881120216827733
	pesos_i(2534) := b"0000000000000000_0000000000000000_0000000101111101_1111111111000011"; -- 0.005828843193687843
	pesos_i(2535) := b"1111111111111111_1111111111111111_1110011101000101_1011110110011001"; -- -0.09659209275404981
	pesos_i(2536) := b"0000000000000000_0000000000000000_0000001010010110_1010011011000000"; -- 0.010111257435013288
	pesos_i(2537) := b"0000000000000000_0000000000000000_0000110010100010_0000111101110011"; -- 0.049347844756081144
	pesos_i(2538) := b"0000000000000000_0000000000000000_0010011011101111_1100001010000111"; -- 0.15209594526176737
	pesos_i(2539) := b"0000000000000000_0000000000000000_0000101101001001_1110001010100101"; -- 0.04409615058374345
	pesos_i(2540) := b"0000000000000000_0000000000000000_0010110111001111_0110011111110110"; -- 0.17894601584607414
	pesos_i(2541) := b"1111111111111111_1111111111111111_1111111000111111_0001000011001000"; -- -0.006850196111737164
	pesos_i(2542) := b"0000000000000000_0000000000000000_0000100110010101_1111011100010000"; -- 0.03744453573386541
	pesos_i(2543) := b"1111111111111111_1111111111111111_1101110000011011_0110100001100111"; -- -0.140206789742107
	pesos_i(2544) := b"0000000000000000_0000000000000000_0010001000000100_1011111100101000"; -- 0.13288492902016005
	pesos_i(2545) := b"0000000000000000_0000000000000000_0000100101101101_1101110111110101"; -- 0.03683268768669667
	pesos_i(2546) := b"1111111111111111_1111111111111111_1101000011001010_0110110111001001"; -- -0.18441118081000865
	pesos_i(2547) := b"1111111111111111_1111111111111111_1110100001100101_0000101010101001"; -- -0.0922082269917498
	pesos_i(2548) := b"0000000000000000_0000000000000000_0000000101011110_0101101001111010"; -- 0.005345968949491051
	pesos_i(2549) := b"0000000000000000_0000000000000000_0000110100010011_1110000000011100"; -- 0.05108452498847293
	pesos_i(2550) := b"0000000000000000_0000000000000000_0000110001110101_1011000100110010"; -- 0.0486708400071104
	pesos_i(2551) := b"0000000000000000_0000000000000000_0010000010110001_0101001010001100"; -- 0.12770572593443538
	pesos_i(2552) := b"0000000000000000_0000000000000000_0010001100000100_1100100001011010"; -- 0.13679172704222622
	pesos_i(2553) := b"1111111111111111_1111111111111111_1111110011100101_0100001111011010"; -- -0.01212669306276624
	pesos_i(2554) := b"1111111111111111_1111111111111111_1101111001111011_1001110011010011"; -- -0.13092632155236836
	pesos_i(2555) := b"1111111111111111_1111111111111111_1111010101110100_1010110111000010"; -- -0.04118837370885071
	pesos_i(2556) := b"1111111111111111_1111111111111111_1101111010100110_1001001000110111"; -- -0.13027082592477346
	pesos_i(2557) := b"0000000000000000_0000000000000000_0010010100100000_0111110001110010"; -- 0.14502694872289748
	pesos_i(2558) := b"0000000000000000_0000000000000000_0000001111000010_1000110111001110"; -- 0.014687407382342806
	pesos_i(2559) := b"1111111111111111_1111111111111111_1110010011110001_1000000010101010"; -- -0.10568996279253705
	pesos_i(2560) := b"0000000000000000_0000000000000000_0000001001101000_0111110010100001"; -- 0.00940684245716164
	pesos_i(2561) := b"0000000000000000_0000000000000000_0010100111000001_0101011000011111"; -- 0.1631063295697748
	pesos_i(2562) := b"1111111111111111_1111111111111111_1111111010111001_0000001000100001"; -- -0.004989497111599878
	pesos_i(2563) := b"0000000000000000_0000000000000000_0010101011101100_1101101100011100"; -- 0.1676766342419172
	pesos_i(2564) := b"0000000000000000_0000000000000000_0010011100011001_0100010000100100"; -- 0.15272928113080758
	pesos_i(2565) := b"0000000000000000_0000000000000000_0000001010101111_1010110001011011"; -- 0.0104930611864309
	pesos_i(2566) := b"1111111111111111_1111111111111111_1101001111110100_1100000011110111"; -- -0.17204660396154814
	pesos_i(2567) := b"1111111111111111_1111111111111111_1111000100010100_0110111101100001"; -- -0.05828193546688405
	pesos_i(2568) := b"1111111111111111_1111111111111111_1110100011100000_1011100101110010"; -- -0.09032097777303204
	pesos_i(2569) := b"0000000000000000_0000000000000000_0000000011010111_1100101001100001"; -- 0.003292702327900055
	pesos_i(2570) := b"0000000000000000_0000000000000000_0010100110111000_1111110101110100"; -- 0.16297897413105933
	pesos_i(2571) := b"1111111111111111_1111111111111111_1110110010011111_0111010000110110"; -- -0.0756919259227572
	pesos_i(2572) := b"0000000000000000_0000000000000000_0010101111010000_0000010100000101"; -- 0.1711428773774871
	pesos_i(2573) := b"1111111111111111_1111111111111111_1101010110011000_0001101100010110"; -- -0.16564779962749435
	pesos_i(2574) := b"0000000000000000_0000000000000000_0000001111101100_1101000001100011"; -- 0.015332244967250837
	pesos_i(2575) := b"0000000000000000_0000000000000000_0000111100110011_0100000101110100"; -- 0.059375849605837486
	pesos_i(2576) := b"1111111111111111_1111111111111111_1110011100000010_0010101101001100"; -- -0.09762315177030448
	pesos_i(2577) := b"1111111111111111_1111111111111111_1111101110011011_0000001010111111"; -- -0.01716597405464089
	pesos_i(2578) := b"1111111111111111_1111111111111111_1110000100000110_0111100000111001"; -- -0.12099503153321438
	pesos_i(2579) := b"0000000000000000_0000000000000000_0001000000001111_1100101110110111"; -- 0.06274102427967572
	pesos_i(2580) := b"0000000000000000_0000000000000000_0000111101100100_0001100010000101"; -- 0.060121090285878885
	pesos_i(2581) := b"1111111111111111_1111111111111111_1110100010110010_1101101110110001"; -- -0.09102084093748755
	pesos_i(2582) := b"0000000000000000_0000000000000000_0010000000000011_1001100001000111"; -- 0.12505485271071642
	pesos_i(2583) := b"1111111111111111_1111111111111111_1111000111001010_0100110000101001"; -- -0.05550693509390005
	pesos_i(2584) := b"1111111111111111_1111111111111111_1111100101001001_1010000011110010"; -- -0.026220265269762913
	pesos_i(2585) := b"1111111111111111_1111111111111111_1111001101000111_0011110100001010"; -- -0.04969423765204799
	pesos_i(2586) := b"1111111111111111_1111111111111111_1101010011101001_0101111101000001"; -- -0.16831402458340675
	pesos_i(2587) := b"1111111111111111_1111111111111111_1110001011101001_0100001111101110"; -- -0.11362815327903585
	pesos_i(2588) := b"0000000000000000_0000000000000000_0010010000010001_1011111011010001"; -- 0.14089577296020453
	pesos_i(2589) := b"1111111111111111_1111111111111111_1111111011110001_1100111111101101"; -- -0.00412273847152059
	pesos_i(2590) := b"1111111111111111_1111111111111111_1110111110000001_1011001111111000"; -- -0.06442713928374928
	pesos_i(2591) := b"1111111111111111_1111111111111111_1110000001001010_1010011000011110"; -- -0.12386094833291167
	pesos_i(2592) := b"0000000000000000_0000000000000000_0010001000111001_0010010100011011"; -- 0.13368446257658453
	pesos_i(2593) := b"1111111111111111_1111111111111111_1111101010101010_0110000101100010"; -- -0.020837701305303925
	pesos_i(2594) := b"1111111111111111_1111111111111111_1111001000000101_1111000010110010"; -- -0.05459685938990033
	pesos_i(2595) := b"1111111111111111_1111111111111111_1101011110011110_1010000100100010"; -- -0.15773575711976945
	pesos_i(2596) := b"1111111111111111_1111111111111111_1111011010010111_1110101111001110"; -- -0.03674436783837462
	pesos_i(2597) := b"1111111111111111_1111111111111111_1111101001101001_1001110000000101"; -- -0.021826027595610604
	pesos_i(2598) := b"1111111111111111_1111111111111111_1111111110010111_1010010110000110"; -- -0.0015923068855067616
	pesos_i(2599) := b"0000000000000000_0000000000000000_0010001001000011_1000111111100110"; -- 0.1338434159306305
	pesos_i(2600) := b"0000000000000000_0000000000000000_0001000011100101_1011000110000111"; -- 0.06600484404087073
	pesos_i(2601) := b"0000000000000000_0000000000000000_0000100111010111_0000001001000000"; -- 0.038437023735854114
	pesos_i(2602) := b"1111111111111111_1111111111111111_1111111011110010_1010101101000011"; -- -0.004109665077542594
	pesos_i(2603) := b"0000000000000000_0000000000000000_0001111010110100_1111101100000011"; -- 0.11994904354228489
	pesos_i(2604) := b"1111111111111111_1111111111111111_1110011010010110_1111001011111101"; -- -0.09925919835993996
	pesos_i(2605) := b"1111111111111111_1111111111111111_1110001000001010_0110000011001110"; -- -0.1170291419854784
	pesos_i(2606) := b"0000000000000000_0000000000000000_0000110000100111_0011100100011000"; -- 0.04747349577091848
	pesos_i(2607) := b"1111111111111111_1111111111111111_1100101000001100_0010011101000010"; -- -0.21075205454477547
	pesos_i(2608) := b"1111111111111111_1111111111111111_1111111000001000_0100101101100110"; -- -0.007685935564091445
	pesos_i(2609) := b"1111111111111111_1111111111111111_1111010010111000_1001100100110111"; -- -0.04405825046238452
	pesos_i(2610) := b"1111111111111111_1111111111111111_1111000111101001_1001101011000100"; -- -0.055029227403319315
	pesos_i(2611) := b"1111111111111111_1111111111111111_1101101011000111_0111101111010101"; -- -0.14539361996733602
	pesos_i(2612) := b"0000000000000000_0000000000000000_0001010110110110_0011011101000100"; -- 0.0848116438034632
	pesos_i(2613) := b"1111111111111111_1111111111111111_1101010010111011_0100010101010000"; -- -0.16901747520655108
	pesos_i(2614) := b"0000000000000000_0000000000000000_0001110000001011_1111010011111010"; -- 0.10955744835315719
	pesos_i(2615) := b"1111111111111111_1111111111111111_1101101010101100_0001101011100111"; -- -0.1458113848602272
	pesos_i(2616) := b"1111111111111111_1111111111111111_1110111000110101_1101010100110001"; -- -0.06949107695128169
	pesos_i(2617) := b"0000000000000000_0000000000000000_0001101011000010_0010001100101011"; -- 0.10452480118922626
	pesos_i(2618) := b"0000000000000000_0000000000000000_0000111001101111_0010001111001010"; -- 0.05638335877421591
	pesos_i(2619) := b"0000000000000000_0000000000000000_0010001100111011_0111011010010001"; -- 0.1376260857542559
	pesos_i(2620) := b"1111111111111111_1111111111111111_1110110100110010_1000010001100111"; -- -0.07344791868659044
	pesos_i(2621) := b"0000000000000000_0000000000000000_0000101111011010_0011100001110110"; -- 0.04629853138578569
	pesos_i(2622) := b"0000000000000000_0000000000000000_0000101101001010_1001010101001011"; -- 0.04410679884120725
	pesos_i(2623) := b"0000000000000000_0000000000000000_0000011100101101_0101000110001101"; -- 0.02803525622428033
	pesos_i(2624) := b"0000000000000000_0000000000000000_0010000100110101_0000110000000101"; -- 0.12971568216902332
	pesos_i(2625) := b"1111111111111111_1111111111111111_1111100001001001_0101000110011010"; -- -0.030131244679252378
	pesos_i(2626) := b"0000000000000000_0000000000000000_0010000001010000_1000111100101100"; -- 0.1262292369425829
	pesos_i(2627) := b"1111111111111111_1111111111111111_1110001010111101_1101000000100111"; -- -0.1142911820150595
	pesos_i(2628) := b"1111111111111111_1111111111111111_1110100000001011_0000001111110110"; -- -0.0935819172439266
	pesos_i(2629) := b"1111111111111111_1111111111111111_1101100000011111_0001000011011110"; -- -0.15577597226932824
	pesos_i(2630) := b"1111111111111111_1111111111111111_1111111111101001_0100111010000001"; -- -0.0003462729955173817
	pesos_i(2631) := b"1111111111111111_1111111111111111_1101101111000010_1001111101110110"; -- -0.14156154035948024
	pesos_i(2632) := b"1111111111111111_1111111111111111_1101111010100111_1100000110000110"; -- -0.13025274729606584
	pesos_i(2633) := b"1111111111111111_1111111111111111_1110010101010101_1110001011000101"; -- -0.1041582364490439
	pesos_i(2634) := b"1111111111111111_1111111111111111_1110010011101101_1101011010101001"; -- -0.10574587229265373
	pesos_i(2635) := b"0000000000000000_0000000000000000_0000110100101110_1101110000011110"; -- 0.05149627424305581
	pesos_i(2636) := b"1111111111111111_1111111111111111_1111011011000101_1101000011001111"; -- -0.03604407268374549
	pesos_i(2637) := b"1111111111111111_1111111111111111_1110100001100001_0101111010110000"; -- -0.09226425360668018
	pesos_i(2638) := b"1111111111111111_1111111111111111_1110000010001111_1100010110101010"; -- -0.12280621144881569
	pesos_i(2639) := b"1111111111111111_1111111111111111_1110101010000001_0110000101110110"; -- -0.08396330710384227
	pesos_i(2640) := b"0000000000000000_0000000000000000_0000010100010011_1100011100111100"; -- 0.019833042270133827
	pesos_i(2641) := b"1111111111111111_1111111111111111_1111111110000111_1000011011001001"; -- -0.0018382795934965943
	pesos_i(2642) := b"0000000000000000_0000000000000000_0001000110000001_1101000111011100"; -- 0.06838714249837329
	pesos_i(2643) := b"1111111111111111_1111111111111111_1110000110110111_1001101100011010"; -- -0.1182921467120504
	pesos_i(2644) := b"0000000000000000_0000000000000000_0001101010101010_1110001101110100"; -- 0.10417005150526092
	pesos_i(2645) := b"1111111111111111_1111111111111111_1111110111101100_1111000011010110"; -- -0.008103320829158876
	pesos_i(2646) := b"0000000000000000_0000000000000000_0010001001111100_0111001001011001"; -- 0.13471140547617746
	pesos_i(2647) := b"1111111111111111_1111111111111111_1110001101100110_1100011110010010"; -- -0.11171295810212972
	pesos_i(2648) := b"1111111111111111_1111111111111111_1111001011100000_0100100100001010"; -- -0.051265177860870655
	pesos_i(2649) := b"1111111111111111_1111111111111111_1101001100110000_0100110011010111"; -- -0.17504424805245652
	pesos_i(2650) := b"1111111111111111_1111111111111111_1110001100100111_1010000001110011"; -- -0.11267659374439497
	pesos_i(2651) := b"1111111111111111_1111111111111111_1101101001111011_1100100000111001"; -- -0.14654873469467344
	pesos_i(2652) := b"1111111111111111_1111111111111111_1101100100011100_1111101100001011"; -- -0.15190154066369907
	pesos_i(2653) := b"1111111111111111_1111111111111111_1101101011000100_0001011100011100"; -- -0.14544539994955935
	pesos_i(2654) := b"1111111111111111_1111111111111111_1111001111111110_1011110010101100"; -- -0.04689427187240377
	pesos_i(2655) := b"0000000000000000_0000000000000000_0000011101011111_1011100101101100"; -- 0.028804386976651802
	pesos_i(2656) := b"0000000000000000_0000000000000000_0010110011000111_1101001111010010"; -- 0.17492412451718334
	pesos_i(2657) := b"0000000000000000_0000000000000000_0010000111110001_0010110010101001"; -- 0.1325862801623112
	pesos_i(2658) := b"1111111111111111_1111111111111111_1110101110101110_0000110110111010"; -- -0.07937540259683755
	pesos_i(2659) := b"1111111111111111_1111111111111111_1111111111011010_0010101000011101"; -- -0.0005773238441105484
	pesos_i(2660) := b"1111111111111111_1111111111111111_1101011100001111_0000010111000111"; -- -0.1599270239178277
	pesos_i(2661) := b"1111111111111111_1111111111111111_1111110010100110_0101010110101001"; -- -0.013086935192990168
	pesos_i(2662) := b"0000000000000000_0000000000000000_0000000110001110_0001000101001001"; -- 0.006074028209514578
	pesos_i(2663) := b"1111111111111111_1111111111111111_1111000100001000_1110110001111011"; -- -0.0584575844488192
	pesos_i(2664) := b"0000000000000000_0000000000000000_0000010011000101_0001001100100001"; -- 0.018632121713277966
	pesos_i(2665) := b"0000000000000000_0000000000000000_0000011000101000_1000110101000011"; -- 0.02405627133009034
	pesos_i(2666) := b"1111111111111111_1111111111111111_1101110110010000_0100001111000111"; -- -0.13451744458461118
	pesos_i(2667) := b"0000000000000000_0000000000000000_0010001011111110_1110110111101011"; -- 0.13670241345170256
	pesos_i(2668) := b"0000000000000000_0000000000000000_0000100010011111_1111011001110011"; -- 0.033690837056373955
	pesos_i(2669) := b"1111111111111111_1111111111111111_1101101001011111_1010110101000111"; -- -0.14697758699896424
	pesos_i(2670) := b"0000000000000000_0000000000000000_0000001111100011_0001011111110110"; -- 0.015183923216969696
	pesos_i(2671) := b"0000000000000000_0000000000000000_0000111010000001_1000010011010100"; -- 0.05666380105590227
	pesos_i(2672) := b"1111111111111111_1111111111111111_1110001101110111_0111001100100110"; -- -0.11145859073148409
	pesos_i(2673) := b"0000000000000000_0000000000000000_0000101010101100_1001001011000111"; -- 0.041695760366990214
	pesos_i(2674) := b"0000000000000000_0000000000000000_0001001100100111_1011111011110111"; -- 0.07482522519858391
	pesos_i(2675) := b"1111111111111111_1111111111111111_1111010100010011_1101101010101111"; -- -0.04266579833393983
	pesos_i(2676) := b"1111111111111111_1111111111111111_1111000111100011_0011100101101111"; -- -0.05512658148190285
	pesos_i(2677) := b"0000000000000000_0000000000000000_0001000101010101_1111000011001011"; -- 0.06771759938176661
	pesos_i(2678) := b"1111111111111111_1111111111111111_1110010001010001_0001000111010110"; -- -0.10813797509496365
	pesos_i(2679) := b"1111111111111111_1111111111111111_1111111001011110_0101110111101001"; -- -0.00637257624088276
	pesos_i(2680) := b"1111111111111111_1111111111111111_1111110011101100_1101100001100010"; -- -0.012011028305624366
	pesos_i(2681) := b"1111111111111111_1111111111111111_1111100000110100_0001101010011010"; -- -0.030454957465879978
	pesos_i(2682) := b"1111111111111111_1111111111111111_1111011110110101_1100110110100011"; -- -0.03238215230075182
	pesos_i(2683) := b"0000000000000000_0000000000000000_0001110101101001_0100000000111110"; -- 0.11488725195483566
	pesos_i(2684) := b"1111111111111111_1111111111111111_1111010001110111_0101100001010100"; -- -0.0450539393522789
	pesos_i(2685) := b"1111111111111111_1111111111111111_1110110011110111_1110011110111110"; -- -0.0743422661170587
	pesos_i(2686) := b"0000000000000000_0000000000000000_0010011100111100_1101100011011001"; -- 0.1532722024515137
	pesos_i(2687) := b"0000000000000000_0000000000000000_0000101000100001_1111111000010001"; -- 0.03958118355846939
	pesos_i(2688) := b"0000000000000000_0000000000000000_0000001100110011_1111110011110100"; -- 0.012512025511838859
	pesos_i(2689) := b"1111111111111111_1111111111111111_1110011000101011_1001110001011110"; -- -0.10089705191115525
	pesos_i(2690) := b"1111111111111111_1111111111111111_1101110100000000_0100010001101000"; -- -0.13671467273382762
	pesos_i(2691) := b"1111111111111111_1111111111111111_1101101010000010_1111000101011010"; -- -0.14643947185591438
	pesos_i(2692) := b"0000000000000000_0000000000000000_0000011110111100_1111100001111011"; -- 0.030227212867277586
	pesos_i(2693) := b"0000000000000000_0000000000000000_0000100100110110_1000000001010100"; -- 0.035987873553904925
	pesos_i(2694) := b"0000000000000000_0000000000000000_0001101010000101_1011110110011111"; -- 0.10360322123897299
	pesos_i(2695) := b"1111111111111111_1111111111111111_1111110100111100_1001100001111111"; -- -0.010794133169870816
	pesos_i(2696) := b"0000000000000000_0000000000000000_0001101110000111_1001100000010110"; -- 0.1075377516010025
	pesos_i(2697) := b"1111111111111111_1111111111111111_1101011011011110_0010110111100100"; -- -0.16067231363435336
	pesos_i(2698) := b"1111111111111111_1111111111111111_1101010101000111_1100001010110010"; -- -0.16687377112757498
	pesos_i(2699) := b"1111111111111111_1111111111111111_1111110001011110_0001111111101111"; -- -0.014188770386174806
	pesos_i(2700) := b"0000000000000000_0000000000000000_0001110000000001_0100011111100001"; -- 0.10939454312118344
	pesos_i(2701) := b"0000000000000000_0000000000000000_0001110101111001_0111110110100101"; -- 0.11513505251434951
	pesos_i(2702) := b"0000000000000000_0000000000000000_0000010101101110_0100010010110101"; -- 0.02121381197228651
	pesos_i(2703) := b"1111111111111111_1111111111111111_1101101110111000_1100011101000110"; -- -0.1417117552173094
	pesos_i(2704) := b"1111111111111111_1111111111111111_1101011011111111_1110010111000000"; -- -0.1601578146947883
	pesos_i(2705) := b"1111111111111111_1111111111111111_1111011110110001_0000110010110101"; -- -0.03245468691955259
	pesos_i(2706) := b"0000000000000000_0000000000000000_0001011100001110_1001100010010011"; -- 0.09006646727699513
	pesos_i(2707) := b"0000000000000000_0000000000000000_0010101001110100_0001101000100101"; -- 0.16583407796975272
	pesos_i(2708) := b"0000000000000000_0000000000000000_0000000001100010_1100000010111011"; -- 0.0015068489634183276
	pesos_i(2709) := b"1111111111111111_1111111111111111_1101100100010000_1110010000011011"; -- -0.15208601322846854
	pesos_i(2710) := b"0000000000000000_0000000000000000_0001110111001010_1001110001110111"; -- 0.11637285149239326
	pesos_i(2711) := b"1111111111111111_1111111111111111_1110101011001100_0111011111100110"; -- -0.08281756050971316
	pesos_i(2712) := b"0000000000000000_0000000000000000_0001110110011100_0111100110011000"; -- 0.11566886872973403
	pesos_i(2713) := b"1111111111111111_1111111111111111_1111111101100111_0100110011110111"; -- -0.0023300073255781892
	pesos_i(2714) := b"0000000000000000_0000000000000000_0000111010011000_1101000101111111"; -- 0.05701932284881705
	pesos_i(2715) := b"1111111111111111_1111111111111111_1110010000111000_0001110011010101"; -- -0.10851878937902161
	pesos_i(2716) := b"1111111111111111_1111111111111111_1111110000100000_0011110000111001"; -- -0.015133129208480697
	pesos_i(2717) := b"1111111111111111_1111111111111111_1111011110110010_1101111101000000"; -- -0.03242687879338731
	pesos_i(2718) := b"0000000000000000_0000000000000000_0000000010111011_0000111001001100"; -- 0.0028542456685323524
	pesos_i(2719) := b"1111111111111111_1111111111111111_1110000101100001_1010011110110011"; -- -0.11960365189959814
	pesos_i(2720) := b"0000000000000000_0000000000000000_0010011001001010_0010101101001100"; -- 0.14956923115431456
	pesos_i(2721) := b"0000000000000000_0000000000000000_0001111011100001_0110000011000010"; -- 0.1206264947199018
	pesos_i(2722) := b"1111111111111111_1111111111111111_1110100011111010_0101001010010100"; -- -0.08993038061928908
	pesos_i(2723) := b"1111111111111111_1111111111111111_1110111010100000_0110100101001010"; -- -0.06786481802350673
	pesos_i(2724) := b"0000000000000000_0000000000000000_0000101110000001_1101010011010111"; -- 0.04494981994143466
	pesos_i(2725) := b"1111111111111111_1111111111111111_1110101000010000_0111000110111111"; -- -0.08568657948631514
	pesos_i(2726) := b"1111111111111111_1111111111111111_1111011100000100_0111101011010011"; -- -0.03508789392740833
	pesos_i(2727) := b"1111111111111111_1111111111111111_1101010010010011_0010100001111101"; -- -0.1696295447796503
	pesos_i(2728) := b"0000000000000000_0000000000000000_0010010001000111_1100000000011110"; -- 0.14171982510973238
	pesos_i(2729) := b"0000000000000000_0000000000000000_0010000100110000_1101010000111100"; -- 0.12965132202487917
	pesos_i(2730) := b"0000000000000000_0000000000000000_0000001111110011_1101001111010110"; -- 0.015439262207807896
	pesos_i(2731) := b"1111111111111111_1111111111111111_1111100001110100_0100001001011100"; -- -0.0294760250894409
	pesos_i(2732) := b"1111111111111111_1111111111111111_1110101000011010_0010111101010011"; -- -0.08553795078943312
	pesos_i(2733) := b"0000000000000000_0000000000000000_0001100100101010_1010010100010101"; -- 0.09830695876559727
	pesos_i(2734) := b"0000000000000000_0000000000000000_0001011000101101_0011111100111110"; -- 0.08662791504287078
	pesos_i(2735) := b"1111111111111111_1111111111111111_1111000001100111_0001010001100011"; -- -0.06092712955137978
	pesos_i(2736) := b"0000000000000000_0000000000000000_0000001101010111_0010110011011101"; -- 0.013048938714391306
	pesos_i(2737) := b"1111111111111111_1111111111111111_1101011010011111_1100111001101010"; -- -0.16162404935355193
	pesos_i(2738) := b"0000000000000000_0000000000000000_0010000010111000_1100100100110101"; -- 0.1278196100707952
	pesos_i(2739) := b"1111111111111111_1111111111111111_1110101110110010_0011111100101110"; -- -0.07931141975398973
	pesos_i(2740) := b"1111111111111111_1111111111111111_1111110110000000_0101011101011001"; -- -0.009760418707331162
	pesos_i(2741) := b"1111111111111111_1111111111111111_1101011011110010_0011100100001001"; -- -0.16036647349252184
	pesos_i(2742) := b"0000000000000000_0000000000000000_0010100101100001_1011101011110110"; -- 0.16164749623691851
	pesos_i(2743) := b"1111111111111111_1111111111111111_1110101011111101_1011000110101101"; -- -0.08206643601220724
	pesos_i(2744) := b"1111111111111111_1111111111111111_1101100110010010_1100101110100111"; -- -0.150103828151429
	pesos_i(2745) := b"0000000000000000_0000000000000000_0001110100000111_1010101000111110"; -- 0.11339820875735462
	pesos_i(2746) := b"0000000000000000_0000000000000000_0010010010010100_1011100110010001"; -- 0.1428943613524545
	pesos_i(2747) := b"0000000000000000_0000000000000000_0000101111010000_0101111011110111"; -- 0.04614823847247986
	pesos_i(2748) := b"1111111111111111_1111111111111111_1110111110010000_1000111110111101"; -- -0.06420041694532543
	pesos_i(2749) := b"1111111111111111_1111111111111111_1110100110001001_0111001110100110"; -- -0.0877464027719013
	pesos_i(2750) := b"0000000000000000_0000000000000000_0000000011000100_1100111110111111"; -- 0.0030031053115922458
	pesos_i(2751) := b"0000000000000000_0000000000000000_0010101101010000_1010110010100111"; -- 0.16919974410271837
	pesos_i(2752) := b"0000000000000000_0000000000000000_0001011101000011_1100100010110010"; -- 0.09087805129703044
	pesos_i(2753) := b"0000000000000000_0000000000000000_0000000000101010_1000010000110100"; -- 0.0006487490197798908
	pesos_i(2754) := b"1111111111111111_1111111111111111_1101100100011110_1101000010101010"; -- -0.15187354889720847
	pesos_i(2755) := b"1111111111111111_1111111111111111_1111011001010110_0000110110011110"; -- -0.03774943257941761
	pesos_i(2756) := b"1111111111111111_1111111111111111_1101111101000101_1111101001100011"; -- -0.1278384694192543
	pesos_i(2757) := b"0000000000000000_0000000000000000_0000101111110010_0100111010101010"; -- 0.046666065640600815
	pesos_i(2758) := b"1111111111111111_1111111111111111_1111000011100010_0101001100100111"; -- -0.05904655735204573
	pesos_i(2759) := b"1111111111111111_1111111111111111_1101110011000010_1011011010101000"; -- -0.13765390781722248
	pesos_i(2760) := b"1111111111111111_1111111111111111_1110111110111001_1000111011100111"; -- -0.06357485645347687
	pesos_i(2761) := b"0000000000000000_0000000000000000_0000111001011001_1111101010010111"; -- 0.05606046864997989
	pesos_i(2762) := b"1111111111111111_1111111111111111_1111100101111100_0100001011111100"; -- -0.0254476676238492
	pesos_i(2763) := b"0000000000000000_0000000000000000_0010000001000011_1111001111001001"; -- 0.1260368695522482
	pesos_i(2764) := b"0000000000000000_0000000000000000_0001101011001101_0010000111011101"; -- 0.10469257006921423
	pesos_i(2765) := b"1111111111111111_1111111111111111_1111010101110111_0110000110101110"; -- -0.041147131857189476
	pesos_i(2766) := b"1111111111111111_1111111111111111_1101010010001101_1011000100011111"; -- -0.1697129534919399
	pesos_i(2767) := b"1111111111111111_1111111111111111_1110111110100001_1110100000101001"; -- -0.06393574712589073
	pesos_i(2768) := b"1111111111111111_1111111111111111_1111110110111101_1111101110101010"; -- -0.008819838420660642
	pesos_i(2769) := b"1111111111111111_1111111111111111_1110100010101100_1000010100111110"; -- -0.09111754646212572
	pesos_i(2770) := b"0000000000000000_0000000000000000_0010010011011111_1010110010100010"; -- 0.14403799967902486
	pesos_i(2771) := b"0000000000000000_0000000000000000_0000011100000110_1111101000110011"; -- 0.027450215703191838
	pesos_i(2772) := b"1111111111111111_1111111111111111_1110010100001011_1111001001001110"; -- -0.10528646085521123
	pesos_i(2773) := b"0000000000000000_0000000000000000_0001010011101100_1000000111111001"; -- 0.0817338211344116
	pesos_i(2774) := b"0000000000000000_0000000000000000_0000000110111001_1111010101110011"; -- 0.006743755996553319
	pesos_i(2775) := b"0000000000000000_0000000000000000_0001011000110110_0100110001001101"; -- 0.0867660225286448
	pesos_i(2776) := b"1111111111111111_1111111111111111_1101110101110100_1011101111111000"; -- -0.1349375265623887
	pesos_i(2777) := b"0000000000000000_0000000000000000_0010001111011111_0110100000110010"; -- 0.14012767056445677
	pesos_i(2778) := b"0000000000000000_0000000000000000_0010100000110001_0001111100011100"; -- 0.1569995348628522
	pesos_i(2779) := b"0000000000000000_0000000000000000_0000100100011111_0111010011100011"; -- 0.03563623953944284
	pesos_i(2780) := b"1111111111111111_1111111111111111_1111011001011010_0110111010000010"; -- -0.03768262218238733
	pesos_i(2781) := b"1111111111111111_1111111111111111_1111100110101100_0011111100000111"; -- -0.02471548155962449
	pesos_i(2782) := b"1111111111111111_1111111111111111_1111101000101101_0001001101100101"; -- -0.02274969859795366
	pesos_i(2783) := b"0000000000000000_0000000000000000_0000111111001011_0101010011001111"; -- 0.06169633913092046
	pesos_i(2784) := b"0000000000000000_0000000000000000_0001001110101011_0000100110000110"; -- 0.07682857066197127
	pesos_i(2785) := b"1111111111111111_1111111111111111_1110100000100100_0000100010000011"; -- -0.09320017617993898
	pesos_i(2786) := b"1111111111111111_1111111111111111_1101011111100010_0100011010101101"; -- -0.1567035510840621
	pesos_i(2787) := b"1111111111111111_1111111111111111_1111100111110110_1001011101000110"; -- -0.023581071248889657
	pesos_i(2788) := b"0000000000000000_0000000000000000_0001000111000010_1010111000011111"; -- 0.06937683353209512
	pesos_i(2789) := b"0000000000000000_0000000000000000_0000100001101001_1111101110001010"; -- 0.03286716567825254
	pesos_i(2790) := b"1111111111111111_1111111111111111_1110110011101000_0111110101010100"; -- -0.07457749086657965
	pesos_i(2791) := b"0000000000000000_0000000000000000_0010101011101110_0001100011111110"; -- 0.1676955814312269
	pesos_i(2792) := b"1111111111111111_1111111111111111_1111111001010001_1110001101010011"; -- -0.006562988538330955
	pesos_i(2793) := b"1111111111111111_1111111111111111_1101111111100110_1100010101110100"; -- -0.12538495946153053
	pesos_i(2794) := b"0000000000000000_0000000000000000_0010000011001110_0001110111010101"; -- 0.1281450886485254
	pesos_i(2795) := b"0000000000000000_0000000000000000_0010010000011111_1000110110010010"; -- 0.14110646082040945
	pesos_i(2796) := b"1111111111111111_1111111111111111_1111001101011100_1110011011110011"; -- -0.049363675705852074
	pesos_i(2797) := b"1111111111111111_1111111111111111_1111101000000001_1100101010110101"; -- -0.023410158916311527
	pesos_i(2798) := b"0000000000000000_0000000000000000_0000001011101011_1111011000101100"; -- 0.011412988483640134
	pesos_i(2799) := b"1111111111111111_1111111111111111_1110001111101000_1010010100100110"; -- -0.10973136729993224
	pesos_i(2800) := b"1111111111111111_1111111111111111_1101110100011001_1011110101011111"; -- -0.13632599286143365
	pesos_i(2801) := b"1111111111111111_1111111111111111_1111001010110001_1110110101110101"; -- -0.05197254068302777
	pesos_i(2802) := b"1111111111111111_1111111111111111_1110101001001100_1001000110001010"; -- -0.08476915720646469
	pesos_i(2803) := b"1111111111111111_1111111111111111_1111100011011110_1110110001000010"; -- -0.02784846665108609
	pesos_i(2804) := b"1111111111111111_1111111111111111_1101110110001111_0111111111110100"; -- -0.13452911651776567
	pesos_i(2805) := b"1111111111111111_1111111111111111_1110101001111101_1001011110111000"; -- -0.08402110818526203
	pesos_i(2806) := b"1111111111111111_1111111111111111_1101111000110000_1110101100110110"; -- -0.13206605841767688
	pesos_i(2807) := b"0000000000000000_0000000000000000_0001110100010011_0101101110000001"; -- 0.11357662103842144
	pesos_i(2808) := b"1111111111111111_1111111111111111_1111000010011101_0011110001001011"; -- -0.06010077648980408
	pesos_i(2809) := b"0000000000000000_0000000000000000_0000001000100010_0101000000010010"; -- 0.008336071486268028
	pesos_i(2810) := b"0000000000000000_0000000000000000_0001111110100111_1011010011101111"; -- 0.12365275216868311
	pesos_i(2811) := b"1111111111111111_1111111111111111_1110000100010001_1101011011001001"; -- -0.12082154849675261
	pesos_i(2812) := b"0000000000000000_0000000000000000_0000111101011101_1000100001101010"; -- 0.06002094835506136
	pesos_i(2813) := b"0000000000000000_0000000000000000_0000111111110010_1110010010000010"; -- 0.06229999710224113
	pesos_i(2814) := b"0000000000000000_0000000000000000_0001101011011010_0000110110101101"; -- 0.10488973121097815
	pesos_i(2815) := b"0000000000000000_0000000000000000_0001011010001111_0110000010001011"; -- 0.08812526115816993
	pesos_i(2816) := b"0000000000000000_0000000000000000_0010110010101000_0111011110010010"; -- 0.17444560360937186
	pesos_i(2817) := b"0000000000000000_0000000000000000_0001101000010111_1011010110010000"; -- 0.10192427400226516
	pesos_i(2818) := b"1111111111111111_1111111111111111_1101000110010110_1010000111100001"; -- -0.1812952829751957
	pesos_i(2819) := b"0000000000000000_0000000000000000_0000011010100111_1111000110101000"; -- 0.02600012158798036
	pesos_i(2820) := b"0000000000000000_0000000000000000_0001001111100111_0010011001011111"; -- 0.07774581728531575
	pesos_i(2821) := b"0000000000000000_0000000000000000_0001010010001101_1100111000011111"; -- 0.08028877496273751
	pesos_i(2822) := b"1111111111111111_1111111111111111_1101111111001111_0101100110101111"; -- -0.12574233499175824
	pesos_i(2823) := b"0000000000000000_0000000000000000_0000100001001110_0010101100001000"; -- 0.03244275036066918
	pesos_i(2824) := b"1111111111111111_1111111111111111_1111111100101100_0001110110100011"; -- -0.003233096888148693
	pesos_i(2825) := b"1111111111111111_1111111111111111_1111001001001101_0101110100011100"; -- -0.05350702352943085
	pesos_i(2826) := b"0000000000000000_0000000000000000_0000101111100000_0000101001110111"; -- 0.046387342443137594
	pesos_i(2827) := b"1111111111111111_1111111111111111_1111111111111011_1000010101011111"; -- -6.834433449574716e-05
	pesos_i(2828) := b"1111111111111111_1111111111111111_1111001000100110_0010100011101000"; -- -0.054105227862207325
	pesos_i(2829) := b"0000000000000000_0000000000000000_0010101000101110_1100101100011010"; -- 0.16477651013726854
	pesos_i(2830) := b"0000000000000000_0000000000000000_0010000100001110_1100010011101000"; -- 0.12913160952256206
	pesos_i(2831) := b"1111111111111111_1111111111111111_1111110110001110_0000101111111010"; -- -0.009551288049258446
	pesos_i(2832) := b"1111111111111111_1111111111111111_1101100011001001_1111101001101110"; -- -0.15316805651636814
	pesos_i(2833) := b"1111111111111111_1111111111111111_1111000000101111_1110000001011110"; -- -0.06176946354164776
	pesos_i(2834) := b"1111111111111111_1111111111111111_1110100111011000_1000011010010100"; -- -0.08653983016249792
	pesos_i(2835) := b"0000000000000000_0000000000000000_0001011110101000_0101110100010001"; -- 0.09241277378641673
	pesos_i(2836) := b"0000000000000000_0000000000000000_0001000010001010_0000010011010010"; -- 0.06460600025761833
	pesos_i(2837) := b"0000000000000000_0000000000000000_0000110110000011_0010101111001101"; -- 0.05278276219296256
	pesos_i(2838) := b"1111111111111111_1111111111111111_1110001000101010_1101110010100010"; -- -0.11653348001531766
	pesos_i(2839) := b"1111111111111111_1111111111111111_1110110001010101_0000001100000000"; -- -0.07682782407517155
	pesos_i(2840) := b"1111111111111111_1111111111111111_1100011100011110_1101001001000001"; -- -0.22218595411744171
	pesos_i(2841) := b"0000000000000000_0000000000000000_0010000010010000_1110111000000001"; -- 0.12721145175459095
	pesos_i(2842) := b"1111111111111111_1111111111111111_1111101011101010_1001001010000001"; -- -0.01985821102239637
	pesos_i(2843) := b"1111111111111111_1111111111111111_1111101110110101_1000101010110110"; -- -0.01676114140520226
	pesos_i(2844) := b"1111111111111111_1111111111111111_1111001110111101_0100001111010010"; -- -0.04789329651213095
	pesos_i(2845) := b"0000000000000000_0000000000000000_0001001110111010_0101110110100110"; -- 0.0770624665903193
	pesos_i(2846) := b"0000000000000000_0000000000000000_0000011011111001_1100100101010111"; -- 0.027248939156192174
	pesos_i(2847) := b"0000000000000000_0000000000000000_0010101100001100_1011011011110010"; -- 0.16816275996220562
	pesos_i(2848) := b"1111111111111111_1111111111111111_1111000101111011_1000110110100010"; -- -0.056708476906872474
	pesos_i(2849) := b"1111111111111111_1111111111111111_1111001000110100_1100010101011110"; -- -0.05388227892270983
	pesos_i(2850) := b"0000000000000000_0000000000000000_0010010000011001_0101111011011001"; -- 0.14101212310689484
	pesos_i(2851) := b"1111111111111111_1111111111111111_1111100111100110_0110000010001100"; -- -0.023828473898288172
	pesos_i(2852) := b"1111111111111111_1111111111111111_1111101100010010_1011100100010010"; -- -0.019245560835550603
	pesos_i(2853) := b"0000000000000000_0000000000000000_0000011100010000_1100000111011001"; -- 0.027599444825333986
	pesos_i(2854) := b"1111111111111111_1111111111111111_1111010011111100_0100000111110100"; -- -0.043025854039046026
	pesos_i(2855) := b"1111111111111111_1111111111111111_1110011100000000_0100011011110100"; -- -0.09765202097910253
	pesos_i(2856) := b"1111111111111111_1111111111111111_1110001111100010_1010000011011001"; -- -0.10982317645907848
	pesos_i(2857) := b"1111111111111111_1111111111111111_1110111000011111_1001010000010001"; -- -0.06983065215293303
	pesos_i(2858) := b"0000000000000000_0000000000000000_0010000010101001_1000010100100010"; -- 0.12758667069640078
	pesos_i(2859) := b"0000000000000000_0000000000000000_0000100001101100_0111100100110111"; -- 0.03290517408401251
	pesos_i(2860) := b"1111111111111111_1111111111111111_1110010100000011_0111100000111011"; -- -0.10541580737643144
	pesos_i(2861) := b"0000000000000000_0000000000000000_0001000101111010_0111101010101011"; -- 0.06827513392480689
	pesos_i(2862) := b"1111111111111111_1111111111111111_1111101101100100_0000001111000010"; -- -0.01800514710838588
	pesos_i(2863) := b"1111111111111111_1111111111111111_1101101101110110_0000110011000010"; -- -0.14272995255248921
	pesos_i(2864) := b"0000000000000000_0000000000000000_0000000101110000_1100011000110000"; -- 0.005627047324300499
	pesos_i(2865) := b"0000000000000000_0000000000000000_0000100100110111_0010100011110010"; -- 0.03599792387801481
	pesos_i(2866) := b"1111111111111111_1111111111111111_1101111001001110_1000010101101000"; -- -0.13161436291291911
	pesos_i(2867) := b"0000000000000000_0000000000000000_0010010010111010_1001000100101001"; -- 0.14347178705661118
	pesos_i(2868) := b"0000000000000000_0000000000000000_0000100000101000_1110101001000110"; -- 0.03187431526609526
	pesos_i(2869) := b"1111111111111111_1111111111111111_1110100100111010_1010010111100110"; -- -0.08894885197833564
	pesos_i(2870) := b"1111111111111111_1111111111111111_1110111001000011_1011010100001000"; -- -0.06927937083643518
	pesos_i(2871) := b"0000000000000000_0000000000000000_0000010111001100_1101010100011001"; -- 0.02265674463041658
	pesos_i(2872) := b"1111111111111111_1111111111111111_1110010100110000_0001011011111110"; -- -0.10473495775112779
	pesos_i(2873) := b"0000000000000000_0000000000000000_0001001101001111_0001111101000011"; -- 0.07542605767433765
	pesos_i(2874) := b"1111111111111111_1111111111111111_1110000111011110_0101001101000001"; -- -0.11770133647469523
	pesos_i(2875) := b"1111111111111111_1111111111111111_1111111010000110_1101110010000010"; -- -0.005754679032338951
	pesos_i(2876) := b"1111111111111111_1111111111111111_1101001001101101_1001101100000001"; -- -0.17801505297720654
	pesos_i(2877) := b"1111111111111111_1111111111111111_1110011100000000_1110001101000000"; -- -0.0976427048755889
	pesos_i(2878) := b"1111111111111111_1111111111111111_1111101010101111_1011110111101110"; -- -0.020755891313696574
	pesos_i(2879) := b"0000000000000000_0000000000000000_0000101011100100_1110000010010100"; -- 0.042554889778036585
	pesos_i(2880) := b"1111111111111111_1111111111111111_1110101001000111_0110000100010011"; -- -0.0848483399465306
	pesos_i(2881) := b"1111111111111111_1111111111111111_1101110010011000_0001100100011110"; -- -0.13830416707619417
	pesos_i(2882) := b"0000000000000000_0000000000000000_0010010010110001_0110001001010100"; -- 0.14333166649604703
	pesos_i(2883) := b"1111111111111111_1111111111111111_1101111110001101_1000001001100010"; -- -0.1267469892890572
	pesos_i(2884) := b"0000000000000000_0000000000000000_0001101100011001_0000100101010111"; -- 0.10585077647979982
	pesos_i(2885) := b"1111111111111111_1111111111111111_1110001110011100_1010010101011011"; -- -0.11089102285533603
	pesos_i(2886) := b"1111111111111111_1111111111111111_1111111110000001_1111101111101111"; -- -0.0019228498706773758
	pesos_i(2887) := b"1111111111111111_1111111111111111_1101110011010000_0000111110000001"; -- -0.13745024784939675
	pesos_i(2888) := b"1111111111111111_1111111111111111_1110110100011100_0111110101010010"; -- -0.07378403425800376
	pesos_i(2889) := b"0000000000000000_0000000000000000_0010001110100100_1110011010010110"; -- 0.13923493529975375
	pesos_i(2890) := b"1111111111111111_1111111111111111_1111011100111110_0101010001000100"; -- -0.034205182527422745
	pesos_i(2891) := b"0000000000000000_0000000000000000_0001110000101010_1100101010001100"; -- 0.1100279418379223
	pesos_i(2892) := b"0000000000000000_0000000000000000_0000011101100111_0010100000110111"; -- 0.028917802362717016
	pesos_i(2893) := b"1111111111111111_1111111111111111_1111000010111001_1110111010101110"; -- -0.059662897593360686
	pesos_i(2894) := b"0000000000000000_0000000000000000_0010000110100011_1000101001101101"; -- 0.13140168342722533
	pesos_i(2895) := b"1111111111111111_1111111111111111_1111101001011100_1010011001110100"; -- -0.022023769916794247
	pesos_i(2896) := b"1111111111111111_1111111111111111_1111010011101101_0110101011100100"; -- -0.04325229583779752
	pesos_i(2897) := b"1111111111111111_1111111111111111_1110001100000001_0010011011011010"; -- -0.11326367547647398
	pesos_i(2898) := b"0000000000000000_0000000000000000_0010100011000010_0001011110011100"; -- 0.1592116123478211
	pesos_i(2899) := b"1111111111111111_1111111111111111_1111001001101111_1000011101011111"; -- -0.05298570562157436
	pesos_i(2900) := b"0000000000000000_0000000000000000_0010001100100010_0001010010101110"; -- 0.13723878145270751
	pesos_i(2901) := b"1111111111111111_1111111111111111_1111101011111101_0101001001111001"; -- -0.019572110568996607
	pesos_i(2902) := b"1111111111111111_1111111111111111_1111101100011010_1101000111100011"; -- -0.01912201125036712
	pesos_i(2903) := b"0000000000000000_0000000000000000_0001001011010111_0111000110010111"; -- 0.07359991014167527
	pesos_i(2904) := b"1111111111111111_1111111111111111_1110001000000110_1000111011111111"; -- -0.11708742397202551
	pesos_i(2905) := b"0000000000000000_0000000000000000_0001010101111101_0111011110101110"; -- 0.08394573200249061
	pesos_i(2906) := b"0000000000000000_0000000000000000_0001001110111110_1110100111001111"; -- 0.07713185610180523
	pesos_i(2907) := b"0000000000000000_0000000000000000_0010001011010011_1101011100010001"; -- 0.13604492342956193
	pesos_i(2908) := b"0000000000000000_0000000000000000_0000110110011010_1010001000111110"; -- 0.05314077399683289
	pesos_i(2909) := b"1111111111111111_1111111111111111_1110000011001111_1010011010110000"; -- -0.12183149537645396
	pesos_i(2910) := b"0000000000000000_0000000000000000_0000111000001110_0000000111010110"; -- 0.05490123241421827
	pesos_i(2911) := b"1111111111111111_1111111111111111_1101101111010111_1101100111111110"; -- -0.1412376169648894
	pesos_i(2912) := b"0000000000000000_0000000000000000_0010000100001101_0010011000110111"; -- 0.1291068920880928
	pesos_i(2913) := b"0000000000000000_0000000000000000_0001100100010000_1011010100100000"; -- 0.09791118655831016
	pesos_i(2914) := b"0000000000000000_0000000000000000_0000111110111000_0101001100011011"; -- 0.061406320629533426
	pesos_i(2915) := b"0000000000000000_0000000000000000_0001000110000101_1010110101011000"; -- 0.06844600097563386
	pesos_i(2916) := b"0000000000000000_0000000000000000_0000100011010111_1001010100110000"; -- 0.03453953189364819
	pesos_i(2917) := b"0000000000000000_0000000000000000_0001111001000111_0100001000101100"; -- 0.11827481824462695
	pesos_i(2918) := b"1111111111111111_1111111111111111_1110100101100110_0101110100010101"; -- -0.0882818053325227
	pesos_i(2919) := b"1111111111111111_1111111111111111_1111011010010000_1111011110101001"; -- -0.03685047257493526
	pesos_i(2920) := b"0000000000000000_0000000000000000_0000110100001001_1011001000110001"; -- 0.05092920010475577
	pesos_i(2921) := b"0000000000000000_0000000000000000_0010001110001001_0111000101010011"; -- 0.13881595876850306
	pesos_i(2922) := b"1111111111111111_1111111111111111_1110001001001101_1000010111010000"; -- -0.11600459744887064
	pesos_i(2923) := b"1111111111111111_1111111111111111_1101100011111000_0001100110111010"; -- -0.15246428695582045
	pesos_i(2924) := b"1111111111111111_1111111111111111_1111111000101000_0100111010100010"; -- -0.007197461526234888
	pesos_i(2925) := b"0000000000000000_0000000000000000_0010100111111010_0001101101100110"; -- 0.16397258027478964
	pesos_i(2926) := b"1111111111111111_1111111111111111_1111010111110011_0010110010110011"; -- -0.03925820004934258
	pesos_i(2927) := b"1111111111111111_1111111111111111_1111000101001101_1110110101011100"; -- -0.057404675479129856
	pesos_i(2928) := b"0000000000000000_0000000000000000_0001010001011010_0011100011111110"; -- 0.07950168800209254
	pesos_i(2929) := b"1111111111111111_1111111111111111_1111011001010011_0000001011010011"; -- -0.03779585212589216
	pesos_i(2930) := b"1111111111111111_1111111111111111_1110011011011010_0001010110110110"; -- -0.09823478997726798
	pesos_i(2931) := b"1111111111111111_1111111111111111_1111110000011100_0101010111010100"; -- -0.015192638048284598
	pesos_i(2932) := b"1111111111111111_1111111111111111_1101101110000111_1111000111001101"; -- -0.14245690110385983
	pesos_i(2933) := b"0000000000000000_0000000000000000_0000100111000011_1011001000010011"; -- 0.03814232788093169
	pesos_i(2934) := b"0000000000000000_0000000000000000_0001011011101110_1101010011111011"; -- 0.089581786408238
	pesos_i(2935) := b"0000000000000000_0000000000000000_0001001010010001_1000100101011000"; -- 0.07253321084950176
	pesos_i(2936) := b"0000000000000000_0000000000000000_0000101100100011_0111110001011111"; -- 0.0435102207536302
	pesos_i(2937) := b"0000000000000000_0000000000000000_0000000010100101_0011100110111011"; -- 0.0025211411731128758
	pesos_i(2938) := b"1111111111111111_1111111111111111_1110011001010000_1110100010111100"; -- -0.10032792480473607
	pesos_i(2939) := b"1111111111111111_1111111111111111_1110001101010011_1101011100110110"; -- -0.11200194286298551
	pesos_i(2940) := b"0000000000000000_0000000000000000_0001110110001010_0111010000100011"; -- 0.11539388509724897
	pesos_i(2941) := b"1111111111111111_1111111111111111_1111110000001110_0010000001111111"; -- -0.015409440076125068
	pesos_i(2942) := b"1111111111111111_1111111111111111_1110010111111111_1100101001100001"; -- -0.10156569605182245
	pesos_i(2943) := b"1111111111111111_1111111111111111_1101000010111010_0001100011101000"; -- -0.18466038059031997
	pesos_i(2944) := b"1111111111111111_1111111111111111_1111000010111100_1111111001110110"; -- -0.05961618058501193
	pesos_i(2945) := b"1111111111111111_1111111111111111_1111011011010110_1100010111111010"; -- -0.035785318716689524
	pesos_i(2946) := b"0000000000000000_0000000000000000_0000111111000011_1001101101101101"; -- 0.06157847792174139
	pesos_i(2947) := b"0000000000000000_0000000000000000_0000000110001001_0001011110000110"; -- 0.005998106225511403
	pesos_i(2948) := b"0000000000000000_0000000000000000_0001101100010001_0010010000110111"; -- 0.10573030807785683
	pesos_i(2949) := b"0000000000000000_0000000000000000_0001101001101100_1111011101000111"; -- 0.10322518800498345
	pesos_i(2950) := b"0000000000000000_0000000000000000_0001001101101101_0010100110001111"; -- 0.07588443516799157
	pesos_i(2951) := b"0000000000000000_0000000000000000_0000110011001110_0010100110001001"; -- 0.050020786125895604
	pesos_i(2952) := b"0000000000000000_0000000000000000_0001011010110000_0111111100011001"; -- 0.08863062251966455
	pesos_i(2953) := b"0000000000000000_0000000000000000_0001011010110010_0111011011111101"; -- 0.08866065666565141
	pesos_i(2954) := b"0000000000000000_0000000000000000_0001010110010100_1100000101110100"; -- 0.08430108143106368
	pesos_i(2955) := b"1111111111111111_1111111111111111_1110111111000101_1010010000111110"; -- -0.06339047898373192
	pesos_i(2956) := b"1111111111111111_1111111111111111_1110000101001110_0010011010011111"; -- -0.11990126236026959
	pesos_i(2957) := b"0000000000000000_0000000000000000_0001101000110111_0111010101100001"; -- 0.10240872981646337
	pesos_i(2958) := b"0000000000000000_0000000000000000_0000001101010110_1101001000110011"; -- 0.013043534697720145
	pesos_i(2959) := b"1111111111111111_1111111111111111_1110010011011110_0100010100011000"; -- -0.10598343061679028
	pesos_i(2960) := b"1111111111111111_1111111111111111_1111010011111101_0001000011100010"; -- -0.04301351997503294
	pesos_i(2961) := b"1111111111111111_1111111111111111_1111010101110011_1101100010101010"; -- -0.04120107511018473
	pesos_i(2962) := b"1111111111111111_1111111111111111_1101110111001000_0101001111101010"; -- -0.13366199059119316
	pesos_i(2963) := b"1111111111111111_1111111111111111_1110000001111100_0000100010110100"; -- -0.12310739129682007
	pesos_i(2964) := b"1111111111111111_1111111111111111_1111001011001001_0101010100110010"; -- -0.05161540545919529
	pesos_i(2965) := b"1111111111111111_1111111111111111_1111001011100111_1100000001101100"; -- -0.051151250512719196
	pesos_i(2966) := b"1111111111111111_1111111111111111_1110110101101011_1001110000001001"; -- -0.07257675907262537
	pesos_i(2967) := b"1111111111111111_1111111111111111_1111000010111001_0000011011111001"; -- -0.059676708449467396
	pesos_i(2968) := b"1111111111111111_1111111111111111_1111111111001110_1010111000101010"; -- -0.0007525585154242239
	pesos_i(2969) := b"0000000000000000_0000000000000000_0010100010010100_1110000110111100"; -- 0.15852175555848697
	pesos_i(2970) := b"0000000000000000_0000000000000000_0010001100101111_0111111101110011"; -- 0.13744350968056163
	pesos_i(2971) := b"0000000000000000_0000000000000000_0000111110001101_1010001010110110"; -- 0.060754937620119645
	pesos_i(2972) := b"0000000000000000_0000000000000000_0000110100101100_0001010110011110"; -- 0.05145392520740647
	pesos_i(2973) := b"1111111111111111_1111111111111111_1111001000110100_1100111010000001"; -- -0.05388173435021811
	pesos_i(2974) := b"1111111111111111_1111111111111111_1111111100001110_0010000100010101"; -- -0.003690655205953567
	pesos_i(2975) := b"1111111111111111_1111111111111111_1101111000101000_0101000101010101"; -- -0.13219730062995816
	pesos_i(2976) := b"1111111111111111_1111111111111111_1110100001010101_0000110110000101"; -- -0.09245219706673274
	pesos_i(2977) := b"0000000000000000_0000000000000000_0010001001101110_1010000000110100"; -- 0.1345005155635028
	pesos_i(2978) := b"0000000000000000_0000000000000000_0010100001010001_1000010010111100"; -- 0.15749387344984853
	pesos_i(2979) := b"0000000000000000_0000000000000000_0001110001011111_1110011000000000"; -- 0.11083829394485219
	pesos_i(2980) := b"1111111111111111_1111111111111111_1111101101010110_1110101111110001"; -- -0.01820493086547407
	pesos_i(2981) := b"0000000000000000_0000000000000000_0000110100010101_1111100100110001"; -- 0.05111653762186401
	pesos_i(2982) := b"0000000000000000_0000000000000000_0001000000110000_1110110010101111"; -- 0.06324652935079068
	pesos_i(2983) := b"0000000000000000_0000000000000000_0001010100111100_1100101011100011"; -- 0.08295887025098617
	pesos_i(2984) := b"0000000000000000_0000000000000000_0010101000010100_0101000011001011"; -- 0.1643724913200794
	pesos_i(2985) := b"1111111111111111_1111111111111111_1101011011000010_1000111110011100"; -- -0.1610937351914458
	pesos_i(2986) := b"0000000000000000_0000000000000000_0000110010101110_1100110101101100"; -- 0.04954227335557256
	pesos_i(2987) := b"0000000000000000_0000000000000000_0000001001001111_1111010111000100"; -- 0.009032593161943712
	pesos_i(2988) := b"1111111111111111_1111111111111111_1110010111011010_0100010111011100"; -- -0.10213816997656064
	pesos_i(2989) := b"0000000000000000_0000000000000000_0000000110000001_0000100001001101"; -- 0.0058751284458087505
	pesos_i(2990) := b"0000000000000000_0000000000000000_0000111101100110_0101101110111101"; -- 0.06015561450862097
	pesos_i(2991) := b"1111111111111111_1111111111111111_1111000100010100_1100001011101000"; -- -0.05827695697147095
	pesos_i(2992) := b"1111111111111111_1111111111111111_1110000001001101_0011000000001011"; -- -0.12382220968181089
	pesos_i(2993) := b"0000000000000000_0000000000000000_0010001011011000_0110001001011111"; -- 0.13611426170172397
	pesos_i(2994) := b"0000000000000000_0000000000000000_0010011000110010_1000011110010011"; -- 0.14920852026639247
	pesos_i(2995) := b"0000000000000000_0000000000000000_0010011101011011_0101100110100111"; -- 0.15373764360336772
	pesos_i(2996) := b"1111111111111111_1111111111111111_1111000011000000_0111111100111100"; -- -0.05956272870683896
	pesos_i(2997) := b"0000000000000000_0000000000000000_0010011100011110_0110000110001110"; -- 0.15280732844242442
	pesos_i(2998) := b"1111111111111111_1111111111111111_1111000001010001_0111000000111101"; -- -0.061257348252735905
	pesos_i(2999) := b"0000000000000000_0000000000000000_0000100100000111_1100101000101001"; -- 0.03527511117097817
	pesos_i(3000) := b"1111111111111111_1111111111111111_1110110101111011_1110101111011101"; -- -0.07232786048699164
	pesos_i(3001) := b"1111111111111111_1111111111111111_1110011111001101_1000111011111011"; -- -0.09451967584139652
	pesos_i(3002) := b"1111111111111111_1111111111111111_1110101010000000_1000000100111011"; -- -0.08397667220325856
	pesos_i(3003) := b"0000000000000000_0000000000000000_0000010111100101_0101011001011111"; -- 0.023030660889887613
	pesos_i(3004) := b"0000000000000000_0000000000000000_0001100010001111_1001000111000111"; -- 0.09594069584100098
	pesos_i(3005) := b"0000000000000000_0000000000000000_0001101010111111_1001101010110001"; -- 0.10448614893867321
	pesos_i(3006) := b"1111111111111111_1111111111111111_1110110001001010_1010100100001000"; -- -0.07698577452970307
	pesos_i(3007) := b"1111111111111111_1111111111111111_1111010111111111_1110011010100011"; -- -0.03906401185540841
	pesos_i(3008) := b"0000000000000000_0000000000000000_0010011010101001_1001001001011110"; -- 0.15102495942653435
	pesos_i(3009) := b"0000000000000000_0000000000000000_0000101110001000_1010010001000111"; -- 0.045053737089776696
	pesos_i(3010) := b"0000000000000000_0000000000000000_0001001101100100_0110100011011011"; -- 0.07575087884941147
	pesos_i(3011) := b"0000000000000000_0000000000000000_0001100111101001_1111110010011001"; -- 0.1012266037699969
	pesos_i(3012) := b"0000000000000000_0000000000000000_0000001111111000_1001011000011001"; -- 0.015511876237216216
	pesos_i(3013) := b"0000000000000000_0000000000000000_0010011011000110_0001101001101010"; -- 0.1514603146390404
	pesos_i(3014) := b"0000000000000000_0000000000000000_0000011101000100_1110011110101001"; -- 0.028395155607789727
	pesos_i(3015) := b"0000000000000000_0000000000000000_0000110000100000_1000100000100110"; -- 0.047371396230286356
	pesos_i(3016) := b"0000000000000000_0000000000000000_0010000100011111_1001000100101100"; -- 0.12938792528605114
	pesos_i(3017) := b"1111111111111111_1111111111111111_1110110101100010_1101000111011101"; -- -0.07271087988173416
	pesos_i(3018) := b"0000000000000000_0000000000000000_0000100101000111_1001111110010000"; -- 0.03624913460175236
	pesos_i(3019) := b"0000000000000000_0000000000000000_0000001011111100_0000001000000110"; -- 0.011657835475752401
	pesos_i(3020) := b"1111111111111111_1111111111111111_1110101011011000_0110111100101010"; -- -0.082634975601689
	pesos_i(3021) := b"1111111111111111_1111111111111111_1111010001101010_0110001010001101"; -- -0.04525169436900684
	pesos_i(3022) := b"1111111111111111_1111111111111111_1111101111001110_0011011111010100"; -- -0.01638461189536695
	pesos_i(3023) := b"1111111111111111_1111111111111111_1111001100100101_0100011101101010"; -- -0.050212418171922506
	pesos_i(3024) := b"1111111111111111_1111111111111111_1101101101110101_0111010011001010"; -- -0.14273901057865324
	pesos_i(3025) := b"0000000000000000_0000000000000000_0001011100000101_0001010100000111"; -- 0.08992129736152421
	pesos_i(3026) := b"1111111111111111_1111111111111111_1110111001101101_1110000011011001"; -- -0.06863588992598009
	pesos_i(3027) := b"0000000000000000_0000000000000000_0000000000000011_0100101011011001"; -- 5.0237580812902256e-05
	pesos_i(3028) := b"0000000000000000_0000000000000000_0000101001100100_0110111000100000"; -- 0.040594942959563396
	pesos_i(3029) := b"0000000000000000_0000000000000000_0001101011011011_1101100100110010"; -- 0.10491712068847178
	pesos_i(3030) := b"1111111111111111_1111111111111111_1111010111111110_1101010000010100"; -- -0.039080376823993755
	pesos_i(3031) := b"1111111111111111_1111111111111111_1110111001100001_1100010110010111"; -- -0.06882062018901772
	pesos_i(3032) := b"1111111111111111_1111111111111111_1111000101010011_1110000111111101"; -- -0.05731380058443362
	pesos_i(3033) := b"1111111111111111_1111111111111111_1111000110110011_0001011100100101"; -- -0.05586104713247537
	pesos_i(3034) := b"1111111111111111_1111111111111111_1110010010000001_0111101001111000"; -- -0.1073993165904229
	pesos_i(3035) := b"0000000000000000_0000000000000000_0000100110101111_0010001101111010"; -- 0.03782865275032291
	pesos_i(3036) := b"0000000000000000_0000000000000000_0000100100001011_1110111011010010"; -- 0.035338331553652826
	pesos_i(3037) := b"1111111111111111_1111111111111111_1111111101000001_1010100011011010"; -- -0.0029043644390614803
	pesos_i(3038) := b"0000000000000000_0000000000000000_0001010101000010_0111001011110010"; -- 0.08304518126452623
	pesos_i(3039) := b"0000000000000000_0000000000000000_0000111010010101_1000111101010100"; -- 0.05696960264919873
	pesos_i(3040) := b"1111111111111111_1111111111111111_1101100000001001_0100110101101010"; -- -0.1561080567691706
	pesos_i(3041) := b"1111111111111111_1111111111111111_1110000000100010_1010000110001000"; -- -0.12447157320834894
	pesos_i(3042) := b"0000000000000000_0000000000000000_0010001010111110_0001110111001101"; -- 0.1357134461334215
	pesos_i(3043) := b"0000000000000000_0000000000000000_0001101100000100_0001101001011010"; -- 0.10553135576616064
	pesos_i(3044) := b"0000000000000000_0000000000000000_0001110100111100_1001010011110001"; -- 0.11420565487041778
	pesos_i(3045) := b"0000000000000000_0000000000000000_0010010001100000_0100011010010101"; -- 0.14209405083566343
	pesos_i(3046) := b"1111111111111111_1111111111111111_1110011010000111_0001001110101101"; -- -0.0995013908086887
	pesos_i(3047) := b"1111111111111111_1111111111111111_1110101101001101_0101101000100110"; -- -0.08085095006491605
	pesos_i(3048) := b"1111111111111111_1111111111111111_1101100101100111_0000001101111011"; -- -0.15077188718082496
	pesos_i(3049) := b"0000000000000000_0000000000000000_0010000111111101_0101001000110000"; -- 0.13277162246057295
	pesos_i(3050) := b"0000000000000000_0000000000000000_0001101011001110_0000001011010001"; -- 0.10470597851715135
	pesos_i(3051) := b"0000000000000000_0000000000000000_0000011000000100_0011111110100100"; -- 0.023502328414338327
	pesos_i(3052) := b"1111111111111111_1111111111111111_1101011111100011_0100100111001101"; -- -0.1566881059512423
	pesos_i(3053) := b"1111111111111111_1111111111111111_1101011010110011_0101001011111010"; -- -0.16132623108010907
	pesos_i(3054) := b"0000000000000000_0000000000000000_0001100110111000_1110110111100000"; -- 0.10047804570205411
	pesos_i(3055) := b"1111111111111111_1111111111111111_1111000000111111_0001101000111100"; -- -0.06153713264352133
	pesos_i(3056) := b"1111111111111111_1111111111111111_1110110000001000_1100001011011001"; -- -0.07799131589623125
	pesos_i(3057) := b"1111111111111111_1111111111111111_1111100100110111_0011011001110001"; -- -0.026501271560284777
	pesos_i(3058) := b"0000000000000000_0000000000000000_0001111101110010_0010010111111111"; -- 0.12283551680528748
	pesos_i(3059) := b"0000000000000000_0000000000000000_0000010100001110_0101010011110011"; -- 0.019749936394046024
	pesos_i(3060) := b"1111111111111111_1111111111111111_1111100001000010_0100001110011000"; -- -0.030238891002838032
	pesos_i(3061) := b"0000000000000000_0000000000000000_0000011100000011_1010101101111110"; -- 0.02739974818243361
	pesos_i(3062) := b"0000000000000000_0000000000000000_0001001001000100_1100011111110111"; -- 0.0713620165343526
	pesos_i(3063) := b"1111111111111111_1111111111111111_1111110100111111_0100110001111011"; -- -0.010752887660153787
	pesos_i(3064) := b"1111111111111111_1111111111111111_1111110111001101_1110111111110011"; -- -0.008576396233465816
	pesos_i(3065) := b"1111111111111111_1111111111111111_1111000111111000_1100000001010011"; -- -0.05479810700301039
	pesos_i(3066) := b"1111111111111111_1111111111111111_1111100010000100_0010000101000111"; -- -0.02923385643315877
	pesos_i(3067) := b"0000000000000000_0000000000000000_0010110000101000_0010010101100110"; -- 0.1724875807128791
	pesos_i(3068) := b"1111111111111111_1111111111111111_1101110000101111_0100000001111110"; -- -0.13990399280383115
	pesos_i(3069) := b"1111111111111111_1111111111111111_1111001110001100_0011100111011000"; -- -0.04864157168203476
	pesos_i(3070) := b"1111111111111111_1111111111111111_1111101110101000_1000010001111001"; -- -0.01695987753651389
	pesos_i(3071) := b"0000000000000000_0000000000000000_0001100100010111_1101000101011001"; -- 0.09801968024200369
	pesos_i(3072) := b"1111111111111111_1111111111111111_1101110111111100_1100110010001001"; -- -0.13286134384992682
	pesos_i(3073) := b"1111111111111111_1111111111111111_1110000101101010_1111010001010000"; -- -0.11946175625900173
	pesos_i(3074) := b"1111111111111111_1111111111111111_1111110011000111_0100101110001111"; -- -0.012583997375867226
	pesos_i(3075) := b"1111111111111111_1111111111111111_1110100100011011_1000110001000011"; -- -0.08942340254003299
	pesos_i(3076) := b"1111111111111111_1111111111111111_1101011111110001_1111000100000010"; -- -0.15646451657367066
	pesos_i(3077) := b"0000000000000000_0000000000000000_0001001111101101_1001110000000111"; -- 0.07784438286622074
	pesos_i(3078) := b"1111111111111111_1111111111111111_1111110000000111_1010011000111000"; -- -0.015508281050129373
	pesos_i(3079) := b"0000000000000000_0000000000000000_0001001000001000_1001000111100010"; -- 0.07044326565360223
	pesos_i(3080) := b"1111111111111111_1111111111111111_1111001101010101_0101010111100001"; -- -0.0494791341368818
	pesos_i(3081) := b"0000000000000000_0000000000000000_0010001010110111_0011110001111001"; -- 0.13560846295510162
	pesos_i(3082) := b"0000000000000000_0000000000000000_0001101111001000_0100001010010011"; -- 0.10852447586401993
	pesos_i(3083) := b"0000000000000000_0000000000000000_0001010100011001_0111011111000010"; -- 0.08241985774024455
	pesos_i(3084) := b"1111111111111111_1111111111111111_1101110010101101_0010011111101110"; -- -0.13798284949784695
	pesos_i(3085) := b"0000000000000000_0000000000000000_0000001111010010_1001101001101100"; -- 0.014932299971117871
	pesos_i(3086) := b"1111111111111111_1111111111111111_1111010100101110_0001001000101110"; -- -0.042265762134611265
	pesos_i(3087) := b"0000000000000000_0000000000000000_0000101111101111_0101100011011110"; -- 0.046620897436863096
	pesos_i(3088) := b"0000000000000000_0000000000000000_0000111011101001_1100000100111001"; -- 0.058254314721051886
	pesos_i(3089) := b"1111111111111111_1111111111111111_1110101110010110_1111010100000000"; -- -0.07972782857280639
	pesos_i(3090) := b"0000000000000000_0000000000000000_0001000100001101_0101001001001010"; -- 0.06660951915101887
	pesos_i(3091) := b"1111111111111111_1111111111111111_1101101000110000_0011000001011001"; -- -0.14770219637980678
	pesos_i(3092) := b"1111111111111111_1111111111111111_1110010111010101_1001100111001110"; -- -0.10220946052645928
	pesos_i(3093) := b"1111111111111111_1111111111111111_1101010111001101_0001110000011111"; -- -0.1648390220998571
	pesos_i(3094) := b"0000000000000000_0000000000000000_0000100000011101_0001100110010011"; -- 0.031694029188989954
	pesos_i(3095) := b"0000000000000000_0000000000000000_0010010011011001_1111010110000101"; -- 0.14395079144507858
	pesos_i(3096) := b"0000000000000000_0000000000000000_0000110001100100_1010011010001001"; -- 0.048410805166554605
	pesos_i(3097) := b"1111111111111111_1111111111111111_1111001010001111_1111001100110110"; -- -0.05249099671406138
	pesos_i(3098) := b"0000000000000000_0000000000000000_0000000110011010_1010011001011010"; -- 0.006266018837511673
	pesos_i(3099) := b"0000000000000000_0000000000000000_0010110000000101_0001101010000010"; -- 0.17195287388712732
	pesos_i(3100) := b"0000000000000000_0000000000000000_0010100000101000_1001010011010111"; -- 0.15686922320790997
	pesos_i(3101) := b"1111111111111111_1111111111111111_1101110010000000_1010000001010100"; -- -0.1386623186939553
	pesos_i(3102) := b"0000000000000000_0000000000000000_0000010110000010_0101111111011100"; -- 0.021520606176890677
	pesos_i(3103) := b"1111111111111111_1111111111111111_1101010010011001_0110001001101010"; -- -0.1695345392794804
	pesos_i(3104) := b"0000000000000000_0000000000000000_0001101001100110_1110011000010011"; -- 0.1031326100136569
	pesos_i(3105) := b"0000000000000000_0000000000000000_0001000010101101_0010101100000101"; -- 0.06514233458681927
	pesos_i(3106) := b"1111111111111111_1111111111111111_1101011011010100_1101010000011010"; -- -0.16081499445767808
	pesos_i(3107) := b"1111111111111111_1111111111111111_1111010101110010_0111111001000100"; -- -0.04122172205001494
	pesos_i(3108) := b"0000000000000000_0000000000000000_0000001100010000_1000110000110110"; -- 0.011971247876272706
	pesos_i(3109) := b"0000000000000000_0000000000000000_0010001110100111_0100111011000011"; -- 0.1392716623240406
	pesos_i(3110) := b"0000000000000000_0000000000000000_0000100000001011_1001011011000111"; -- 0.031426833712912654
	pesos_i(3111) := b"1111111111111111_1111111111111111_1110011101100010_0110010001011101"; -- -0.09615490649506382
	pesos_i(3112) := b"0000000000000000_0000000000000000_0000111101110100_0001010011111011"; -- 0.06036502015230852
	pesos_i(3113) := b"0000000000000000_0000000000000000_0001110111101010_1110100010000101"; -- 0.116865665892067
	pesos_i(3114) := b"0000000000000000_0000000000000000_0001100001011101_1100001110000001"; -- 0.09518072022021568
	pesos_i(3115) := b"1111111111111111_1111111111111111_1101110011101111_0010001101010010"; -- -0.13697604420977322
	pesos_i(3116) := b"0000000000000000_0000000000000000_0001011000101110_1111110010100110"; -- 0.08665446321297887
	pesos_i(3117) := b"0000000000000000_0000000000000000_0001000110001101_0000001011001000"; -- 0.06855790514772825
	pesos_i(3118) := b"0000000000000000_0000000000000000_0001111101100000_1001010110010100"; -- 0.12256750919424511
	pesos_i(3119) := b"1111111111111111_1111111111111111_1101110000001101_1111001000010000"; -- -0.14041220780481287
	pesos_i(3120) := b"0000000000000000_0000000000000000_0000000100011110_0010011100011001"; -- 0.004366343984214122
	pesos_i(3121) := b"0000000000000000_0000000000000000_0010101110001110_1001011010100100"; -- 0.17014447701741964
	pesos_i(3122) := b"1111111111111111_1111111111111111_1110011100010010_1110000001110001"; -- -0.09736821394592443
	pesos_i(3123) := b"0000000000000000_0000000000000000_0001000100101001_1110101111100011"; -- 0.06704592028847733
	pesos_i(3124) := b"0000000000000000_0000000000000000_0001110101101011_1001001111010001"; -- 0.11492275096082606
	pesos_i(3125) := b"1111111111111111_1111111111111111_1110001001100101_0011100000100000"; -- -0.11564301705947444
	pesos_i(3126) := b"1111111111111111_1111111111111111_1101010110001000_0110001100100101"; -- -0.16588764526997404
	pesos_i(3127) := b"0000000000000000_0000000000000000_0000100011001101_1110110110011000"; -- 0.03439221339485256
	pesos_i(3128) := b"0000000000000000_0000000000000000_0001011000101101_1110001010001100"; -- 0.08663764877390709
	pesos_i(3129) := b"0000000000000000_0000000000000000_0001010011001111_1110011100011000"; -- 0.08129734353684662
	pesos_i(3130) := b"1111111111111111_1111111111111111_1110101000010101_0101100111010011"; -- -0.08561171146391815
	pesos_i(3131) := b"1111111111111111_1111111111111111_1110000010111010_1100100001100000"; -- -0.12214992188567152
	pesos_i(3132) := b"1111111111111111_1111111111111111_1110101000011100_1111011011110111"; -- -0.08549553359779248
	pesos_i(3133) := b"1111111111111111_1111111111111111_1110010101101111_0010000111101101"; -- -0.10377300217867974
	pesos_i(3134) := b"1111111111111111_1111111111111111_1111001100010000_1100110001001010"; -- -0.05052493287229749
	pesos_i(3135) := b"1111111111111111_1111111111111111_1110111000000000_0010001000001001"; -- -0.07031047123179396
	pesos_i(3136) := b"1111111111111111_1111111111111111_1101100101101111_1101101010100111"; -- -0.1506369916129833
	pesos_i(3137) := b"1111111111111111_1111111111111111_1111100001101100_1110110100010010"; -- -0.029587920336840746
	pesos_i(3138) := b"1111111111111111_1111111111111111_1101111011100010_0011010111001001"; -- -0.12936080787836346
	pesos_i(3139) := b"0000000000000000_0000000000000000_0010011001000011_0110010011111000"; -- 0.14946585718090316
	pesos_i(3140) := b"1111111111111111_1111111111111111_1110101101011100_0100110000010110"; -- -0.08062290628303156
	pesos_i(3141) := b"1111111111111111_1111111111111111_1110101010011011_0110000101111101"; -- -0.0835665769724423
	pesos_i(3142) := b"0000000000000000_0000000000000000_0001001110000101_0010001110010000"; -- 0.07625028870051141
	pesos_i(3143) := b"1111111111111111_1111111111111111_1101101000100111_1010100010011001"; -- -0.1478323579096264
	pesos_i(3144) := b"0000000000000000_0000000000000000_0000110111001011_0100001111101000"; -- 0.0538828318157127
	pesos_i(3145) := b"0000000000000000_0000000000000000_0000110101101110_0000001000111100"; -- 0.05245985007578849
	pesos_i(3146) := b"0000000000000000_0000000000000000_0001000100111001_0110110010001111"; -- 0.0672824716364495
	pesos_i(3147) := b"0000000000000000_0000000000000000_0010001100010010_1001001001001001"; -- 0.1370021273645306
	pesos_i(3148) := b"1111111111111111_1111111111111111_1110001000000100_1001100001110111"; -- -0.11711737711744642
	pesos_i(3149) := b"0000000000000000_0000000000000000_0000110011111101_0011000101100100"; -- 0.05073841744355387
	pesos_i(3150) := b"1111111111111111_1111111111111111_1101110111101010_1101101000101000"; -- -0.13313519013370342
	pesos_i(3151) := b"1111111111111111_1111111111111111_1110100111010101_1000111000001001"; -- -0.08658516204966019
	pesos_i(3152) := b"1111111111111111_1111111111111111_1101011111000000_0110010000100100"; -- -0.1572205936676747
	pesos_i(3153) := b"1111111111111111_1111111111111111_1111001101011001_0011011001110001"; -- -0.04941997270140066
	pesos_i(3154) := b"0000000000000000_0000000000000000_0000000011101100_1101110001010111"; -- 0.0036142074924667604
	pesos_i(3155) := b"1111111111111111_1111111111111111_1110001011010100_0010111010110101"; -- -0.11394985280168278
	pesos_i(3156) := b"1111111111111111_1111111111111111_1101100101110000_1100110010000101"; -- -0.15062257542369165
	pesos_i(3157) := b"0000000000000000_0000000000000000_0000011001100111_1010011010110110"; -- 0.025019091984405953
	pesos_i(3158) := b"0000000000000000_0000000000000000_0010001101011111_0110001001001010"; -- 0.1381741934341831
	pesos_i(3159) := b"0000000000000000_0000000000000000_0000110001010111_1100011111001001"; -- 0.04821442287535075
	pesos_i(3160) := b"0000000000000000_0000000000000000_0000000000000100_1001101000111101"; -- 7.02284929738426e-05
	pesos_i(3161) := b"0000000000000000_0000000000000000_0000010111010010_1001011110000110"; -- 0.02274462727572193
	pesos_i(3162) := b"0000000000000000_0000000000000000_0010011111000110_1011000110001100"; -- 0.15537557275082528
	pesos_i(3163) := b"0000000000000000_0000000000000000_0000100011110011_0110100010010000"; -- 0.034964118235868175
	pesos_i(3164) := b"1111111111111111_1111111111111111_1111010010110001_1010100010011010"; -- -0.04416414483764398
	pesos_i(3165) := b"1111111111111111_1111111111111111_1101111010011110_1101000101011110"; -- -0.13038913200015675
	pesos_i(3166) := b"1111111111111111_1111111111111111_1101110011000101_0001001110101000"; -- -0.13761784690491763
	pesos_i(3167) := b"1111111111111111_1111111111111111_1111110010010011_0001101000001010"; -- -0.01338040602941079
	pesos_i(3168) := b"0000000000000000_0000000000000000_0001001001000001_1101010001100001"; -- 0.07131698011650611
	pesos_i(3169) := b"1111111111111111_1111111111111111_1110000110100101_0101110000110110"; -- -0.11857055369602358
	pesos_i(3170) := b"1111111111111111_1111111111111111_1111100110101010_0110000100100101"; -- -0.024743965496233335
	pesos_i(3171) := b"1111111111111111_1111111111111111_1110101001000110_1111110001000010"; -- -0.08485434906100461
	pesos_i(3172) := b"1111111111111111_1111111111111111_1111010111110101_0101010111011111"; -- -0.03922522842507899
	pesos_i(3173) := b"0000000000000000_0000000000000000_0000011001100011_0101110101011110"; -- 0.024953685299908216
	pesos_i(3174) := b"0000000000000000_0000000000000000_0001010001110100_0101010100000000"; -- 0.07990008597229874
	pesos_i(3175) := b"0000000000000000_0000000000000000_0000010011000100_0111110001101111"; -- 0.01862313946430441
	pesos_i(3176) := b"0000000000000000_0000000000000000_0010100110010010_1011001001010000"; -- 0.16239466136070127
	pesos_i(3177) := b"0000000000000000_0000000000000000_0001010001101100_0100111011111111"; -- 0.07977765782418733
	pesos_i(3178) := b"1111111111111111_1111111111111111_1110101010000111_0010001000000100"; -- -0.08387553594687566
	pesos_i(3179) := b"0000000000000000_0000000000000000_0001110001010111_0111110010010100"; -- 0.11070994007992307
	pesos_i(3180) := b"1111111111111111_1111111111111111_1110000000010000_1000101011010110"; -- -0.12474758417374747
	pesos_i(3181) := b"1111111111111111_1111111111111111_1110000100000111_0110111110100000"; -- -0.12098028512774184
	pesos_i(3182) := b"0000000000000000_0000000000000000_0001001110111010_0011100100000101"; -- 0.0770602833009957
	pesos_i(3183) := b"0000000000000000_0000000000000000_0001010000100001_0110001000011010"; -- 0.07863438728102898
	pesos_i(3184) := b"1111111111111111_1111111111111111_1111010110001100_1111111011000000"; -- -0.040817335259899695
	pesos_i(3185) := b"0000000000000000_0000000000000000_0010001010001101_1100111100010001"; -- 0.13497633147017885
	pesos_i(3186) := b"0000000000000000_0000000000000000_0000010010101010_0000010001001111"; -- 0.01821925103778363
	pesos_i(3187) := b"1111111111111111_1111111111111111_1110010001101011_0011001101010000"; -- -0.10773925101270568
	pesos_i(3188) := b"0000000000000000_0000000000000000_0010100000100010_1010100100111100"; -- 0.15677888603698623
	pesos_i(3189) := b"0000000000000000_0000000000000000_0000101101000011_0101100100101000"; -- 0.043996402930667054
	pesos_i(3190) := b"0000000000000000_0000000000000000_0001111101001001_1110011000011011"; -- 0.12222135690329362
	pesos_i(3191) := b"1111111111111111_1111111111111111_1101101011001001_0001101110001000"; -- -0.14536884233481795
	pesos_i(3192) := b"1111111111111111_1111111111111111_1111000000110101_0100110100010101"; -- -0.06168668962324715
	pesos_i(3193) := b"1111111111111111_1111111111111111_1101110111110100_1111111000101010"; -- -0.13298045622627933
	pesos_i(3194) := b"1111111111111111_1111111111111111_1110111100011000_1010110111010001"; -- -0.0660296787650842
	pesos_i(3195) := b"0000000000000000_0000000000000000_0001000011111101_0101100011010001"; -- 0.0663657674007142
	pesos_i(3196) := b"0000000000000000_0000000000000000_0010100011000001_1000100100001001"; -- 0.15920311414074714
	pesos_i(3197) := b"1111111111111111_1111111111111111_1110010100011111_1000011110010101"; -- -0.10498764615425649
	pesos_i(3198) := b"0000000000000000_0000000000000000_0001100000100111_0100011010101011"; -- 0.09434930486899294
	pesos_i(3199) := b"0000000000000000_0000000000000000_0000010101001001_1111110010010101"; -- 0.020660196647171957
	pesos_i(3200) := b"0000000000000000_0000000000000000_0010101001001111_1000101000011000"; -- 0.16527617543404824
	pesos_i(3201) := b"0000000000000000_0000000000000000_0000101000111111_1001011001101001"; -- 0.04003276894715709
	pesos_i(3202) := b"0000000000000000_0000000000000000_0010010101110011_1000101010010001"; -- 0.14629427004950848
	pesos_i(3203) := b"1111111111111111_1111111111111111_1101111101000000_1100100000001101"; -- -0.12791776357224252
	pesos_i(3204) := b"0000000000000000_0000000000000000_0001100010110101_1010000101110000"; -- 0.09652146322602406
	pesos_i(3205) := b"1111111111111111_1111111111111111_1111101111100111_0110110011111110"; -- -0.015999973232773263
	pesos_i(3206) := b"0000000000000000_0000000000000000_0000100000010110_1011011111111111"; -- 0.031596660486877495
	pesos_i(3207) := b"1111111111111111_1111111111111111_1110001010000011_1001001000110000"; -- -0.1151798852251048
	pesos_i(3208) := b"1111111111111111_1111111111111111_1111101100011000_0111100111111010"; -- -0.019157768641790304
	pesos_i(3209) := b"1111111111111111_1111111111111111_1110011011001000_1101001010011010"; -- -0.09849818936444239
	pesos_i(3210) := b"0000000000000000_0000000000000000_0010101001111001_0111110101000101"; -- 0.16591628015296195
	pesos_i(3211) := b"0000000000000000_0000000000000000_0000110101010011_1010100111100111"; -- 0.052057856522832555
	pesos_i(3212) := b"1111111111111111_1111111111111111_1110110111100010_1000001000000111"; -- -0.07076251339548327
	pesos_i(3213) := b"1111111111111111_1111111111111111_1110011101001000_0100101011001011"; -- -0.09655315916376148
	pesos_i(3214) := b"1111111111111111_1111111111111111_1101101011110001_1000000001011101"; -- -0.14475248074398514
	pesos_i(3215) := b"0000000000000000_0000000000000000_0010001001000011_1101110011101110"; -- 0.13384800736633398
	pesos_i(3216) := b"1111111111111111_1111111111111111_1101011010111001_1101011101110100"; -- -0.1612267820528988
	pesos_i(3217) := b"1111111111111111_1111111111111111_1110100100100010_1011011100101001"; -- -0.0893140338594438
	pesos_i(3218) := b"0000000000000000_0000000000000000_0010110000011111_0100000111111000"; -- 0.17235195457685304
	pesos_i(3219) := b"1111111111111111_1111111111111111_1101100010010101_0100000011001011"; -- -0.15397257843724935
	pesos_i(3220) := b"0000000000000000_0000000000000000_0000011000101000_1011000111100011"; -- 0.0240584543711764
	pesos_i(3221) := b"0000000000000000_0000000000000000_0010001001001110_1100000000010100"; -- 0.1340141342365671
	pesos_i(3222) := b"1111111111111111_1111111111111111_1100111011111011_0000100001100011"; -- -0.19148204412619868
	pesos_i(3223) := b"1111111111111111_1111111111111111_1110111110011010_1011110100101011"; -- -0.06404512118783283
	pesos_i(3224) := b"1111111111111111_1111111111111111_1111100111010000_1110100110101001"; -- -0.024155994575022943
	pesos_i(3225) := b"0000000000000000_0000000000000000_0000000001110001_0000111001000110"; -- 0.0017250939296529805
	pesos_i(3226) := b"1111111111111111_1111111111111111_1111000110001111_1011000100111000"; -- -0.05640118021069393
	pesos_i(3227) := b"0000000000000000_0000000000000000_0010101101001010_1011111111011011"; -- 0.1691093357869754
	pesos_i(3228) := b"0000000000000000_0000000000000000_0001011110011010_1011010011111100"; -- 0.0922043909091568
	pesos_i(3229) := b"0000000000000000_0000000000000000_0001011010111010_0011110110001111"; -- 0.08877930401045782
	pesos_i(3230) := b"1111111111111111_1111111111111111_1110000100001110_1110011010111010"; -- -0.12086637464322308
	pesos_i(3231) := b"0000000000000000_0000000000000000_0001101011011001_0111010111110111"; -- 0.10488068838249784
	pesos_i(3232) := b"0000000000000000_0000000000000000_0010011111100100_0101010101101000"; -- 0.15582784448790862
	pesos_i(3233) := b"1111111111111111_1111111111111111_1101011000100100_0101010101001100"; -- -0.16350809940101776
	pesos_i(3234) := b"0000000000000000_0000000000000000_0000111111110111_1110101001010000"; -- 0.06237663708118535
	pesos_i(3235) := b"1111111111111111_1111111111111111_1110011001110110_0010011100000010"; -- -0.0997596379205973
	pesos_i(3236) := b"1111111111111111_1111111111111111_1110111010100011_1101100011001111"; -- -0.06781239461465831
	pesos_i(3237) := b"0000000000000000_0000000000000000_0010011100011100_1100110101101101"; -- 0.15278324042649385
	pesos_i(3238) := b"1111111111111111_1111111111111111_1110110001100101_1001000001110010"; -- -0.07657525269146545
	pesos_i(3239) := b"1111111111111111_1111111111111111_1110100111001010_0110101101011111"; -- -0.08675507483607382
	pesos_i(3240) := b"1111111111111111_1111111111111111_1111001001101101_0010100010100001"; -- -0.053021870384515044
	pesos_i(3241) := b"1111111111111111_1111111111111111_1111011000111000_1100010100110101"; -- -0.03819625340433387
	pesos_i(3242) := b"1111111111111111_1111111111111111_1111110000000000_1110000000011101"; -- -0.01561164182756953
	pesos_i(3243) := b"0000000000000000_0000000000000000_0000001001110101_0000100010100110"; -- 0.009598293698557662
	pesos_i(3244) := b"0000000000000000_0000000000000000_0000110001010011_0101001101100010"; -- 0.0481464494527638
	pesos_i(3245) := b"1111111111111111_1111111111111111_1101100010110011_1001111010001101"; -- -0.15350922637010128
	pesos_i(3246) := b"1111111111111111_1111111111111111_1111011001101010_1101110001000010"; -- -0.037431939964416405
	pesos_i(3247) := b"0000000000000000_0000000000000000_0001011111011001_1111111111011010"; -- 0.09317015708531506
	pesos_i(3248) := b"0000000000000000_0000000000000000_0000010100100110_0101101011011111"; -- 0.020116500278951344
	pesos_i(3249) := b"1111111111111111_1111111111111111_1101110110000111_0100001100111010"; -- -0.13465480635177507
	pesos_i(3250) := b"1111111111111111_1111111111111111_1111101010011001_0111111111010011"; -- -0.021095286465270688
	pesos_i(3251) := b"1111111111111111_1111111111111111_1110000111000111_0000010011101111"; -- -0.11805695698517635
	pesos_i(3252) := b"0000000000000000_0000000000000000_0001001100111010_1011100110010111"; -- 0.07511482187174778
	pesos_i(3253) := b"1111111111111111_1111111111111111_1111111110011000_0000000000110011"; -- -0.0015869022698759155
	pesos_i(3254) := b"0000000000000000_0000000000000000_0000011110101010_0100010000001111"; -- 0.029941800723873153
	pesos_i(3255) := b"1111111111111111_1111111111111111_1111001010000100_0010000000001001"; -- -0.05267143039587606
	pesos_i(3256) := b"0000000000000000_0000000000000000_0000010000011010_0000101110000110"; -- 0.01602241544839439
	pesos_i(3257) := b"1111111111111111_1111111111111111_1110100001010101_1010100111100011"; -- -0.09244287696207643
	pesos_i(3258) := b"0000000000000000_0000000000000000_0001110101110000_1100110010100110"; -- 0.11500243248393448
	pesos_i(3259) := b"0000000000000000_0000000000000000_0010010001011100_1001000100001111"; -- 0.1420374547625796
	pesos_i(3260) := b"0000000000000000_0000000000000000_0001011010111010_1101001001010000"; -- 0.08878817034645399
	pesos_i(3261) := b"0000000000000000_0000000000000000_0010011000101011_0111010000011001"; -- 0.1491005478400922
	pesos_i(3262) := b"0000000000000000_0000000000000000_0010110101000111_1110101110111111"; -- 0.17687867562748055
	pesos_i(3263) := b"1111111111111111_1111111111111111_1110000001111011_1100001100011111"; -- -0.12311153881178966
	pesos_i(3264) := b"0000000000000000_0000000000000000_0000000111110101_0110011010010101"; -- 0.007650767773648509
	pesos_i(3265) := b"1111111111111111_1111111111111111_1101011010101010_1111100001100000"; -- -0.16145370166862194
	pesos_i(3266) := b"1111111111111111_1111111111111111_1101001011011111_1011000101000100"; -- -0.1762742242518934
	pesos_i(3267) := b"0000000000000000_0000000000000000_0001001110110010_1110100011101001"; -- 0.07694869706523547
	pesos_i(3268) := b"0000000000000000_0000000000000000_0010011101000010_0100010001100000"; -- 0.15335490560064993
	pesos_i(3269) := b"0000000000000000_0000000000000000_0000100000100010_1100100000110101"; -- 0.03178073206519929
	pesos_i(3270) := b"0000000000000000_0000000000000000_0010000101011011_0010010110110111"; -- 0.13029704781408444
	pesos_i(3271) := b"1111111111111111_1111111111111111_1111011011011011_1100111101100001"; -- -0.03570846439384947
	pesos_i(3272) := b"0000000000000000_0000000000000000_0001101101100110_1110010001010011"; -- 0.10703875571588128
	pesos_i(3273) := b"0000000000000000_0000000000000000_0010000101001110_1011111101010111"; -- 0.13010784036329673
	pesos_i(3274) := b"0000000000000000_0000000000000000_0001101100101011_0010100101010010"; -- 0.1061273408590425
	pesos_i(3275) := b"0000000000000000_0000000000000000_0000001000010001_1100010000011101"; -- 0.008083588728472738
	pesos_i(3276) := b"0000000000000000_0000000000000000_0000000000010100_0101001110111001"; -- 0.00031016613627802875
	pesos_i(3277) := b"1111111111111111_1111111111111111_1111000111111111_0001001011010001"; -- -0.05470163735178332
	pesos_i(3278) := b"1111111111111111_1111111111111111_1110000111010111_1111101111111100"; -- -0.11779809094557636
	pesos_i(3279) := b"0000000000000000_0000000000000000_0001000001110100_1111110011010100"; -- 0.06428508917435374
	pesos_i(3280) := b"0000000000000000_0000000000000000_0001101010111111_0111101101011011"; -- 0.10448428120356132
	pesos_i(3281) := b"0000000000000000_0000000000000000_0010001101110101_0111101111010010"; -- 0.1385114086063874
	pesos_i(3282) := b"1111111111111111_1111111111111111_1101111011111101_0000110111110001"; -- -0.12895119541258127
	pesos_i(3283) := b"1111111111111111_1111111111111111_1110110111001111_1100101010000110"; -- -0.07104810939451077
	pesos_i(3284) := b"0000000000000000_0000000000000000_0010001011011110_0111101001001011"; -- 0.13620724030435954
	pesos_i(3285) := b"1111111111111111_1111111111111111_1110001000100010_0010001110001101"; -- -0.11666658229276458
	pesos_i(3286) := b"1111111111111111_1111111111111111_1111101001001111_0100000010101100"; -- -0.022228200857824523
	pesos_i(3287) := b"0000000000000000_0000000000000000_0000011010001001_1100111010000011"; -- 0.025540263059523515
	pesos_i(3288) := b"0000000000000000_0000000000000000_0000110010111001_0111100101011011"; -- 0.0497051093092324
	pesos_i(3289) := b"1111111111111111_1111111111111111_1110001100111010_1010001110000011"; -- -0.11238649415610605
	pesos_i(3290) := b"0000000000000000_0000000000000000_0001010100010001_1100000010100111"; -- 0.08230213229865793
	pesos_i(3291) := b"0000000000000000_0000000000000000_0001010010010110_1000100000100101"; -- 0.08042193310791267
	pesos_i(3292) := b"0000000000000000_0000000000000000_0001110110011001_1101111100011110"; -- 0.11562914352533167
	pesos_i(3293) := b"1111111111111111_1111111111111111_1111100111100001_1010101011111010"; -- -0.023900331532692578
	pesos_i(3294) := b"1111111111111111_1111111111111111_1110000001011000_0011000101000101"; -- -0.12365428976305093
	pesos_i(3295) := b"1111111111111111_1111111111111111_1111000010111001_1010001010111101"; -- -0.0596674239965161
	pesos_i(3296) := b"0000000000000000_0000000000000000_0000110001111111_0000110010001110"; -- 0.04881361456017316
	pesos_i(3297) := b"1111111111111111_1111111111111111_1110101111000100_0100110000011100"; -- -0.07903599080722941
	pesos_i(3298) := b"0000000000000000_0000000000000000_0000110111110111_1010100111110100"; -- 0.05456030086140196
	pesos_i(3299) := b"1111111111111111_1111111111111111_1111110110011100_0010100100111010"; -- -0.009335921677759785
	pesos_i(3300) := b"1111111111111111_1111111111111111_1111000001010111_1111000100111001"; -- -0.0611581073264527
	pesos_i(3301) := b"1111111111111111_1111111111111111_1101100100001011_0111001101110000"; -- -0.1521690228202402
	pesos_i(3302) := b"0000000000000000_0000000000000000_0001000010010111_1011010101100000"; -- 0.06481488798668289
	pesos_i(3303) := b"0000000000000000_0000000000000000_0000100100110001_1011111001111001"; -- 0.035915283803222925
	pesos_i(3304) := b"0000000000000000_0000000000000000_0010100111111011_1100100001001101"; -- 0.16399814491897105
	pesos_i(3305) := b"1111111111111111_1111111111111111_1101111111001111_0001000000011100"; -- -0.12574672044756258
	pesos_i(3306) := b"1111111111111111_1111111111111111_1111000111001001_0001101011000110"; -- -0.05552513761118263
	pesos_i(3307) := b"0000000000000000_0000000000000000_0010101111111000_1110101110001110"; -- 0.17176696980578557
	pesos_i(3308) := b"0000000000000000_0000000000000000_0001110101111100_0111000101101100"; -- 0.1151801003151782
	pesos_i(3309) := b"0000000000000000_0000000000000000_0010001010010111_1101010001111101"; -- 0.13512924246194696
	pesos_i(3310) := b"1111111111111111_1111111111111111_1111001110100000_1010011010111110"; -- -0.04832990522321448
	pesos_i(3311) := b"0000000000000000_0000000000000000_0000000000011110_0101000000011111"; -- 0.00046253934913575284
	pesos_i(3312) := b"1111111111111111_1111111111111111_1101011100100111_0101111101110001"; -- -0.15955546856952904
	pesos_i(3313) := b"1111111111111111_1111111111111111_1110101110100111_0001100100001000"; -- -0.07948154022994751
	pesos_i(3314) := b"1111111111111111_1111111111111111_1111001110111011_1100111000001111"; -- -0.04791557450281724
	pesos_i(3315) := b"0000000000000000_0000000000000000_0001110111110110_1011001101111111"; -- 0.1170456109688631
	pesos_i(3316) := b"0000000000000000_0000000000000000_0010100000011010_1100000100010110"; -- 0.15665823728534173
	pesos_i(3317) := b"0000000000000000_0000000000000000_0000011000110010_1100011111000011"; -- 0.024212346088845482
	pesos_i(3318) := b"0000000000000000_0000000000000000_0001011111101111_1110110000000011"; -- 0.09350466806914116
	pesos_i(3319) := b"1111111111111111_1111111111111111_1110011101111100_1100010010100001"; -- -0.09575244016992954
	pesos_i(3320) := b"1111111111111111_1111111111111111_1101110111000101_1000011011011111"; -- -0.13370472962462532
	pesos_i(3321) := b"1111111111111111_1111111111111111_1110110011100001_0001011010100001"; -- -0.07469042368831129
	pesos_i(3322) := b"1111111111111111_1111111111111111_1101100010110111_1111000000011111"; -- -0.15344332933646446
	pesos_i(3323) := b"1111111111111111_1111111111111111_1101001001011011_1010110100111011"; -- -0.17828862488149677
	pesos_i(3324) := b"0000000000000000_0000000000000000_0000011110110101_0100011111000001"; -- 0.03010986778416947
	pesos_i(3325) := b"1111111111111111_1111111111111111_1110001110000101_0111100010111001"; -- -0.11124463538782257
	pesos_i(3326) := b"1111111111111111_1111111111111111_1110110101010011_0111110010111111"; -- -0.07294483511609871
	pesos_i(3327) := b"1111111111111111_1111111111111111_1110010110011010_0100000001110100"; -- -0.10311505468679613
	pesos_i(3328) := b"0000000000000000_0000000000000000_0000111101100111_1100010110100011"; -- 0.06017718527644467
	pesos_i(3329) := b"0000000000000000_0000000000000000_0010000101001100_1100100011111001"; -- 0.1300778968622303
	pesos_i(3330) := b"0000000000000000_0000000000000000_0001010010111010_1011101101111100"; -- 0.08097430971326895
	pesos_i(3331) := b"1111111111111111_1111111111111111_1101010101100000_0101010000010110"; -- -0.16649889442002025
	pesos_i(3332) := b"0000000000000000_0000000000000000_0000100010001100_0011000001110001"; -- 0.03338911779352271
	pesos_i(3333) := b"1111111111111111_1111111111111111_1110011011001011_1101111111100100"; -- -0.09845162098829725
	pesos_i(3334) := b"0000000000000000_0000000000000000_0001010100100000_1100000011000100"; -- 0.08253102095417007
	pesos_i(3335) := b"0000000000000000_0000000000000000_0010100011000110_1001110000100000"; -- 0.159280546068907
	pesos_i(3336) := b"1111111111111111_1111111111111111_1111100111111111_1000011111101110"; -- -0.02344465682937466
	pesos_i(3337) := b"1111111111111111_1111111111111111_1110000001011100_0011000101100001"; -- -0.12359324819703105
	pesos_i(3338) := b"0000000000000000_0000000000000000_0010011101110000_1011000011010100"; -- 0.15406327408687365
	pesos_i(3339) := b"1111111111111111_1111111111111111_1101010101011101_1100011010100010"; -- -0.16653784327957752
	pesos_i(3340) := b"0000000000000000_0000000000000000_0001000011010011_1101000011101100"; -- 0.06573205717576383
	pesos_i(3341) := b"1111111111111111_1111111111111111_1101101110101101_1111000010001110"; -- -0.1418771414193581
	pesos_i(3342) := b"1111111111111111_1111111111111111_1111100100001111_0100011001010110"; -- -0.027110675746093688
	pesos_i(3343) := b"0000000000000000_0000000000000000_0001000110000000_0000110011110100"; -- 0.06836014702080798
	pesos_i(3344) := b"1111111111111111_1111111111111111_1111001000100001_1011110000110101"; -- -0.054172741970378774
	pesos_i(3345) := b"0000000000000000_0000000000000000_0010101001011100_0101011111010000"; -- 0.1654715427213548
	pesos_i(3346) := b"1111111111111111_1111111111111111_1111101111001001_0101001011001001"; -- -0.016459299036383487
	pesos_i(3347) := b"1111111111111111_1111111111111111_1101110010001110_0011110111101011"; -- -0.138454561294941
	pesos_i(3348) := b"1111111111111111_1111111111111111_1111101110101001_0110010110001000"; -- -0.016946462851172312
	pesos_i(3349) := b"1111111111111111_1111111111111111_1110100001010111_1101110111111011"; -- -0.09240925439428387
	pesos_i(3350) := b"0000000000000000_0000000000000000_0001000000001010_1100011100000000"; -- 0.06266444922209986
	pesos_i(3351) := b"1111111111111111_1111111111111111_1110011011110000_1101100111010011"; -- -0.09788740730833312
	pesos_i(3352) := b"1111111111111111_1111111111111111_1100110111000000_0010011000111100"; -- -0.19628678346430575
	pesos_i(3353) := b"0000000000000000_0000000000000000_0000101110101000_1110111101011111"; -- 0.045546494205655756
	pesos_i(3354) := b"0000000000000000_0000000000000000_0001000001100000_1001000011110011"; -- 0.06397348335689186
	pesos_i(3355) := b"0000000000000000_0000000000000000_0010110001100111_0111000000001010"; -- 0.1734533332203408
	pesos_i(3356) := b"0000000000000000_0000000000000000_0001011010000001_0101100111001011"; -- 0.08791123590214082
	pesos_i(3357) := b"0000000000000000_0000000000000000_0000011110111000_0111000101100001"; -- 0.030158125073422807
	pesos_i(3358) := b"1111111111111111_1111111111111111_1111010010001100_0100011001101011"; -- -0.04473457240088617
	pesos_i(3359) := b"1111111111111111_1111111111111111_1101101101000001_1100011000010100"; -- -0.1435276222418898
	pesos_i(3360) := b"0000000000000000_0000000000000000_0000111111010101_0001110110000011"; -- 0.06184563101285975
	pesos_i(3361) := b"0000000000000000_0000000000000000_0010000101010001_0011100111000111"; -- 0.13014565573843834
	pesos_i(3362) := b"0000000000000000_0000000000000000_0010010000011010_1011110000010101"; -- 0.14103293913921114
	pesos_i(3363) := b"0000000000000000_0000000000000000_0001110100010000_0110110000001111"; -- 0.11353183136622165
	pesos_i(3364) := b"1111111111111111_1111111111111111_1101101111001100_1101100110010011"; -- -0.14140548850693568
	pesos_i(3365) := b"1111111111111111_1111111111111111_1111110011010010_1101000111100100"; -- -0.012408143940235265
	pesos_i(3366) := b"1111111111111111_1111111111111111_1101011000111000_0011100111011111"; -- -0.1632045584273981
	pesos_i(3367) := b"0000000000000000_0000000000000000_0000001010111111_0010010100000101"; -- 0.010729135356616737
	pesos_i(3368) := b"0000000000000000_0000000000000000_0000001111100010_1111010111011100"; -- 0.015181890702161
	pesos_i(3369) := b"0000000000000000_0000000000000000_0010001100101111_1000110001001111"; -- 0.13744427609136706
	pesos_i(3370) := b"1111111111111111_1111111111111111_1111010000101011_0111100010100000"; -- -0.04621168229277903
	pesos_i(3371) := b"0000000000000000_0000000000000000_0000100011000110_0100000111101111"; -- 0.034275170263169695
	pesos_i(3372) := b"1111111111111111_1111111111111111_1101110000111111_1011100110011010"; -- -0.13965263365428604
	pesos_i(3373) := b"1111111111111111_1111111111111111_1110100010100010_0010010100111100"; -- -0.09127585675164501
	pesos_i(3374) := b"0000000000000000_0000000000000000_0000101111001000_0000000010010001"; -- 0.04602054147898547
	pesos_i(3375) := b"0000000000000000_0000000000000000_0000010111010010_0110110011101101"; -- 0.022742088198762826
	pesos_i(3376) := b"1111111111111111_1111111111111111_1111110000100111_1001100010110011"; -- -0.01502080562696878
	pesos_i(3377) := b"1111111111111111_1111111111111111_1111100001000111_1101001001000001"; -- -0.030154093807827152
	pesos_i(3378) := b"0000000000000000_0000000000000000_0001011011111110_1010101011101110"; -- 0.0898234205304048
	pesos_i(3379) := b"1111111111111111_1111111111111111_1101110001110110_1110001010101101"; -- -0.13881095201014768
	pesos_i(3380) := b"1111111111111111_1111111111111111_1101111111000110_1110110000101001"; -- -0.12587093354443257
	pesos_i(3381) := b"1111111111111111_1111111111111111_1111011001100111_0001011001101111"; -- -0.037489507590944986
	pesos_i(3382) := b"1111111111111111_1111111111111111_1110111011101100_1110111001011010"; -- -0.0666972189313316
	pesos_i(3383) := b"1111111111111111_1111111111111111_1110110011111011_1011111011010000"; -- -0.07428367068451244
	pesos_i(3384) := b"0000000000000000_0000000000000000_0001110001101011_1000011111111011"; -- 0.11101579544515691
	pesos_i(3385) := b"1111111111111111_1111111111111111_1110011101000010_1111110001011010"; -- -0.09663412859597362
	pesos_i(3386) := b"1111111111111111_1111111111111111_1110101100110010_1111101110101011"; -- -0.08125331005641875
	pesos_i(3387) := b"1111111111111111_1111111111111111_1110101001101000_1101101101101100"; -- -0.08433750727592387
	pesos_i(3388) := b"1111111111111111_1111111111111111_1111001010101101_1110010111010101"; -- -0.052034030394833695
	pesos_i(3389) := b"1111111111111111_1111111111111111_1110011000110010_1000111111001010"; -- -0.10079098993624011
	pesos_i(3390) := b"0000000000000000_0000000000000000_0000110000010110_1111010000100011"; -- 0.04722524512355132
	pesos_i(3391) := b"0000000000000000_0000000000000000_0000010111001110_1100100100001101"; -- 0.022686544160883747
	pesos_i(3392) := b"0000000000000000_0000000000000000_0000111001010001_1110101011000110"; -- 0.05593745551644566
	pesos_i(3393) := b"1111111111111111_1111111111111111_1110011011001010_1110000011001101"; -- -0.09846682540503796
	pesos_i(3394) := b"1111111111111111_1111111111111111_1110111001111010_1101111011110011"; -- -0.06843763898063593
	pesos_i(3395) := b"0000000000000000_0000000000000000_0010111011101001_0111011010111111"; -- 0.18324987573678664
	pesos_i(3396) := b"0000000000000000_0000000000000000_0000101111001000_0000110000001011"; -- 0.04602122567816621
	pesos_i(3397) := b"0000000000000000_0000000000000000_0010001111010110_0000010001100001"; -- 0.1399843918570705
	pesos_i(3398) := b"1111111111111111_1111111111111111_1111010110001011_1000010100111010"; -- -0.04083983743916889
	pesos_i(3399) := b"0000000000000000_0000000000000000_0001011001100011_0100000000000010"; -- 0.08745193519996862
	pesos_i(3400) := b"0000000000000000_0000000000000000_0010000000011110_1010111000011111"; -- 0.12546814200722517
	pesos_i(3401) := b"1111111111111111_1111111111111111_1101100011010111_0110110010110100"; -- -0.15296288104148736
	pesos_i(3402) := b"0000000000000000_0000000000000000_0010101101010101_1011001111001101"; -- 0.16927646395011
	pesos_i(3403) := b"1111111111111111_1111111111111111_1101001111100100_1111011101010001"; -- -0.17228750485038588
	pesos_i(3404) := b"0000000000000000_0000000000000000_0000001101010010_1111011101010100"; -- 0.012984712536907942
	pesos_i(3405) := b"0000000000000000_0000000000000000_0001100011000100_1011010111011100"; -- 0.0967515622500255
	pesos_i(3406) := b"0000000000000000_0000000000000000_0000111100011111_1001000110010111"; -- 0.05907545024716791
	pesos_i(3407) := b"0000000000000000_0000000000000000_0010011101110100_1000101101110000"; -- 0.15412208062076346
	pesos_i(3408) := b"1111111111111111_1111111111111111_1111101011110100_1001100010010010"; -- -0.019705261567484228
	pesos_i(3409) := b"0000000000000000_0000000000000000_0010111011011010_0001110001100010"; -- 0.18301560772197561
	pesos_i(3410) := b"1111111111111111_1111111111111111_1110001100011010_1010010011100010"; -- -0.1128746936043989
	pesos_i(3411) := b"0000000000000000_0000000000000000_0001001001000011_0001111001111111"; -- 0.07133665649683574
	pesos_i(3412) := b"1111111111111111_1111111111111111_1101011111001001_0010110101110101"; -- -0.15708652388311448
	pesos_i(3413) := b"1111111111111111_1111111111111111_1101101100011010_0011011101001111"; -- -0.14413122489340882
	pesos_i(3414) := b"1111111111111111_1111111111111111_1110110110001100_1100011101100001"; -- -0.07207063556286408
	pesos_i(3415) := b"0000000000000000_0000000000000000_0001110101100110_1011111000011100"; -- 0.11484897785760517
	pesos_i(3416) := b"1111111111111111_1111111111111111_1111010011011010_0001010110101110"; -- -0.043547291758866534
	pesos_i(3417) := b"1111111111111111_1111111111111111_1101110010000111_0101111010101111"; -- -0.13855941981306735
	pesos_i(3418) := b"1111111111111111_1111111111111111_1110110101100010_1101110000111101"; -- -0.07271026156288764
	pesos_i(3419) := b"0000000000000000_0000000000000000_0000011101100111_0010001011001111"; -- 0.02891748009392512
	pesos_i(3420) := b"1111111111111111_1111111111111111_1110100001111001_0110010001110110"; -- -0.09189769847642001
	pesos_i(3421) := b"0000000000000000_0000000000000000_0010100101110110_1111000100000000"; -- 0.1619711519143306
	pesos_i(3422) := b"0000000000000000_0000000000000000_0001110010001110_1100001101010101"; -- 0.11155339066690156
	pesos_i(3423) := b"0000000000000000_0000000000000000_0010110011011001_1101000000101100"; -- 0.17519856526612335
	pesos_i(3424) := b"0000000000000000_0000000000000000_0010011000100100_0100000000110101"; -- 0.14899064347001298
	pesos_i(3425) := b"0000000000000000_0000000000000000_0000010011001011_1101100010110110"; -- 0.0187354512457765
	pesos_i(3426) := b"0000000000000000_0000000000000000_0000000011010100_0100000001111010"; -- 0.0032387064407041126
	pesos_i(3427) := b"1111111111111111_1111111111111111_1110100001010011_0000110010101110"; -- -0.09248276464812347
	pesos_i(3428) := b"1111111111111111_1111111111111111_1101001101001011_1001000110111111"; -- -0.1746281536959505
	pesos_i(3429) := b"1111111111111111_1111111111111111_1110000001111110_0110110110011110"; -- -0.12307085883341003
	pesos_i(3430) := b"1111111111111111_1111111111111111_1111000100001001_0111011001111000"; -- -0.05844935971940309
	pesos_i(3431) := b"0000000000000000_0000000000000000_0001101101111101_1100011001111100"; -- 0.10738792931666633
	pesos_i(3432) := b"0000000000000000_0000000000000000_0001001110000100_1011111011100100"; -- 0.07624428814850784
	pesos_i(3433) := b"0000000000000000_0000000000000000_0001001110101100_0100110100100010"; -- 0.07684785926109483
	pesos_i(3434) := b"1111111111111111_1111111111111111_1101101011010111_0110010100000010"; -- -0.14515083990206773
	pesos_i(3435) := b"0000000000000000_0000000000000000_0010011001101100_1110101100101011"; -- 0.15009946632819857
	pesos_i(3436) := b"1111111111111111_1111111111111111_1111111101110101_0000111110101101"; -- -0.0021200374215994185
	pesos_i(3437) := b"1111111111111111_1111111111111111_1111011011011100_0110000011000000"; -- -0.035699799759558185
	pesos_i(3438) := b"0000000000000000_0000000000000000_0001110000100111_1011100100101100"; -- 0.10998112988581317
	pesos_i(3439) := b"0000000000000000_0000000000000000_0000001110111111_1001101110101110"; -- 0.014642457978484015
	pesos_i(3440) := b"0000000000000000_0000000000000000_0001001011111010_1010100000011111"; -- 0.07413721812108218
	pesos_i(3441) := b"0000000000000000_0000000000000000_0000110001000111_1001110111000100"; -- 0.0479677776909065
	pesos_i(3442) := b"0000000000000000_0000000000000000_0000000000110100_1110100101101110"; -- 0.000807370545740925
	pesos_i(3443) := b"0000000000000000_0000000000000000_0010000101000110_0111101110110011"; -- 0.12998173836107077
	pesos_i(3444) := b"0000000000000000_0000000000000000_0001010011110000_1110100100111010"; -- 0.08180101085941009
	pesos_i(3445) := b"1111111111111111_1111111111111111_1111001010111010_0101001101110001"; -- -0.051844391784735974
	pesos_i(3446) := b"0000000000000000_0000000000000000_0001001000110111_0111011110110110"; -- 0.0711588686864903
	pesos_i(3447) := b"1111111111111111_1111111111111111_1111000001000100_1010101100111011"; -- -0.061452196231139476
	pesos_i(3448) := b"1111111111111111_1111111111111111_1110010101011100_1000100010101011"; -- -0.10405679535916369
	pesos_i(3449) := b"1111111111111111_1111111111111111_1111011111110111_0100101110111101"; -- -0.0313828147983379
	pesos_i(3450) := b"0000000000000000_0000000000000000_0000001110010001_0101110110000001"; -- 0.013936847636875032
	pesos_i(3451) := b"1111111111111111_1111111111111111_1101111001010110_0010011011010010"; -- -0.13149793025153747
	pesos_i(3452) := b"0000000000000000_0000000000000000_0001101111110100_0110011001001101"; -- 0.10919799206872997
	pesos_i(3453) := b"1111111111111111_1111111111111111_1110100000010000_1110111001101010"; -- -0.09349164883625904
	pesos_i(3454) := b"1111111111111111_1111111111111111_1110010000001100_1100111101100000"; -- -0.10917953410596991
	pesos_i(3455) := b"1111111111111111_1111111111111111_1111001001101010_1010100110011010"; -- -0.05305995926295267
	pesos_i(3456) := b"0000000000000000_0000000000000000_0000101101001110_0110110011100101"; -- 0.04416542606494167
	pesos_i(3457) := b"0000000000000000_0000000000000000_0010011111001010_1111100001101001"; -- 0.15544083169030362
	pesos_i(3458) := b"0000000000000000_0000000000000000_0001011101110010_0100101000011011"; -- 0.09158766890529167
	pesos_i(3459) := b"1111111111111111_1111111111111111_1111011110110110_1001111011000011"; -- -0.03236968738074186
	pesos_i(3460) := b"1111111111111111_1111111111111111_1101001010100111_0011001001100000"; -- -0.1771362795923456
	pesos_i(3461) := b"0000000000000000_0000000000000000_0000000111011101_1101111010110110"; -- 0.00729171704732239
	pesos_i(3462) := b"1111111111111111_1111111111111111_1111001101011000_1011010110011000"; -- -0.0494276528271087
	pesos_i(3463) := b"0000000000000000_0000000000000000_0000110111111101_0100001010100101"; -- 0.05464569585540404
	pesos_i(3464) := b"0000000000000000_0000000000000000_0011011011000111_1100110101011100"; -- 0.21398623942862227
	pesos_i(3465) := b"0000000000000000_0000000000000000_0000001110110111_0001110001101000"; -- 0.014512801594480942
	pesos_i(3466) := b"0000000000000000_0000000000000000_0000110111010000_1110011011101010"; -- 0.05396884171551514
	pesos_i(3467) := b"1111111111111111_1111111111111111_1110000011110110_0100011100100001"; -- -0.12124209839265224
	pesos_i(3468) := b"1111111111111111_1111111111111111_1110001111101111_1111111000110001"; -- -0.10961924847580777
	pesos_i(3469) := b"0000000000000000_0000000000000000_0000100011110011_0110100011011101"; -- 0.0349641360817772
	pesos_i(3470) := b"1111111111111111_1111111111111111_1111001110010111_1101011000001011"; -- -0.048464414927226994
	pesos_i(3471) := b"1111111111111111_1111111111111111_1111010101000110_1001101011100100"; -- -0.04189140246270023
	pesos_i(3472) := b"0000000000000000_0000000000000000_0000100110111101_0010110100000110"; -- 0.03804284478207329
	pesos_i(3473) := b"1111111111111111_1111111111111111_1111010100101000_1101011010001100"; -- -0.042345610415380514
	pesos_i(3474) := b"0000000000000000_0000000000000000_0000110001100001_1100010101011101"; -- 0.048366866228877474
	pesos_i(3475) := b"0000000000000000_0000000000000000_0010100001011101_1101001001101001"; -- 0.15768160871993242
	pesos_i(3476) := b"0000000000000000_0000000000000000_0000010011110101_1110000001010001"; -- 0.019376773593822276
	pesos_i(3477) := b"0000000000000000_0000000000000000_0010000100010110_1101001101000111"; -- 0.12925453647791948
	pesos_i(3478) := b"0000000000000000_0000000000000000_0000111100100011_1111001000000011"; -- 0.05914223253508089
	pesos_i(3479) := b"1111111111111111_1111111111111111_1110110111101001_1010110010011100"; -- -0.07065316385158284
	pesos_i(3480) := b"0000000000000000_0000000000000000_0000000010101000_1111100100110010"; -- 0.002578329762504054
	pesos_i(3481) := b"1111111111111111_1111111111111111_1111001011110111_1001111010101011"; -- -0.050909121803860896
	pesos_i(3482) := b"0000000000000000_0000000000000000_0000100110110110_0001001010000000"; -- 0.037934452300338706
	pesos_i(3483) := b"0000000000000000_0000000000000000_0001110111010000_0111011110000001"; -- 0.11646220111267848
	pesos_i(3484) := b"1111111111111111_1111111111111111_1110110100111100_1000011100010001"; -- -0.07329517208310408
	pesos_i(3485) := b"1111111111111111_1111111111111111_1101101011011001_1010100111101000"; -- -0.14511621563963847
	pesos_i(3486) := b"1111111111111111_1111111111111111_1110001010011001_1110100000001000"; -- -0.11483907503533561
	pesos_i(3487) := b"1111111111111111_1111111111111111_1110001001000100_1001011000100111"; -- -0.1161409526787113
	pesos_i(3488) := b"0000000000000000_0000000000000000_0000111001001001_0011101010111011"; -- 0.0558048921587648
	pesos_i(3489) := b"1111111111111111_1111111111111111_1101101101010010_1000000011101100"; -- -0.14327234496875918
	pesos_i(3490) := b"1111111111111111_1111111111111111_1110111000110100_1010001111100000"; -- -0.06950927529736016
	pesos_i(3491) := b"1111111111111111_1111111111111111_1111101011101010_1111110001110001"; -- -0.01985189672805704
	pesos_i(3492) := b"0000000000000000_0000000000000000_0000001100110011_0001001011001001"; -- 0.012498067826898138
	pesos_i(3493) := b"1111111111111111_1111111111111111_1110011110101101_0010100110100001"; -- -0.09501399818995235
	pesos_i(3494) := b"0000000000000000_0000000000000000_0000101101010001_0110011100111010"; -- 0.044210864652275986
	pesos_i(3495) := b"0000000000000000_0000000000000000_0000011101111001_0011110010000101"; -- 0.029193670746984868
	pesos_i(3496) := b"1111111111111111_1111111111111111_1111001111111111_0011011100100010"; -- -0.04688697260650049
	pesos_i(3497) := b"0000000000000000_0000000000000000_0010001011011011_0000001101110000"; -- 0.13615437971090105
	pesos_i(3498) := b"1111111111111111_1111111111111111_1101100101100000_0001100001010011"; -- -0.15087745638106054
	pesos_i(3499) := b"0000000000000000_0000000000000000_0001001010101010_1011011101111110"; -- 0.07291743109708823
	pesos_i(3500) := b"1111111111111111_1111111111111111_1111110111011110_1101010101001011"; -- -0.008318585586986045
	pesos_i(3501) := b"0000000000000000_0000000000000000_0000001100001011_1111100001011101"; -- 0.011901400242123765
	pesos_i(3502) := b"1111111111111111_1111111111111111_1101001011100101_0000001101101101"; -- -0.17619303306138753
	pesos_i(3503) := b"0000000000000000_0000000000000000_0010001110110010_1011011101001011"; -- 0.13944573947487454
	pesos_i(3504) := b"0000000000000000_0000000000000000_0000000001111111_1110001111110101"; -- 0.0019514534143386941
	pesos_i(3505) := b"1111111111111111_1111111111111111_1110001101101101_0111100110000010"; -- -0.11161079959366797
	pesos_i(3506) := b"1111111111111111_1111111111111111_1111001100100111_0111110100001011"; -- -0.05017870399927885
	pesos_i(3507) := b"1111111111111111_1111111111111111_1111010100110000_0110000100111111"; -- -0.04223053190374911
	pesos_i(3508) := b"1111111111111111_1111111111111111_1110010110001101_1110101001000001"; -- -0.10330329813279496
	pesos_i(3509) := b"0000000000000000_0000000000000000_0000111010110001_1100011001100100"; -- 0.05740013061762983
	pesos_i(3510) := b"1111111111111111_1111111111111111_1111100001100110_0110001011001100"; -- -0.029687714845758918
	pesos_i(3511) := b"0000000000000000_0000000000000000_0010001111101110_1111000011110111"; -- 0.14036470453089436
	pesos_i(3512) := b"0000000000000000_0000000000000000_0010011010001110_0000001110001111"; -- 0.1506044600459496
	pesos_i(3513) := b"0000000000000000_0000000000000000_0000101001100100_1100001101001000"; -- 0.04060001847691672
	pesos_i(3514) := b"1111111111111111_1111111111111111_1111010110100110_0111001001110101"; -- -0.0404289688276123
	pesos_i(3515) := b"0000000000000000_0000000000000000_0001101111010100_0011001000010011"; -- 0.10870659785423444
	pesos_i(3516) := b"1111111111111111_1111111111111111_1110111010111111_0011001011011100"; -- -0.06739503981298163
	pesos_i(3517) := b"0000000000000000_0000000000000000_0001110101110100_0111100000100101"; -- 0.11505843059446802
	pesos_i(3518) := b"1111111111111111_1111111111111111_1110001001010101_1110100111101110"; -- -0.11587655969517159
	pesos_i(3519) := b"1111111111111111_1111111111111111_1111001110000101_1100010101101100"; -- -0.048740063877816785
	pesos_i(3520) := b"0000000000000000_0000000000000000_0010001110110110_1010011000100110"; -- 0.13950575272603152
	pesos_i(3521) := b"0000000000000000_0000000000000000_0000110100001111_1000111101001101"; -- 0.05101867312517988
	pesos_i(3522) := b"0000000000000000_0000000000000000_0000011001101001_0110001110000010"; -- 0.025045604032630644
	pesos_i(3523) := b"1111111111111111_1111111111111111_1110011001111101_1011011010100001"; -- -0.0996442658432755
	pesos_i(3524) := b"0000000000000000_0000000000000000_0001001000101101_0001010101011011"; -- 0.07100041844390428
	pesos_i(3525) := b"0000000000000000_0000000000000000_0000010001100101_0001001000001110"; -- 0.01716721376797514
	pesos_i(3526) := b"0000000000000000_0000000000000000_0001111100000110_0010001100110100"; -- 0.12118740109323282
	pesos_i(3527) := b"0000000000000000_0000000000000000_0010101111011100_1110010011110001"; -- 0.1713393294926571
	pesos_i(3528) := b"1111111111111111_1111111111111111_1110000110101110_1001010011101111"; -- -0.1184298435131826
	pesos_i(3529) := b"1111111111111111_1111111111111111_1111011010001111_1011111111010001"; -- -0.03686906001912072
	pesos_i(3530) := b"0000000000000000_0000000000000000_0000111000110101_1001000110110110"; -- 0.05550490082621728
	pesos_i(3531) := b"1111111111111111_1111111111111111_1101010100001011_0110001001010001"; -- -0.16779504326071668
	pesos_i(3532) := b"0000000000000000_0000000000000000_0001001001011000_1100000101000101"; -- 0.07166679318919489
	pesos_i(3533) := b"1111111111111111_1111111111111111_1101101001010111_1110011011001010"; -- -0.14709622924314922
	pesos_i(3534) := b"1111111111111111_1111111111111111_1101110111001000_1011010001011110"; -- -0.13365624148322525
	pesos_i(3535) := b"0000000000000000_0000000000000000_0001010111100101_1110100100001111"; -- 0.08553940408672171
	pesos_i(3536) := b"1111111111111111_1111111111111111_1111110010001111_1000011100011111"; -- -0.013434939210652336
	pesos_i(3537) := b"0000000000000000_0000000000000000_0001110011110000_1100001011111010"; -- 0.11304873092830378
	pesos_i(3538) := b"0000000000000000_0000000000000000_0000101000111010_1111110000111010"; -- 0.03996254362697462
	pesos_i(3539) := b"1111111111111111_1111111111111111_1110000110101101_0101000100111001"; -- -0.1184491382263761
	pesos_i(3540) := b"1111111111111111_1111111111111111_1110111101110101_1000001000101110"; -- -0.06461321232442686
	pesos_i(3541) := b"1111111111111111_1111111111111111_1101011111000110_1011111011111010"; -- -0.15712362657139797
	pesos_i(3542) := b"0000000000000000_0000000000000000_0000100111011101_0101000000011110"; -- 0.03853321774886698
	pesos_i(3543) := b"1111111111111111_1111111111111111_1111011110111010_1011001000001011"; -- -0.032307502959469755
	pesos_i(3544) := b"1111111111111111_1111111111111111_1110000100101101_1001111101110011"; -- -0.12039760061781607
	pesos_i(3545) := b"0000000000000000_0000000000000000_0001111010011010_1000110100101111"; -- 0.11954576869954874
	pesos_i(3546) := b"1111111111111111_1111111111111111_1101111010100001_0100101101001010"; -- -0.13035134739650622
	pesos_i(3547) := b"0000000000000000_0000000000000000_0000101111001011_0100000100111001"; -- 0.04607017168821107
	pesos_i(3548) := b"0000000000000000_0000000000000000_0010111010110100_0010000111111011"; -- 0.1824361074926381
	pesos_i(3549) := b"1111111111111111_1111111111111111_1111000010101100_0101000001011000"; -- -0.05987069932723272
	pesos_i(3550) := b"0000000000000000_0000000000000000_0010100111011110_0011111000101000"; -- 0.1635474058807211
	pesos_i(3551) := b"1111111111111111_1111111111111111_1110000100110011_0111110001111100"; -- -0.12030813185294464
	pesos_i(3552) := b"0000000000000000_0000000000000000_0010000011010010_1011001001100110"; -- 0.12821497913170352
	pesos_i(3553) := b"0000000000000000_0000000000000000_0000110001110100_1011100010101111"; -- 0.04865602750567461
	pesos_i(3554) := b"1111111111111111_1111111111111111_1111001111111101_1101010001111011"; -- -0.04690811152326231
	pesos_i(3555) := b"1111111111111111_1111111111111111_1110000000011001_1100011101010011"; -- -0.12460664959847838
	pesos_i(3556) := b"0000000000000000_0000000000000000_0010000110100100_1110001000011100"; -- 0.1314221684898239
	pesos_i(3557) := b"0000000000000000_0000000000000000_0000000000100010_0000100101010000"; -- 0.0005193539634364608
	pesos_i(3558) := b"1111111111111111_1111111111111111_1101100110101011_0100101110110110"; -- -0.14972998426993325
	pesos_i(3559) := b"0000000000000000_0000000000000000_0010000101000001_0010001110010101"; -- 0.12990019211430473
	pesos_i(3560) := b"1111111111111111_1111111111111111_1111010010010101_0100000001011110"; -- -0.04459760378397595
	pesos_i(3561) := b"0000000000000000_0000000000000000_0001100011100010_0111110010101011"; -- 0.09720591703083821
	pesos_i(3562) := b"1111111111111111_1111111111111111_1110001011100000_1110010111100101"; -- -0.11375582854725814
	pesos_i(3563) := b"1111111111111111_1111111111111111_1101010101111001_1100001011011001"; -- -0.16611082281200332
	pesos_i(3564) := b"0000000000000000_0000000000000000_0001100010001000_0001010101010101"; -- 0.09582646684530584
	pesos_i(3565) := b"1111111111111111_1111111111111111_1111101101110110_1010111000011000"; -- -0.017720336008334468
	pesos_i(3566) := b"0000000000000000_0000000000000000_0001100101000101_1011111011101001"; -- 0.09872048552621854
	pesos_i(3567) := b"0000000000000000_0000000000000000_0001000100011001_0010000010001100"; -- 0.06678965974403742
	pesos_i(3568) := b"1111111111111111_1111111111111111_1111000010100010_1000010010010000"; -- -0.06002017477578643
	pesos_i(3569) := b"1111111111111111_1111111111111111_1110101101011110_1011100101011001"; -- -0.08058587627904794
	pesos_i(3570) := b"0000000000000000_0000000000000000_0010011101011110_1010011011010100"; -- 0.15378801981485493
	pesos_i(3571) := b"0000000000000000_0000000000000000_0001101111001110_1110100001001001"; -- 0.10862590578170818
	pesos_i(3572) := b"1111111111111111_1111111111111111_1111010100110000_0010010100110000"; -- -0.04223411158543155
	pesos_i(3573) := b"1111111111111111_1111111111111111_1101101000010101_1110010010001100"; -- -0.14810344304412906
	pesos_i(3574) := b"0000000000000000_0000000000000000_0010110101011100_1101001101010110"; -- 0.17719765514945307
	pesos_i(3575) := b"1111111111111111_1111111111111111_1111001110000001_1111001011011001"; -- -0.04879839142728612
	pesos_i(3576) := b"1111111111111111_1111111111111111_1111101010010101_1001000000110000"; -- -0.021155346140642906
	pesos_i(3577) := b"1111111111111111_1111111111111111_1101110000010111_1101010010010010"; -- -0.14026137763062202
	pesos_i(3578) := b"1111111111111111_1111111111111111_1110110011011100_0011111000100100"; -- -0.07476436261723729
	pesos_i(3579) := b"0000000000000000_0000000000000000_0001011001101110_1000011100001111"; -- 0.08762401691818364
	pesos_i(3580) := b"0000000000000000_0000000000000000_0001000111100110_0111010011010010"; -- 0.06992273454843091
	pesos_i(3581) := b"1111111111111111_1111111111111111_1110011000011110_0001000101010010"; -- -0.10110370398371835
	pesos_i(3582) := b"0000000000000000_0000000000000000_0000110011010011_1110000111101001"; -- 0.05010806975738218
	pesos_i(3583) := b"1111111111111111_1111111111111111_1110100110011111_1001100110100100"; -- -0.08740844478484545
	pesos_i(3584) := b"0000000000000000_0000000000000000_0010010010001100_0101000000111101"; -- 0.14276601295623778
	pesos_i(3585) := b"1111111111111111_1111111111111111_1111011000100111_1011000011000100"; -- -0.038456871286871766
	pesos_i(3586) := b"1111111111111111_1111111111111111_1110111110111100_0101100101001000"; -- -0.06353227614989392
	pesos_i(3587) := b"0000000000000000_0000000000000000_0001011011001000_1110001110000111"; -- 0.08900281950421139
	pesos_i(3588) := b"1111111111111111_1111111111111111_1110110010001100_0100011011110111"; -- -0.07598453972200013
	pesos_i(3589) := b"1111111111111111_1111111111111111_1101100111011101_1110101011001101"; -- -0.1489575624132207
	pesos_i(3590) := b"0000000000000000_0000000000000000_0000001010001110_1010001100110111"; -- 0.009988976395812713
	pesos_i(3591) := b"1111111111111111_1111111111111111_1111000101000100_0010000001101111"; -- -0.05755421914815824
	pesos_i(3592) := b"0000000000000000_0000000000000000_0010000011101111_1001000101101100"; -- 0.12865551843250708
	pesos_i(3593) := b"0000000000000000_0000000000000000_0001100100001101_0100001011011010"; -- 0.09785859884521929
	pesos_i(3594) := b"1111111111111111_1111111111111111_1111010111111001_0100111001010001"; -- -0.039164643389865694
	pesos_i(3595) := b"1111111111111111_1111111111111111_1111100100111110_1101100101110001"; -- -0.02638474462962706
	pesos_i(3596) := b"0000000000000000_0000000000000000_0000111111001101_0011010000000010"; -- 0.06172490171240791
	pesos_i(3597) := b"0000000000000000_0000000000000000_0000010101000000_1010010010101010"; -- 0.020517627351699444
	pesos_i(3598) := b"0000000000000000_0000000000000000_0000101111001001_1100110100000111"; -- 0.0460479872832877
	pesos_i(3599) := b"0000000000000000_0000000000000000_0001111101010101_0010110101100010"; -- 0.12239345204207644
	pesos_i(3600) := b"0000000000000000_0000000000000000_0000100101101010_0110001100100110"; -- 0.036779591264044315
	pesos_i(3601) := b"0000000000000000_0000000000000000_0000011110101000_1110100001100000"; -- 0.029921077292865896
	pesos_i(3602) := b"0000000000000000_0000000000000000_0001010001111011_0111011110100010"; -- 0.08000896175582146
	pesos_i(3603) := b"1111111111111111_1111111111111111_1101100101001011_1011010000011011"; -- -0.1511886056145076
	pesos_i(3604) := b"0000000000000000_0000000000000000_0001111000001110_0010011011000000"; -- 0.11740343261363541
	pesos_i(3605) := b"1111111111111111_1111111111111111_1111100100101111_0001001001100100"; -- -0.026625490773897847
	pesos_i(3606) := b"1111111111111111_1111111111111111_1110100000010010_0100011001000000"; -- -0.09347115458897767
	pesos_i(3607) := b"0000000000000000_0000000000000000_0010101001101000_1001011100110000"; -- 0.16565842563292832
	pesos_i(3608) := b"0000000000000000_0000000000000000_0000000100100011_1100100011100101"; -- 0.00445228178439031
	pesos_i(3609) := b"0000000000000000_0000000000000000_0001011000000011_0011111100111000"; -- 0.08598704443094338
	pesos_i(3610) := b"1111111111111111_1111111111111111_1111001101110011_1101010011010100"; -- -0.04901380376110271
	pesos_i(3611) := b"0000000000000000_0000000000000000_0000001000010100_1000000110100000"; -- 0.008125402114245577
	pesos_i(3612) := b"0000000000000000_0000000000000000_0000001100000111_0001001100001001"; -- 0.011826696027752244
	pesos_i(3613) := b"0000000000000000_0000000000000000_0000110010010111_0100111011001101"; -- 0.049183773994789584
	pesos_i(3614) := b"1111111111111111_1111111111111111_1101100001110110_0110011101011111"; -- -0.15444330150078683
	pesos_i(3615) := b"0000000000000000_0000000000000000_0001010101111000_0101110011111101"; -- 0.0838678471253839
	pesos_i(3616) := b"0000000000000000_0000000000000000_0001111111000111_1000101011110100"; -- 0.12413853133357253
	pesos_i(3617) := b"0000000000000000_0000000000000000_0000101110011010_0000010001011101"; -- 0.045318863474940685
	pesos_i(3618) := b"1111111111111111_1111111111111111_1110110011000110_1111110100110000"; -- -0.07508866863859821
	pesos_i(3619) := b"0000000000000000_0000000000000000_0010011101101011_0100001111100110"; -- 0.15398048746591916
	pesos_i(3620) := b"0000000000000000_0000000000000000_0000111001101100_1001111111101110"; -- 0.05634498188635324
	pesos_i(3621) := b"1111111111111111_1111111111111111_1110011010110010_0001001011011100"; -- -0.09884531154734039
	pesos_i(3622) := b"1111111111111111_1111111111111111_1111111110010110_1011100001101111"; -- -0.0016064386127809568
	pesos_i(3623) := b"0000000000000000_0000000000000000_0001011010000010_0010111110001110"; -- 0.08792397715842046
	pesos_i(3624) := b"0000000000000000_0000000000000000_0000101011010000_0011011100010010"; -- 0.04223961050693095
	pesos_i(3625) := b"1111111111111111_1111111111111111_1110100111011011_1100000101000101"; -- -0.08649055549296997
	pesos_i(3626) := b"1111111111111111_1111111111111111_1101100100110111_1000011111011010"; -- -0.15149641920702353
	pesos_i(3627) := b"0000000000000000_0000000000000000_0000000000001110_0011100100100011"; -- 0.0002170286742056121
	pesos_i(3628) := b"1111111111111111_1111111111111111_1111010100100100_1110110011101100"; -- -0.04240531198197727
	pesos_i(3629) := b"0000000000000000_0000000000000000_0010010110011100_1011110010110010"; -- 0.14692286822601547
	pesos_i(3630) := b"0000000000000000_0000000000000000_0001100011010001_0000011100110001"; -- 0.09693951558663301
	pesos_i(3631) := b"1111111111111111_1111111111111111_1111000010011001_1001111000010011"; -- -0.06015598321491492
	pesos_i(3632) := b"1111111111111111_1111111111111111_1110111001010010_0100110010011000"; -- -0.06905671387914392
	pesos_i(3633) := b"0000000000000000_0000000000000000_0010001001100111_1011101110101011"; -- 0.13439534108021395
	pesos_i(3634) := b"1111111111111111_1111111111111111_1101100101100001_0101000100000101"; -- -0.1508588184268454
	pesos_i(3635) := b"0000000000000000_0000000000000000_0001111111111101_0100010111111000"; -- 0.12495839416119556
	pesos_i(3636) := b"0000000000000000_0000000000000000_0001000000101100_0101011100110100"; -- 0.06317658452129804
	pesos_i(3637) := b"0000000000000000_0000000000000000_0010110100001000_0000101100000010"; -- 0.17590397636068433
	pesos_i(3638) := b"0000000000000000_0000000000000000_0010000100110001_0111011000011111"; -- 0.12966097133958565
	pesos_i(3639) := b"0000000000000000_0000000000000000_0000100100010100_1101110110110111"; -- 0.035474640954712616
	pesos_i(3640) := b"1111111111111111_1111111111111111_1111100111000101_0011011110000000"; -- -0.024334460458731944
	pesos_i(3641) := b"1111111111111111_1111111111111111_1101110111101100_1110000110110100"; -- -0.13310422293771437
	pesos_i(3642) := b"0000000000000000_0000000000000000_0001100101001110_0000011000001011"; -- 0.09884679576786864
	pesos_i(3643) := b"0000000000000000_0000000000000000_0001111011101010_0000100101111111"; -- 0.12075862265563371
	pesos_i(3644) := b"0000000000000000_0000000000000000_0001100111011111_0101101101010110"; -- 0.10106440401442299
	pesos_i(3645) := b"1111111111111111_1111111111111111_1110001011100100_1101100000100010"; -- -0.11369561348185814
	pesos_i(3646) := b"0000000000000000_0000000000000000_0010011111101001_0101110100010100"; -- 0.15590459571714255
	pesos_i(3647) := b"0000000000000000_0000000000000000_0001010111011011_1000011111001011"; -- 0.08538101876921668
	pesos_i(3648) := b"1111111111111111_1111111111111111_1111100010010111_1111110101110111"; -- -0.028930815141779587
	pesos_i(3649) := b"1111111111111111_1111111111111111_1110010001111000_1000100100111010"; -- -0.10753576599878618
	pesos_i(3650) := b"1111111111111111_1111111111111111_1110011110011001_1010111010010111"; -- -0.09531124895092166
	pesos_i(3651) := b"1111111111111111_1111111111111111_1111101001011110_1110111011101101"; -- -0.021988932821970515
	pesos_i(3652) := b"0000000000000000_0000000000000000_0000000110101000_1111010011000100"; -- 0.006484315645047183
	pesos_i(3653) := b"0000000000000000_0000000000000000_0000100111101101_1001000000110110"; -- 0.03878117868268587
	pesos_i(3654) := b"1111111111111111_1111111111111111_1101100100100100_0000001110010010"; -- -0.15179422074448934
	pesos_i(3655) := b"0000000000000000_0000000000000000_0001111010100000_0010111110000000"; -- 0.11963173743359135
	pesos_i(3656) := b"1111111111111111_1111111111111111_1110001000001101_1101100111100010"; -- -0.11697614885889747
	pesos_i(3657) := b"0000000000000000_0000000000000000_0001100000111101_1010111000100000"; -- 0.09469116486084167
	pesos_i(3658) := b"1111111111111111_1111111111111111_1111111000100010_1011001001100110"; -- -0.007283067825632711
	pesos_i(3659) := b"0000000000000000_0000000000000000_0000111101111010_0000001001110100"; -- 0.06045546839761695
	pesos_i(3660) := b"0000000000000000_0000000000000000_0001111110001000_1011101000000001"; -- 0.12318003197214808
	pesos_i(3661) := b"1111111111111111_1111111111111111_1101111101000101_1000011001111100"; -- -0.12784537768081353
	pesos_i(3662) := b"1111111111111111_1111111111111111_1101011110010011_0101001111110000"; -- -0.15790820488610097
	pesos_i(3663) := b"0000000000000000_0000000000000000_0000110100011010_0001101001100100"; -- 0.05117955144006986
	pesos_i(3664) := b"1111111111111111_1111111111111111_1110111111110010_1010110111111001"; -- -0.0627032535043067
	pesos_i(3665) := b"0000000000000000_0000000000000000_0001110000100011_1001110001001000"; -- 0.1099183727826899
	pesos_i(3666) := b"1111111111111111_1111111111111111_1111001100100101_0110110100100111"; -- -0.05021016879341928
	pesos_i(3667) := b"0000000000000000_0000000000000000_0001011000101000_1101111001100101"; -- 0.08656110730050709
	pesos_i(3668) := b"1111111111111111_1111111111111111_1101100011000001_0101000011101010"; -- -0.15330023081653765
	pesos_i(3669) := b"1111111111111111_1111111111111111_1111100001001011_1011101001101010"; -- -0.030094479565185652
	pesos_i(3670) := b"1111111111111111_1111111111111111_1101011010010000_1010111010110100"; -- -0.16185482123511977
	pesos_i(3671) := b"0000000000000000_0000000000000000_0001101000110010_0111001011010100"; -- 0.10233228374998751
	pesos_i(3672) := b"0000000000000000_0000000000000000_0010100110011110_0000110010110111"; -- 0.1625678964641075
	pesos_i(3673) := b"1111111111111111_1111111111111111_1111001010110010_0111101100011001"; -- -0.051964098243941007
	pesos_i(3674) := b"1111111111111111_1111111111111111_1111101001000010_0010111101010110"; -- -0.022427598579196947
	pesos_i(3675) := b"1111111111111111_1111111111111111_1111101011100100_1101000000001111"; -- -0.0199460948918793
	pesos_i(3676) := b"0000000000000000_0000000000000000_0010100110101100_1111111010001101"; -- 0.16279593407641338
	pesos_i(3677) := b"0000000000000000_0000000000000000_0001011001110000_0111101101000010"; -- 0.08765383101423332
	pesos_i(3678) := b"0000000000000000_0000000000000000_0000001011101101_1100110010100111"; -- 0.011441031230324238
	pesos_i(3679) := b"0000000000000000_0000000000000000_0000010000010000_1001001100010100"; -- 0.015877907279852888
	pesos_i(3680) := b"0000000000000000_0000000000000000_0010011101011000_0001000001000110"; -- 0.1536874933190124
	pesos_i(3681) := b"0000000000000000_0000000000000000_0010001000001000_1100111010000110"; -- 0.13294687995690438
	pesos_i(3682) := b"1111111111111111_1111111111111111_1111100010011111_0000111000111111"; -- -0.02882300332922209
	pesos_i(3683) := b"0000000000000000_0000000000000000_0010000010000101_0000111010001011"; -- 0.127030285875705
	pesos_i(3684) := b"1111111111111111_1111111111111111_1110011010001000_1000110011000001"; -- -0.09947891504927361
	pesos_i(3685) := b"0000000000000000_0000000000000000_0001110100001010_0001110111111100"; -- 0.11343562510827114
	pesos_i(3686) := b"1111111111111111_1111111111111111_1101100111001000_1101011010011110"; -- -0.14927919990211191
	pesos_i(3687) := b"0000000000000000_0000000000000000_0000101100111110_1001111100001110"; -- 0.043924275340270685
	pesos_i(3688) := b"1111111111111111_1111111111111111_1111110101010100_0101100110101101"; -- -0.0104316667154849
	pesos_i(3689) := b"1111111111111111_1111111111111111_1101110110110111_1011100010000000"; -- -0.13391539446725895
	pesos_i(3690) := b"1111111111111111_1111111111111111_1111010001001001_1000101100001010"; -- -0.045752821053852706
	pesos_i(3691) := b"0000000000000000_0000000000000000_0010011111010110_0011100011111100"; -- 0.15561252732254288
	pesos_i(3692) := b"0000000000000000_0000000000000000_0001101010001101_1010111010100100"; -- 0.10372439862486972
	pesos_i(3693) := b"1111111111111111_1111111111111111_1110000101101101_1010010111000100"; -- -0.1194206615291647
	pesos_i(3694) := b"0000000000000000_0000000000000000_0010000001100011_0001011110000101"; -- 0.126512022050425
	pesos_i(3695) := b"0000000000000000_0000000000000000_0010000011110111_0110110000101111"; -- 0.12877536903355968
	pesos_i(3696) := b"0000000000000000_0000000000000000_0001110111001110_0010001010100000"; -- 0.11642662430421444
	pesos_i(3697) := b"0000000000000000_0000000000000000_0001000110000111_1110000001000001"; -- 0.06847955308788622
	pesos_i(3698) := b"1111111111111111_1111111111111111_1110001010011001_0000001001001101"; -- -0.11485276815092078
	pesos_i(3699) := b"1111111111111111_1111111111111111_1111110001111001_1000100001101101"; -- -0.013770554913844732
	pesos_i(3700) := b"1111111111111111_1111111111111111_1110111001100100_1110100100010111"; -- -0.06877272786840631
	pesos_i(3701) := b"1111111111111111_1111111111111111_1111010011001000_1101111000001110"; -- -0.04381000669573639
	pesos_i(3702) := b"0000000000000000_0000000000000000_0000110110011100_0110100111100111"; -- 0.05316793325291069
	pesos_i(3703) := b"1111111111111111_1111111111111111_1110001101000101_1101011101011010"; -- -0.1122155574991831
	pesos_i(3704) := b"0000000000000000_0000000000000000_0001111000010000_1111110010101011"; -- 0.1174467007163871
	pesos_i(3705) := b"0000000000000000_0000000000000000_0000111100100110_0011101001011010"; -- 0.05917706191789359
	pesos_i(3706) := b"1111111111111111_1111111111111111_1111010011100000_0010101001010010"; -- -0.043454508798575646
	pesos_i(3707) := b"0000000000000000_0000000000000000_0000000000011000_0101110001010111"; -- 0.0003717147739316714
	pesos_i(3708) := b"0000000000000000_0000000000000000_0001110000101100_0110100011111001"; -- 0.11005264354694894
	pesos_i(3709) := b"1111111111111111_1111111111111111_1111010000101100_1111101101101011"; -- -0.046188627675956904
	pesos_i(3710) := b"0000000000000000_0000000000000000_0010101100010111_1101011010100000"; -- 0.1683324947627561
	pesos_i(3711) := b"0000000000000000_0000000000000000_0010111111111100_1111000110100001"; -- 0.18745336699446694
	pesos_i(3712) := b"0000000000000000_0000000000000000_0000101110010110_0000001100011001"; -- 0.04525775303003182
	pesos_i(3713) := b"1111111111111111_1111111111111111_1110101001101001_0011010000000110"; -- -0.08433222622928584
	pesos_i(3714) := b"1111111111111111_1111111111111111_1111111101010100_0000101100010000"; -- -0.0026238523150159338
	pesos_i(3715) := b"1111111111111111_1111111111111111_1110001111010010_1110101101101101"; -- -0.11006287190342642
	pesos_i(3716) := b"1111111111111111_1111111111111111_1110011010011000_0111010000100110"; -- -0.09923624116940936
	pesos_i(3717) := b"1111111111111111_1111111111111111_1111100100110011_0011100111011000"; -- -0.026562103954025192
	pesos_i(3718) := b"1111111111111111_1111111111111111_1111011101100010_0100110100110000"; -- -0.03365628801324214
	pesos_i(3719) := b"1111111111111111_1111111111111111_1110100110100101_1110011100001010"; -- -0.08731227875151787
	pesos_i(3720) := b"1111111111111111_1111111111111111_1110001010111011_0011011011101100"; -- -0.11433083274018069
	pesos_i(3721) := b"0000000000000000_0000000000000000_0001101101010001_0101111101000011"; -- 0.10671038995606935
	pesos_i(3722) := b"1111111111111111_1111111111111111_1101010100100010_1100101111011010"; -- -0.16743780056292565
	pesos_i(3723) := b"1111111111111111_1111111111111111_1110111011111101_0101011110101101"; -- -0.06644680054940592
	pesos_i(3724) := b"0000000000000000_0000000000000000_0001001110111110_0011000100000000"; -- 0.07712084057154814
	pesos_i(3725) := b"1111111111111111_1111111111111111_1110000111100100_0011110101011010"; -- -0.11761108919459198
	pesos_i(3726) := b"1111111111111111_1111111111111111_1101101000010000_1000010010010001"; -- -0.1481854579143684
	pesos_i(3727) := b"0000000000000000_0000000000000000_0001111110111001_0001001110000010"; -- 0.12391778870369863
	pesos_i(3728) := b"0000000000000000_0000000000000000_0000010111011111_0100101110101101"; -- 0.022938470478104295
	pesos_i(3729) := b"0000000000000000_0000000000000000_0010010011111111_0110011010100001"; -- 0.14452210839361515
	pesos_i(3730) := b"0000000000000000_0000000000000000_0000110000110011_0001100000110101"; -- 0.04765464115960538
	pesos_i(3731) := b"0000000000000000_0000000000000000_0010101001000010_1010111000000001"; -- 0.16507995144481313
	pesos_i(3732) := b"0000000000000000_0000000000000000_0000001001010101_0100001001011000"; -- 0.00911345135423001
	pesos_i(3733) := b"1111111111111111_1111111111111111_1111010101000110_1010111111100111"; -- -0.04189015021621766
	pesos_i(3734) := b"0000000000000000_0000000000000000_0000110000101110_0011001111001000"; -- 0.04757999077301513
	pesos_i(3735) := b"0000000000000000_0000000000000000_0001001001010000_0001011001110111"; -- 0.07153454202360385
	pesos_i(3736) := b"0000000000000000_0000000000000000_0000100111111011_1000000110001000"; -- 0.038993926624999876
	pesos_i(3737) := b"0000000000000000_0000000000000000_0000011001111111_1011010101101001"; -- 0.025386179198333178
	pesos_i(3738) := b"1111111111111111_1111111111111111_1101001110111101_0001100000111001"; -- -0.17289589497335445
	pesos_i(3739) := b"1111111111111111_1111111111111111_1101110100111101_0000101000101000"; -- -0.13578735860606564
	pesos_i(3740) := b"0000000000000000_0000000000000000_0000101110111101_0001010111011100"; -- 0.04585396416121319
	pesos_i(3741) := b"0000000000000000_0000000000000000_0010010111011001_1111000110111100"; -- 0.14785681573254092
	pesos_i(3742) := b"1111111111111111_1111111111111111_1110011100101100_1011111011110101"; -- -0.09697348131784606
	pesos_i(3743) := b"1111111111111111_1111111111111111_1111111001100011_0111011000010001"; -- -0.006294842530679912
	pesos_i(3744) := b"0000000000000000_0000000000000000_0001101000010111_0100100000111001"; -- 0.10191775695129388
	pesos_i(3745) := b"0000000000000000_0000000000000000_0000110110001110_1001100110110011"; -- 0.05295715920575689
	pesos_i(3746) := b"0000000000000000_0000000000000000_0001100001101101_1111001001111111"; -- 0.09542766192693684
	pesos_i(3747) := b"0000000000000000_0000000000000000_0000000111011101_0000101000111110"; -- 0.007279052756410409
	pesos_i(3748) := b"1111111111111111_1111111111111111_1111111100111000_1000010110011100"; -- -0.003043794016343227
	pesos_i(3749) := b"0000000000000000_0000000000000000_0010100110101111_1011000011111010"; -- 0.16283708677649328
	pesos_i(3750) := b"1111111111111111_1111111111111111_1110101001011010_1010011110011111"; -- -0.08455421803647485
	pesos_i(3751) := b"0000000000000000_0000000000000000_0001000101000111_0111110110000110"; -- 0.06749710576208726
	pesos_i(3752) := b"1111111111111111_1111111111111111_1101101100100110_0011011010100111"; -- -0.14394815856899945
	pesos_i(3753) := b"1111111111111111_1111111111111111_1101001001011111_1001101111001011"; -- -0.17822862901414044
	pesos_i(3754) := b"0000000000000000_0000000000000000_0010000111001010_1011110100100010"; -- 0.1319997986974912
	pesos_i(3755) := b"1111111111111111_1111111111111111_1101011001110101_1000001001011100"; -- -0.16226945173441712
	pesos_i(3756) := b"1111111111111111_1111111111111111_1101011111001110_1011101000000111"; -- -0.15700185125507407
	pesos_i(3757) := b"0000000000000000_0000000000000000_0000101111011100_1010001111000111"; -- 0.04633544551247091
	pesos_i(3758) := b"0000000000000000_0000000000000000_0010110101110111_1000101000100010"; -- 0.17760527919273253
	pesos_i(3759) := b"0000000000000000_0000000000000000_0010000010001111_1010001001110010"; -- 0.12719168937601172
	pesos_i(3760) := b"1111111111111111_1111111111111111_1110101010011001_0111000010011011"; -- -0.08359619353465067
	pesos_i(3761) := b"1111111111111111_1111111111111111_1111000010001011_0001101011101000"; -- -0.060377424557801075
	pesos_i(3762) := b"0000000000000000_0000000000000000_0000001110101100_0011101100111000"; -- 0.014346791370603811
	pesos_i(3763) := b"0000000000000000_0000000000000000_0000000110100111_1101110100011010"; -- 0.006467646560301427
	pesos_i(3764) := b"0000000000000000_0000000000000000_0000110000100010_0101101011110101"; -- 0.04739922025005927
	pesos_i(3765) := b"0000000000000000_0000000000000000_0000011110010001_0101110110000110"; -- 0.029561848901518323
	pesos_i(3766) := b"0000000000000000_0000000000000000_0010011111011000_1000011111111100"; -- 0.1556477538512906
	pesos_i(3767) := b"1111111111111111_1111111111111111_1111110010001101_1001011100011100"; -- -0.013464503829899471
	pesos_i(3768) := b"1111111111111111_1111111111111111_1111111001000001_1100001000000111"; -- -0.006809113817287965
	pesos_i(3769) := b"0000000000000000_0000000000000000_0001111111010011_1011010100001101"; -- 0.12432414594449148
	pesos_i(3770) := b"1111111111111111_1111111111111111_1110100111100001_0010011011000110"; -- -0.08640821138892096
	pesos_i(3771) := b"1111111111111111_1111111111111111_1111000101010011_0111100001000001"; -- -0.05732010271828087
	pesos_i(3772) := b"1111111111111111_1111111111111111_1110111111110101_0001110000100110"; -- -0.06266616883425301
	pesos_i(3773) := b"1111111111111111_1111111111111111_1110001010010101_1000100110100011"; -- -0.11490573672720547
	pesos_i(3774) := b"0000000000000000_0000000000000000_0000010101011000_0000000110101010"; -- 0.02087412253265412
	pesos_i(3775) := b"0000000000000000_0000000000000000_0001000100011111_1010100001100111"; -- 0.06688930992368308
	pesos_i(3776) := b"0000000000000000_0000000000000000_0000000111100110_1111010110010000"; -- 0.007430408224128798
	pesos_i(3777) := b"0000000000000000_0000000000000000_0000001010111101_1110100001110010"; -- 0.010710266024506341
	pesos_i(3778) := b"0000000000000000_0000000000000000_0010000100101011_1100101010000001"; -- 0.12957444808337445
	pesos_i(3779) := b"1111111111111111_1111111111111111_1111101111001110_0001110010001010"; -- -0.016386238325543742
	pesos_i(3780) := b"0000000000000000_0000000000000000_0010000110100100_0011110000010101"; -- 0.1314122726874334
	pesos_i(3781) := b"1111111111111111_1111111111111111_1110110101101010_0010000010101000"; -- -0.07259937190788157
	pesos_i(3782) := b"0000000000000000_0000000000000000_0001001111100010_1000000100000111"; -- 0.07767492692365537
	pesos_i(3783) := b"1111111111111111_1111111111111111_1101010010110000_1110011110011111"; -- -0.16917564748327799
	pesos_i(3784) := b"1111111111111111_1111111111111111_1111011011000100_0100000110001100"; -- -0.03606787036060706
	pesos_i(3785) := b"1111111111111111_1111111111111111_1101100101000111_0110010010010100"; -- -0.15125438116575227
	pesos_i(3786) := b"0000000000000000_0000000000000000_0001001100010100_1100010000101110"; -- 0.07453561903548035
	pesos_i(3787) := b"1111111111111111_1111111111111111_1110100100011001_1011101001110000"; -- -0.0894511677827555
	pesos_i(3788) := b"0000000000000000_0000000000000000_0001100111011010_0011110011101010"; -- 0.10098629673798028
	pesos_i(3789) := b"0000000000000000_0000000000000000_0001010011011000_0111001110000100"; -- 0.08142778361234047
	pesos_i(3790) := b"1111111111111111_1111111111111111_1101101100111100_1111111110111101"; -- -0.1436004794778537
	pesos_i(3791) := b"1111111111111111_1111111111111111_1101101000101011_0010000100000110"; -- -0.14777940375135895
	pesos_i(3792) := b"0000000000000000_0000000000000000_0000010101000101_1111000010111000"; -- 0.020598454475821287
	pesos_i(3793) := b"0000000000000000_0000000000000000_0000100000011010_0010101000110010"; -- 0.03164924362857196
	pesos_i(3794) := b"1111111111111111_1111111111111111_1111010001110000_0101111111110001"; -- -0.04516029702381751
	pesos_i(3795) := b"1111111111111111_1111111111111111_1110000011111110_1110011110110101"; -- -0.12111045680129047
	pesos_i(3796) := b"0000000000000000_0000000000000000_0010100010101100_0010000011001111"; -- 0.15887646718870865
	pesos_i(3797) := b"0000000000000000_0000000000000000_0010011011101001_0011001001101001"; -- 0.15199580263402823
	pesos_i(3798) := b"0000000000000000_0000000000000000_0010011010010011_0110110100110001"; -- 0.15068705021292428
	pesos_i(3799) := b"0000000000000000_0000000000000000_0000110110010000_1101111101000010"; -- 0.05299182293468066
	pesos_i(3800) := b"1111111111111111_1111111111111111_1110011001010011_0011100000101111"; -- -0.1002926716859211
	pesos_i(3801) := b"0000000000000000_0000000000000000_0000101111000111_0010101101011001"; -- 0.04600783278909568
	pesos_i(3802) := b"1111111111111111_1111111111111111_1111000110000011_0110010101001001"; -- -0.05658881154003921
	pesos_i(3803) := b"1111111111111111_1111111111111111_1111001101111110_1001111011101011"; -- -0.048849170269415494
	pesos_i(3804) := b"0000000000000000_0000000000000000_0010010011100110_1111100001010110"; -- 0.14414932355627694
	pesos_i(3805) := b"1111111111111111_1111111111111111_1111011000101000_0010011110110010"; -- -0.03844978239642496
	pesos_i(3806) := b"0000000000000000_0000000000000000_0000010101101010_1011110000100011"; -- 0.021159895471470794
	pesos_i(3807) := b"0000000000000000_0000000000000000_0001000101100110_0100001001000001"; -- 0.06796659544664901
	pesos_i(3808) := b"0000000000000000_0000000000000000_0001100110100010_0000000111011001"; -- 0.10012828387670955
	pesos_i(3809) := b"0000000000000000_0000000000000000_0001110001100100_1001011111010101"; -- 0.11090992876744833
	pesos_i(3810) := b"1111111111111111_1111111111111111_1110011101111000_1001011011001010"; -- -0.0958162075041
	pesos_i(3811) := b"1111111111111111_1111111111111111_1111011001111100_0011100101101110"; -- -0.03716698716699179
	pesos_i(3812) := b"0000000000000000_0000000000000000_0010001100100000_0100010001000101"; -- 0.13721110032759934
	pesos_i(3813) := b"1111111111111111_1111111111111111_1101111011000110_0000010000111010"; -- -0.1297910079080779
	pesos_i(3814) := b"1111111111111111_1111111111111111_1110110111100001_0110111100011101"; -- -0.07077889955247768
	pesos_i(3815) := b"0000000000000000_0000000000000000_0000100110010110_1111001111100000"; -- 0.03745960449502733
	pesos_i(3816) := b"1111111111111111_1111111111111111_1111101011010001_0111110000001110"; -- -0.02024101895417954
	pesos_i(3817) := b"1111111111111111_1111111111111111_1110001001010001_1001111011001110"; -- -0.11594207263207956
	pesos_i(3818) := b"0000000000000000_0000000000000000_0001111011101010_1110110010100100"; -- 0.12077216141235866
	pesos_i(3819) := b"1111111111111111_1111111111111111_1110000100110111_1101011101110111"; -- -0.12024167383867189
	pesos_i(3820) := b"1111111111111111_1111111111111111_1111011000101100_1100011001000011"; -- -0.038379295962209514
	pesos_i(3821) := b"0000000000000000_0000000000000000_0000011101000101_0110101010010111"; -- 0.028402959707679202
	pesos_i(3822) := b"0000000000000000_0000000000000000_0000001101100100_1010101110110110"; -- 0.01325486371815899
	pesos_i(3823) := b"0000000000000000_0000000000000000_0001101101000100_1101100111110100"; -- 0.10651933874860589
	pesos_i(3824) := b"1111111111111111_1111111111111111_1101111000111110_0011000000010001"; -- -0.1318635900945704
	pesos_i(3825) := b"0000000000000000_0000000000000000_0001001011000010_1100000001110100"; -- 0.07328417617093465
	pesos_i(3826) := b"0000000000000000_0000000000000000_0010001010010111_0101001000110111"; -- 0.13512147742023747
	pesos_i(3827) := b"0000000000000000_0000000000000000_0001101110001111_0111100001100000"; -- 0.1076579317162667
	pesos_i(3828) := b"1111111111111111_1111111111111111_1110011101001101_0110100111100111"; -- -0.09647501089602485
	pesos_i(3829) := b"0000000000000000_0000000000000000_0010100101100000_0101101011111110"; -- 0.16162651721337565
	pesos_i(3830) := b"1111111111111111_1111111111111111_1110001010101000_0010110111010100"; -- -0.11462129185903719
	pesos_i(3831) := b"0000000000000000_0000000000000000_0000001010100000_0100101111111010"; -- 0.010258434868348413
	pesos_i(3832) := b"0000000000000000_0000000000000000_0000001111100010_1011100010000001"; -- 0.015178233619249248
	pesos_i(3833) := b"1111111111111111_1111111111111111_1101001101111001_1000011111000100"; -- -0.17392684420831717
	pesos_i(3834) := b"1111111111111111_1111111111111111_1110001000110011_0000100000000001"; -- -0.11640882478621928
	pesos_i(3835) := b"1111111111111111_1111111111111111_1111100111100100_0101000111100011"; -- -0.023859865307527785
	pesos_i(3836) := b"0000000000000000_0000000000000000_0001011001000000_1101100111010110"; -- 0.08692704646959101
	pesos_i(3837) := b"1111111111111111_1111111111111111_1101100010111111_1001101110111111"; -- -0.1533262880847079
	pesos_i(3838) := b"0000000000000000_0000000000000000_0010000011001110_0100100111001100"; -- 0.12814770929230798
	pesos_i(3839) := b"1111111111111111_1111111111111111_1110001001110001_0100100001101110"; -- -0.11545893976266305
	pesos_i(3840) := b"0000000000000000_0000000000000000_0010100111101100_0110110110010001"; -- 0.16376385482364683
	pesos_i(3841) := b"1111111111111111_1111111111111111_1110100001111001_1010101011100110"; -- -0.0918935002015409
	pesos_i(3842) := b"0000000000000000_0000000000000000_0010001001010110_1100110110000110"; -- 0.13413700606917753
	pesos_i(3843) := b"0000000000000000_0000000000000000_0010010100010000_0001000011111110"; -- 0.14477640339976441
	pesos_i(3844) := b"0000000000000000_0000000000000000_0010011100110011_1110110101001000"; -- 0.15313609136918457
	pesos_i(3845) := b"0000000000000000_0000000000000000_0010000101010000_1010111110100011"; -- 0.1301374218191907
	pesos_i(3846) := b"1111111111111111_1111111111111111_1111110111100110_0110000011001100"; -- -0.00820345888428753
	pesos_i(3847) := b"0000000000000000_0000000000000000_0001111110110001_0000011111101001"; -- 0.12379502725752037
	pesos_i(3848) := b"0000000000000000_0000000000000000_0000100110110010_1001110110000100"; -- 0.037881703003825144
	pesos_i(3849) := b"0000000000000000_0000000000000000_0010010100101011_0000100111110000"; -- 0.145187970221518
	pesos_i(3850) := b"0000000000000000_0000000000000000_0000111110000000_0101000000111100"; -- 0.06055165723572622
	pesos_i(3851) := b"0000000000000000_0000000000000000_0010101110010110_1000100111111111"; -- 0.17026579353151558
	pesos_i(3852) := b"1111111111111111_1111111111111111_1110111110000100_1101011111011010"; -- -0.06437922410536544
	pesos_i(3853) := b"0000000000000000_0000000000000000_0010011001101001_0000001000011101"; -- 0.1500397987034533
	pesos_i(3854) := b"1111111111111111_1111111111111111_1101001100010011_0011001110100010"; -- -0.1754882554458725
	pesos_i(3855) := b"0000000000000000_0000000000000000_0001111100101100_1100010001110000"; -- 0.12177684532830528
	pesos_i(3856) := b"1111111111111111_1111111111111111_1101110100101001_1011111100011011"; -- -0.1360817489000329
	pesos_i(3857) := b"1111111111111111_1111111111111111_1111000111110001_1100000001011100"; -- -0.05490491624662875
	pesos_i(3858) := b"0000000000000000_0000000000000000_0000101011110111_0111101001001001"; -- 0.04283870976446808
	pesos_i(3859) := b"0000000000000000_0000000000000000_0010011011000011_1101111010111101"; -- 0.15142624016890321
	pesos_i(3860) := b"1111111111111111_1111111111111111_1101101001100100_1101100110101101"; -- -0.14689864664021077
	pesos_i(3861) := b"0000000000000000_0000000000000000_0001110001111111_0000100010101001"; -- 0.11131338235629222
	pesos_i(3862) := b"1111111111111111_1111111111111111_1110000000110001_1011010110011000"; -- -0.12424149556675157
	pesos_i(3863) := b"0000000000000000_0000000000000000_0010001100001010_1100001000010011"; -- 0.13688290555477398
	pesos_i(3864) := b"1111111111111111_1111111111111111_1111000110111011_0011100011111110"; -- -0.05573695948612044
	pesos_i(3865) := b"0000000000000000_0000000000000000_0000111000001011_0110111101100111"; -- 0.054861986769218114
	pesos_i(3866) := b"1111111111111111_1111111111111111_1110011000000000_0010111101000011"; -- -0.10155968307653868
	pesos_i(3867) := b"0000000000000000_0000000000000000_0001100001011100_0011100100110010"; -- 0.09515721770095491
	pesos_i(3868) := b"1111111111111111_1111111111111111_1111001100110100_0001100011000100"; -- -0.049986316812432034
	pesos_i(3869) := b"0000000000000000_0000000000000000_0010101010100000_1001110000000111"; -- 0.16651320609178186
	pesos_i(3870) := b"1111111111111111_1111111111111111_1110110111111111_1110011101101111"; -- -0.07031396418551562
	pesos_i(3871) := b"1111111111111111_1111111111111111_1111001100000010_0100110111110101"; -- -0.050746085728022056
	pesos_i(3872) := b"0000000000000000_0000000000000000_0000001110011011_0011000010001111"; -- 0.014086756510398396
	pesos_i(3873) := b"1111111111111111_1111111111111111_1101110000011011_1110000101011011"; -- -0.14019958057552764
	pesos_i(3874) := b"0000000000000000_0000000000000000_0010100000101011_1011000111101001"; -- 0.15691673209090914
	pesos_i(3875) := b"0000000000000000_0000000000000000_0001011001101100_1010010100101010"; -- 0.08759529379432253
	pesos_i(3876) := b"0000000000000000_0000000000000000_0001100011101000_1101110111100101"; -- 0.09730326501283436
	pesos_i(3877) := b"1111111111111111_1111111111111111_1110110110111111_1011100100101101"; -- -0.07129328402429869
	pesos_i(3878) := b"1111111111111111_1111111111111111_1111011000110010_0111000000110011"; -- -0.03829287295008024
	pesos_i(3879) := b"1111111111111111_1111111111111111_1110010100100110_0000011110100100"; -- -0.10488846067915353
	pesos_i(3880) := b"1111111111111111_1111111111111111_1110011010110001_0011101101011011"; -- -0.09885815639507275
	pesos_i(3881) := b"1111111111111111_1111111111111111_1101110011100101_1000100100010111"; -- -0.1371225660395859
	pesos_i(3882) := b"0000000000000000_0000000000000000_0000100100110100_0001100111011101"; -- 0.03595124857891489
	pesos_i(3883) := b"0000000000000000_0000000000000000_0001101001000101_1101111011100001"; -- 0.10262864102009109
	pesos_i(3884) := b"1111111111111111_1111111111111111_1110000001110101_0101100011110111"; -- -0.12320941905997694
	pesos_i(3885) := b"0000000000000000_0000000000000000_0010001111001001_1010110111111110"; -- 0.1397961372526705
	pesos_i(3886) := b"0000000000000000_0000000000000000_0000111001100011_0110000011010101"; -- 0.056203891752033004
	pesos_i(3887) := b"0000000000000000_0000000000000000_0001011101100101_1110111001111111"; -- 0.09139910323203508
	pesos_i(3888) := b"0000000000000000_0000000000000000_0000110010011111_1111011101110000"; -- 0.04931589578246012
	pesos_i(3889) := b"1111111111111111_1111111111111111_1101111000110010_1000110110011001"; -- -0.13204112061197962
	pesos_i(3890) := b"1111111111111111_1111111111111111_1111000001000100_0011011110100011"; -- -0.06145908609472168
	pesos_i(3891) := b"0000000000000000_0000000000000000_0001101111010100_0100011100011100"; -- 0.1087078516702922
	pesos_i(3892) := b"1111111111111111_1111111111111111_1101010101100110_0010010000010100"; -- -0.1664102032037121
	pesos_i(3893) := b"0000000000000000_0000000000000000_0001101001111011_1100111111010001"; -- 0.10345171784379824
	pesos_i(3894) := b"1111111111111111_1111111111111111_1111100000010011_0011011011110101"; -- -0.03095680738084414
	pesos_i(3895) := b"1111111111111111_1111111111111111_1111111010100111_1111010000011000"; -- -0.0052497332161208525
	pesos_i(3896) := b"0000000000000000_0000000000000000_0000011101000000_1100011001011000"; -- 0.02833213469496143
	pesos_i(3897) := b"1111111111111111_1111111111111111_1111111101001011_1101010010111101"; -- -0.002749160547172643
	pesos_i(3898) := b"0000000000000000_0000000000000000_0001000101101111_1101001101110000"; -- 0.06811257813645422
	pesos_i(3899) := b"0000000000000000_0000000000000000_0000001011001001_1111111101111111"; -- 0.01089474542306722
	pesos_i(3900) := b"1111111111111111_1111111111111111_1111110110001011_0000110011100001"; -- -0.009597010705826164
	pesos_i(3901) := b"1111111111111111_1111111111111111_1110100101000110_1010111001101100"; -- -0.08876523839434568
	pesos_i(3902) := b"1111111111111111_1111111111111111_1110101000000000_1000010001111010"; -- -0.08592960386358954
	pesos_i(3903) := b"1111111111111111_1111111111111111_1110000000110110_0001010101011101"; -- -0.12417475214393561
	pesos_i(3904) := b"0000000000000000_0000000000000000_0000010010000101_0010110010110010"; -- 0.017657082969675802
	pesos_i(3905) := b"1111111111111111_1111111111111111_1101111100000001_0011101110011001"; -- -0.12888743884693435
	pesos_i(3906) := b"0000000000000000_0000000000000000_0001010100100011_0101010010110101"; -- 0.08257035660838276
	pesos_i(3907) := b"0000000000000000_0000000000000000_0010000011111000_1100111000011110"; -- 0.12879646522144336
	pesos_i(3908) := b"0000000000000000_0000000000000000_0001111001011000_0101011110010001"; -- 0.11853549291125079
	pesos_i(3909) := b"0000000000000000_0000000000000000_0001011010111000_1110111010001101"; -- 0.08875933593952719
	pesos_i(3910) := b"0000000000000000_0000000000000000_0011000111010111_0100111000111001"; -- 0.1946915521791288
	pesos_i(3911) := b"0000000000000000_0000000000000000_0000000101001000_0010100000110100"; -- 0.00500727919190757
	pesos_i(3912) := b"1111111111111111_1111111111111111_1111000000110111_1000100111101101"; -- -0.06165254565666456
	pesos_i(3913) := b"0000000000000000_0000000000000000_0010100001000011_1001011111011000"; -- 0.15728138956318413
	pesos_i(3914) := b"1111111111111111_1111111111111111_1111111000000100_0110100110111111"; -- -0.0077451617761768645
	pesos_i(3915) := b"1111111111111111_1111111111111111_1111100001010111_1011111111100110"; -- -0.029911047303819483
	pesos_i(3916) := b"0000000000000000_0000000000000000_0001100111101010_1010111101001111"; -- 0.10123725591678272
	pesos_i(3917) := b"1111111111111111_1111111111111111_1110100000011111_0111101110100010"; -- -0.09326960848824824
	pesos_i(3918) := b"1111111111111111_1111111111111111_1110010100111000_0000111000100101"; -- -0.10461341462493316
	pesos_i(3919) := b"1111111111111111_1111111111111111_1111101000111000_1101111111010010"; -- -0.02256966716235517
	pesos_i(3920) := b"1111111111111111_1111111111111111_1110110011001001_1100100010100001"; -- -0.07504602502370841
	pesos_i(3921) := b"1111111111111111_1111111111111111_1110010011001101_1000011111100111"; -- -0.10623884775532995
	pesos_i(3922) := b"0000000000000000_0000000000000000_0001011000000011_1011101011001000"; -- 0.08599440935880996
	pesos_i(3923) := b"0000000000000000_0000000000000000_0000100000101100_1011110111111111"; -- 0.03193271144099888
	pesos_i(3924) := b"0000000000000000_0000000000000000_0010011011011011_0011000101101111"; -- 0.15178212116404008
	pesos_i(3925) := b"0000000000000000_0000000000000000_0010010011010101_0111000010010100"; -- 0.14388183226362877
	pesos_i(3926) := b"0000000000000000_0000000000000000_0010101100011110_1011001011000100"; -- 0.16843716901312364
	pesos_i(3927) := b"0000000000000000_0000000000000000_0011011001001111_0011110000111010"; -- 0.21214653419800744
	pesos_i(3928) := b"0000000000000000_0000000000000000_0000110010010000_1000001101101110"; -- 0.049080099503606506
	pesos_i(3929) := b"0000000000000000_0000000000000000_0001000111010111_0011110100001101"; -- 0.06969052860332588
	pesos_i(3930) := b"1111111111111111_1111111111111111_1110010001101001_0110110011111111"; -- -0.10776633036530418
	pesos_i(3931) := b"0000000000000000_0000000000000000_0000111001010011_1101110011011110"; -- 0.05596714418781857
	pesos_i(3932) := b"1111111111111111_1111111111111111_1111000010101010_1100110101100101"; -- -0.05989376348945504
	pesos_i(3933) := b"0000000000000000_0000000000000000_0000000001111010_1110111101100110"; -- 0.0018758414397102249
	pesos_i(3934) := b"0000000000000000_0000000000000000_0001000111011001_1101010100000100"; -- 0.0697301039492905
	pesos_i(3935) := b"1111111111111111_1111111111111111_1110110101001110_0110010001111101"; -- -0.07302257495479152
	pesos_i(3936) := b"0000000000000000_0000000000000000_0010000010010111_1000110000001011"; -- 0.12731242432870285
	pesos_i(3937) := b"1111111111111111_1111111111111111_1101110110000110_1101011111010010"; -- -0.1346612083950401
	pesos_i(3938) := b"1111111111111111_1111111111111111_1110110100011110_0010110010100000"; -- -0.0737583264484874
	pesos_i(3939) := b"1111111111111111_1111111111111111_1111001001001110_0101100001001010"; -- -0.05349205207919153
	pesos_i(3940) := b"0000000000000000_0000000000000000_0001001001010010_1011001111110001"; -- 0.07157444609928817
	pesos_i(3941) := b"1111111111111111_1111111111111111_1110001001110011_0111000110010001"; -- -0.11542597006181303
	pesos_i(3942) := b"0000000000000000_0000000000000000_0010000011001100_1101100110010011"; -- 0.12812576128646036
	pesos_i(3943) := b"1111111111111111_1111111111111111_1101111111110010_1100100010110000"; -- -0.12520166110059466
	pesos_i(3944) := b"0000000000000000_0000000000000000_0000000011000110_1101001001010110"; -- 0.0030337771471787567
	pesos_i(3945) := b"0000000000000000_0000000000000000_0000110110101111_1110100001101000"; -- 0.05346539057699166
	pesos_i(3946) := b"0000000000000000_0000000000000000_0001101111000111_1111011110011000"; -- 0.10852000677668239
	pesos_i(3947) := b"1111111111111111_1111111111111111_1110101101100110_1000010101111101"; -- -0.08046689692099666
	pesos_i(3948) := b"1111111111111111_1111111111111111_1101111010000010_1111100000000110"; -- -0.1308140741374903
	pesos_i(3949) := b"0000000000000000_0000000000000000_0000111001111011_0110011101111011"; -- 0.056570499031202315
	pesos_i(3950) := b"0000000000000000_0000000000000000_0000110100010001_0110101011111111"; -- 0.05104702682919691
	pesos_i(3951) := b"0000000000000000_0000000000000000_0001001110000101_0000110010110000"; -- 0.07624892517403163
	pesos_i(3952) := b"1111111111111111_1111111111111111_1101011010111101_1000100000110100"; -- -0.1611704705084123
	pesos_i(3953) := b"1111111111111111_1111111111111111_1110101000010110_0001101001000100"; -- -0.08560024117635036
	pesos_i(3954) := b"0000000000000000_0000000000000000_0000110110101101_0000111001110010"; -- 0.053421881555513445
	pesos_i(3955) := b"0000000000000000_0000000000000000_0000001101001011_0111100011000100"; -- 0.012870357267317382
	pesos_i(3956) := b"1111111111111111_1111111111111111_1101111101011100_1011000010110111"; -- -0.1274919084717092
	pesos_i(3957) := b"1111111111111111_1111111111111111_1110101111100101_0100000100101111"; -- -0.07853310202844246
	pesos_i(3958) := b"0000000000000000_0000000000000000_0001110111010000_1000101001011011"; -- 0.11646332466115455
	pesos_i(3959) := b"1111111111111111_1111111111111111_1101010000101010_1100000001101111"; -- -0.17122266093022984
	pesos_i(3960) := b"0000000000000000_0000000000000000_0000110011000101_1100011100100111"; -- 0.04989285196522375
	pesos_i(3961) := b"1111111111111111_1111111111111111_1101111111000111_0111101000011110"; -- -0.12586247215517546
	pesos_i(3962) := b"0000000000000000_0000000000000000_0000111111000111_0100001100000010"; -- 0.0616342430656891
	pesos_i(3963) := b"1111111111111111_1111111111111111_1101110011100001_1110001110010110"; -- -0.1371782072229682
	pesos_i(3964) := b"0000000000000000_0000000000000000_0001110100000010_0000011011111111"; -- 0.11331218452803006
	pesos_i(3965) := b"1111111111111111_1111111111111111_1101100001010000_1110001110000001"; -- -0.1550157365788449
	pesos_i(3966) := b"1111111111111111_1111111111111111_1101011111111110_0011110111101101"; -- -0.15627682656572925
	pesos_i(3967) := b"0000000000000000_0000000000000000_0000010111110111_1001001100011000"; -- 0.023308938324598474
	pesos_i(3968) := b"0000000000000000_0000000000000000_0001011111110101_1011111010011111"; -- 0.09359351523570295
	pesos_i(3969) := b"0000000000000000_0000000000000000_0011001010010001_1010000110101101"; -- 0.19753466094605301
	pesos_i(3970) := b"0000000000000000_0000000000000000_0001011010011110_1101010110001101"; -- 0.08836111730177579
	pesos_i(3971) := b"0000000000000000_0000000000000000_0010000000010111_1100110001001100"; -- 0.1253631291398008
	pesos_i(3972) := b"0000000000000000_0000000000000000_0010100001001100_1100000001011000"; -- 0.15742113249075226
	pesos_i(3973) := b"1111111111111111_1111111111111111_1111000101110000_0111010110100100"; -- -0.056877753619723775
	pesos_i(3974) := b"0000000000000000_0000000000000000_0001010001101001_0100100100101111"; -- 0.07973153488108697
	pesos_i(3975) := b"1111111111111111_1111111111111111_1111100010111010_1100001001010101"; -- -0.02840028221676804
	pesos_i(3976) := b"1111111111111111_1111111111111111_1110011101101101_1010010010101011"; -- -0.09598322692926263
	pesos_i(3977) := b"1111111111111111_1111111111111111_1101110001101101_1010010000000111"; -- -0.1389520151780506
	pesos_i(3978) := b"1111111111111111_1111111111111111_1111010111110111_0000000110001101"; -- -0.039199736746531016
	pesos_i(3979) := b"0000000000000000_0000000000000000_0000111100100111_0011010011100101"; -- 0.059191995633166065
	pesos_i(3980) := b"0000000000000000_0000000000000000_0001100101101101_1001011001101000"; -- 0.09932842294620908
	pesos_i(3981) := b"0000000000000000_0000000000000000_0010111000011111_0000100101000111"; -- 0.18016107548545562
	pesos_i(3982) := b"1111111111111111_1111111111111111_1111110010110000_0010011110000011"; -- -0.01293709802028404
	pesos_i(3983) := b"1111111111111111_1111111111111111_1110101111000011_1001101111001101"; -- -0.07904649978149525
	pesos_i(3984) := b"1111111111111111_1111111111111111_1101111001011010_0111111111000101"; -- -0.13143159334711987
	pesos_i(3985) := b"0000000000000000_0000000000000000_0000100101010101_1100100101110111"; -- 0.03646525541306484
	pesos_i(3986) := b"0000000000000000_0000000000000000_0000101000001110_0101010100101000"; -- 0.03928119867562835
	pesos_i(3987) := b"0000000000000000_0000000000000000_0001001001100100_0000001000000100"; -- 0.07183849899254627
	pesos_i(3988) := b"0000000000000000_0000000000000000_0001110101011111_0111010011101101"; -- 0.11473780433580727
	pesos_i(3989) := b"0000000000000000_0000000000000000_0010011010101010_0110001100111101"; -- 0.1510374091374901
	pesos_i(3990) := b"1111111111111111_1111111111111111_1111110100001001_1110010110000011"; -- -0.011567740878727086
	pesos_i(3991) := b"0000000000000000_0000000000000000_0001010111100110_0001000001111110"; -- 0.08554175449851069
	pesos_i(3992) := b"0000000000000000_0000000000000000_0010001011111011_1101110110011011"; -- 0.13665566468330684
	pesos_i(3993) := b"1111111111111111_1111111111111111_1111001110110001_1111101110001110"; -- -0.048065450488810724
	pesos_i(3994) := b"1111111111111111_1111111111111111_1110011111101110_0100010101001100"; -- -0.09402052768202605
	pesos_i(3995) := b"1111111111111111_1111111111111111_1101111011000001_1101100011001100"; -- -0.12985463164908242
	pesos_i(3996) := b"0000000000000000_0000000000000000_0000000100101101_1011110011000010"; -- 0.00460414642792646
	pesos_i(3997) := b"1111111111111111_1111111111111111_1101010101100100_0111011000100100"; -- -0.1664358294298727
	pesos_i(3998) := b"1111111111111111_1111111111111111_1110100111010100_1001110010110111"; -- -0.08659954578233214
	pesos_i(3999) := b"1111111111111111_1111111111111111_1111110100111110_1010110011000001"; -- -0.010762408076698815
	pesos_i(4000) := b"1111111111111111_1111111111111111_1101001101111111_0111110110111010"; -- -0.1738358898407172
	pesos_i(4001) := b"0000000000000000_0000000000000000_0001101100101111_0001001011101100"; -- 0.10618704099012156
	pesos_i(4002) := b"0000000000000000_0000000000000000_0010110000000011_1011110000011000"; -- 0.17193198757273218
	pesos_i(4003) := b"1111111111111111_1111111111111111_1101111011110110_0110101011101010"; -- -0.12905246530545772
	pesos_i(4004) := b"0000000000000000_0000000000000000_0001000101011011_1101001011110110"; -- 0.06780737409025099
	pesos_i(4005) := b"1111111111111111_1111111111111111_1110001100111110_1100000000000101"; -- -0.11232375972162299
	pesos_i(4006) := b"0000000000000000_0000000000000000_0000010001110000_1101010010110001"; -- 0.01734666167592165
	pesos_i(4007) := b"0000000000000000_0000000000000000_0001100011001010_1101000100101111"; -- 0.09684474362544629
	pesos_i(4008) := b"1111111111111111_1111111111111111_1101111100001111_1000101101010010"; -- -0.12866906413847606
	pesos_i(4009) := b"0000000000000000_0000000000000000_0000111111000101_0110111111110100"; -- 0.06160640448475139
	pesos_i(4010) := b"1111111111111111_1111111111111111_1110111000100000_0011111101000111"; -- -0.06982044702395686
	pesos_i(4011) := b"0000000000000000_0000000000000000_0010100111101011_1100101111111101"; -- 0.1637542241813606
	pesos_i(4012) := b"1111111111111111_1111111111111111_1110110001010001_1101011010110000"; -- -0.07687624168197844
	pesos_i(4013) := b"1111111111111111_1111111111111111_1101101111001001_0011110111000011"; -- -0.14146055213708467
	pesos_i(4014) := b"0000000000000000_0000000000000000_0001001101010101_1010101000111110"; -- 0.07552589426667429
	pesos_i(4015) := b"0000000000000000_0000000000000000_0000110100011011_0100100100100100"; -- 0.051197596821704515
	pesos_i(4016) := b"1111111111111111_1111111111111111_1101100110000101_0010101100111100"; -- -0.15031175412560552
	pesos_i(4017) := b"0000000000000000_0000000000000000_0001111010110111_0111100010000100"; -- 0.11998704178289131
	pesos_i(4018) := b"1111111111111111_1111111111111111_1110010111001000_1100000001000100"; -- -0.10240553223847733
	pesos_i(4019) := b"1111111111111111_1111111111111111_1110001100001010_1101011110111100"; -- -0.11311580331197506
	pesos_i(4020) := b"0000000000000000_0000000000000000_0000101001011111_1101100011001001"; -- 0.040525006290989804
	pesos_i(4021) := b"1111111111111111_1111111111111111_1111010111011010_1100010110110110"; -- -0.03963054959849357
	pesos_i(4022) := b"1111111111111111_1111111111111111_1110010111101001_0111001000100101"; -- -0.10190664856402203
	pesos_i(4023) := b"1111111111111111_1111111111111111_1101100111101000_1111000011000100"; -- -0.1487893602733674
	pesos_i(4024) := b"1111111111111111_1111111111111111_1111010111100111_1101001110001111"; -- -0.03943135984542567
	pesos_i(4025) := b"0000000000000000_0000000000000000_0000111001010001_0110110110111010"; -- 0.055930002114418405
	pesos_i(4026) := b"1111111111111111_1111111111111111_1101010100011110_0011011111000000"; -- -0.16750766329526837
	pesos_i(4027) := b"1111111111111111_1111111111111111_1111010001000010_0101010000000000"; -- -0.04586291320000522
	pesos_i(4028) := b"1111111111111111_1111111111111111_1101001111001101_0010001000000001"; -- -0.17265117153472706
	pesos_i(4029) := b"0000000000000000_0000000000000000_0010101101000100_1011101000101000"; -- 0.1690174434973309
	pesos_i(4030) := b"0000000000000000_0000000000000000_0000111011001110_1011111110111010"; -- 0.0578422384039884
	pesos_i(4031) := b"0000000000000000_0000000000000000_0000000111010011_0010001110011010"; -- 0.007127976474409874
	pesos_i(4032) := b"1111111111111111_1111111111111111_1101001110001110_0110100100010010"; -- -0.1736082392610771
	pesos_i(4033) := b"0000000000000000_0000000000000000_0001111011000000_0101011000110010"; -- 0.12012232515647392
	pesos_i(4034) := b"1111111111111111_1111111111111111_1110001100011101_0100110111100011"; -- -0.11283410278655523
	pesos_i(4035) := b"1111111111111111_1111111111111111_1101010011000000_1000101101101011"; -- -0.16893700264646386
	pesos_i(4036) := b"1111111111111111_1111111111111111_1110001101010010_1101100010010001"; -- -0.11201712095358547
	pesos_i(4037) := b"0000000000000000_0000000000000000_0001011010010000_0010010011001001"; -- 0.08813695823993342
	pesos_i(4038) := b"1111111111111111_1111111111111111_1111100100001011_0100111100010000"; -- -0.02717119084279127
	pesos_i(4039) := b"0000000000000000_0000000000000000_0001001001110110_0100001101011110"; -- 0.07211705259444084
	pesos_i(4040) := b"0000000000000000_0000000000000000_0000010011010000_0000111100100110"; -- 0.018799731132637092
	pesos_i(4041) := b"0000000000000000_0000000000000000_0000000100110101_1001011111111000"; -- 0.004724023865228633
	pesos_i(4042) := b"0000000000000000_0000000000000000_0001101100011101_0000001011001011"; -- 0.10591142132604503
	pesos_i(4043) := b"1111111111111111_1111111111111111_1101101010111100_1100101010100110"; -- -0.14555676884203556
	pesos_i(4044) := b"1111111111111111_1111111111111111_1110101101000100_1001010101011110"; -- -0.08098474933628318
	pesos_i(4045) := b"1111111111111111_1111111111111111_1111011111011001_1110110000000100"; -- -0.03183102521311638
	pesos_i(4046) := b"0000000000000000_0000000000000000_0010010011100111_0111111110111000"; -- 0.1441573928413776
	pesos_i(4047) := b"0000000000000000_0000000000000000_0000001111100011_1110011010110011"; -- 0.015196245969192081
	pesos_i(4048) := b"0000000000000000_0000000000000000_0010001001011111_0100111110000010"; -- 0.13426682399798737
	pesos_i(4049) := b"0000000000000000_0000000000000000_0010111000010000_1001110001100100"; -- 0.17994096222708586
	pesos_i(4050) := b"1111111111111111_1111111111111111_1101010100010100_1011011101011011"; -- -0.16765264541486105
	pesos_i(4051) := b"1111111111111111_1111111111111111_1101110000100111_0000101101000010"; -- -0.14002923615924553
	pesos_i(4052) := b"0000000000000000_0000000000000000_0000100101001101_0100111011110000"; -- 0.03633588183050843
	pesos_i(4053) := b"0000000000000000_0000000000000000_0000100001011010_0010111101111101"; -- 0.03262612147324428
	pesos_i(4054) := b"0000000000000000_0000000000000000_0001000011011000_1101011001100010"; -- 0.06580867658688301
	pesos_i(4055) := b"0000000000000000_0000000000000000_0000011000100001_0001110100000010"; -- 0.02394276909334498
	pesos_i(4056) := b"0000000000000000_0000000000000000_0000100101110101_1111111100000010"; -- 0.03695672803513313
	pesos_i(4057) := b"1111111111111111_1111111111111111_1111110101110011_1101101001010010"; -- -0.009950976258332798
	pesos_i(4058) := b"1111111111111111_1111111111111111_1110110000110000_1000001011100010"; -- -0.07738477699261534
	pesos_i(4059) := b"0000000000000000_0000000000000000_0010001011101011_1100011001110011"; -- 0.13641014386533343
	pesos_i(4060) := b"1111111111111111_1111111111111111_1101101000011000_0000101001001000"; -- -0.14807067630840348
	pesos_i(4061) := b"0000000000000000_0000000000000000_0000010010110100_0000000101000011"; -- 0.018371657316491898
	pesos_i(4062) := b"1111111111111111_1111111111111111_1101000110100010_0010011110101010"; -- -0.1811194620355277
	pesos_i(4063) := b"1111111111111111_1111111111111111_1110011110100001_0011010101010100"; -- -0.09519640637478874
	pesos_i(4064) := b"1111111111111111_1111111111111111_1110010100011011_1101111010010011"; -- -0.10504349633276044
	pesos_i(4065) := b"1111111111111111_1111111111111111_1111001010010000_0110000000001111"; -- -0.05248450876295946
	pesos_i(4066) := b"1111111111111111_1111111111111111_1110100001110110_1101000110111111"; -- -0.09193696100502315
	pesos_i(4067) := b"0000000000000000_0000000000000000_0001101000111111_1111111000010000"; -- 0.10253894694006335
	pesos_i(4068) := b"1111111111111111_1111111111111111_1110100001000001_1111001011101100"; -- -0.0927436994668215
	pesos_i(4069) := b"0000000000000000_0000000000000000_0000100111100001_1001101010101110"; -- 0.03859869709333215
	pesos_i(4070) := b"1111111111111111_1111111111111111_1111001001001111_1101100101001011"; -- -0.05346910399440965
	pesos_i(4071) := b"1111111111111111_1111111111111111_1101011111000110_1100001010101001"; -- -0.15712340704295935
	pesos_i(4072) := b"1111111111111111_1111111111111111_1101001110010101_1011100111100010"; -- -0.1734966109601313
	pesos_i(4073) := b"1111111111111111_1111111111111111_1111100010111001_0010011010001101"; -- -0.028424826266266592
	pesos_i(4074) := b"0000000000000000_0000000000000000_0000110101001110_1011010001010010"; -- 0.05198218348485722
	pesos_i(4075) := b"0000000000000000_0000000000000000_0000101001111110_1000100000110100"; -- 0.040993225719870005
	pesos_i(4076) := b"0000000000000000_0000000000000000_0010000110000010_0100000101100110"; -- 0.13089379073800994
	pesos_i(4077) := b"1111111111111111_1111111111111111_1110101100000001_1110110011100111"; -- -0.08200187075668142
	pesos_i(4078) := b"0000000000000000_0000000000000000_0010011101011011_0010100010001011"; -- 0.1537347163025036
	pesos_i(4079) := b"1111111111111111_1111111111111111_1110110001011011_0100101011000000"; -- -0.07673199474411194
	pesos_i(4080) := b"0000000000000000_0000000000000000_0000100000011000_0101001011100010"; -- 0.03162115107018615
	pesos_i(4081) := b"1111111111111111_1111111111111111_1110101110000011_1100100100101101"; -- -0.08002035757518537
	pesos_i(4082) := b"0000000000000000_0000000000000000_0000111010010101_1001000101011011"; -- 0.056969723376917705
	pesos_i(4083) := b"1111111111111111_1111111111111111_1111011011101101_0101010100011111"; -- -0.035441093411895
	pesos_i(4084) := b"1111111111111111_1111111111111111_1111011001110110_1001101111000111"; -- -0.037252677935712394
	pesos_i(4085) := b"1111111111111111_1111111111111111_1111101110111111_0110110011001110"; -- -0.016610335921833384
	pesos_i(4086) := b"0000000000000000_0000000000000000_0000110010100011_1001101001001100"; -- 0.04937137943676177
	pesos_i(4087) := b"0000000000000000_0000000000000000_0001001111110111_0010010010001010"; -- 0.07798984882755917
	pesos_i(4088) := b"0000000000000000_0000000000000000_0010000010010101_0111010111111110"; -- 0.12728059236898834
	pesos_i(4089) := b"1111111111111111_1111111111111111_1101110000000110_1011100111100111"; -- -0.1405223666749926
	pesos_i(4090) := b"0000000000000000_0000000000000000_0010011100000110_1101010001000100"; -- 0.15244795477999654
	pesos_i(4091) := b"0000000000000000_0000000000000000_0001010100110010_0001000110000001"; -- 0.08279523269498712
	pesos_i(4092) := b"0000000000000000_0000000000000000_0000111101110011_1001100111110101"; -- 0.06035768732933884
	pesos_i(4093) := b"0000000000000000_0000000000000000_0010101011111101_0000111010001000"; -- 0.1679238397408533
	pesos_i(4094) := b"1111111111111111_1111111111111111_1111011110111110_1111111111001010"; -- -0.03224183395135335
	pesos_i(4095) := b"1111111111111111_1111111111111111_1101111000010110_0001111101101110"; -- -0.13247493334522617
	pesos_i(4096) := b"1111111111111111_1111111111111111_1111001001010001_1101111011000001"; -- -0.05343826101898069
	pesos_i(4097) := b"1111111111111111_1111111111111111_1111111000100000_0111111010101110"; -- -0.007316668047729192
	pesos_i(4098) := b"0000000000000000_0000000000000000_0010101110110110_0001010100000111"; -- 0.17074710287225345
	pesos_i(4099) := b"0000000000000000_0000000000000000_0000001100111100_1111000101111011"; -- 0.012648670700597102
	pesos_i(4100) := b"0000000000000000_0000000000000000_0001100010101011_0000111110110011"; -- 0.09636018859929063
	pesos_i(4101) := b"0000000000000000_0000000000000000_0001100111000110_0010110011100101"; -- 0.10068016620638916
	pesos_i(4102) := b"1111111111111111_1111111111111111_1111010011001111_1001100111011000"; -- -0.04370726074836702
	pesos_i(4103) := b"1111111111111111_1111111111111111_1111001001001111_0110101000100010"; -- -0.05347572973733664
	pesos_i(4104) := b"0000000000000000_0000000000000000_0001010011111100_0000011001010100"; -- 0.08197059200186708
	pesos_i(4105) := b"1111111111111111_1111111111111111_1110110011110001_0001001101001111"; -- -0.07444648103735331
	pesos_i(4106) := b"1111111111111111_1111111111111111_1111000001110011_0100000111111111"; -- -0.06074130554657592
	pesos_i(4107) := b"0000000000000000_0000000000000000_0000110010101111_1100111001001001"; -- 0.049557583530656854
	pesos_i(4108) := b"0000000000000000_0000000000000000_0010011101010000_1111001100111100"; -- 0.15357895108975314
	pesos_i(4109) := b"1111111111111111_1111111111111111_1111000010110111_0001111000000110"; -- -0.05970585213887934
	pesos_i(4110) := b"1111111111111111_1111111111111111_1110010001010011_0111100010001010"; -- -0.10810133581666574
	pesos_i(4111) := b"0000000000000000_0000000000000000_0001010011001011_0100000101011110"; -- 0.08122643032878894
	pesos_i(4112) := b"1111111111111111_1111111111111111_1110110110000000_0010000100110000"; -- -0.07226364692951918
	pesos_i(4113) := b"1111111111111111_1111111111111111_1101111010011001_1010011011101111"; -- -0.1304679551476232
	pesos_i(4114) := b"0000000000000000_0000000000000000_0001110001001000_0001100011001101"; -- 0.11047511111530559
	pesos_i(4115) := b"0000000000000000_0000000000000000_0001100000001101_1111001100000001"; -- 0.09396284839487705
	pesos_i(4116) := b"1111111111111111_1111111111111111_1110100101110110_0111100110110111"; -- -0.08803595805978694
	pesos_i(4117) := b"0000000000000000_0000000000000000_0001001010111000_0111100100011100"; -- 0.07312733581852944
	pesos_i(4118) := b"1111111111111111_1111111111111111_1110001010110111_1010000101000100"; -- -0.11438552943543635
	pesos_i(4119) := b"1111111111111111_1111111111111111_1111011110111010_0100001101011000"; -- -0.03231410114620415
	pesos_i(4120) := b"0000000000000000_0000000000000000_0000000000001000_0100111100111000"; -- 0.00012679222646219888
	pesos_i(4121) := b"1111111111111111_1111111111111111_1111101000001011_1001001011100011"; -- -0.023260898187620394
	pesos_i(4122) := b"0000000000000000_0000000000000000_0001000100001011_1000110010111100"; -- 0.06658248509105062
	pesos_i(4123) := b"0000000000000000_0000000000000000_0000111001010011_0001011010010100"; -- 0.055955325262541225
	pesos_i(4124) := b"1111111111111111_1111111111111111_1110001111011000_0100000111000101"; -- -0.1099814313930244
	pesos_i(4125) := b"0000000000000000_0000000000000000_0001000111110010_1111101010011010"; -- 0.07011381407211977
	pesos_i(4126) := b"1111111111111111_1111111111111111_1111100001101010_0001100010111011"; -- -0.029631094371180687
	pesos_i(4127) := b"1111111111111111_1111111111111111_1110100010100100_0011100100110010"; -- -0.09124414957921825
	pesos_i(4128) := b"1111111111111111_1111111111111111_1111110111001001_1100100100000011"; -- -0.008639752132469591
	pesos_i(4129) := b"1111111111111111_1111111111111111_1101011000100100_1001001010100101"; -- -0.16350444282961304
	pesos_i(4130) := b"0000000000000000_0000000000000000_0001000011000000_0001101111010100"; -- 0.06543134607635873
	pesos_i(4131) := b"0000000000000000_0000000000000000_0000100110001110_1101111100001001"; -- 0.03733629208271382
	pesos_i(4132) := b"1111111111111111_1111111111111111_1111100010010110_0101010000101110"; -- -0.028956164211497343
	pesos_i(4133) := b"1111111111111111_1111111111111111_1111000111110100_1101000100011101"; -- -0.05485814132505463
	pesos_i(4134) := b"0000000000000000_0000000000000000_0010010010110000_1111000110100101"; -- 0.14332495002524892
	pesos_i(4135) := b"1111111111111111_1111111111111111_1111110100101110_1011011101110101"; -- -0.011005910802600077
	pesos_i(4136) := b"1111111111111111_1111111111111111_1111110000110010_0011000101001111"; -- -0.014859121543753573
	pesos_i(4137) := b"0000000000000000_0000000000000000_0001011011000110_1110011000000010"; -- 0.08897244979643695
	pesos_i(4138) := b"0000000000000000_0000000000000000_0000000011001011_0111011010001100"; -- 0.0031046000209347903
	pesos_i(4139) := b"0000000000000000_0000000000000000_0000101011101011_0000100101000010"; -- 0.04264886718097806
	pesos_i(4140) := b"0000000000000000_0000000000000000_0010010011111000_1011010001010001"; -- 0.1444199274027844
	pesos_i(4141) := b"0000000000000000_0000000000000000_0001101011101000_1111001110111100"; -- 0.10511706676666223
	pesos_i(4142) := b"1111111111111111_1111111111111111_1110001001001101_1111100000100010"; -- -0.11599778328617164
	pesos_i(4143) := b"1111111111111111_1111111111111111_1100110111000110_1110101001100110"; -- -0.19618353847031636
	pesos_i(4144) := b"0000000000000000_0000000000000000_0001011111101001_1000100000000111"; -- 0.09340715567033828
	pesos_i(4145) := b"1111111111111111_1111111111111111_1110010111111011_1100101001000101"; -- -0.10162673778733912
	pesos_i(4146) := b"0000000000000000_0000000000000000_0001001001011111_1011101101011001"; -- 0.07177325168110611
	pesos_i(4147) := b"0000000000000000_0000000000000000_0001100001100100_0111101011111000"; -- 0.09528320849237142
	pesos_i(4148) := b"1111111111111111_1111111111111111_1110101110101011_1100100111000111"; -- -0.07940997014333502
	pesos_i(4149) := b"0000000000000000_0000000000000000_0001010100001001_1111010011000110"; -- 0.08218316882870998
	pesos_i(4150) := b"1111111111111111_1111111111111111_1110101010000010_0100010111110101"; -- -0.08394968761238153
	pesos_i(4151) := b"0000000000000000_0000000000000000_0000010100101101_0110111001110011"; -- 0.020224478848428463
	pesos_i(4152) := b"1111111111111111_1111111111111111_1101001011001101_0011001011010000"; -- -0.17655641954439805
	pesos_i(4153) := b"1111111111111111_1111111111111111_1110000000101001_1011001111101100"; -- -0.12436366538089651
	pesos_i(4154) := b"1111111111111111_1111111111111111_1111100000101000_0101100101001000"; -- -0.030634326817627917
	pesos_i(4155) := b"1111111111111111_1111111111111111_1101010011101111_0101000111101011"; -- -0.16822326664119863
	pesos_i(4156) := b"0000000000000000_0000000000000000_0000100000100100_1101101101110011"; -- 0.03181239664675819
	pesos_i(4157) := b"1111111111111111_1111111111111111_1110110011101000_1110110111100011"; -- -0.07457078181882719
	pesos_i(4158) := b"0000000000000000_0000000000000000_0001101001011110_0000111000010000"; -- 0.10299766425227136
	pesos_i(4159) := b"1111111111111111_1111111111111111_1110111111001001_1111110001110010"; -- -0.06332418641133687
	pesos_i(4160) := b"0000000000000000_0000000000000000_0000101010000000_1000000111110110"; -- 0.041023371186030916
	pesos_i(4161) := b"0000000000000000_0000000000000000_0000111000101011_0101010101111000"; -- 0.055348722222586286
	pesos_i(4162) := b"1111111111111111_1111111111111111_1111111001100111_0101101101000000"; -- -0.006235405824499738
	pesos_i(4163) := b"1111111111111111_1111111111111111_1110000111010111_1101011000010011"; -- -0.11780035060027338
	pesos_i(4164) := b"1111111111111111_1111111111111111_1101110100011010_1010001111010000"; -- -0.13631225759044674
	pesos_i(4165) := b"0000000000000000_0000000000000000_0000111110010001_1101000011011010"; -- 0.06081872287233677
	pesos_i(4166) := b"1111111111111111_1111111111111111_1101101111010101_1000100101011100"; -- -0.14127294062856946
	pesos_i(4167) := b"0000000000000000_0000000000000000_0000010000011111_0011011000000001"; -- 0.016101241277387733
	pesos_i(4168) := b"0000000000000000_0000000000000000_0000001000100101_0001000010111101"; -- 0.008378072897234674
	pesos_i(4169) := b"1111111111111111_1111111111111111_1111011110100000_1110000101011000"; -- -0.032701412131747244
	pesos_i(4170) := b"0000000000000000_0000000000000000_0001110010111001_1101111111000110"; -- 0.11221121397016555
	pesos_i(4171) := b"1111111111111111_1111111111111111_1110001001001010_0000111101001010"; -- -0.11605743820127198
	pesos_i(4172) := b"1111111111111111_1111111111111111_1111001111111010_0001011010100100"; -- -0.046965203197591156
	pesos_i(4173) := b"0000000000000000_0000000000000000_0001111000001001_0101010110110011"; -- 0.117329937264755
	pesos_i(4174) := b"1111111111111111_1111111111111111_1110001010100000_0101010111111101"; -- -0.11474096838102119
	pesos_i(4175) := b"1111111111111111_1111111111111111_1110010101000001_1101010011100010"; -- -0.10446424000816827
	pesos_i(4176) := b"0000000000000000_0000000000000000_0001000001100110_0001110100100001"; -- 0.06405813267236513
	pesos_i(4177) := b"1111111111111111_1111111111111111_1101001111101001_0111111111101110"; -- -0.17221832697221515
	pesos_i(4178) := b"0000000000000000_0000000000000000_0000011111001110_1110000001101111"; -- 0.030500437871855548
	pesos_i(4179) := b"0000000000000000_0000000000000000_0010000101001010_1111010100110111"; -- 0.13005001636171945
	pesos_i(4180) := b"0000000000000000_0000000000000000_0010000100100101_0011100000111100"; -- 0.12947417707690578
	pesos_i(4181) := b"1111111111111111_1111111111111111_1111111010000010_1110011110000110"; -- -0.00581505757175316
	pesos_i(4182) := b"0000000000000000_0000000000000000_0010100001100011_0010110111110101"; -- 0.157763359450552
	pesos_i(4183) := b"1111111111111111_1111111111111111_1111010011000110_0010111010010010"; -- -0.04385098400772659
	pesos_i(4184) := b"0000000000000000_0000000000000000_0001001010111110_1010010011000000"; -- 0.07322148990176323
	pesos_i(4185) := b"0000000000000000_0000000000000000_0010011011000010_0110001100011000"; -- 0.1514036114827386
	pesos_i(4186) := b"0000000000000000_0000000000000000_0000110001010101_1010010001101100"; -- 0.04818179732540834
	pesos_i(4187) := b"1111111111111111_1111111111111111_1110000000110001_0100111100000010"; -- -0.12424761009196608
	pesos_i(4188) := b"1111111111111111_1111111111111111_1111100111000101_0110110001111011"; -- -0.024331302672216042
	pesos_i(4189) := b"1111111111111111_1111111111111111_1111101111010110_1011000000110110"; -- -0.016255366062361255
	pesos_i(4190) := b"1111111111111111_1111111111111111_1110101010011001_0111100011111001"; -- -0.08359569479777913
	pesos_i(4191) := b"0000000000000000_0000000000000000_0001011101001111_0100100111010100"; -- 0.09105359487742423
	pesos_i(4192) := b"0000000000000000_0000000000000000_0000111001000100_0001010001010010"; -- 0.0557263088661733
	pesos_i(4193) := b"1111111111111111_1111111111111111_1101101010101100_0110011010000111"; -- -0.1458068772242391
	pesos_i(4194) := b"1111111111111111_1111111111111111_1110000011010101_1101100010101100"; -- -0.12173696328464047
	pesos_i(4195) := b"0000000000000000_0000000000000000_0010100000101000_1000001111100000"; -- 0.15686821189422348
	pesos_i(4196) := b"0000000000000000_0000000000000000_0001110011101011_0101010011011010"; -- 0.11296587288353031
	pesos_i(4197) := b"1111111111111111_1111111111111111_1101010101110000_1000100001000110"; -- -0.16625164302436826
	pesos_i(4198) := b"0000000000000000_0000000000000000_0000010010111110_1101010101110111"; -- 0.01853689350969331
	pesos_i(4199) := b"1111111111111111_1111111111111111_1110110111000000_0111101001111010"; -- -0.07128176232148255
	pesos_i(4200) := b"1111111111111111_1111111111111111_1111001110011011_0100011010001010"; -- -0.04841193316227485
	pesos_i(4201) := b"0000000000000000_0000000000000000_0001110010110111_0110101110100101"; -- 0.11217377461557612
	pesos_i(4202) := b"1111111111111111_1111111111111111_1101001001110101_0111110011011010"; -- -0.1778947800531564
	pesos_i(4203) := b"1111111111111111_1111111111111111_1111001111101001_0010011101101111"; -- -0.04722360182572565
	pesos_i(4204) := b"0000000000000000_0000000000000000_0010101110000110_1111110111101011"; -- 0.1700285624812253
	pesos_i(4205) := b"1111111111111111_1111111111111111_1110101100100010_1010000100001011"; -- -0.08150285233592171
	pesos_i(4206) := b"1111111111111111_1111111111111111_1110001001001010_1110010010000011"; -- -0.1160447291735952
	pesos_i(4207) := b"1111111111111111_1111111111111111_1110110101000100_1000001000111011"; -- -0.07317339010243162
	pesos_i(4208) := b"1111111111111111_1111111111111111_1101101111101001_1101001100101101"; -- -0.14096336519648062
	pesos_i(4209) := b"0000000000000000_0000000000000000_0000000011001011_0000011010011111"; -- 0.003097928930280939
	pesos_i(4210) := b"0000000000000000_0000000000000000_0001110000000101_1111101000011000"; -- 0.10946620058722246
	pesos_i(4211) := b"0000000000000000_0000000000000000_0001010001000011_0111100011000010"; -- 0.07915453667863835
	pesos_i(4212) := b"0000000000000000_0000000000000000_0010001011010111_1010111110010011"; -- 0.13610360460458745
	pesos_i(4213) := b"0000000000000000_0000000000000000_0010001011011010_0001010011011111"; -- 0.1361401600359823
	pesos_i(4214) := b"0000000000000000_0000000000000000_0001000010100000_1000100001101001"; -- 0.06494953703136909
	pesos_i(4215) := b"0000000000000000_0000000000000000_0010000010100110_0010010011111101"; -- 0.12753516374194432
	pesos_i(4216) := b"1111111111111111_1111111111111111_1111110111011101_1101110110101110"; -- -0.00833334446611636
	pesos_i(4217) := b"0000000000000000_0000000000000000_0001000101100001_0000100000000000"; -- 0.06788682940501242
	pesos_i(4218) := b"0000000000000000_0000000000000000_0010110100101111_0001111100111111"; -- 0.17650027555186135
	pesos_i(4219) := b"1111111111111111_1111111111111111_1110101010100101_1000111101110001"; -- -0.08341125012102091
	pesos_i(4220) := b"1111111111111111_1111111111111111_1110011100100000_0110110000011101"; -- -0.09716152465089914
	pesos_i(4221) := b"1111111111111111_1111111111111111_1101011000000010_0011100100000010"; -- -0.16402858452234478
	pesos_i(4222) := b"0000000000000000_0000000000000000_0001110100101100_0100110001110001"; -- 0.11395719295929113
	pesos_i(4223) := b"0000000000000000_0000000000000000_0010110001100110_0011101011100100"; -- 0.1734349065335276
	pesos_i(4224) := b"0000000000000000_0000000000000000_0001110010111001_0101011110010000"; -- 0.1122030951042153
	pesos_i(4225) := b"1111111111111111_1111111111111111_1101101110000100_0110011001111011"; -- -0.1425109816093785
	pesos_i(4226) := b"0000000000000000_0000000000000000_0010010101100000_1000110011011111"; -- 0.14600449032501495
	pesos_i(4227) := b"1111111111111111_1111111111111111_1101011010001110_1100100001101010"; -- -0.16188380626555196
	pesos_i(4228) := b"1111111111111111_1111111111111111_1111011111101010_1111010110000100"; -- -0.03157105957333669
	pesos_i(4229) := b"1111111111111111_1111111111111111_1110110011111001_0011000001111101"; -- -0.07432267143275748
	pesos_i(4230) := b"0000000000000000_0000000000000000_0000001010010000_0001100110110011"; -- 0.01001129744414336
	pesos_i(4231) := b"1111111111111111_1111111111111111_1111011100001100_1101011010100100"; -- -0.03496035105457492
	pesos_i(4232) := b"0000000000000000_0000000000000000_0000011111101100_0111001001110001"; -- 0.030951645361197707
	pesos_i(4233) := b"1111111111111111_1111111111111111_1101100111000000_1111000111101100"; -- -0.14939964288576596
	pesos_i(4234) := b"0000000000000000_0000000000000000_0000000111011111_1100001111100111"; -- 0.007320636623206926
	pesos_i(4235) := b"1111111111111111_1111111111111111_1111110101010011_1110101101010000"; -- -0.010438244785798472
	pesos_i(4236) := b"1111111111111111_1111111111111111_1110000100001010_1100011010000111"; -- -0.12092932887479282
	pesos_i(4237) := b"1111111111111111_1111111111111111_1101111110001011_1000000001011001"; -- -0.12677762830287928
	pesos_i(4238) := b"0000000000000000_0000000000000000_0000111110001111_1111101101111100"; -- 0.06079074652074148
	pesos_i(4239) := b"0000000000000000_0000000000000000_0000010101000100_1111011100000101"; -- 0.020583571181591508
	pesos_i(4240) := b"0000000000000000_0000000000000000_0001111000011000_1000100101111010"; -- 0.11756190509677192
	pesos_i(4241) := b"1111111111111111_1111111111111111_1101001101011111_1110000001100100"; -- -0.17431829039516444
	pesos_i(4242) := b"1111111111111111_1111111111111111_1110001110101010_1001000000101010"; -- -0.11067866292384299
	pesos_i(4243) := b"1111111111111111_1111111111111111_1111100101111010_0010100010011110"; -- -0.025479756814787296
	pesos_i(4244) := b"1111111111111111_1111111111111111_1101001000101110_0011010001010101"; -- -0.1789824765286594
	pesos_i(4245) := b"1111111111111111_1111111111111111_1101010011111100_0000110100101100"; -- -0.16802900000682786
	pesos_i(4246) := b"1111111111111111_1111111111111111_1110110001100011_1011001100100101"; -- -0.07660370215287855
	pesos_i(4247) := b"0000000000000000_0000000000000000_0001110100110001_1001101001001110"; -- 0.1140381278908619
	pesos_i(4248) := b"0000000000000000_0000000000000000_0001111010010011_0010100111111110"; -- 0.11943304500046102
	pesos_i(4249) := b"1111111111111111_1111111111111111_1111101010110000_1111111100100001"; -- -0.02073674637353395
	pesos_i(4250) := b"0000000000000000_0000000000000000_0001000011110000_0101011001001101"; -- 0.06616725326709029
	pesos_i(4251) := b"0000000000000000_0000000000000000_0010100101001000_0101110010110000"; -- 0.16126040734463126
	pesos_i(4252) := b"1111111111111111_1111111111111111_1110101011000011_1101011100010110"; -- -0.08294921600018003
	pesos_i(4253) := b"1111111111111111_1111111111111111_1101100010011010_0010111101010100"; -- -0.15389732545997578
	pesos_i(4254) := b"0000000000000000_0000000000000000_0010011001100011_1110101110010010"; -- 0.14996216126382614
	pesos_i(4255) := b"0000000000000000_0000000000000000_0001111001000101_1011011100011000"; -- 0.11825126968177227
	pesos_i(4256) := b"0000000000000000_0000000000000000_0010001101010111_1110011001000010"; -- 0.13805998897339858
	pesos_i(4257) := b"0000000000000000_0000000000000000_0001001010010010_1011000011100000"; -- 0.0725508258191112
	pesos_i(4258) := b"0000000000000000_0000000000000000_0000001100111110_1111011001010001"; -- 0.012679476622095787
	pesos_i(4259) := b"0000000000000000_0000000000000000_0001101110101101_1001001101111100"; -- 0.10811731132133699
	pesos_i(4260) := b"1111111111111111_1111111111111111_1110000101101100_0001111000011010"; -- -0.11944400661607234
	pesos_i(4261) := b"0000000000000000_0000000000000000_0000110111111011_0110000110100111"; -- 0.05461702647590051
	pesos_i(4262) := b"1111111111111111_1111111111111111_1111011101101011_1001101001001100"; -- -0.0335143626668688
	pesos_i(4263) := b"0000000000000000_0000000000000000_0000111110010001_0001001100001100"; -- 0.060807409649238614
	pesos_i(4264) := b"0000000000000000_0000000000000000_0000100100110111_0110111110101101"; -- 0.036002139714686104
	pesos_i(4265) := b"0000000000000000_0000000000000000_0010101000010011_0100011001110110"; -- 0.16435661686418307
	pesos_i(4266) := b"1111111111111111_1111111111111111_1111111000111000_1000010011011101"; -- -0.006950088497107892
	pesos_i(4267) := b"0000000000000000_0000000000000000_0000101110110101_1110111000110011"; -- 0.04574478857997583
	pesos_i(4268) := b"0000000000000000_0000000000000000_0001011111000000_1110001110111010"; -- 0.0927870110442662
	pesos_i(4269) := b"0000000000000000_0000000000000000_0001010010110110_0101101001011011"; -- 0.08090748514708748
	pesos_i(4270) := b"0000000000000000_0000000000000000_0010000110010100_1000110001100101"; -- 0.13117291890695043
	pesos_i(4271) := b"1111111111111111_1111111111111111_1111111111001010_1001000100010111"; -- -0.0008153266018345089
	pesos_i(4272) := b"0000000000000000_0000000000000000_0000100101111111_1101100000100101"; -- 0.0371069993235951
	pesos_i(4273) := b"0000000000000000_0000000000000000_0001000101001100_1001010010110000"; -- 0.0675747804607965
	pesos_i(4274) := b"1111111111111111_1111111111111111_1111101101001110_0101101101101010"; -- -0.018335615829775977
	pesos_i(4275) := b"0000000000000000_0000000000000000_0001001010100000_0101111100010101"; -- 0.07275957347982227
	pesos_i(4276) := b"0000000000000000_0000000000000000_0010100010101100_0101001001010110"; -- 0.15887941925546956
	pesos_i(4277) := b"0000000000000000_0000000000000000_0001011001101001_0101110000000110"; -- 0.08754515782546056
	pesos_i(4278) := b"1111111111111111_1111111111111111_1111001100001010_1101111011100010"; -- -0.05061537719903093
	pesos_i(4279) := b"1111111111111111_1111111111111111_1111110110001111_0010101000101001"; -- -0.00953423026130145
	pesos_i(4280) := b"1111111111111111_1111111111111111_1111001101011001_1001000000101011"; -- -0.04941462462881391
	pesos_i(4281) := b"0000000000000000_0000000000000000_0001011010000001_0111110110100001"; -- 0.08791337193274862
	pesos_i(4282) := b"1111111111111111_1111111111111111_1111000001101001_1011110001010001"; -- -0.060886602620867564
	pesos_i(4283) := b"0000000000000000_0000000000000000_0010000111110101_1010111100101001"; -- 0.13265509378718032
	pesos_i(4284) := b"1111111111111111_1111111111111111_1111101011011100_1101111101101101"; -- -0.02006724915773854
	pesos_i(4285) := b"1111111111111111_1111111111111111_1110010011011000_0011100010101110"; -- -0.10607572314182898
	pesos_i(4286) := b"1111111111111111_1111111111111111_1101100010110111_1010001110100010"; -- -0.15344788834333656
	pesos_i(4287) := b"0000000000000000_0000000000000000_0010001111001100_1101010010011001"; -- 0.13984421468620345
	pesos_i(4288) := b"0000000000000000_0000000000000000_0001010101000111_1000101000001010"; -- 0.08312285189962146
	pesos_i(4289) := b"1111111111111111_1111111111111111_1111000110010001_0001010001110101"; -- -0.056380006166480326
	pesos_i(4290) := b"1111111111111111_1111111111111111_1101100110010111_1010110001110010"; -- -0.1500293942110825
	pesos_i(4291) := b"1111111111111111_1111111111111111_1110000100110011_1001100101010101"; -- -0.12030641256719687
	pesos_i(4292) := b"1111111111111111_1111111111111111_1101011011110100_0100001000111001"; -- -0.16033540831489412
	pesos_i(4293) := b"1111111111111111_1111111111111111_1111110111101101_0111110110100000"; -- -0.008094929249807415
	pesos_i(4294) := b"1111111111111111_1111111111111111_1110010111001101_1111011101101101"; -- -0.10232595052773898
	pesos_i(4295) := b"0000000000000000_0000000000000000_0010000000100000_0110011010111000"; -- 0.12549440372902268
	pesos_i(4296) := b"1111111111111111_1111111111111111_1101101101100001_0111011101110100"; -- -0.14304402740648214
	pesos_i(4297) := b"0000000000000000_0000000000000000_0000000001100001_0111000100010100"; -- 0.0014868424523124286
	pesos_i(4298) := b"1111111111111111_1111111111111111_1110101001001010_1011110100000111"; -- -0.08479708278404904
	pesos_i(4299) := b"1111111111111111_1111111111111111_1110010100011111_0000110111110010"; -- -0.10499489632272642
	pesos_i(4300) := b"1111111111111111_1111111111111111_1111001011001001_1000100101100011"; -- -0.05161229445272138
	pesos_i(4301) := b"0000000000000000_0000000000000000_0000011100111101_0001100011000011"; -- 0.028276012006485312
	pesos_i(4302) := b"1111111111111111_1111111111111111_1110111101110010_0101010010010111"; -- -0.06466170609242365
	pesos_i(4303) := b"1111111111111111_1111111111111111_1101100001000011_0000001100000111"; -- -0.15522748077913748
	pesos_i(4304) := b"1111111111111111_1111111111111111_1111010111001000_0010000001110010"; -- -0.039915058231735495
	pesos_i(4305) := b"1111111111111111_1111111111111111_1110111100010011_1010010101110101"; -- -0.06610647092345595
	pesos_i(4306) := b"0000000000000000_0000000000000000_0000100011110001_0101001000011010"; -- 0.03493226175304913
	pesos_i(4307) := b"0000000000000000_0000000000000000_0000011111110101_1101011101100110"; -- 0.031094992162967173
	pesos_i(4308) := b"1111111111111111_1111111111111111_1110010110011111_0100111110001110"; -- -0.10303786076763928
	pesos_i(4309) := b"0000000000000000_0000000000000000_0001001000101111_1110011001011011"; -- 0.0710433932952863
	pesos_i(4310) := b"0000000000000000_0000000000000000_0010100010110001_0001110101111011"; -- 0.1589525629127513
	pesos_i(4311) := b"1111111111111111_1111111111111111_1100101010111100_1110011001010110"; -- -0.20805511855397815
	pesos_i(4312) := b"1111111111111111_1111111111111111_1101000001010011_1011010111100010"; -- -0.18622267950942842
	pesos_i(4313) := b"1111111111111111_1111111111111111_1111000101010101_0000001000011010"; -- -0.05729662765767996
	pesos_i(4314) := b"1111111111111111_1111111111111111_1111110110111100_0010011011001111"; -- -0.008847784391983278
	pesos_i(4315) := b"1111111111111111_1111111111111111_1110011110101110_0111101101100101"; -- -0.09499386580933059
	pesos_i(4316) := b"0000000000000000_0000000000000000_0000100110010000_0000010101110110"; -- 0.03735384111512976
	pesos_i(4317) := b"1111111111111111_1111111111111111_1110110010001110_1111101000001001"; -- -0.07594334861994047
	pesos_i(4318) := b"1111111111111111_1111111111111111_1110011111110011_0111001000111111"; -- -0.09394155458322913
	pesos_i(4319) := b"0000000000000000_0000000000000000_0000100000111111_1110111011100100"; -- 0.03222554270706329
	pesos_i(4320) := b"0000000000000000_0000000000000000_0001100100011110_1101000001001010"; -- 0.09812642869681545
	pesos_i(4321) := b"1111111111111111_1111111111111111_1111100101001011_0011101110010100"; -- -0.026195789802903956
	pesos_i(4322) := b"0000000000000000_0000000000000000_0001111101110011_1001001001011101"; -- 0.12285723459963743
	pesos_i(4323) := b"0000000000000000_0000000000000000_0001010100111100_1111110000010101"; -- 0.08296180264952074
	pesos_i(4324) := b"0000000000000000_0000000000000000_0010010100111100_0010101111001100"; -- 0.14544938790939238
	pesos_i(4325) := b"0000000000000000_0000000000000000_0000100101000110_1010001010000111"; -- 0.03623405265896755
	pesos_i(4326) := b"1111111111111111_1111111111111111_1111101000101001_0000111011001001"; -- -0.022811008497773108
	pesos_i(4327) := b"0000000000000000_0000000000000000_0010110011110000_0010100000101001"; -- 0.17553950300888918
	pesos_i(4328) := b"0000000000000000_0000000000000000_0001100011100001_1011110101001101"; -- 0.09719451074703625
	pesos_i(4329) := b"1111111111111111_1111111111111111_1110010111110110_0101100010000111"; -- -0.10170981128618795
	pesos_i(4330) := b"1111111111111111_1111111111111111_1101111110010011_0101000101010101"; -- -0.12665836019636484
	pesos_i(4331) := b"1111111111111111_1111111111111111_1101100110000010_1000111110110101"; -- -0.15035154191864966
	pesos_i(4332) := b"1111111111111111_1111111111111111_1101100101011100_0110101000011000"; -- -0.15093361777144904
	pesos_i(4333) := b"0000000000000000_0000000000000000_0000011101111000_1001111110010000"; -- 0.029184315363332932
	pesos_i(4334) := b"0000000000000000_0000000000000000_0001001010010101_0010110101000001"; -- 0.07258875685417573
	pesos_i(4335) := b"1111111111111111_1111111111111111_1101110000100000_1110110011010100"; -- -0.1401226027396492
	pesos_i(4336) := b"1111111111111111_1111111111111111_1110111101011101_1010110010000000"; -- -0.06497690092476356
	pesos_i(4337) := b"1111111111111111_1111111111111111_1111110011011011_1110001010011000"; -- -0.012269819179581021
	pesos_i(4338) := b"1111111111111111_1111111111111111_1110000001001100_1110011000000111"; -- -0.12382662131898203
	pesos_i(4339) := b"0000000000000000_0000000000000000_0001110001100010_1000111011000000"; -- 0.11087886997739758
	pesos_i(4340) := b"1111111111111111_1111111111111111_1110010010001011_0010010111010000"; -- -0.10725177460084367
	pesos_i(4341) := b"0000000000000000_0000000000000000_0001001010011110_1110101110011000"; -- 0.07273743124934948
	pesos_i(4342) := b"1111111111111111_1111111111111111_1110111110001110_0010111110110001"; -- -0.06423665936090463
	pesos_i(4343) := b"1111111111111111_1111111111111111_1110011000000010_1000001111101111"; -- -0.10152411858476469
	pesos_i(4344) := b"1111111111111111_1111111111111111_1101111101010010_1001110101001100"; -- -0.1276456537734459
	pesos_i(4345) := b"0000000000000000_0000000000000000_0000000111110110_1100101000001111"; -- 0.0076719557691287184
	pesos_i(4346) := b"0000000000000000_0000000000000000_0010011100001010_0110101010110011"; -- 0.1525026975680945
	pesos_i(4347) := b"1111111111111111_1111111111111111_1101010111010010_0100001100000111"; -- -0.16476040906321052
	pesos_i(4348) := b"1111111111111111_1111111111111111_1110001011010101_1110000101001010"; -- -0.11392394973848882
	pesos_i(4349) := b"1111111111111111_1111111111111111_1101110000100100_0011111100010000"; -- -0.14007192481906106
	pesos_i(4350) := b"1111111111111111_1111111111111111_1111110110101000_0001111110101110"; -- -0.009153385116945224
	pesos_i(4351) := b"1111111111111111_1111111111111111_1111111001010001_0000000111010000"; -- -0.006576430058435691
	pesos_i(4352) := b"0000000000000000_0000000000000000_0010101100111100_0111011101111110"; -- 0.16889139966914432
	pesos_i(4353) := b"0000000000000000_0000000000000000_0000101010000000_0001110110010110"; -- 0.04101738847337719
	pesos_i(4354) := b"1111111111111111_1111111111111111_1110001110010101_1111110111101110"; -- -0.11099255498673241
	pesos_i(4355) := b"0000000000000000_0000000000000000_0001001010001011_1101101000000010"; -- 0.07244646589965827
	pesos_i(4356) := b"1111111111111111_1111111111111111_1110001111110111_1110101011001100"; -- -0.10949833403822783
	pesos_i(4357) := b"0000000000000000_0000000000000000_0000111110111100_1000100010000001"; -- 0.06147053852302459
	pesos_i(4358) := b"1111111111111111_1111111111111111_1111010011010001_0010101111111110"; -- -0.043683290881445506
	pesos_i(4359) := b"1111111111111111_1111111111111111_1111011111001001_0110001011111101"; -- -0.03208333332977972
	pesos_i(4360) := b"1111111111111111_1111111111111111_1101100010010100_0000111111101011"; -- -0.15399075037357784
	pesos_i(4361) := b"1111111111111111_1111111111111111_1110001011010111_1100011111100000"; -- -0.11389494693896605
	pesos_i(4362) := b"1111111111111111_1111111111111111_1111010111000010_1111011011111101"; -- -0.039993823309824594
	pesos_i(4363) := b"0000000000000000_0000000000000000_0000001101010010_0011000000101010"; -- 0.01297284142348218
	pesos_i(4364) := b"0000000000000000_0000000000000000_0001110101101010_0001010001001000"; -- 0.11489989038956334
	pesos_i(4365) := b"1111111111111111_1111111111111111_1101001001001000_1010101001010110"; -- -0.17857871444917003
	pesos_i(4366) := b"0000000000000000_0000000000000000_0000011100001010_0100011011111011"; -- 0.027500568754096125
	pesos_i(4367) := b"0000000000000000_0000000000000000_0001000010011010_1110000011001100"; -- 0.06486325242005321
	pesos_i(4368) := b"0000000000000000_0000000000000000_0001111101000101_1110111001111111"; -- 0.12216082191448283
	pesos_i(4369) := b"0000000000000000_0000000000000000_0000010111111010_0101101010101000"; -- 0.023351350846876257
	pesos_i(4370) := b"0000000000000000_0000000000000000_0010101111110000_0001010011100010"; -- 0.17163210404521348
	pesos_i(4371) := b"0000000000000000_0000000000000000_0001110011100111_1101011000101100"; -- 0.11291254595474459
	pesos_i(4372) := b"1111111111111111_1111111111111111_1111001011001001_1111110001100001"; -- -0.05160544050059638
	pesos_i(4373) := b"0000000000000000_0000000000000000_0001111001001111_1100011110100011"; -- 0.11840484361149298
	pesos_i(4374) := b"1111111111111111_1111111111111111_1110101111101101_0001000010000101"; -- -0.0784139324281022
	pesos_i(4375) := b"0000000000000000_0000000000000000_0010001111001101_0100000000100011"; -- 0.1398506245783121
	pesos_i(4376) := b"0000000000000000_0000000000000000_0011101011111000_0101111100010111"; -- 0.2303523474398287
	pesos_i(4377) := b"1111111111111111_1111111111111111_1111111001010011_1000110001110100"; -- -0.006537648779458719
	pesos_i(4378) := b"1111111111111111_1111111111111111_1101011100011001_1001000010001110"; -- -0.15976616405717534
	pesos_i(4379) := b"1111111111111111_1111111111111111_1101110100101110_1111100000000110"; -- -0.13600206227241243
	pesos_i(4380) := b"0000000000000000_0000000000000000_0001100100100010_0011001110000110"; -- 0.0981781198406905
	pesos_i(4381) := b"1111111111111111_1111111111111111_1111100100010110_1100100000010101"; -- -0.026996130891090587
	pesos_i(4382) := b"1111111111111111_1111111111111111_1110110111101101_1001110100110101"; -- -0.07059304677640087
	pesos_i(4383) := b"0000000000000000_0000000000000000_0001110110001111_0110011011111011"; -- 0.11546939496790662
	pesos_i(4384) := b"0000000000000000_0000000000000000_0010110001010100_0000101010111100"; -- 0.17315737803889744
	pesos_i(4385) := b"1111111111111111_1111111111111111_1111111000011000_1111100010011101"; -- -0.007431470519902248
	pesos_i(4386) := b"1111111111111111_1111111111111111_1111000011010100_0001011000110001"; -- -0.05926381399698023
	pesos_i(4387) := b"0000000000000000_0000000000000000_0000000111100101_1101000110011011"; -- 0.007413006266695686
	pesos_i(4388) := b"1111111111111111_1111111111111111_1111010011001101_0101011010011000"; -- -0.043741786790063596
	pesos_i(4389) := b"0000000000000000_0000000000000000_0000001111110001_0001010010100001"; -- 0.01539734767319473
	pesos_i(4390) := b"1111111111111111_1111111111111111_1101111010100111_0000100100101010"; -- -0.13026373610028652
	pesos_i(4391) := b"0000000000000000_0000000000000000_0010110011000101_0001011100111110"; -- 0.17488236686182038
	pesos_i(4392) := b"0000000000000000_0000000000000000_0000100100011111_1000110101101000"; -- 0.035637701032313895
	pesos_i(4393) := b"0000000000000000_0000000000000000_0001101011100111_1000010100111100"; -- 0.10509522173782113
	pesos_i(4394) := b"1111111111111111_1111111111111111_1101110001101111_0000101111110100"; -- -0.13893056192001968
	pesos_i(4395) := b"0000000000000000_0000000000000000_0001101111001011_1100101101100100"; -- 0.10857840723549858
	pesos_i(4396) := b"1111111111111111_1111111111111111_1101010010000001_0101001000000101"; -- -0.16990172738412257
	pesos_i(4397) := b"0000000000000000_0000000000000000_0000111100111100_1001010111110100"; -- 0.05951821532948907
	pesos_i(4398) := b"0000000000000000_0000000000000000_0000011100101110_1010100111010011"; -- 0.028055776621235477
	pesos_i(4399) := b"1111111111111111_1111111111111111_1111111101110000_1001100000111001"; -- -0.0021881924054027585
	pesos_i(4400) := b"0000000000000000_0000000000000000_0000100010110000_1100001110000011"; -- 0.033947200358533686
	pesos_i(4401) := b"1111111111111111_1111111111111111_1111111111011010_1100101000011110"; -- -0.0005677868340799865
	pesos_i(4402) := b"1111111111111111_1111111111111111_1111001001010010_0110010110011111"; -- -0.053430222301542055
	pesos_i(4403) := b"1111111111111111_1111111111111111_1111111100010101_0100101110010101"; -- -0.0035813105048155226
	pesos_i(4404) := b"1111111111111111_1111111111111111_1110010011010010_0011101010011001"; -- -0.10616716157846248
	pesos_i(4405) := b"1111111111111111_1111111111111111_1110011101111001_0011111101111100"; -- -0.09580615266373668
	pesos_i(4406) := b"0000000000000000_0000000000000000_0001101101110000_0100110111011001"; -- 0.10718237444944424
	pesos_i(4407) := b"1111111111111111_1111111111111111_1111000010010111_0111000111010011"; -- -0.060189138467415845
	pesos_i(4408) := b"0000000000000000_0000000000000000_0001011010011000_0100010000111011"; -- 0.08826090267966943
	pesos_i(4409) := b"1111111111111111_1111111111111111_1111011110101110_0000001111001110"; -- -0.03250099397280358
	pesos_i(4410) := b"1111111111111111_1111111111111111_1110101100001011_0001100110011110"; -- -0.08186187650650578
	pesos_i(4411) := b"0000000000000000_0000000000000000_0000001101101000_1111001101111101"; -- 0.01332017707548152
	pesos_i(4412) := b"1111111111111111_1111111111111111_1110000110011110_1100101100010000"; -- -0.11867075779777121
	pesos_i(4413) := b"1111111111111111_1111111111111111_1111110100010011_1101100010011010"; -- -0.011415922531983307
	pesos_i(4414) := b"0000000000000000_0000000000000000_0000001011010100_1100010011011100"; -- 0.01105909694331059
	pesos_i(4415) := b"0000000000000000_0000000000000000_0001100111001011_0011110111011110"; -- 0.10075747183488068
	pesos_i(4416) := b"0000000000000000_0000000000000000_0010100000000001_1000100110001110"; -- 0.15627345762753217
	pesos_i(4417) := b"1111111111111111_1111111111111111_1110111001111010_1011011010011010"; -- -0.06844004372401136
	pesos_i(4418) := b"0000000000000000_0000000000000000_0010000000001001_0001000000101110"; -- 0.12513829340678417
	pesos_i(4419) := b"1111111111111111_1111111111111111_1111111101000010_1111011000001001"; -- -0.0028845051147556875
	pesos_i(4420) := b"1111111111111111_1111111111111111_1110100011000001_0111000101101110"; -- -0.09079829285738689
	pesos_i(4421) := b"1111111111111111_1111111111111111_1110101000011100_1011100010110010"; -- -0.08549924513755497
	pesos_i(4422) := b"1111111111111111_1111111111111111_1111010010001110_0011011011100011"; -- -0.0447049803997883
	pesos_i(4423) := b"0000000000000000_0000000000000000_0001101001011001_1101001110000100"; -- 0.10293313964284452
	pesos_i(4424) := b"1111111111111111_1111111111111111_1100101010001101_1111101000000001"; -- -0.20877110929140408
	pesos_i(4425) := b"0000000000000000_0000000000000000_0000001000101001_0100101000010110"; -- 0.008442526254242516
	pesos_i(4426) := b"1111111111111111_1111111111111111_1101111101100100_1101011000111011"; -- -0.12736760190469593
	pesos_i(4427) := b"0000000000000000_0000000000000000_0000101010001001_1011100011010001"; -- 0.04116397003935495
	pesos_i(4428) := b"0000000000000000_0000000000000000_0001101011110010_0001100111011001"; -- 0.10525666767054563
	pesos_i(4429) := b"0000000000000000_0000000000000000_0010011011011110_1111001011111101"; -- 0.15183943444335013
	pesos_i(4430) := b"0000000000000000_0000000000000000_0000010101000000_0000110010110000"; -- 0.02050856873031814
	pesos_i(4431) := b"1111111111111111_1111111111111111_1111010000011111_0101100010110011"; -- -0.04639669057802088
	pesos_i(4432) := b"0000000000000000_0000000000000000_0000010001101111_1111001110011111"; -- 0.017333246431593508
	pesos_i(4433) := b"1111111111111111_1111111111111111_1111101010010011_1111101110010111"; -- -0.02117946204769738
	pesos_i(4434) := b"1111111111111111_1111111111111111_1110011010011011_0100110110001101"; -- -0.09919276525045141
	pesos_i(4435) := b"1111111111111111_1111111111111111_1111100100100101_0110011101001010"; -- -0.026773018274858375
	pesos_i(4436) := b"1111111111111111_1111111111111111_1110000001100000_1110111101000101"; -- -0.12352089466911832
	pesos_i(4437) := b"1111111111111111_1111111111111111_1111011000011010_0010110101101000"; -- -0.03866306503294024
	pesos_i(4438) := b"1111111111111111_1111111111111111_1111010010111100_0111011100011101"; -- -0.04399924797475312
	pesos_i(4439) := b"0000000000000000_0000000000000000_0001000110000001_1000001011011100"; -- 0.06838243350551647
	pesos_i(4440) := b"0000000000000000_0000000000000000_0001011001000100_1111110111000000"; -- 0.08699022222814877
	pesos_i(4441) := b"1111111111111111_1111111111111111_1110110100110111_0101111011111110"; -- -0.07337385451536935
	pesos_i(4442) := b"1111111111111111_1111111111111111_1111011001111001_1100111100010011"; -- -0.03720384400566176
	pesos_i(4443) := b"1111111111111111_1111111111111111_1101001100010011_0111100100001001"; -- -0.17548411881566786
	pesos_i(4444) := b"0000000000000000_0000000000000000_0000110101011001_1110010100001101"; -- 0.05215293473715128
	pesos_i(4445) := b"1111111111111111_1111111111111111_1111110101000001_0101000011100110"; -- -0.010722106712995725
	pesos_i(4446) := b"0000000000000000_0000000000000000_0001110000110011_1100001111110011"; -- 0.11016487780358196
	pesos_i(4447) := b"1111111111111111_1111111111111111_1111110101000011_0110001001111001"; -- -0.010690541681907167
	pesos_i(4448) := b"1111111111111111_1111111111111111_1111101100001111_1101010110000110"; -- -0.019289641121435358
	pesos_i(4449) := b"0000000000000000_0000000000000000_0000101001101000_1001111101111110"; -- 0.04065892061639372
	pesos_i(4450) := b"1111111111111111_1111111111111111_1110110011001010_1111000001111101"; -- -0.07502839047793086
	pesos_i(4451) := b"0000000000000000_0000000000000000_0010100000101001_0011110001010011"; -- 0.15687920592098273
	pesos_i(4452) := b"0000000000000000_0000000000000000_0000000111110000_1001101101001001"; -- 0.007577614994121112
	pesos_i(4453) := b"1111111111111111_1111111111111111_1111001101011011_1011110001001011"; -- -0.04938147715812793
	pesos_i(4454) := b"0000000000000000_0000000000000000_0000101110011011_0010010011000011"; -- 0.04533605340947595
	pesos_i(4455) := b"0000000000000000_0000000000000000_0010011011010001_0011100000110011"; -- 0.15162993658702925
	pesos_i(4456) := b"0000000000000000_0000000000000000_0010110100100011_1101110010000110"; -- 0.17632845192995603
	pesos_i(4457) := b"1111111111111111_1111111111111111_1101100011101101_1111100001000010"; -- -0.152618869650595
	pesos_i(4458) := b"0000000000000000_0000000000000000_0000000001101110_1100000001011101"; -- 0.0016899325807144695
	pesos_i(4459) := b"0000000000000000_0000000000000000_0010011010010110_0001000011101011"; -- 0.15072732670491737
	pesos_i(4460) := b"1111111111111111_1111111111111111_1110100111100010_1100110010010001"; -- -0.08638307053347645
	pesos_i(4461) := b"1111111111111111_1111111111111111_1110111111100100_0101001110001110"; -- -0.062922265922355
	pesos_i(4462) := b"0000000000000000_0000000000000000_0000001000111011_0011101001011110"; -- 0.008716247554425193
	pesos_i(4463) := b"1111111111111111_1111111111111111_1110010111001101_1111111011010001"; -- -0.10232551006863075
	pesos_i(4464) := b"0000000000000000_0000000000000000_0001100010011011_0001010111101010"; -- 0.09611641859444361
	pesos_i(4465) := b"0000000000000000_0000000000000000_0001011110101001_0010000011001101"; -- 0.09242444038766778
	pesos_i(4466) := b"0000000000000000_0000000000000000_0010011000111100_0101011111000110"; -- 0.14935825906506175
	pesos_i(4467) := b"1111111111111111_1111111111111111_1101110000011110_1011010010100010"; -- -0.14015646983062932
	pesos_i(4468) := b"0000000000000000_0000000000000000_0010011011111001_1101111011010001"; -- 0.15225021933237246
	pesos_i(4469) := b"0000000000000000_0000000000000000_0000110100100101_1001011011011101"; -- 0.05135481743968176
	pesos_i(4470) := b"1111111111111111_1111111111111111_1111010001001100_0011101001110110"; -- -0.04571184739003312
	pesos_i(4471) := b"1111111111111111_1111111111111111_1111101100011010_1101000110101110"; -- -0.01912202353590779
	pesos_i(4472) := b"0000000000000000_0000000000000000_0010110010101101_1101000100010110"; -- 0.1745272329586494
	pesos_i(4473) := b"1111111111111111_1111111111111111_1111000111100100_0000010001001110"; -- -0.05511448945532653
	pesos_i(4474) := b"1111111111111111_1111111111111111_1110011011000111_1110010100010010"; -- -0.09851234734291629
	pesos_i(4475) := b"1111111111111111_1111111111111111_1111100010000101_0101011010110000"; -- -0.029215413981047367
	pesos_i(4476) := b"0000000000000000_0000000000000000_0010001000110001_0111100100101110"; -- 0.13356740363328637
	pesos_i(4477) := b"0000000000000000_0000000000000000_0010000110101110_1110011010000010"; -- 0.13157501858994958
	pesos_i(4478) := b"0000000000000000_0000000000000000_0001010010101011_1101011000011001"; -- 0.08074701423103554
	pesos_i(4479) := b"0000000000000000_0000000000000000_0001011010001000_1011000001000101"; -- 0.08802320169844466
	pesos_i(4480) := b"0000000000000000_0000000000000000_0000110101111011_1011111100110111"; -- 0.05266947837994018
	pesos_i(4481) := b"1111111111111111_1111111111111111_1111100000110100_0111111110011000"; -- -0.030448937841326126
	pesos_i(4482) := b"0000000000000000_0000000000000000_0001010110100000_0001000110100011"; -- 0.08447370743838287
	pesos_i(4483) := b"0000000000000000_0000000000000000_0000011000010001_1011010110100010"; -- 0.023707725477080784
	pesos_i(4484) := b"1111111111111111_1111111111111111_1110111101001001_0001011000001101"; -- -0.06529104409568802
	pesos_i(4485) := b"0000000000000000_0000000000000000_0001011010011101_0011110111000111"; -- 0.08833681206019559
	pesos_i(4486) := b"1111111111111111_1111111111111111_1101101100110011_1011000000110000"; -- -0.14374255007502457
	pesos_i(4487) := b"1111111111111111_1111111111111111_1111110011010111_0100110000011111"; -- -0.01233982317928063
	pesos_i(4488) := b"1111111111111111_1111111111111111_1011101110111100_0000011001001001"; -- -0.2666622230007831
	pesos_i(4489) := b"1111111111111111_1111111111111111_1110101010000011_1100101010011011"; -- -0.08392652250448625
	pesos_i(4490) := b"1111111111111111_1111111111111111_1111000111101000_0011111000110011"; -- -0.05505000347002218
	pesos_i(4491) := b"0000000000000000_0000000000000000_0000011100101000_0100010011101101"; -- 0.02795820991877643
	pesos_i(4492) := b"1111111111111111_1111111111111111_1101111111010011_0001101110001001"; -- -0.1256850041792752
	pesos_i(4493) := b"1111111111111111_1111111111111111_1101010100111010_1101100000101000"; -- -0.1670708563235478
	pesos_i(4494) := b"0000000000000000_0000000000000000_0001101000111101_0011000010100010"; -- 0.10249618484551222
	pesos_i(4495) := b"1111111111111111_1111111111111111_1101000011110111_1001010101110010"; -- -0.18372217139181216
	pesos_i(4496) := b"1111111111111111_1111111111111111_1111001010011011_0000110011111101"; -- -0.0523216135520415
	pesos_i(4497) := b"0000000000000000_0000000000000000_0010101111010101_0000000001010000"; -- 0.17121889081159616
	pesos_i(4498) := b"1111111111111111_1111111111111111_1110111101011101_1111011110101000"; -- -0.06497242115697899
	pesos_i(4499) := b"0000000000000000_0000000000000000_0001111110101000_0001000000100100"; -- 0.12365818853726074
	pesos_i(4500) := b"1111111111111111_1111111111111111_1110100010010011_1111001010111100"; -- -0.09149248999894724
	pesos_i(4501) := b"0000000000000000_0000000000000000_0010010101100100_0101010100011011"; -- 0.146062201624207
	pesos_i(4502) := b"0000000000000000_0000000000000000_0010100101010101_1000011111010111"; -- 0.16146134369382997
	pesos_i(4503) := b"1111111111111111_1111111111111111_1110010011110100_1101110101111010"; -- -0.10563865437605412
	pesos_i(4504) := b"1111111111111111_1111111111111111_1111010011011000_1100110001000111"; -- -0.043566925689924214
	pesos_i(4505) := b"1111111111111111_1111111111111111_1110111011100000_1100011100110110"; -- -0.06688265734869667
	pesos_i(4506) := b"0000000000000000_0000000000000000_0000101000101010_1110010101011000"; -- 0.039717039041569216
	pesos_i(4507) := b"1111111111111111_1111111111111111_1110100100110101_1100001101000000"; -- -0.08902339640461675
	pesos_i(4508) := b"1111111111111111_1111111111111111_1111001111010110_0101000011000011"; -- -0.04751105527427291
	pesos_i(4509) := b"0000000000000000_0000000000000000_0001000110011110_0100000100011010"; -- 0.06882101896538982
	pesos_i(4510) := b"0000000000000000_0000000000000000_0001101100000110_0011101111001100"; -- 0.1055638670023112
	pesos_i(4511) := b"1111111111111111_1111111111111111_1111110110101100_0000010110011101"; -- -0.009093903811644044
	pesos_i(4512) := b"1111111111111111_1111111111111111_1110011100000101_0110110111011111"; -- -0.09757340718321089
	pesos_i(4513) := b"1111111111111111_1111111111111111_1111111111010111_1011001001110000"; -- -0.0006149746965194634
	pesos_i(4514) := b"0000000000000000_0000000000000000_0010101001100110_0011111001010000"; -- 0.1656226106715746
	pesos_i(4515) := b"0000000000000000_0000000000000000_0000101001111000_1011111100110100"; -- 0.04090495130428522
	pesos_i(4516) := b"0000000000000000_0000000000000000_0000011001001010_0111010111010011"; -- 0.024573673208351382
	pesos_i(4517) := b"1111111111111111_1111111111111111_1110101010101001_0101011011011100"; -- -0.08335358734521152
	pesos_i(4518) := b"0000000000000000_0000000000000000_0000000100011100_0100111010101010"; -- 0.004338184733112812
	pesos_i(4519) := b"1111111111111111_1111111111111111_1110101101011010_0010011100000000"; -- -0.08065563442469709
	pesos_i(4520) := b"1111111111111111_1111111111111111_1111101110101101_0011010101110110"; -- -0.016888292913445235
	pesos_i(4521) := b"0000000000000000_0000000000000000_0001100011010100_0001010110110110"; -- 0.09698615730091716
	pesos_i(4522) := b"1111111111111111_1111111111111111_1111011100110010_0011100010000000"; -- -0.03438994289834129
	pesos_i(4523) := b"0000000000000000_0000000000000000_0001001110000010_1100100100101001"; -- 0.07621438266311399
	pesos_i(4524) := b"0000000000000000_0000000000000000_0001001100100000_1010110100111000"; -- 0.07471735594782154
	pesos_i(4525) := b"0000000000000000_0000000000000000_0010010100100010_0101010000010001"; -- 0.14505505961739143
	pesos_i(4526) := b"0000000000000000_0000000000000000_0010100001110100_1110010110001010"; -- 0.15803370113553042
	pesos_i(4527) := b"1111111111111111_1111111111111111_1110110001000001_0001101101010100"; -- -0.07713154975577807
	pesos_i(4528) := b"1111111111111111_1111111111111111_1110111000001011_1100111011010001"; -- -0.0701323261554796
	pesos_i(4529) := b"1111111111111111_1111111111111111_1111111100111100_0010101101101001"; -- -0.002988135271425915
	pesos_i(4530) := b"1111111111111111_1111111111111111_1111111000011110_0001001011110011"; -- -0.007353606951364958
	pesos_i(4531) := b"1111111111111111_1111111111111111_1110001100100000_1111001000110111"; -- -0.11277853162857614
	pesos_i(4532) := b"0000000000000000_0000000000000000_0001010000101110_0010001100011111"; -- 0.07882899757289798
	pesos_i(4533) := b"0000000000000000_0000000000000000_0000010101110000_0000101011100100"; -- 0.02124088339954264
	pesos_i(4534) := b"1111111111111111_1111111111111111_1111101110100100_0100010010111010"; -- -0.01702471227016838
	pesos_i(4535) := b"1111111111111111_1111111111111111_1111110000010011_1010010000011001"; -- -0.015325301925794167
	pesos_i(4536) := b"0000000000000000_0000000000000000_0000000100001111_0000000101001010"; -- 0.004135208728471063
	pesos_i(4537) := b"1111111111111111_1111111111111111_1110101001110010_1000101011111000"; -- -0.08418971495925076
	pesos_i(4538) := b"1111111111111111_1111111111111111_1111110010000100_0011000010111001"; -- -0.013607935796535757
	pesos_i(4539) := b"1111111111111111_1111111111111111_1111100101110000_1100101101101010"; -- -0.025622641150091597
	pesos_i(4540) := b"1111111111111111_1111111111111111_1101011101111110_0101000000110000"; -- -0.1582288631314048
	pesos_i(4541) := b"1111111111111111_1111111111111111_1110100100010011_1110000001001001"; -- -0.08954046467429626
	pesos_i(4542) := b"0000000000000000_0000000000000000_0001101010110011_0011000011110110"; -- 0.10429674155541961
	pesos_i(4543) := b"0000000000000000_0000000000000000_0000110010101110_1101010110111101"; -- 0.049542769141950875
	pesos_i(4544) := b"1111111111111111_1111111111111111_1111101111110100_0010010100010111"; -- -0.01580589465697302
	pesos_i(4545) := b"1111111111111111_1111111111111111_1111101100110000_0101111011011001"; -- -0.018793174653809582
	pesos_i(4546) := b"1111111111111111_1111111111111111_1101101111101001_1111001110111011"; -- -0.14096142461905237
	pesos_i(4547) := b"0000000000000000_0000000000000000_0001101100111011_0001101101110101"; -- 0.10637065511664404
	pesos_i(4548) := b"1111111111111111_1111111111111111_1101110011000100_1011010100011000"; -- -0.13762348335157454
	pesos_i(4549) := b"0000000000000000_0000000000000000_0001001110111010_1111101100111110"; -- 0.07707185999657393
	pesos_i(4550) := b"1111111111111111_1111111111111111_1111010100100111_1110111001100000"; -- -0.04235944890405383
	pesos_i(4551) := b"1111111111111111_1111111111111111_1110010000111010_1011011000011000"; -- -0.10847913660539683
	pesos_i(4552) := b"1111111111111111_1111111111111111_1101110101010111_0001111011001100"; -- -0.13538939977027142
	pesos_i(4553) := b"0000000000000000_0000000000000000_0001101110001111_1100111101101111"; -- 0.1076631207536472
	pesos_i(4554) := b"1111111111111111_1111111111111111_1101101110011111_0000011110101101"; -- -0.14210464511752285
	pesos_i(4555) := b"1111111111111111_1111111111111111_1110010011100011_0111110010110000"; -- -0.1059038228874573
	pesos_i(4556) := b"1111111111111111_1111111111111111_1110101110001001_1111101010110101"; -- -0.07992585262876438
	pesos_i(4557) := b"1111111111111111_1111111111111111_1110000011011011_1110010101101000"; -- -0.12164465158347237
	pesos_i(4558) := b"0000000000000000_0000000000000000_0001111001111000_0000000100010100"; -- 0.11901861900668279
	pesos_i(4559) := b"1111111111111111_1111111111111111_1101101101101000_1001011011110010"; -- -0.14293533896142574
	pesos_i(4560) := b"1111111111111111_1111111111111111_1101101110011010_0010000000111100"; -- -0.14217947513178422
	pesos_i(4561) := b"1111111111111111_1111111111111111_1110110000001001_0010110000000000"; -- -0.07798504838129948
	pesos_i(4562) := b"0000000000000000_0000000000000000_0001000101111011_1111011101000010"; -- 0.06829781881765862
	pesos_i(4563) := b"0000000000000000_0000000000000000_0010001111111110_0111000010001100"; -- 0.14060119076117947
	pesos_i(4564) := b"0000000000000000_0000000000000000_0000001001111101_1000001001000000"; -- 0.00972761223761414
	pesos_i(4565) := b"0000000000000000_0000000000000000_0000111101010101_1000010111100011"; -- 0.05989872742832342
	pesos_i(4566) := b"1111111111111111_1111111111111111_1101100000000110_1111011000001001"; -- -0.156143782352257
	pesos_i(4567) := b"0000000000000000_0000000000000000_0010111100000001_1110100011101001"; -- 0.18362289141285723
	pesos_i(4568) := b"0000000000000000_0000000000000000_0001001001100000_0101000001011011"; -- 0.07178213333281831
	pesos_i(4569) := b"0000000000000000_0000000000000000_0000101110010100_1010111110000100"; -- 0.04523751238555337
	pesos_i(4570) := b"1111111111111111_1111111111111111_1101110110000101_1100111001111100"; -- -0.1346770235839781
	pesos_i(4571) := b"0000000000000000_0000000000000000_0000111001111011_0010000011010011"; -- 0.056566287510634285
	pesos_i(4572) := b"1111111111111111_1111111111111111_1101110101011100_1001001100011010"; -- -0.13530617339868356
	pesos_i(4573) := b"1111111111111111_1111111111111111_1111111100001110_0011001001101101"; -- -0.00368962145429355
	pesos_i(4574) := b"0000000000000000_0000000000000000_0001100101100000_1010110000100001"; -- 0.09913135333544651
	pesos_i(4575) := b"1111111111111111_1111111111111111_1110001111000110_0010111100111000"; -- -0.11025719537027939
	pesos_i(4576) := b"1111111111111111_1111111111111111_1101010001100000_0100001011011101"; -- -0.17040617099245764
	pesos_i(4577) := b"0000000000000000_0000000000000000_0010100000111111_0101101001001110"; -- 0.15721668629885155
	pesos_i(4578) := b"0000000000000000_0000000000000000_0010001110010110_1000001111011111"; -- 0.13901542850033732
	pesos_i(4579) := b"1111111111111111_1111111111111111_1111111011010011_0101011110111000"; -- -0.004587667120342853
	pesos_i(4580) := b"0000000000000000_0000000000000000_0000000111100001_0110101001110100"; -- 0.007345822678088715
	pesos_i(4581) := b"1111111111111111_1111111111111111_1101011100010101_1001111010110111"; -- -0.1598263552865969
	pesos_i(4582) := b"0000000000000000_0000000000000000_0001100001101001_1000000111010100"; -- 0.09535991113041917
	pesos_i(4583) := b"0000000000000000_0000000000000000_0010001000010011_1011100111101100"; -- 0.13311349886652232
	pesos_i(4584) := b"0000000000000000_0000000000000000_0010011111010000_0000000110010101"; -- 0.1555176725149117
	pesos_i(4585) := b"0000000000000000_0000000000000000_0010001011000010_1011100011111111"; -- 0.13578373173807626
	pesos_i(4586) := b"1111111111111111_1111111111111111_1111100110100001_1101101100111000"; -- -0.02487401852458598
	pesos_i(4587) := b"0000000000000000_0000000000000000_0010010010110110_1100101100010111"; -- 0.14341420470788682
	pesos_i(4588) := b"1111111111111111_1111111111111111_1110101100010101_0011110100111000"; -- -0.081707166544519
	pesos_i(4589) := b"1111111111111111_1111111111111111_1101011001110100_1101100001001000"; -- -0.16227958898720493
	pesos_i(4590) := b"0000000000000000_0000000000000000_0000001010101111_1111010101010001"; -- 0.01049741005518659
	pesos_i(4591) := b"1111111111111111_1111111111111111_1101011100010001_1000010100010010"; -- -0.15988891897926885
	pesos_i(4592) := b"1111111111111111_1111111111111111_1111101110010001_0100100011100011"; -- -0.01731438112232292
	pesos_i(4593) := b"1111111111111111_1111111111111111_1110101011111101_0100111010010110"; -- -0.08207234220885297
	pesos_i(4594) := b"1111111111111111_1111111111111111_1101110010010101_1011110000001110"; -- -0.13834023147842736
	pesos_i(4595) := b"0000000000000000_0000000000000000_0000100111101010_1110011101000111"; -- 0.03874059178892123
	pesos_i(4596) := b"1111111111111111_1111111111111111_1111111011011010_1011011110100101"; -- -0.004475137939586669
	pesos_i(4597) := b"1111111111111111_1111111111111111_1111111000010101_0011010010111111"; -- -0.007488921420023271
	pesos_i(4598) := b"0000000000000000_0000000000000000_0001110000101000_0110010001110100"; -- 0.10999133910142023
	pesos_i(4599) := b"0000000000000000_0000000000000000_0001100000101001_0101001010101000"; -- 0.09438053696592226
	pesos_i(4600) := b"0000000000000000_0000000000000000_0010100011101010_0010010100001011"; -- 0.15982276455453645
	pesos_i(4601) := b"1111111111111111_1111111111111111_1110111101100101_1111110110011010"; -- -0.0648499965084788
	pesos_i(4602) := b"1111111111111111_1111111111111111_1111110100100010_1000001110001011"; -- -0.011192110656552748
	pesos_i(4603) := b"1111111111111111_1111111111111111_1110011010011000_1000010111000000"; -- -0.09923519193572196
	pesos_i(4604) := b"0000000000000000_0000000000000000_0001111000010001_1011110111011100"; -- 0.11745821592839725
	pesos_i(4605) := b"0000000000000000_0000000000000000_0010010001100000_0111000100110001"; -- 0.14209659044408637
	pesos_i(4606) := b"1111111111111111_1111111111111111_1110100000110101_1110011110000001"; -- -0.09292748535832
	pesos_i(4607) := b"0000000000000000_0000000000000000_0000010111111100_0110100111000101"; -- 0.02338276924512921
	pesos_i(4608) := b"1111111111111111_1111111111111111_1101100011101011_1010111111010001"; -- -0.15265370517441282
	pesos_i(4609) := b"0000000000000000_0000000000000000_0010000000101000_1010011011101101"; -- 0.1256203012027827
	pesos_i(4610) := b"1111111111111111_1111111111111111_1110101010010000_0111000011110010"; -- -0.0837335022002133
	pesos_i(4611) := b"0000000000000000_0000000000000000_0001010101011011_0001001010110111"; -- 0.08342091537556089
	pesos_i(4612) := b"0000000000000000_0000000000000000_0001111001111010_1110110110000110"; -- 0.11906322979554865
	pesos_i(4613) := b"0000000000000000_0000000000000000_0010100010100100_1000110010100100"; -- 0.15876082414145057
	pesos_i(4614) := b"1111111111111111_1111111111111111_1101101101101110_1000010111100100"; -- -0.14284480259974824
	pesos_i(4615) := b"1111111111111111_1111111111111111_1101100100110101_0101000110010101"; -- -0.1515301716099157
	pesos_i(4616) := b"0000000000000000_0000000000000000_0000001100111010_1001110001100001"; -- 0.012613080664071453
	pesos_i(4617) := b"1111111111111111_1111111111111111_1111110011111110_1000100001010110"; -- -0.011741141294155908
	pesos_i(4618) := b"0000000000000000_0000000000000000_0010000000000100_0110011011101001"; -- 0.12506716907667048
	pesos_i(4619) := b"0000000000000000_0000000000000000_0010100000111100_0011111110011000"; -- 0.15716931789425206
	pesos_i(4620) := b"0000000000000000_0000000000000000_0010100111010010_0101011100101000"; -- 0.16336579056145692
	pesos_i(4621) := b"1111111111111111_1111111111111111_1110001101011001_1110111110000011"; -- -0.11190894167326998
	pesos_i(4622) := b"0000000000000000_0000000000000000_0001111101111111_0111001000111001"; -- 0.12303842445527484
	pesos_i(4623) := b"1111111111111111_1111111111111111_1111011110000101_0100111110001100"; -- -0.03312208978037151
	pesos_i(4624) := b"0000000000000000_0000000000000000_0000110100111100_1010011111111011"; -- 0.05170678984479482
	pesos_i(4625) := b"0000000000000000_0000000000000000_0010010000010100_0001011111010101"; -- 0.14093159633504598
	pesos_i(4626) := b"1111111111111111_1111111111111111_1111011101100011_1101100001111111"; -- -0.03363272577763082
	pesos_i(4627) := b"1111111111111111_1111111111111111_1101001100101111_0100011011111011"; -- -0.1750598561389139
	pesos_i(4628) := b"1111111111111111_1111111111111111_1110000010011010_0000000101110100"; -- -0.1226500598012654
	pesos_i(4629) := b"1111111111111111_1111111111111111_1111001000010010_0101001000010010"; -- -0.054407950088540415
	pesos_i(4630) := b"1111111111111111_1111111111111111_1110011010101001_0111101010011100"; -- -0.0989764565919543
	pesos_i(4631) := b"0000000000000000_0000000000000000_0011111111101111_0001000110011010"; -- 0.24974164961230166
	pesos_i(4632) := b"1111111111111111_1111111111111111_1110000101001101_1110110110000011"; -- -0.11990466654099873
	pesos_i(4633) := b"0000000000000000_0000000000000000_0000101111111001_1001101001100110"; -- 0.046777391235208375
	pesos_i(4634) := b"1111111111111111_1111111111111111_1110000110101000_0110010111101000"; -- -0.11852419927114698
	pesos_i(4635) := b"1111111111111111_1111111111111111_1101100000111111_1001100100110010"; -- -0.15527956512797086
	pesos_i(4636) := b"0000000000000000_0000000000000000_0010001111000000_0001110110010010"; -- 0.1396502000572939
	pesos_i(4637) := b"1111111111111111_1111111111111111_1101000110110101_0100000100001110"; -- -0.18082803157523758
	pesos_i(4638) := b"1111111111111111_1111111111111111_1110000010110010_1000001011010101"; -- -0.12227613743867334
	pesos_i(4639) := b"0000000000000000_0000000000000000_0010101101010110_1101110000100100"; -- 0.16929412729889684
	pesos_i(4640) := b"1111111111111111_1111111111111111_1101111010010011_0011011011101001"; -- -0.1305661851708152
	pesos_i(4641) := b"0000000000000000_0000000000000000_0010001000111101_1000000100001101"; -- 0.1337509781296137
	pesos_i(4642) := b"1111111111111111_1111111111111111_1111011101100001_1001010110001001"; -- -0.033667234537231396
	pesos_i(4643) := b"1111111111111111_1111111111111111_1111011100111010_1110100001110101"; -- -0.034257384661798014
	pesos_i(4644) := b"1111111111111111_1111111111111111_1111011000010110_0100011110011000"; -- -0.0387225393311148
	pesos_i(4645) := b"1111111111111111_1111111111111111_1111011101101101_1100110011000010"; -- -0.033480837391992695
	pesos_i(4646) := b"1111111111111111_1111111111111111_1101100110101010_0011001101111010"; -- -0.14974668762583895
	pesos_i(4647) := b"0000000000000000_0000000000000000_0001100111100000_0011000001000100"; -- 0.1010770955193642
	pesos_i(4648) := b"1111111111111111_1111111111111111_1110101111000111_0001100011010110"; -- -0.07899327059091604
	pesos_i(4649) := b"1111111111111111_1111111111111111_1101001100111100_1110000111011010"; -- -0.1748522609513582
	pesos_i(4650) := b"1111111111111111_1111111111111111_1110101101111000_1101001100001111"; -- -0.08018761523160495
	pesos_i(4651) := b"1111111111111111_1111111111111111_1111111010101001_1010101110000000"; -- -0.005223542441994021
	pesos_i(4652) := b"0000000000000000_0000000000000000_0010001100111100_1100111000011010"; -- 0.13764656184052568
	pesos_i(4653) := b"0000000000000000_0000000000000000_0010011110010100_0110011101100101"; -- 0.15460821357626053
	pesos_i(4654) := b"1111111111111111_1111111111111111_1101111010010101_1100100111010110"; -- -0.1305269101630323
	pesos_i(4655) := b"0000000000000000_0000000000000000_0010110010110011_0010101010101001"; -- 0.17460886601433767
	pesos_i(4656) := b"0000000000000000_0000000000000000_0010100100000110_0000100101001011"; -- 0.1602483565319223
	pesos_i(4657) := b"0000000000000000_0000000000000000_0000100000000011_0111011001000111"; -- 0.03130282618110983
	pesos_i(4658) := b"0000000000000000_0000000000000000_0001101010000000_1000000110101101"; -- 0.10352335427078849
	pesos_i(4659) := b"0000000000000000_0000000000000000_0000111110111001_0101111110010110"; -- 0.061422323448913456
	pesos_i(4660) := b"0000000000000000_0000000000000000_0010010011010001_1001001001101100"; -- 0.14382281426439783
	pesos_i(4661) := b"1111111111111111_1111111111111111_1110011000111100_1100101101000011"; -- -0.10063485740100266
	pesos_i(4662) := b"0000000000000000_0000000000000000_0000000110100000_1110000111001100"; -- 0.006361114721987685
	pesos_i(4663) := b"1111111111111111_1111111111111111_1110010101111110_0001001110000001"; -- -0.1035449800473184
	pesos_i(4664) := b"0000000000000000_0000000000000000_0010001010101101_0000100010011000"; -- 0.13545278268643093
	pesos_i(4665) := b"0000000000000000_0000000000000000_0001001011001011_1110111010001101"; -- 0.07342425281018314
	pesos_i(4666) := b"0000000000000000_0000000000000000_0010010000001000_1100100110001001"; -- 0.1407590828233445
	pesos_i(4667) := b"1111111111111111_1111111111111111_1110100110100000_0100100110000110"; -- -0.08739796143227263
	pesos_i(4668) := b"0000000000000000_0000000000000000_0000111101111010_1000110111100001"; -- 0.0604637788076539
	pesos_i(4669) := b"1111111111111111_1111111111111111_1110110011100010_1100000111011011"; -- -0.07466495888836688
	pesos_i(4670) := b"1111111111111111_1111111111111111_1111100000111011_0110010011001110"; -- -0.030343722999651195
	pesos_i(4671) := b"1111111111111111_1111111111111111_1110111100001111_0010001010011000"; -- -0.06617530617046483
	pesos_i(4672) := b"1111111111111111_1111111111111111_1110011000001101_1011101110010001"; -- -0.10135295599847474
	pesos_i(4673) := b"0000000000000000_0000000000000000_0001010000111011_1111110011100011"; -- 0.07904034186853896
	pesos_i(4674) := b"0000000000000000_0000000000000000_0001111100001101_0100110001100100"; -- 0.12129666740336659
	pesos_i(4675) := b"1111111111111111_1111111111111111_1110100111011111_0100100110011011"; -- -0.08643665285625331
	pesos_i(4676) := b"0000000000000000_0000000000000000_0001100011000010_1010011010111101"; -- 0.09672014355680544
	pesos_i(4677) := b"1111111111111111_1111111111111111_1110011110010010_0110101010101101"; -- -0.09542210837235938
	pesos_i(4678) := b"1111111111111111_1111111111111111_1111100001011011_0100111001001011"; -- -0.029856783620877174
	pesos_i(4679) := b"1111111111111111_1111111111111111_1101010000101100_1100100000110011"; -- -0.1711916804483558
	pesos_i(4680) := b"0000000000000000_0000000000000000_0010110010110010_0011000110110110"; -- 0.17459402747713407
	pesos_i(4681) := b"0000000000000000_0000000000000000_0001011000110100_1000011101111001"; -- 0.08673903177730162
	pesos_i(4682) := b"1111111111111111_1111111111111111_1110000110111111_1101100001011110"; -- -0.11816642471278309
	pesos_i(4683) := b"1111111111111111_1111111111111111_1111011000010100_0010101100100010"; -- -0.03875475334145909
	pesos_i(4684) := b"0000000000000000_0000000000000000_0000011110110101_1010101011100010"; -- 0.030115776179340012
	pesos_i(4685) := b"1111111111111111_1111111111111111_1110110010100000_1011111100001100"; -- -0.07567220641909775
	pesos_i(4686) := b"0000000000000000_0000000000000000_0010010010111101_0011010001011111"; -- 0.14351203263108062
	pesos_i(4687) := b"1111111111111111_1111111111111111_1110001000011111_1000101000010110"; -- -0.1167062470144463
	pesos_i(4688) := b"1111111111111111_1111111111111111_1101100001011011_1010111100111100"; -- -0.15485100530295406
	pesos_i(4689) := b"0000000000000000_0000000000000000_0000101010000111_1000101110111001"; -- 0.041130764729985565
	pesos_i(4690) := b"1111111111111111_1111111111111111_1101100101001111_1110011100011011"; -- -0.15112453067242554
	pesos_i(4691) := b"1111111111111111_1111111111111111_1101110000001010_1010100110000100"; -- -0.14046230829828224
	pesos_i(4692) := b"0000000000000000_0000000000000000_0000110011011101_1101110110111101"; -- 0.050260409126155
	pesos_i(4693) := b"1111111111111111_1111111111111111_1110111110001110_1101010001011001"; -- -0.06422684503588767
	pesos_i(4694) := b"0000000000000000_0000000000000000_0000001000101001_1000100101011001"; -- 0.008446296809270075
	pesos_i(4695) := b"0000000000000000_0000000000000000_0010010100100011_1010010111110110"; -- 0.14507519964529164
	pesos_i(4696) := b"0000000000000000_0000000000000000_0010101011111000_0000001010011001"; -- 0.16784683455163066
	pesos_i(4697) := b"0000000000000000_0000000000000000_0010010101101010_1011000010011001"; -- 0.14615920769240823
	pesos_i(4698) := b"1111111111111111_1111111111111111_1111001100001101_0001010100101111"; -- -0.05058162299675561
	pesos_i(4699) := b"1111111111111111_1111111111111111_1101110101101011_0010101111010111"; -- -0.13508344642112743
	pesos_i(4700) := b"1111111111111111_1111111111111111_1101111011110010_1101001110010110"; -- -0.12910726153531152
	pesos_i(4701) := b"1111111111111111_1111111111111111_1111110100010111_1011011101110111"; -- -0.011356862582738648
	pesos_i(4702) := b"0000000000000000_0000000000000000_0000000001101100_0111001101110110"; -- 0.0016548311209015362
	pesos_i(4703) := b"1111111111111111_1111111111111111_1110111010111000_1010001101111010"; -- -0.06749513877028625
	pesos_i(4704) := b"1111111111111111_1111111111111111_1101010100100100_0001110001111110"; -- -0.16741773530745757
	pesos_i(4705) := b"0000000000000000_0000000000000000_0010011100100101_0100101011011011"; -- 0.15291278692397112
	pesos_i(4706) := b"1111111111111111_1111111111111111_1110110001110101_0110010001001111"; -- -0.07633374293376982
	pesos_i(4707) := b"1111111111111111_1111111111111111_1110100110010111_1111011100000001"; -- -0.08752495032587908
	pesos_i(4708) := b"1111111111111111_1111111111111111_1110000110011110_0110001100001101"; -- -0.11867695737085235
	pesos_i(4709) := b"0000000000000000_0000000000000000_0000110110001010_1111101000011101"; -- 0.05290187073016792
	pesos_i(4710) := b"1111111111111111_1111111111111111_1110011111011100_0111000111111110"; -- -0.09429252205301157
	pesos_i(4711) := b"1111111111111111_1111111111111111_1111101111000101_0110110000011111"; -- -0.01651882396166779
	pesos_i(4712) := b"0000000000000000_0000000000000000_0000100000111000_0100110001010101"; -- 0.032109041910112296
	pesos_i(4713) := b"1111111111111111_1111111111111111_1110011101001001_1110000110111011"; -- -0.09652890379540652
	pesos_i(4714) := b"0000000000000000_0000000000000000_0000000000011011_1110111110010101"; -- 0.0004262675841864796
	pesos_i(4715) := b"0000000000000000_0000000000000000_0000011110110000_1101001001101100"; -- 0.0300418389640602
	pesos_i(4716) := b"0000000000000000_0000000000000000_0000011110000101_0011100100010110"; -- 0.02937657143199239
	pesos_i(4717) := b"0000000000000000_0000000000000000_0001000100110101_1101100010001111"; -- 0.06722787370993014
	pesos_i(4718) := b"1111111111111111_1111111111111111_1101110100100111_0111001000110101"; -- -0.1361168499150716
	pesos_i(4719) := b"1111111111111111_1111111111111111_1111110101111011_1101010110110100"; -- -0.009829181190207899
	pesos_i(4720) := b"0000000000000000_0000000000000000_0010011110010101_1001011001010011"; -- 0.15462626965079843
	pesos_i(4721) := b"1111111111111111_1111111111111111_1110101001111001_0110001101001110"; -- -0.08408526744414839
	pesos_i(4722) := b"1111111111111111_1111111111111111_1110110010111010_0001010000010000"; -- -0.07528566950576307
	pesos_i(4723) := b"0000000000000000_0000000000000000_0010010001001000_0011110101110011"; -- 0.1417272955595422
	pesos_i(4724) := b"0000000000000000_0000000000000000_0000010100000011_0100000110000111"; -- 0.019580932022067888
	pesos_i(4725) := b"1111111111111111_1111111111111111_1111101011110100_0110000000001101"; -- -0.019708630415659623
	pesos_i(4726) := b"0000000000000000_0000000000000000_0001101011101100_0011010000010000"; -- 0.10516667736517417
	pesos_i(4727) := b"1111111111111111_1111111111111111_1110000111010111_0000110010010111"; -- -0.11781235990142906
	pesos_i(4728) := b"0000000000000000_0000000000000000_0000111000111000_1111111001110100"; -- 0.055557158805450424
	pesos_i(4729) := b"0000000000000000_0000000000000000_0000011011100110_0111101010100010"; -- 0.02695433090079886
	pesos_i(4730) := b"0000000000000000_0000000000000000_0000111010001011_1011111110101001"; -- 0.05681989548937032
	pesos_i(4731) := b"0000000000000000_0000000000000000_0001010101101110_0011100001001001"; -- 0.08371307168492638
	pesos_i(4732) := b"1111111111111111_1111111111111111_1111001000100001_0100111110001011"; -- -0.05417921882074122
	pesos_i(4733) := b"1111111111111111_1111111111111111_1110001000011111_1011000010100101"; -- -0.11670394865663727
	pesos_i(4734) := b"1111111111111111_1111111111111111_1111010000111100_1001000101001010"; -- -0.045950812802530265
	pesos_i(4735) := b"0000000000000000_0000000000000000_0001010111101010_1010001110011011"; -- 0.08561155823593594
	pesos_i(4736) := b"0000000000000000_0000000000000000_0010100101011111_0001001111011111"; -- 0.16160701929175544
	pesos_i(4737) := b"0000000000000000_0000000000000000_0001100001010011_1001011100010100"; -- 0.09502548454723803
	pesos_i(4738) := b"0000000000000000_0000000000000000_0001001101000110_1101001000110111"; -- 0.0752993950225239
	pesos_i(4739) := b"0000000000000000_0000000000000000_0010100111010010_0010001000100010"; -- 0.1633626302193313
	pesos_i(4740) := b"0000000000000000_0000000000000000_0001001010110001_0010000001000000"; -- 0.07301522786187456
	pesos_i(4741) := b"0000000000000000_0000000000000000_0010001100110010_1001010000101000"; -- 0.13749052029243605
	pesos_i(4742) := b"1111111111111111_1111111111111111_1101111000010110_1110100101010101"; -- -0.13246289905519537
	pesos_i(4743) := b"1111111111111111_1111111111111111_1111111010000100_1010010001111110"; -- -0.0057885354157704285
	pesos_i(4744) := b"0000000000000000_0000000000000000_0000101001001000_1100010110001001"; -- 0.04017290672471124
	pesos_i(4745) := b"1111111111111111_1111111111111111_1110100011101011_0100100001111001"; -- -0.0901598649709397
	pesos_i(4746) := b"0000000000000000_0000000000000000_0010100110011001_1100000011011000"; -- 0.1625023391812109
	pesos_i(4747) := b"1111111111111111_1111111111111111_1110111011100111_1011001100110001"; -- -0.06677703907005283
	pesos_i(4748) := b"1111111111111111_1111111111111111_1110011001100110_0111110000111110"; -- -0.0999986980840781
	pesos_i(4749) := b"0000000000000000_0000000000000000_0000111001001000_1000101101100111"; -- 0.05579444177707601
	pesos_i(4750) := b"0000000000000000_0000000000000000_0001111000110101_0100111111011001"; -- 0.11800097500509328
	pesos_i(4751) := b"0000000000000000_0000000000000000_0001010011111101_1000100011100001"; -- 0.08199363228646304
	pesos_i(4752) := b"1111111111111111_1111111111111111_1111111000010111_0101001110001101"; -- -0.0074565678154139
	pesos_i(4753) := b"1111111111111111_1111111111111111_1111011111000011_1110101110110110"; -- -0.03216673661858794
	pesos_i(4754) := b"0000000000000000_0000000000000000_0010000110110100_1001110110011101"; -- 0.13166222644430267
	pesos_i(4755) := b"1111111111111111_1111111111111111_1110110100111001_0100001001011010"; -- -0.07334504414418166
	pesos_i(4756) := b"1111111111111111_1111111111111111_1110001000100110_1110100000000100"; -- -0.11659383676902814
	pesos_i(4757) := b"0000000000000000_0000000000000000_0010001100000001_0111111010101010"; -- 0.13674155864104803
	pesos_i(4758) := b"0000000000000000_0000000000000000_0001101000110111_1001000000100110"; -- 0.10241032538126824
	pesos_i(4759) := b"0000000000000000_0000000000000000_0001011000000010_0011111001100110"; -- 0.08597173688173022
	pesos_i(4760) := b"0000000000000000_0000000000000000_0000100111110101_1011110101110101"; -- 0.038905945873443114
	pesos_i(4761) := b"0000000000000000_0000000000000000_0010000000011010_1111110111110111"; -- 0.1254118660514932
	pesos_i(4762) := b"1111111111111111_1111111111111111_1101111100100101_0111011111001001"; -- -0.12833453512586868
	pesos_i(4763) := b"1111111111111111_1111111111111111_1101001000010001_0010000010011000"; -- -0.17942615779059476
	pesos_i(4764) := b"0000000000000000_0000000000000000_0001001101001110_1110000100000101"; -- 0.07542234768388854
	pesos_i(4765) := b"1111111111111111_1111111111111111_1101101111001101_1101100110001011"; -- -0.14139023171888734
	pesos_i(4766) := b"1111111111111111_1111111111111111_1101101001010110_0001111100100110"; -- -0.14712338761239113
	pesos_i(4767) := b"0000000000000000_0000000000000000_0010000101110101_0000100111011011"; -- 0.1306921157356922
	pesos_i(4768) := b"1111111111111111_1111111111111111_1111011100010110_1011110001101110"; -- -0.03480932527083663
	pesos_i(4769) := b"0000000000000000_0000000000000000_0000100011100111_1110100001001011"; -- 0.03478862591244446
	pesos_i(4770) := b"0000000000000000_0000000000000000_0010101010111011_1101011000010101"; -- 0.16692865388594735
	pesos_i(4771) := b"1111111111111111_1111111111111111_1110110101101111_1101110111001100"; -- -0.07251180423127705
	pesos_i(4772) := b"1111111111111111_1111111111111111_1111000011101111_1011111000100001"; -- -0.05884181685858914
	pesos_i(4773) := b"1111111111111111_1111111111111111_1111111111011011_0010010000011010"; -- -0.0005624233839681802
	pesos_i(4774) := b"1111111111111111_1111111111111111_1111011100100100_1111100100011111"; -- -0.03459208470446396
	pesos_i(4775) := b"0000000000000000_0000000000000000_0010011001000000_0111001001101010"; -- 0.14942088214679497
	pesos_i(4776) := b"0000000000000000_0000000000000000_0000000001001000_0101100010001111"; -- 0.0011039114157657404
	pesos_i(4777) := b"1111111111111111_1111111111111111_1110111011001001_0101101010000000"; -- -0.06724008907118283
	pesos_i(4778) := b"0000000000000000_0000000000000000_0010101111111111_1110100000011011"; -- 0.17187357578917287
	pesos_i(4779) := b"0000000000000000_0000000000000000_0001101010010111_0001101110010001"; -- 0.10386822014311214
	pesos_i(4780) := b"1111111111111111_1111111111111111_1111111011001110_1001100101111111"; -- -0.004660040300031891
	pesos_i(4781) := b"0000000000000000_0000000000000000_0001010100110011_0100100010000011"; -- 0.08281377017012297
	pesos_i(4782) := b"0000000000000000_0000000000000000_0001101001010100_0011010110100011"; -- 0.1028474352951361
	pesos_i(4783) := b"1111111111111111_1111111111111111_1110111000011011_0101110100111111"; -- -0.0698949547102013
	pesos_i(4784) := b"1111111111111111_1111111111111111_1101001011110011_1110110100101101"; -- -0.17596547745109897
	pesos_i(4785) := b"1111111111111111_1111111111111111_1111011000000000_1101000111111001"; -- -0.039049984587644866
	pesos_i(4786) := b"0000000000000000_0000000000000000_0001011010111111_1110001011000100"; -- 0.08886544493548224
	pesos_i(4787) := b"1111111111111111_1111111111111111_1110100001100100_1000101101101011"; -- -0.09221581117981996
	pesos_i(4788) := b"0000000000000000_0000000000000000_0010100001110010_1001110010100010"; -- 0.15799883793824834
	pesos_i(4789) := b"0000000000000000_0000000000000000_0000110100000011_0010111100000001"; -- 0.05082982800799485
	pesos_i(4790) := b"0000000000000000_0000000000000000_0001001101000001_1011010100000101"; -- 0.07522136099368125
	pesos_i(4791) := b"1111111111111111_1111111111111111_1101110100111100_1000000101100000"; -- -0.13579551138555618
	pesos_i(4792) := b"1111111111111111_1111111111111111_1110100010010101_0101000100000110"; -- -0.09147161116884377
	pesos_i(4793) := b"1111111111111111_1111111111111111_1111011111101110_0000001011100111"; -- -0.03152448517426139
	pesos_i(4794) := b"0000000000000000_0000000000000000_0010100010011111_0101001100101011"; -- 0.15868110472626448
	pesos_i(4795) := b"1111111111111111_1111111111111111_1111010000011001_1010100111111010"; -- -0.04648339883464944
	pesos_i(4796) := b"1111111111111111_1111111111111111_1101110011011000_1011011110011011"; -- -0.1373181579271746
	pesos_i(4797) := b"1111111111111111_1111111111111111_1101100110010110_0111111011101011"; -- -0.15004736679415154
	pesos_i(4798) := b"0000000000000000_0000000000000000_0010100111111101_1000111000100010"; -- 0.1640251954417713
	pesos_i(4799) := b"0000000000000000_0000000000000000_0000000101011001_0111010001111110"; -- 0.0052712256562644525
	pesos_i(4800) := b"0000000000000000_0000000000000000_0010000000011110_0001010000011101"; -- 0.1254589624049923
	pesos_i(4801) := b"0000000000000000_0000000000000000_0010000100010000_1010010010100101"; -- 0.12916020412907916
	pesos_i(4802) := b"0000000000000000_0000000000000000_0001101000110100_1101100000100111"; -- 0.10236884059963437
	pesos_i(4803) := b"1111111111111111_1111111111111111_1111111010000100_0111011100111101"; -- -0.0057912325944731655
	pesos_i(4804) := b"0000000000000000_0000000000000000_0001010111111000_0100010001001010"; -- 0.08581950012815094
	pesos_i(4805) := b"1111111111111111_1111111111111111_1101010010010100_1000010111010110"; -- -0.1696087219592115
	pesos_i(4806) := b"1111111111111111_1111111111111111_1111100101101010_0011110111110001"; -- -0.02572262629053747
	pesos_i(4807) := b"0000000000000000_0000000000000000_0000111101000001_0111001101111011"; -- 0.05959245441148006
	pesos_i(4808) := b"0000000000000000_0000000000000000_0000100111000011_1001111101001100"; -- 0.038141208593419657
	pesos_i(4809) := b"1111111111111111_1111111111111111_1111001000000001_1100100000011010"; -- -0.054660314248523044
	pesos_i(4810) := b"1111111111111111_1111111111111111_1110100001011010_1111011111010000"; -- -0.09236193831907939
	pesos_i(4811) := b"1111111111111111_1111111111111111_1111111111001101_0010110010111101"; -- -0.000775531642371012
	pesos_i(4812) := b"0000000000000000_0000000000000000_0010000001010000_0100011001101011"; -- 0.12622490031643435
	pesos_i(4813) := b"1111111111111111_1111111111111111_1101110000100011_1100011111100110"; -- -0.14007902761427515
	pesos_i(4814) := b"1111111111111111_1111111111111111_1101110101011000_1111100101111001"; -- -0.13536110674955518
	pesos_i(4815) := b"0000000000000000_0000000000000000_0000110101010011_1001011001011010"; -- 0.052056691036602105
	pesos_i(4816) := b"1111111111111111_1111111111111111_1101010000101101_1000011000000111"; -- -0.1711803657691644
	pesos_i(4817) := b"0000000000000000_0000000000000000_0010000101100011_1111010111110100"; -- 0.1304315300509886
	pesos_i(4818) := b"0000000000000000_0000000000000000_0010110000111000_0101010111110100"; -- 0.17273461534712706
	pesos_i(4819) := b"1111111111111111_1111111111111111_1110011110001100_1110100001000000"; -- -0.09550617644126867
	pesos_i(4820) := b"1111111111111111_1111111111111111_1110011010001010_0100001011000110"; -- -0.09945280709096033
	pesos_i(4821) := b"1111111111111111_1111111111111111_1111110111111011_0001011011100010"; -- -0.00788742995261705
	pesos_i(4822) := b"1111111111111111_1111111111111111_1101110001000010_1101111011101011"; -- -0.13960463292788658
	pesos_i(4823) := b"0000000000000000_0000000000000000_0011001001100110_1011000111110000"; -- 0.19687950231187507
	pesos_i(4824) := b"1111111111111111_1111111111111111_1111000010010110_1001100100010000"; -- -0.06020205844699915
	pesos_i(4825) := b"1111111111111111_1111111111111111_1111100111111000_0000111000001110"; -- -0.023558732682100382
	pesos_i(4826) := b"1111111111111111_1111111111111111_1110010001110110_0111010010110010"; -- -0.10756750733692685
	pesos_i(4827) := b"0000000000000000_0000000000000000_0001111100111001_0010110011111111"; -- 0.12196618295254509
	pesos_i(4828) := b"0000000000000000_0000000000000000_0010101011011100_1011011111001001"; -- 0.16743038811102146
	pesos_i(4829) := b"1111111111111111_1111111111111111_1111010100001000_1011100110000010"; -- -0.04283562261154984
	pesos_i(4830) := b"1111111111111111_1111111111111111_1111101110110011_1100100010011000"; -- -0.01678797048360721
	pesos_i(4831) := b"0000000000000000_0000000000000000_0010001101110001_0010010001000010"; -- 0.13844515430758506
	pesos_i(4832) := b"0000000000000000_0000000000000000_0010000000100100_1111110111111001"; -- 0.12556445442422096
	pesos_i(4833) := b"0000000000000000_0000000000000000_0001001000000110_0110001011100110"; -- 0.07040994746268991
	pesos_i(4834) := b"0000000000000000_0000000000000000_0010011001011011_0111100001001010"; -- 0.1498332195328398
	pesos_i(4835) := b"0000000000000000_0000000000000000_0000101011011110_1011001001011111"; -- 0.042460582921320995
	pesos_i(4836) := b"0000000000000000_0000000000000000_0000100011001000_0101100111101110"; -- 0.0343071180696885
	pesos_i(4837) := b"1111111111111111_1111111111111111_1111000001110101_0101110110111101"; -- -0.060709134547807436
	pesos_i(4838) := b"0000000000000000_0000000000000000_0000101111011000_1100110110010101"; -- 0.046276902007780674
	pesos_i(4839) := b"0000000000000000_0000000000000000_0010001101101111_1011110101011001"; -- 0.13842376166355244
	pesos_i(4840) := b"0000000000000000_0000000000000000_0001100011001101_1000111100111101"; -- 0.0968865893629032
	pesos_i(4841) := b"0000000000000000_0000000000000000_0000000111011110_0100101010000001"; -- 0.007298142020400872
	pesos_i(4842) := b"0000000000000000_0000000000000000_0000101111011100_1000010111010011"; -- 0.04633366015974773
	pesos_i(4843) := b"1111111111111111_1111111111111111_1110011010111001_1011011110001001"; -- -0.09872868444332374
	pesos_i(4844) := b"0000000000000000_0000000000000000_0001011111110101_0101110110001000"; -- 0.09358772820024107
	pesos_i(4845) := b"1111111111111111_1111111111111111_1110001011001111_0111111011010001"; -- -0.11402137190168536
	pesos_i(4846) := b"1111111111111111_1111111111111111_1110111001010110_0001011111010110"; -- -0.0689988233870216
	pesos_i(4847) := b"1111111111111111_1111111111111111_1110010011000001_0000010001001001"; -- -0.10642979826253585
	pesos_i(4848) := b"1111111111111111_1111111111111111_1111110100101100_0010011100111000"; -- -0.011045025761629634
	pesos_i(4849) := b"0000000000000000_0000000000000000_0000000000011111_1011011101110010"; -- 0.00048395673911075655
	pesos_i(4850) := b"0000000000000000_0000000000000000_0010001000101010_0011101001100111"; -- 0.1334568500917844
	pesos_i(4851) := b"1111111111111111_1111111111111111_1101110111100001_0000111101101000"; -- -0.13328460426886138
	pesos_i(4852) := b"1111111111111111_1111111111111111_1110101101000001_1111111101001001"; -- -0.08102421247621261
	pesos_i(4853) := b"0000000000000000_0000000000000000_0001100000011100_0010101000000110"; -- 0.09417975084182796
	pesos_i(4854) := b"0000000000000000_0000000000000000_0010011111000110_1010111010010000"; -- 0.15537539504349748
	pesos_i(4855) := b"1111111111111111_1111111111111111_1110110010001101_1010100111011110"; -- -0.07596338595885836
	pesos_i(4856) := b"0000000000000000_0000000000000000_0010100001010011_1111010101100000"; -- 0.1575311050791842
	pesos_i(4857) := b"0000000000000000_0000000000000000_0001010011001110_1110101110001010"; -- 0.08128234982731422
	pesos_i(4858) := b"1111111111111111_1111111111111111_1110010111001101_0000100110111000"; -- -0.10234011897292969
	pesos_i(4859) := b"0000000000000000_0000000000000000_0001000011110101_1101010010011111"; -- 0.06625107656161937
	pesos_i(4860) := b"0000000000000000_0000000000000000_0001101100100011_0001110101010100"; -- 0.1060045556009841
	pesos_i(4861) := b"1111111111111111_1111111111111111_1110111001100101_0001011011011001"; -- -0.06877000057094974
	pesos_i(4862) := b"1111111111111111_1111111111111111_1110100101000110_0000011001001000"; -- -0.08877526044729615
	pesos_i(4863) := b"0000000000000000_0000000000000000_0000000001010111_0001011001110110"; -- 0.0013288534157173961
	pesos_i(4864) := b"0000000000000000_0000000000000000_0001011101011101_0101111100110011"; -- 0.09126849164473524
	pesos_i(4865) := b"0000000000000000_0000000000000000_0001001100111100_0011101001111101"; -- 0.07513776360684735
	pesos_i(4866) := b"1111111111111111_1111111111111111_1101011000010110_1111111100001101"; -- -0.16371160448846478
	pesos_i(4867) := b"1111111111111111_1111111111111111_1111100001100100_0011100101100010"; -- -0.029720700922274523
	pesos_i(4868) := b"0000000000000000_0000000000000000_0000100001101111_1010011001000000"; -- 0.03295363477103243
	pesos_i(4869) := b"0000000000000000_0000000000000000_0001100100100111_1110100111101010"; -- 0.09826528519430432
	pesos_i(4870) := b"1111111111111111_1111111111111111_1111110100001110_1000001011110100"; -- -0.011497321593689715
	pesos_i(4871) := b"1111111111111111_1111111111111111_1111110000111011_1101101100111000"; -- -0.01471166497734793
	pesos_i(4872) := b"1111111111111111_1111111111111111_1111010100011011_0100110111001101"; -- -0.04255212548501044
	pesos_i(4873) := b"1111111111111111_1111111111111111_1111111111000110_1101110000000001"; -- -0.0008718963964781766
	pesos_i(4874) := b"1111111111111111_1111111111111111_1110000100001100_1111110000100001"; -- -0.12089561656597726
	pesos_i(4875) := b"0000000000000000_0000000000000000_0000111001101001_0010110001111101"; -- 0.056292324511536734
	pesos_i(4876) := b"1111111111111111_1111111111111111_1110011001111000_0001100001111101"; -- -0.09972998573397578
	pesos_i(4877) := b"1111111111111111_1111111111111111_1110011001000010_0110111111010000"; -- -0.10054875532590979
	pesos_i(4878) := b"0000000000000000_0000000000000000_0000011010011011_0111000110001100"; -- 0.02580938024839123
	pesos_i(4879) := b"1111111111111111_1111111111111111_1110111010001100_1011000100100001"; -- -0.06816571175206952
	pesos_i(4880) := b"0000000000000000_0000000000000000_0010110010101111_0000100100001100"; -- 0.17454582723416492
	pesos_i(4881) := b"0000000000000000_0000000000000000_0001111101111101_0100110110111010"; -- 0.1230057314381978
	pesos_i(4882) := b"0000000000000000_0000000000000000_0010000011110001_0100110000111100"; -- 0.1286819121352003
	pesos_i(4883) := b"1111111111111111_1111111111111111_1111000010111010_0111010001001010"; -- -0.059654933912623546
	pesos_i(4884) := b"1111111111111111_1111111111111111_1101110100110100_1000010111011000"; -- -0.13591731518010788
	pesos_i(4885) := b"0000000000000000_0000000000000000_0001010111100111_1010010011000110"; -- 0.08556585163708473
	pesos_i(4886) := b"0000000000000000_0000000000000000_0010100100001110_0010101101100101"; -- 0.16037245960097918
	pesos_i(4887) := b"0000000000000000_0000000000000000_0010000111000101_0010000011010100"; -- 0.13191418804437638
	pesos_i(4888) := b"1111111111111111_1111111111111111_1111010000100001_1101100110010100"; -- -0.04635849131393675
	pesos_i(4889) := b"1111111111111111_1111111111111111_1111010110100110_1000011011110011"; -- -0.04042774732887216
	pesos_i(4890) := b"1111111111111111_1111111111111111_1111011111101101_0101100001110000"; -- -0.031534645766009554
	pesos_i(4891) := b"0000000000000000_0000000000000000_0001010010110010_1011101111000001"; -- 0.08085225546820593
	pesos_i(4892) := b"1111111111111111_1111111111111111_1111110000000010_1000100110110011"; -- -0.01558627488523715
	pesos_i(4893) := b"0000000000000000_0000000000000000_0000110001011000_0010011011100111"; -- 0.0482200920887886
	pesos_i(4894) := b"0000000000000000_0000000000000000_0000011000110001_0101100110110100"; -- 0.024190527424248418
	pesos_i(4895) := b"0000000000000000_0000000000000000_0010000101011010_0110110001001001"; -- 0.13028599530613746
	pesos_i(4896) := b"0000000000000000_0000000000000000_0000011010011001_1101111010100001"; -- 0.025785364559452434
	pesos_i(4897) := b"0000000000000000_0000000000000000_0001001001110000_1011011011010101"; -- 0.07203238190487357
	pesos_i(4898) := b"0000000000000000_0000000000000000_0000010010001100_1100111110100011"; -- 0.017773606686899143
	pesos_i(4899) := b"0000000000000000_0000000000000000_0001001000110110_1010011001001110"; -- 0.07114638718008903
	pesos_i(4900) := b"1111111111111111_1111111111111111_1110100011101000_1100110100110010"; -- -0.09019773037656952
	pesos_i(4901) := b"0000000000000000_0000000000000000_0000000011011100_0010100011001100"; -- 0.0033593652323780695
	pesos_i(4902) := b"1111111111111111_1111111111111111_1110111010010100_0100110000111000"; -- -0.06804965628548597
	pesos_i(4903) := b"0000000000000000_0000000000000000_0001110011000010_1011010110111000"; -- 0.11234603644135835
	pesos_i(4904) := b"0000000000000000_0000000000000000_0001001000100110_0010101001100001"; -- 0.07089485997149741
	pesos_i(4905) := b"1111111111111111_1111111111111111_1111001011100111_0100101110100101"; -- -0.05115821107436995
	pesos_i(4906) := b"0000000000000000_0000000000000000_0001000111000001_1101010000011011"; -- 0.06936383887400267
	pesos_i(4907) := b"1111111111111111_1111111111111111_1111101010110010_1000010100101000"; -- -0.02071349890943056
	pesos_i(4908) := b"1111111111111111_1111111111111111_1101011100101000_0001010011010010"; -- -0.15954465741425963
	pesos_i(4909) := b"0000000000000000_0000000000000000_0001001000000011_1001111110101010"; -- 0.070367793195875
	pesos_i(4910) := b"0000000000000000_0000000000000000_0010111010000111_0001000110100010"; -- 0.1817484876125213
	pesos_i(4911) := b"0000000000000000_0000000000000000_0010101000111111_0110111101010101"; -- 0.16503043963946235
	pesos_i(4912) := b"0000000000000000_0000000000000000_0001011001001111_1001110001000011"; -- 0.08715225819657527
	pesos_i(4913) := b"1111111111111111_1111111111111111_1111111111000001_0101111011001001"; -- -0.0009556540866678719
	pesos_i(4914) := b"1111111111111111_1111111111111111_1110101100110001_1001000111100110"; -- -0.08127487310043974
	pesos_i(4915) := b"0000000000000000_0000000000000000_0001110001101100_0111110110111111"; -- 0.11103044423068245
	pesos_i(4916) := b"0000000000000000_0000000000000000_0001100010001100_1100011011000000"; -- 0.09589807699518424
	pesos_i(4917) := b"0000000000000000_0000000000000000_0000011110010111_1100011111111110"; -- 0.029659747699035163
	pesos_i(4918) := b"1111111111111111_1111111111111111_1110111001110000_0010001010011110"; -- -0.06860145231900094
	pesos_i(4919) := b"1111111111111111_1111111111111111_1110000100001010_1111100101011100"; -- -0.1209262991437335
	pesos_i(4920) := b"0000000000000000_0000000000000000_0010100110010111_1011110101110100"; -- 0.16247161950674868
	pesos_i(4921) := b"1111111111111111_1111111111111111_1111101000110110_1100101110111110"; -- -0.022601381489407484
	pesos_i(4922) := b"1111111111111111_1111111111111111_1111110010100101_1010111101110111"; -- -0.013096841348229365
	pesos_i(4923) := b"1111111111111111_1111111111111111_1111001000000111_0010011011100100"; -- -0.054578370339473964
	pesos_i(4924) := b"0000000000000000_0000000000000000_0001010110010011_1110010000011110"; -- 0.08428788884393604
	pesos_i(4925) := b"0000000000000000_0000000000000000_0000000101110010_0101001011100100"; -- 0.00565069255038287
	pesos_i(4926) := b"0000000000000000_0000000000000000_0001101010100011_1000011011110011"; -- 0.10405772630609347
	pesos_i(4927) := b"0000000000000000_0000000000000000_0000011101101011_1111010101000111"; -- 0.0289910600312234
	pesos_i(4928) := b"0000000000000000_0000000000000000_0001010001111011_1110000011000011"; -- 0.08001522788836726
	pesos_i(4929) := b"0000000000000000_0000000000000000_0001111001001011_0111011000100100"; -- 0.11833895095276367
	pesos_i(4930) := b"0000000000000000_0000000000000000_0000001011010001_0110111111101011"; -- 0.011008257695591848
	pesos_i(4931) := b"0000000000000000_0000000000000000_0001100111011110_0011011111110001"; -- 0.1010470354701203
	pesos_i(4932) := b"1111111111111111_1111111111111111_1101011010110010_1111001011101101"; -- -0.16133195603735018
	pesos_i(4933) := b"1111111111111111_1111111111111111_1101001111001011_0101110111001010"; -- -0.17267812548042205
	pesos_i(4934) := b"0000000000000000_0000000000000000_0001011110100000_0001001101010001"; -- 0.09228630762775153
	pesos_i(4935) := b"0000000000000000_0000000000000000_0010111100000011_0001001001001101"; -- 0.18364061716309413
	pesos_i(4936) := b"0000000000000000_0000000000000000_0010000100000111_0110010100011100"; -- 0.12901908807212523
	pesos_i(4937) := b"1111111111111111_1111111111111111_1110100111101001_0011001010010101"; -- -0.08628543715082918
	pesos_i(4938) := b"1111111111111111_1111111111111111_1111000010000010_1001010100101000"; -- -0.06050746696476905
	pesos_i(4939) := b"0000000000000000_0000000000000000_0010000101100011_1110111010110110"; -- 0.1304310984700201
	pesos_i(4940) := b"0000000000000000_0000000000000000_0001110111100001_0010000001001100"; -- 0.11671640252963289
	pesos_i(4941) := b"0000000000000000_0000000000000000_0000011110101010_0010000010111000"; -- 0.029939694294736897
	pesos_i(4942) := b"0000000000000000_0000000000000000_0000111101111011_0111001110101010"; -- 0.0604774751194021
	pesos_i(4943) := b"1111111111111111_1111111111111111_1110100010101000_1100011110001100"; -- -0.09117462958114093
	pesos_i(4944) := b"1111111111111111_1111111111111111_1110100100111000_1000111011001110"; -- -0.08898074604856293
	pesos_i(4945) := b"1111111111111111_1111111111111111_1110000000010001_0011001001101001"; -- -0.12473759585375793
	pesos_i(4946) := b"0000000000000000_0000000000000000_0000010111010000_1011011011001101"; -- 0.022715973980214493
	pesos_i(4947) := b"0000000000000000_0000000000000000_0001111010000101_0000010001101001"; -- 0.11921718185379714
	pesos_i(4948) := b"0000000000000000_0000000000000000_0010001111000100_0010100110110011"; -- 0.13971195823319998
	pesos_i(4949) := b"1111111111111111_1111111111111111_1110111001111111_1110010111010011"; -- -0.06836093515097974
	pesos_i(4950) := b"1111111111111111_1111111111111111_1101100111000101_0000010111100111"; -- -0.14933741668553993
	pesos_i(4951) := b"0000000000000000_0000000000000000_0010111011010101_1000010101110101"; -- 0.1829455767048513
	pesos_i(4952) := b"1111111111111111_1111111111111111_1111011101111101_1100011001000110"; -- -0.03323708335635258
	pesos_i(4953) := b"1111111111111111_1111111111111111_1101111111011110_0001100110001101"; -- -0.1255172758732767
	pesos_i(4954) := b"0000000000000000_0000000000000000_0001011001011111_0110010101001101"; -- 0.08739312285006232
	pesos_i(4955) := b"0000000000000000_0000000000000000_0000010111110000_1101101000100010"; -- 0.023206361219606304
	pesos_i(4956) := b"1111111111111111_1111111111111111_1111000001101001_0100100100110100"; -- -0.06089346382039851
	pesos_i(4957) := b"0000000000000000_0000000000000000_0010011110011001_1011011111100110"; -- 0.1546893060155349
	pesos_i(4958) := b"0000000000000000_0000000000000000_0001011011101001_0011000111101010"; -- 0.0894957730166891
	pesos_i(4959) := b"1111111111111111_1111111111111111_1111001110100100_0000000101100011"; -- -0.048278725965301555
	pesos_i(4960) := b"1111111111111111_1111111111111111_1111110011100111_1011011111100101"; -- -0.012089258725531654
	pesos_i(4961) := b"0000000000000000_0000000000000000_0001100100011110_1111111010011101"; -- 0.09812918977763563
	pesos_i(4962) := b"1111111111111111_1111111111111111_1111100000011000_0110101100011000"; -- -0.030877405672351855
	pesos_i(4963) := b"1111111111111111_1111111111111111_1110001100100111_0011111000010001"; -- -0.11268245777730258
	pesos_i(4964) := b"1111111111111111_1111111111111111_1101000100000110_1001101011001001"; -- -0.1834929713719282
	pesos_i(4965) := b"1111111111111111_1111111111111111_1111110000100111_0001101111010000"; -- -0.015028249520392908
	pesos_i(4966) := b"0000000000000000_0000000000000000_0000010010101000_1010000110001010"; -- 0.018198104934752872
	pesos_i(4967) := b"0000000000000000_0000000000000000_0001100000101010_1000001101111111"; -- 0.09439870690097604
	pesos_i(4968) := b"1111111111111111_1111111111111111_1101100010110010_1110010111001111"; -- -0.1535202377937216
	pesos_i(4969) := b"0000000000000000_0000000000000000_0000111001111100_1111110011000010"; -- 0.0565946553515827
	pesos_i(4970) := b"1111111111111111_1111111111111111_1101101101000001_0011010011010000"; -- -0.1435362809524617
	pesos_i(4971) := b"1111111111111111_1111111111111111_1111111100011111_1011110110011010"; -- -0.0034219263651873604
	pesos_i(4972) := b"0000000000000000_0000000000000000_0010001100001001_1111011101111111"; -- 0.13687083092647706
	pesos_i(4973) := b"0000000000000000_0000000000000000_0001101110111100_1111010111011101"; -- 0.10835205692052712
	pesos_i(4974) := b"1111111111111111_1111111111111111_1101010110111000_1101101001111000"; -- -0.165148111125546
	pesos_i(4975) := b"1111111111111111_1111111111111111_1110100110001111_0010111000100001"; -- -0.08765899366822093
	pesos_i(4976) := b"0000000000000000_0000000000000000_0000000101100100_0001111011001000"; -- 0.005433963695597788
	pesos_i(4977) := b"1111111111111111_1111111111111111_1110100101100110_0111101111110010"; -- -0.08827996577290326
	pesos_i(4978) := b"1111111111111111_1111111111111111_1101110110101110_1000110010010011"; -- -0.13405534191728047
	pesos_i(4979) := b"1111111111111111_1111111111111111_1101010011010110_0011011000011111"; -- -0.1686063932643649
	pesos_i(4980) := b"0000000000000000_0000000000000000_0010111000001011_1100011001000100"; -- 0.17986716419436274
	pesos_i(4981) := b"1111111111111111_1111111111111111_1110001000101110_0011111100000101"; -- -0.1164818395554079
	pesos_i(4982) := b"1111111111111111_1111111111111111_1110011110111011_1101110001000101"; -- -0.09478972734409716
	pesos_i(4983) := b"1111111111111111_1111111111111111_1101110100010100_0011000110101010"; -- -0.13641061399538126
	pesos_i(4984) := b"0000000000000000_0000000000000000_0010110100101000_1100100010100111"; -- 0.17640356125971193
	pesos_i(4985) := b"0000000000000000_0000000000000000_0000100110100111_1111001100010011"; -- 0.03771895602612451
	pesos_i(4986) := b"0000000000000000_0000000000000000_0001010000100011_1111000110001001"; -- 0.07867345420461831
	pesos_i(4987) := b"0000000000000000_0000000000000000_0010001110110000_1111000010011100"; -- 0.13941863821751488
	pesos_i(4988) := b"1111111111111111_1111111111111111_1111111110000101_0100001000010111"; -- -0.001872891867463783
	pesos_i(4989) := b"1111111111111111_1111111111111111_1110010101101010_0010000110001011"; -- -0.1038493189525032
	pesos_i(4990) := b"0000000000000000_0000000000000000_0010001100001101_0010011101000000"; -- 0.13691945369662206
	pesos_i(4991) := b"1111111111111111_1111111111111111_1110000001011111_1101111100111010"; -- -0.12353710964271614
	pesos_i(4992) := b"1111111111111111_1111111111111111_1111100001010111_1100100000010000"; -- -0.029910560731802788
	pesos_i(4993) := b"0000000000000000_0000000000000000_0011001011010000_1100110100001101"; -- 0.19849855014609644
	pesos_i(4994) := b"1111111111111111_1111111111111111_1111010101101001_1100111011111100"; -- -0.041354239962097035
	pesos_i(4995) := b"1111111111111111_1111111111111111_1101010100111110_0010010111101110"; -- -0.16702044437177102
	pesos_i(4996) := b"0000000000000000_0000000000000000_0010100001100111_0000011110010010"; -- 0.15782210651125156
	pesos_i(4997) := b"0000000000000000_0000000000000000_0001100110100111_1000001000100010"; -- 0.10021222425268954
	pesos_i(4998) := b"1111111111111111_1111111111111111_1111101001110101_0001000100101010"; -- -0.0216511987331603
	pesos_i(4999) := b"0000000000000000_0000000000000000_0000100110001111_1100000101111010"; -- 0.037349789049855045
	pesos_i(5000) := b"1111111111111111_1111111111111111_1110111001010100_1001101101000011"; -- -0.06902150735526788
	pesos_i(5001) := b"0000000000000000_0000000000000000_0000011100110110_1110011011001011"; -- 0.028181480847686076
	pesos_i(5002) := b"0000000000000000_0000000000000000_0001111101001110_0100011111101001"; -- 0.1222882217334806
	pesos_i(5003) := b"1111111111111111_1111111111111111_1101100011101011_1110111010110101"; -- -0.15264995653280475
	pesos_i(5004) := b"1111111111111111_1111111111111111_1111001111110101_0100000101001010"; -- -0.04703895509206437
	pesos_i(5005) := b"0000000000000000_0000000000000000_0010000101111001_0010110111100111"; -- 0.13075529937547103
	pesos_i(5006) := b"1111111111111111_1111111111111111_1111110001010001_0101100001111110"; -- -0.014383763607737562
	pesos_i(5007) := b"1111111111111111_1111111111111111_1110101111011110_0111010001110010"; -- -0.07863685813506975
	pesos_i(5008) := b"1111111111111111_1111111111111111_1101010001010100_0011010110110011"; -- -0.17059006090063025
	pesos_i(5009) := b"0000000000000000_0000000000000000_0001010101011010_1111110010010000"; -- 0.08341959498951601
	pesos_i(5010) := b"1111111111111111_1111111111111111_1111111100000000_1001111110101011"; -- -0.0038967330132580824
	pesos_i(5011) := b"1111111111111111_1111111111111111_1101100010011100_1000111001001110"; -- -0.1538611469772971
	pesos_i(5012) := b"0000000000000000_0000000000000000_0000000100011101_0101001101000110"; -- 0.004353718406386159
	pesos_i(5013) := b"1111111111111111_1111111111111111_1101111101000000_1000110011101100"; -- -0.12792128799487198
	pesos_i(5014) := b"0000000000000000_0000000000000000_0001010111011000_1100000000100000"; -- 0.08533860002677675
	pesos_i(5015) := b"0000000000000000_0000000000000000_0001000100100110_1100101100000101"; -- 0.06699818492666743
	pesos_i(5016) := b"0000000000000000_0000000000000000_0010010011000101_0010101010000100"; -- 0.14363351547954445
	pesos_i(5017) := b"0000000000000000_0000000000000000_0001100001011100_0010001110111100"; -- 0.09515593856091925
	pesos_i(5018) := b"0000000000000000_0000000000000000_0001010000101011_0000100110100101"; -- 0.07878170283137534
	pesos_i(5019) := b"0000000000000000_0000000000000000_0001101100011100_1110001000010001"; -- 0.10590947077664935
	pesos_i(5020) := b"0000000000000000_0000000000000000_0001101100101100_0010101001011111"; -- 0.10614266215920964
	pesos_i(5021) := b"1111111111111111_1111111111111111_1110111101010111_0101001110000111"; -- -0.06507375672848491
	pesos_i(5022) := b"0000000000000000_0000000000000000_0010111001010001_0110001011011010"; -- 0.180929354025038
	pesos_i(5023) := b"1111111111111111_1111111111111111_1110000101011101_1011110001011111"; -- -0.1196634548388012
	pesos_i(5024) := b"1111111111111111_1111111111111111_1110100010000000_1011111101010110"; -- -0.09178547057633148
	pesos_i(5025) := b"0000000000000000_0000000000000000_0001101100110010_1001100101001000"; -- 0.10624082567231607
	pesos_i(5026) := b"0000000000000000_0000000000000000_0010010100010001_0001111010101001"; -- 0.14479247685065313
	pesos_i(5027) := b"0000000000000000_0000000000000000_0000000100010100_0000001011011011"; -- 0.004211595951126428
	pesos_i(5028) := b"1111111111111111_1111111111111111_1110111001110111_1110011101100100"; -- -0.06848291224517396
	pesos_i(5029) := b"0000000000000000_0000000000000000_0010001001011010_0101010001110011"; -- 0.13419082450953757
	pesos_i(5030) := b"1111111111111111_1111111111111111_1111110110111000_0011111101111010"; -- -0.008907349268117643
	pesos_i(5031) := b"1111111111111111_1111111111111111_1101011011001001_1110100100010110"; -- -0.16098159038425122
	pesos_i(5032) := b"1111111111111111_1111111111111111_1111101010101010_0111101010111010"; -- -0.020836190672464866
	pesos_i(5033) := b"1111111111111111_1111111111111111_1111101100011111_0000100011010111"; -- -0.01905770065737281
	pesos_i(5034) := b"1111111111111111_1111111111111111_1110010001010111_0000101110001101"; -- -0.1080467969079158
	pesos_i(5035) := b"1111111111111111_1111111111111111_1110111111001101_0010000000011110"; -- -0.06327628388803444
	pesos_i(5036) := b"0000000000000000_0000000000000000_0000110011000010_0000011000010101"; -- 0.04983556761545876
	pesos_i(5037) := b"0000000000000000_0000000000000000_0010011100110011_1010111110101011"; -- 0.15313241875299446
	pesos_i(5038) := b"0000000000000000_0000000000000000_0000111011000001_0011110000010010"; -- 0.057636026872680955
	pesos_i(5039) := b"0000000000000000_0000000000000000_0001101010001110_1010000101111001"; -- 0.10373887247180273
	pesos_i(5040) := b"0000000000000000_0000000000000000_0001101110001101_1111001101011101"; -- 0.10763474488468991
	pesos_i(5041) := b"1111111111111111_1111111111111111_1111011001101101_1101010001010010"; -- -0.037386636728318864
	pesos_i(5042) := b"0000000000000000_0000000000000000_0001010001000001_0110101011101111"; -- 0.07912319492319095
	pesos_i(5043) := b"1111111111111111_1111111111111111_1111110001010101_0100001101011100"; -- -0.014323988070351073
	pesos_i(5044) := b"1111111111111111_1111111111111111_1111110011011011_0100010101010001"; -- -0.012279193663468852
	pesos_i(5045) := b"1111111111111111_1111111111111111_1110100010111101_1000010111011101"; -- -0.09085810994259716
	pesos_i(5046) := b"1111111111111111_1111111111111111_1110100111110001_0001110100100011"; -- -0.08616464512533098
	pesos_i(5047) := b"1111111111111111_1111111111111111_1111000111110001_1010000100010011"; -- -0.05490678095361051
	pesos_i(5048) := b"1111111111111111_1111111111111111_1111011100011011_1011110101110010"; -- -0.034732970911626804
	pesos_i(5049) := b"1111111111111111_1111111111111111_1110100000111111_0101101110000111"; -- -0.09278324089236571
	pesos_i(5050) := b"1111111111111111_1111111111111111_1110100101101101_1000111110100101"; -- -0.08817198015828924
	pesos_i(5051) := b"0000000000000000_0000000000000000_0010100001110110_0111101110101000"; -- 0.15805790750539936
	pesos_i(5052) := b"0000000000000000_0000000000000000_0001011110011011_1000011110011101"; -- 0.09221694543615837
	pesos_i(5053) := b"1111111111111111_1111111111111111_1111010110110000_0000011010010001"; -- -0.040282811664239505
	pesos_i(5054) := b"1111111111111111_1111111111111111_1111101110011110_1010000110010100"; -- -0.017110730407745457
	pesos_i(5055) := b"0000000000000000_0000000000000000_0001010101101001_1010110101100100"; -- 0.08364375772693372
	pesos_i(5056) := b"0000000000000000_0000000000000000_0001011010000101_0001010111010010"; -- 0.08796821959434473
	pesos_i(5057) := b"1111111111111111_1111111111111111_1111100101001011_0001111001010010"; -- -0.026197533514535517
	pesos_i(5058) := b"0000000000000000_0000000000000000_0001110000101011_1010011010101111"; -- 0.11004106299461586
	pesos_i(5059) := b"1111111111111111_1111111111111111_1111100000111001_1000011011010100"; -- -0.030372212659622425
	pesos_i(5060) := b"1111111111111111_1111111111111111_1111111101111001_1011010011000111"; -- -0.002049161242923107
	pesos_i(5061) := b"0000000000000000_0000000000000000_0001010001000010_1001101001001010"; -- 0.0791412764269623
	pesos_i(5062) := b"0000000000000000_0000000000000000_0001010101001000_0000011011100011"; -- 0.08313029339629785
	pesos_i(5063) := b"0000000000000000_0000000000000000_0001000001001000_1001111100010111"; -- 0.06360811528124277
	pesos_i(5064) := b"0000000000000000_0000000000000000_0001000000101101_0010011001000100"; -- 0.06318892636672255
	pesos_i(5065) := b"1111111111111111_1111111111111111_1110100001111011_1010110011110110"; -- -0.09186285962703374
	pesos_i(5066) := b"0000000000000000_0000000000000000_0000010001101001_0111110010010001"; -- 0.017234597619412276
	pesos_i(5067) := b"0000000000000000_0000000000000000_0001011001110111_1110010100111011"; -- 0.08776695920955238
	pesos_i(5068) := b"1111111111111111_1111111111111111_1110110110101100_1010010101011000"; -- -0.07158438306330064
	pesos_i(5069) := b"1111111111111111_1111111111111111_1110101000100111_1010001011000110"; -- -0.0853327052456208
	pesos_i(5070) := b"1111111111111111_1111111111111111_1110101110010001_0010100110010000"; -- -0.07981624833856676
	pesos_i(5071) := b"1111111111111111_1111111111111111_1101111011011000_0100100000000000"; -- -0.1295123099946403
	pesos_i(5072) := b"0000000000000000_0000000000000000_0010010000100100_0001101011111011"; -- 0.14117592467135712
	pesos_i(5073) := b"1111111111111111_1111111111111111_1111101110111010_1100110111011100"; -- -0.016680845090552135
	pesos_i(5074) := b"1111111111111111_1111111111111111_1111000110101000_0111110000110110"; -- -0.056022869921807425
	pesos_i(5075) := b"0000000000000000_0000000000000000_0010110011101000_1110111101000010"; -- 0.17542929996027137
	pesos_i(5076) := b"1111111111111111_1111111111111111_1110111001001111_1010011101100110"; -- -0.06909707798577472
	pesos_i(5077) := b"1111111111111111_1111111111111111_1110010010111000_0110100101111101"; -- -0.10656109514234366
	pesos_i(5078) := b"1111111111111111_1111111111111111_1110110111011101_1011000111001000"; -- -0.07083596097402417
	pesos_i(5079) := b"1111111111111111_1111111111111111_1110001010110000_0111011111101101"; -- -0.11449480497707093
	pesos_i(5080) := b"0000000000000000_0000000000000000_0010010000100111_1001010001000001"; -- 0.14122892930399458
	pesos_i(5081) := b"1111111111111111_1111111111111111_1111110010100001_1110000000101011"; -- -0.013154973410790827
	pesos_i(5082) := b"1111111111111111_1111111111111111_1101111101110110_1001000001111110"; -- -0.1270971005797037
	pesos_i(5083) := b"0000000000000000_0000000000000000_0001110010001101_1001101000001101"; -- 0.11153567142265444
	pesos_i(5084) := b"0000000000000000_0000000000000000_0001100011001000_0001001011101101"; -- 0.09680288594073942
	pesos_i(5085) := b"1111111111111111_1111111111111111_1111000110011111_0011101110001001"; -- -0.056164053952532954
	pesos_i(5086) := b"0000000000000000_0000000000000000_0001000100000010_1001100010001101"; -- 0.06644586029283199
	pesos_i(5087) := b"0000000000000000_0000000000000000_0001101111011011_1100000101001011"; -- 0.10882194595516262
	pesos_i(5088) := b"0000000000000000_0000000000000000_0010011110101111_1101000100101100"; -- 0.1550265056656309
	pesos_i(5089) := b"0000000000000000_0000000000000000_0000011111100000_0011010001110111"; -- 0.030764845925649403
	pesos_i(5090) := b"1111111111111111_1111111111111111_1110110100000001_1001001101011100"; -- -0.07419470799146265
	pesos_i(5091) := b"0000000000000000_0000000000000000_0000001011001000_1100110000101000"; -- 0.010876426368437726
	pesos_i(5092) := b"0000000000000000_0000000000000000_0000101000100001_1011011000100111"; -- 0.039576897213183464
	pesos_i(5093) := b"1111111111111111_1111111111111111_1111010000010001_0111101001100110"; -- -0.04660830515181695
	pesos_i(5094) := b"0000000000000000_0000000000000000_0001001000000101_0001010011101011"; -- 0.07039004079175226
	pesos_i(5095) := b"1111111111111111_1111111111111111_1110001100010110_0001100110111010"; -- -0.11294402315106417
	pesos_i(5096) := b"1111111111111111_1111111111111111_1111001110010010_1110000111011011"; -- -0.04854000475966949
	pesos_i(5097) := b"0000000000000000_0000000000000000_0010101011101011_0110100011011110"; -- 0.16765456589712316
	pesos_i(5098) := b"1111111111111111_1111111111111111_1111011100111000_1110010011101101"; -- -0.034288112822755526
	pesos_i(5099) := b"1111111111111111_1111111111111111_1101011101000111_1100011011011101"; -- -0.15906102277516612
	pesos_i(5100) := b"0000000000000000_0000000000000000_0000000001100101_0001100100101010"; -- 0.0015426375741124996
	pesos_i(5101) := b"1111111111111111_1111111111111111_1101100101001100_1000000110010111"; -- -0.15117635778498476
	pesos_i(5102) := b"1111111111111111_1111111111111111_1111101101101011_0011001111010000"; -- -0.0178954712486164
	pesos_i(5103) := b"1111111111111111_1111111111111111_1110011011101000_1000001100100110"; -- -0.0980146438143512
	pesos_i(5104) := b"0000000000000000_0000000000000000_0001110100001111_0111000001001100"; -- 0.11351682530635035
	pesos_i(5105) := b"1111111111111111_1111111111111111_1111001100010011_0100110110001110"; -- -0.05048671046652491
	pesos_i(5106) := b"0000000000000000_0000000000000000_0010101110000001_0110010010010100"; -- 0.16994312880610604
	pesos_i(5107) := b"0000000000000000_0000000000000000_0000111001100110_0011010000010001"; -- 0.056246999822870826
	pesos_i(5108) := b"0000000000000000_0000000000000000_0000100100010111_0110011101100111"; -- 0.03551336542952333
	pesos_i(5109) := b"1111111111111111_1111111111111111_1110101010001001_0001011101101110"; -- -0.08384564927803244
	pesos_i(5110) := b"0000000000000000_0000000000000000_0001101110100010_0101101010101110"; -- 0.10794607867416793
	pesos_i(5111) := b"1111111111111111_1111111111111111_1101101000101110_1110001100101110"; -- -0.14772205479172143
	pesos_i(5112) := b"0000000000000000_0000000000000000_0000101100001110_1111001001110101"; -- 0.04319682454853588
	pesos_i(5113) := b"1111111111111111_1111111111111111_1111000000110001_0011111111010000"; -- -0.06174851589714204
	pesos_i(5114) := b"0000000000000000_0000000000000000_0001110011011001_0110101011000011"; -- 0.1126925206862873
	pesos_i(5115) := b"1111111111111111_1111111111111111_1111010100100010_0011010100111110"; -- -0.042446777669693486
	pesos_i(5116) := b"1111111111111111_1111111111111111_1111010101111000_0111111111101110"; -- -0.04113007010891154
	pesos_i(5117) := b"0000000000000000_0000000000000000_0000100110011110_1101100110110000"; -- 0.037580113834344175
	pesos_i(5118) := b"0000000000000000_0000000000000000_0010100011101100_0010111000111111"; -- 0.15985383077044787
	pesos_i(5119) := b"1111111111111111_1111111111111111_1110100000000001_1101100111010010"; -- -0.09372175812047659
	pesos_i(5120) := b"0000000000000000_0000000000000000_0010011010011101_1001010011000001"; -- 0.15084199640221488
	pesos_i(5121) := b"1111111111111111_1111111111111111_1101100000011011_0100010000111001"; -- -0.1558339462967084
	pesos_i(5122) := b"1111111111111111_1111111111111111_1101011001010110_0100001011000110"; -- -0.16274626414997315
	pesos_i(5123) := b"1111111111111111_1111111111111111_1111000111110000_1010000111011110"; -- -0.054921992546527174
	pesos_i(5124) := b"0000000000000000_0000000000000000_0010011100111110_0101100111000011"; -- 0.15329514523894874
	pesos_i(5125) := b"1111111111111111_1111111111111111_1110110110101011_0101000110101100"; -- -0.07160462896554806
	pesos_i(5126) := b"0000000000000000_0000000000000000_0010101001101010_1111010011010100"; -- 0.16569452452753766
	pesos_i(5127) := b"1111111111111111_1111111111111111_1110100110011010_1011010011001010"; -- -0.08748312066857358
	pesos_i(5128) := b"0000000000000000_0000000000000000_0000000001111101_0000111100011001"; -- 0.0019082486065983679
	pesos_i(5129) := b"1111111111111111_1111111111111111_1111100010110110_0111110001110010"; -- -0.028465482856164806
	pesos_i(5130) := b"0000000000000000_0000000000000000_0000011001100010_1011010001000111"; -- 0.02494360672230187
	pesos_i(5131) := b"0000000000000000_0000000000000000_0001001101101010_0111001000101111"; -- 0.0758429875909875
	pesos_i(5132) := b"0000000000000000_0000000000000000_0000100000000010_1111010010111100"; -- 0.03129510477872174
	pesos_i(5133) := b"0000000000000000_0000000000000000_0000011010001011_1110000111100011"; -- 0.0255719354947208
	pesos_i(5134) := b"1111111111111111_1111111111111111_1110001100101111_0011000110110001"; -- -0.11256112512278273
	pesos_i(5135) := b"1111111111111111_1111111111111111_1110011010011110_0010001111101111"; -- -0.09914946957159522
	pesos_i(5136) := b"1111111111111111_1111111111111111_1111000001110101_1011010101000011"; -- -0.06070391763670041
	pesos_i(5137) := b"0000000000000000_0000000000000000_0010000100000001_0000110011101110"; -- 0.128922279568323
	pesos_i(5138) := b"1111111111111111_1111111111111111_1101001111100010_1011010011110100"; -- -0.17232197808870384
	pesos_i(5139) := b"0000000000000000_0000000000000000_0000001001001000_1000001110010101"; -- 0.008918975732054756
	pesos_i(5140) := b"0000000000000000_0000000000000000_0001000111011010_0100101100100001"; -- 0.06973714415572639
	pesos_i(5141) := b"1111111111111111_1111111111111111_1110100010100000_1111010010010000"; -- -0.09129401676218236
	pesos_i(5142) := b"0000000000000000_0000000000000000_0001111100111100_1101010100000001"; -- 0.12202197326316126
	pesos_i(5143) := b"0000000000000000_0000000000000000_0000010010010010_1110110110111111"; -- 0.01786695390756449
	pesos_i(5144) := b"0000000000000000_0000000000000000_0000111001000111_1100010111011111"; -- 0.05578266814043528
	pesos_i(5145) := b"1111111111111111_1111111111111111_1111001010001001_0100000111011110"; -- -0.05259312000330483
	pesos_i(5146) := b"0000000000000000_0000000000000000_0001001010111100_0100110011010010"; -- 0.07318573126345268
	pesos_i(5147) := b"0000000000000000_0000000000000000_0001101101010111_0100011011011100"; -- 0.10680048811733144
	pesos_i(5148) := b"1111111111111111_1111111111111111_1111111011001100_0111110100100110"; -- -0.004692247642313532
	pesos_i(5149) := b"1111111111111111_1111111111111111_1110101101101000_1011000100111010"; -- -0.0804337725055057
	pesos_i(5150) := b"1111111111111111_1111111111111111_1111111101110001_0100010001011010"; -- -0.0021779327343179598
	pesos_i(5151) := b"0000000000000000_0000000000000000_0010010101010011_1010111000011110"; -- 0.1458081077721263
	pesos_i(5152) := b"1111111111111111_1111111111111111_1101010011111110_1100100001111111"; -- -0.16798731697916502
	pesos_i(5153) := b"0000000000000000_0000000000000000_0000100000011110_0110001111001000"; -- 0.03171371119353964
	pesos_i(5154) := b"0000000000000000_0000000000000000_0010000101110110_1000000100101010"; -- 0.13071448589886853
	pesos_i(5155) := b"0000000000000000_0000000000000000_0001101001001101_0101101100001100"; -- 0.10274285349321235
	pesos_i(5156) := b"1111111111111111_1111111111111111_1111110011011111_1000111000111100"; -- -0.012213812217552295
	pesos_i(5157) := b"0000000000000000_0000000000000000_0000101100111010_0110000101111110"; -- 0.04385957082886528
	pesos_i(5158) := b"1111111111111111_1111111111111111_1111011101111001_0010001110111010"; -- -0.033307807034010775
	pesos_i(5159) := b"1111111111111111_1111111111111111_1110111010101000_0010000111110110"; -- -0.06774699923677134
	pesos_i(5160) := b"1111111111111111_1111111111111111_1111100011111011_0010100010000101"; -- -0.027417628698178487
	pesos_i(5161) := b"0000000000000000_0000000000000000_0001010011110110_0101010010000101"; -- 0.08188369988203094
	pesos_i(5162) := b"1111111111111111_1111111111111111_1110011001010010_0101100100101100"; -- -0.10030596428714786
	pesos_i(5163) := b"0000000000000000_0000000000000000_0001101111101111_1011111111100111"; -- 0.10912703884146352
	pesos_i(5164) := b"1111111111111111_1111111111111111_1111101111000101_1011111101110011"; -- -0.016513857325810396
	pesos_i(5165) := b"1111111111111111_1111111111111111_1110100101111000_0101110001110111"; -- -0.08800718403619448
	pesos_i(5166) := b"1111111111111111_1111111111111111_1101101001110111_1110111111101100"; -- -0.14660740362891805
	pesos_i(5167) := b"0000000000000000_0000000000000000_0000000010111001_1001110010010110"; -- 0.002832209138495531
	pesos_i(5168) := b"1111111111111111_1111111111111111_1101101000000100_1010001111001010"; -- -0.1483667022868295
	pesos_i(5169) := b"1111111111111111_1111111111111111_1111101110000000_0100100011000001"; -- -0.017573788441722117
	pesos_i(5170) := b"0000000000000000_0000000000000000_0000101010001101_1011110001011000"; -- 0.04122521550069831
	pesos_i(5171) := b"0000000000000000_0000000000000000_0000111001000000_1001110010001101"; -- 0.05567339370171894
	pesos_i(5172) := b"0000000000000000_0000000000000000_0010100000111011_0110010101111110"; -- 0.15715631787224277
	pesos_i(5173) := b"1111111111111111_1111111111111111_1111111100101101_0001110001111100"; -- -0.003217906655793431
	pesos_i(5174) := b"0000000000000000_0000000000000000_0000001000011111_1101011011100100"; -- 0.008298331018424846
	pesos_i(5175) := b"0000000000000000_0000000000000000_0001101100111011_1111010000110010"; -- 0.10638357368443939
	pesos_i(5176) := b"0000000000000000_0000000000000000_0010110010101101_0101011100011011"; -- 0.17451996250550986
	pesos_i(5177) := b"0000000000000000_0000000000000000_0010011001011111_1001101010000101"; -- 0.1498962949683677
	pesos_i(5178) := b"1111111111111111_1111111111111111_1111100110101000_1100000111111101"; -- -0.0247687107450537
	pesos_i(5179) := b"1111111111111111_1111111111111111_1110101110111111_1010000000011101"; -- -0.07910727783532655
	pesos_i(5180) := b"1111111111111111_1111111111111111_1101101100011001_0110111111100001"; -- -0.14414311168865468
	pesos_i(5181) := b"1111111111111111_1111111111111111_1111110010010110_0000000000100101"; -- -0.013336173080478134
	pesos_i(5182) := b"0000000000000000_0000000000000000_0000011010111110_0011101010000011"; -- 0.026340157566946062
	pesos_i(5183) := b"0000000000000000_0000000000000000_0001011010011001_0011101001111100"; -- 0.08827558058601961
	pesos_i(5184) := b"1111111111111111_1111111111111111_1110001001010100_0011011101110101"; -- -0.1159024562386742
	pesos_i(5185) := b"0000000000000000_0000000000000000_0001011111110111_1001001010010011"; -- 0.09362140745339734
	pesos_i(5186) := b"1111111111111111_1111111111111111_1110000000011001_0011000110100111"; -- -0.12461557081300915
	pesos_i(5187) := b"1111111111111111_1111111111111111_1101111000010001_0101001111101000"; -- -0.13254809927564337
	pesos_i(5188) := b"0000000000000000_0000000000000000_0000100111111101_1000011011111110"; -- 0.03902476974861863
	pesos_i(5189) := b"1111111111111111_1111111111111111_1111010001101000_0010001000111101"; -- -0.045286045080359036
	pesos_i(5190) := b"1111111111111111_1111111111111111_1111000000000101_1110000001100100"; -- -0.06241033126441297
	pesos_i(5191) := b"0000000000000000_0000000000000000_0001010010100000_1011111110011111"; -- 0.08057782775863076
	pesos_i(5192) := b"0000000000000000_0000000000000000_0010100101110010_1101011101001111"; -- 0.16190858531857785
	pesos_i(5193) := b"1111111111111111_1111111111111111_1111011100111111_0000010100111001"; -- -0.034194634992847826
	pesos_i(5194) := b"0000000000000000_0000000000000000_0000101101010010_0011001101110011"; -- 0.044223037317637354
	pesos_i(5195) := b"1111111111111111_1111111111111111_1110000111000001_0011101101000001"; -- -0.11814527188238033
	pesos_i(5196) := b"1111111111111111_1111111111111111_1111011110011100_0100111101001111"; -- -0.032771151725881575
	pesos_i(5197) := b"1111111111111111_1111111111111111_1111101011011101_1111000111011010"; -- -0.020050892102436473
	pesos_i(5198) := b"1111111111111111_1111111111111111_1101011110011001_0110010101010001"; -- -0.15781561641758377
	pesos_i(5199) := b"0000000000000000_0000000000000000_0010011100010110_1111000100001100"; -- 0.15269381077129954
	pesos_i(5200) := b"0000000000000000_0000000000000000_0001000001010000_0011100110110010"; -- 0.06372414195736165
	pesos_i(5201) := b"0000000000000000_0000000000000000_0001111100110110_1110100100111111"; -- 0.12193162714674047
	pesos_i(5202) := b"0000000000000000_0000000000000000_0010011000001110_1000010101101011"; -- 0.14865907543491647
	pesos_i(5203) := b"0000000000000000_0000000000000000_0010001101001110_1010110000110011"; -- 0.13791919931987648
	pesos_i(5204) := b"1111111111111111_1111111111111111_1101100100100001_0011100000110011"; -- -0.1518368601951693
	pesos_i(5205) := b"1111111111111111_1111111111111111_1111011000010111_0101000010001101"; -- -0.03870674665369644
	pesos_i(5206) := b"0000000000000000_0000000000000000_0001011011010110_1100101000001111"; -- 0.08921492456716593
	pesos_i(5207) := b"1111111111111111_1111111111111111_1110111011101000_0010010010000110"; -- -0.06677028401245566
	pesos_i(5208) := b"1111111111111111_1111111111111111_1100101111111000_1011000011101110"; -- -0.20323652451203336
	pesos_i(5209) := b"1111111111111111_1111111111111111_1110011100011011_1111111110110100"; -- -0.09722902150724579
	pesos_i(5210) := b"1111111111111111_1111111111111111_1101010011110100_0100000001000001"; -- -0.1681480256735757
	pesos_i(5211) := b"1111111111111111_1111111111111111_1111100001110101_1111110001100101"; -- -0.02944967787270931
	pesos_i(5212) := b"1111111111111111_1111111111111111_1101101111000100_1100110110010001"; -- -0.14152827464519138
	pesos_i(5213) := b"0000000000000000_0000000000000000_0000110111111101_0111010111100000"; -- 0.05464874964406545
	pesos_i(5214) := b"0000000000000000_0000000000000000_0001100010111101_1101110001110010"; -- 0.09664705074794432
	pesos_i(5215) := b"1111111111111111_1111111111111111_1110011110101110_1101000111100000"; -- -0.09498871107497864
	pesos_i(5216) := b"0000000000000000_0000000000000000_0000110110100011_1100110111110101"; -- 0.053280708710132296
	pesos_i(5217) := b"0000000000000000_0000000000000000_0011000111100001_1100001110001101"; -- 0.19485113324529965
	pesos_i(5218) := b"0000000000000000_0000000000000000_0000110011001111_0001100111110001"; -- 0.05003511546001942
	pesos_i(5219) := b"1111111111111111_1111111111111111_1111011100100101_0101011011100111"; -- -0.034586495047177715
	pesos_i(5220) := b"0000000000000000_0000000000000000_0000100011101111_1001011110000110"; -- 0.034905882163113335
	pesos_i(5221) := b"1111111111111111_1111111111111111_1111000100101100_1100110100001110"; -- -0.057910141151924006
	pesos_i(5222) := b"1111111111111111_1111111111111111_1110001001000110_1101000100111001"; -- -0.11610691421980027
	pesos_i(5223) := b"1111111111111111_1111111111111111_1101011110101001_1100011100011101"; -- -0.1575656466310283
	pesos_i(5224) := b"0000000000000000_0000000000000000_0000010011010100_1100110010010001"; -- 0.01887205644658768
	pesos_i(5225) := b"0000000000000000_0000000000000000_0000000010110000_1110001111100111"; -- 0.0026991309651882914
	pesos_i(5226) := b"1111111111111111_1111111111111111_1110011011100111_1010011110011111"; -- -0.09802772883511122
	pesos_i(5227) := b"1111111111111111_1111111111111111_1101101101000110_1110101011001010"; -- -0.1434491401338086
	pesos_i(5228) := b"1111111111111111_1111111111111111_1111001001101010_1000011000010011"; -- -0.05306207699379549
	pesos_i(5229) := b"0000000000000000_0000000000000000_0000001100110011_0001001100111101"; -- 0.012498094932639089
	pesos_i(5230) := b"0000000000000000_0000000000000000_0001001110000001_1111110111011100"; -- 0.07620226508267577
	pesos_i(5231) := b"0000000000000000_0000000000000000_0001010101100101_1000110010111100"; -- 0.08358077612663943
	pesos_i(5232) := b"0000000000000000_0000000000000000_0000110011110011_0100011101110000"; -- 0.050587143817112074
	pesos_i(5233) := b"0000000000000000_0000000000000000_0001101011110011_1011010100111101"; -- 0.10528118836419148
	pesos_i(5234) := b"0000000000000000_0000000000000000_0010100100110100_1010001001111111"; -- 0.16095939246708696
	pesos_i(5235) := b"1111111111111111_1111111111111111_1111001001000001_1001111101001000"; -- -0.05368618492091082
	pesos_i(5236) := b"1111111111111111_1111111111111111_1111100101000101_0010011101000111"; -- -0.02628855249716306
	pesos_i(5237) := b"0000000000000000_0000000000000000_0000100101111011_0111010110100000"; -- 0.03704009194550813
	pesos_i(5238) := b"1111111111111111_1111111111111111_1110110001000000_0011111111010100"; -- -0.07714463311928725
	pesos_i(5239) := b"1111111111111111_1111111111111111_1110100001011000_1001101011100010"; -- -0.09239799472215574
	pesos_i(5240) := b"1111111111111111_1111111111111111_1110111111010010_0110100000001110"; -- -0.06319570222579166
	pesos_i(5241) := b"0000000000000000_0000000000000000_0000000001100110_0110111100000010"; -- 0.0015630131335341562
	pesos_i(5242) := b"0000000000000000_0000000000000000_0010110110111000_1000000011000110"; -- 0.1785965425743084
	pesos_i(5243) := b"1111111111111111_1111111111111111_1110000100001101_1101100101100000"; -- -0.12088242927961328
	pesos_i(5244) := b"1111111111111111_1111111111111111_1110010110101000_1001101110010100"; -- -0.10289600015235004
	pesos_i(5245) := b"0000000000000000_0000000000000000_0010000001001100_0011010001111011"; -- 0.12616279597826574
	pesos_i(5246) := b"0000000000000000_0000000000000000_0001111001001111_1010101000011101"; -- 0.11840308386162803
	pesos_i(5247) := b"0000000000000000_0000000000000000_0011000000001100_1000100110100000"; -- 0.18769130864479966
	pesos_i(5248) := b"1111111111111111_1111111111111111_1110110111100101_0000101001010111"; -- -0.07072387104739791
	pesos_i(5249) := b"1111111111111111_1111111111111111_1111010111011101_1101010001010100"; -- -0.03958390188923587
	pesos_i(5250) := b"1111111111111111_1111111111111111_1101011001011101_1001000101010010"; -- -0.1626347708826056
	pesos_i(5251) := b"1111111111111111_1111111111111111_1111011101111111_0101110010110011"; -- -0.03321285846577132
	pesos_i(5252) := b"1111111111111111_1111111111111111_1110110001110010_0011110110011101"; -- -0.07638182553974696
	pesos_i(5253) := b"1111111111111111_1111111111111111_1101010100011100_0111110011101001"; -- -0.16753405876316957
	pesos_i(5254) := b"1111111111111111_1111111111111111_1111010110011000_0110101111111100"; -- -0.040642977670365676
	pesos_i(5255) := b"0000000000000000_0000000000000000_0000111100010001_1011010100001010"; -- 0.05886394028042063
	pesos_i(5256) := b"0000000000000000_0000000000000000_0001000110100000_0101000001101001"; -- 0.0688524491147049
	pesos_i(5257) := b"0000000000000000_0000000000000000_0000011000011011_1000001111001010"; -- 0.023857342609548464
	pesos_i(5258) := b"0000000000000000_0000000000000000_0000010100010111_1100001101101010"; -- 0.019893849818911995
	pesos_i(5259) := b"1111111111111111_1111111111111111_1101110111000010_0011101000000010"; -- -0.13375508733662103
	pesos_i(5260) := b"1111111111111111_1111111111111111_1111110000110101_0111101001110110"; -- -0.014808984832543521
	pesos_i(5261) := b"1111111111111111_1111111111111111_1110001101111001_0110010010111110"; -- -0.11142893174625208
	pesos_i(5262) := b"1111111111111111_1111111111111111_1101101101101011_1011001111000011"; -- -0.1428878450495807
	pesos_i(5263) := b"1111111111111111_1111111111111111_1111101001101011_0001111110100110"; -- -0.021802923227384294
	pesos_i(5264) := b"1111111111111111_1111111111111111_1110111100010110_1100010110100111"; -- -0.0660587757296791
	pesos_i(5265) := b"1111111111111111_1111111111111111_1110100101001010_1001011111000110"; -- -0.08870555326783641
	pesos_i(5266) := b"1111111111111111_1111111111111111_1101110110110011_1111000011000111"; -- -0.13397307532222194
	pesos_i(5267) := b"0000000000000000_0000000000000000_0000011001100001_1111001000011101"; -- 0.024932033718299444
	pesos_i(5268) := b"1111111111111111_1111111111111111_1110000100010101_1000111001001001"; -- -0.12076483459145079
	pesos_i(5269) := b"1111111111111111_1111111111111111_1101110000100000_1000110101001110"; -- -0.1401282963801073
	pesos_i(5270) := b"1111111111111111_1111111111111111_1101100101111110_1100000001011000"; -- -0.15040967800955735
	pesos_i(5271) := b"1111111111111111_1111111111111111_1111000110110011_1011110001110010"; -- -0.055851194461193625
	pesos_i(5272) := b"0000000000000000_0000000000000000_0001000010010011_0000000110000000"; -- 0.06474313144434528
	pesos_i(5273) := b"0000000000000000_0000000000000000_0010010110010010_0110000110110011"; -- 0.146764856637134
	pesos_i(5274) := b"1111111111111111_1111111111111111_1110001101010101_1000110110001111"; -- -0.11197581540714957
	pesos_i(5275) := b"1111111111111111_1111111111111111_1111000010100101_1100111100011000"; -- -0.05996995597302743
	pesos_i(5276) := b"1111111111111111_1111111111111111_1111011101001111_0110010000011010"; -- -0.033944839234591184
	pesos_i(5277) := b"0000000000000000_0000000000000000_0000011111110010_0100010100100001"; -- 0.03104049745280002
	pesos_i(5278) := b"1111111111111111_1111111111111111_1101101110010000_0001010111011010"; -- -0.14233268180601322
	pesos_i(5279) := b"1111111111111111_1111111111111111_1111101010010111_1000110010110100"; -- -0.021125036388976892
	pesos_i(5280) := b"1111111111111111_1111111111111111_1110011111010101_0100001000000000"; -- -0.09440219407313186
	pesos_i(5281) := b"0000000000000000_0000000000000000_0010100011111001_1100000000000101"; -- 0.16006088372884367
	pesos_i(5282) := b"0000000000000000_0000000000000000_0000010010110110_1001100001000101"; -- 0.018411175585947147
	pesos_i(5283) := b"0000000000000000_0000000000000000_0000100000100010_0100110101011100"; -- 0.03177340978233159
	pesos_i(5284) := b"0000000000000000_0000000000000000_0000010111100001_0111011011010100"; -- 0.02297156027191096
	pesos_i(5285) := b"0000000000000000_0000000000000000_0010000000111111_1111100010010110"; -- 0.12597612050751814
	pesos_i(5286) := b"0000000000000000_0000000000000000_0010011110110100_1001110000100001"; -- 0.1550996380679907
	pesos_i(5287) := b"1111111111111111_1111111111111111_1111011011110100_1110011010111011"; -- -0.035325602888381324
	pesos_i(5288) := b"0000000000000000_0000000000000000_0010001011101101_0010011001111000"; -- 0.13643112599133364
	pesos_i(5289) := b"0000000000000000_0000000000000000_0001010111110110_1111111010001011"; -- 0.08580008412446385
	pesos_i(5290) := b"1111111111111111_1111111111111111_1111010110011010_1110010110010010"; -- -0.040605213142539495
	pesos_i(5291) := b"1111111111111111_1111111111111111_1111011010010000_0011100101000010"; -- -0.036861821455413606
	pesos_i(5292) := b"0000000000000000_0000000000000000_0001101001000001_1100011000000101"; -- 0.10256612422115162
	pesos_i(5293) := b"1111111111111111_1111111111111111_1110101110111000_1000100110000001"; -- -0.07921543695829766
	pesos_i(5294) := b"1111111111111111_1111111111111111_1110001101101100_1001001000001001"; -- -0.11162459634135409
	pesos_i(5295) := b"0000000000000000_0000000000000000_0010111001101011_1000100100000110"; -- 0.1813283576030918
	pesos_i(5296) := b"1111111111111111_1111111111111111_1111011111100000_0000000011000110"; -- -0.03173823514295379
	pesos_i(5297) := b"1111111111111111_1111111111111111_1111110111000000_1011010110010011"; -- -0.008778239779634716
	pesos_i(5298) := b"1111111111111111_1111111111111111_1110110110000111_1001011100001011"; -- -0.0721498105540759
	pesos_i(5299) := b"0000000000000000_0000000000000000_0000110001011011_1101000110110010"; -- 0.04827604867535666
	pesos_i(5300) := b"1111111111111111_1111111111111111_1101110011011000_1000100101100011"; -- -0.13732091263907223
	pesos_i(5301) := b"0000000000000000_0000000000000000_0001101001110101_0100011100111000"; -- 0.10335202338901331
	pesos_i(5302) := b"1111111111111111_1111111111111111_1101100111100010_1101110101110001"; -- -0.1488820648445191
	pesos_i(5303) := b"1111111111111111_1111111111111111_1101101101110011_1101010001100010"; -- -0.1427638303263591
	pesos_i(5304) := b"1111111111111111_1111111111111111_1101110000000101_1000101110111000"; -- -0.14054037819711737
	pesos_i(5305) := b"1111111111111111_1111111111111111_1111110011101011_0100000000110000"; -- -0.0120353585939762
	pesos_i(5306) := b"1111111111111111_1111111111111111_1111010101101111_1101111100111011"; -- -0.04126171882701938
	pesos_i(5307) := b"0000000000000000_0000000000000000_0000001001100000_1111010010111100"; -- 0.009291931105990853
	pesos_i(5308) := b"0000000000000000_0000000000000000_0010100111011001_1100001010100010"; -- 0.16347900829203263
	pesos_i(5309) := b"0000000000000000_0000000000000000_0010100101011010_0000101010110000"; -- 0.16153017813867887
	pesos_i(5310) := b"0000000000000000_0000000000000000_0010000000010111_0110101010111101"; -- 0.12535731424965685
	pesos_i(5311) := b"1111111111111111_1111111111111111_1111100100111100_1110110111101001"; -- -0.026414042033154422
	pesos_i(5312) := b"1111111111111111_1111111111111111_1110101100010010_1000100011010010"; -- -0.08174843671102586
	pesos_i(5313) := b"1111111111111111_1111111111111111_1110110000101011_1100000101110101"; -- -0.07745734108945208
	pesos_i(5314) := b"1111111111111111_1111111111111111_1101101001000001_1111110000000110"; -- -0.1474306568845766
	pesos_i(5315) := b"0000000000000000_0000000000000000_0010011000111000_0110000100110101"; -- 0.14929778609397823
	pesos_i(5316) := b"1111111111111111_1111111111111111_1110010011111011_1100111011011000"; -- -0.1055327151005643
	pesos_i(5317) := b"0000000000000000_0000000000000000_0001011000100100_1000011000000000"; -- 0.08649480347608347
	pesos_i(5318) := b"1111111111111111_1111111111111111_1101011010110010_1010111010010010"; -- -0.16133603042358396
	pesos_i(5319) := b"1111111111111111_1111111111111111_1110111000010010_0010010111110010"; -- -0.07003558015196018
	pesos_i(5320) := b"0000000000000000_0000000000000000_0000110000000010_1110001111110110"; -- 0.04691910513908871
	pesos_i(5321) := b"0000000000000000_0000000000000000_0010011101001000_1111100110100010"; -- 0.15345726199412457
	pesos_i(5322) := b"1111111111111111_1111111111111111_1110110100001001_0100111110011000"; -- -0.07407667677461176
	pesos_i(5323) := b"1111111111111111_1111111111111111_1101110100100100_1011001010110110"; -- -0.13615878156806682
	pesos_i(5324) := b"1111111111111111_1111111111111111_1111011101011110_1011000110011101"; -- -0.033711337165241065
	pesos_i(5325) := b"1111111111111111_1111111111111111_1111100011000011_0010111001110001"; -- -0.028271768001548025
	pesos_i(5326) := b"1111111111111111_1111111111111111_1101110011111000_1001111000010011"; -- -0.1368313984034368
	pesos_i(5327) := b"0000000000000000_0000000000000000_0000111001001110_1110011111111000"; -- 0.0558915120584868
	pesos_i(5328) := b"0000000000000000_0000000000000000_0000110111110111_1100011011101100"; -- 0.05456202745959138
	pesos_i(5329) := b"1111111111111111_1111111111111111_1111101001011010_1010100001010110"; -- -0.02205417531199962
	pesos_i(5330) := b"1111111111111111_1111111111111111_1101000011101111_1010001111001010"; -- -0.1838433868323061
	pesos_i(5331) := b"1111111111111111_1111111111111111_1110111111000101_1001110011101001"; -- -0.06339091606071494
	pesos_i(5332) := b"1111111111111111_1111111111111111_1110011100010110_0100100001110011"; -- -0.09731623829772225
	pesos_i(5333) := b"0000000000000000_0000000000000000_0010000111010101_1101111100101111"; -- 0.13216967477563993
	pesos_i(5334) := b"1111111111111111_1111111111111111_1101001101000001_1101110100001011"; -- -0.17477625351520468
	pesos_i(5335) := b"1111111111111111_1111111111111111_1111011101110111_1100011001001110"; -- -0.033328634311759926
	pesos_i(5336) := b"0000000000000000_0000000000000000_0010001000000101_0010111111001101"; -- 0.13289164310884466
	pesos_i(5337) := b"0000000000000000_0000000000000000_0000111110101011_0100000010100101"; -- 0.06120685601608032
	pesos_i(5338) := b"0000000000000000_0000000000000000_0010010110100000_0101100110111111"; -- 0.14697800562544716
	pesos_i(5339) := b"1111111111111111_1111111111111111_1110010010011010_1110111011110011"; -- -0.10701090406986005
	pesos_i(5340) := b"1111111111111111_1111111111111111_1111000100001000_1110001011001111"; -- -0.0584581607521351
	pesos_i(5341) := b"1111111111111111_1111111111111111_1111110111011001_0101000100000111"; -- -0.00840276309485928
	pesos_i(5342) := b"0000000000000000_0000000000000000_0010110000100000_0010101101110011"; -- 0.17236587107717088
	pesos_i(5343) := b"1111111111111111_1111111111111111_1111101001111010_0110111000100010"; -- -0.021569363270143582
	pesos_i(5344) := b"1111111111111111_1111111111111111_1101101000011100_0010001110011111"; -- -0.1480081306720514
	pesos_i(5345) := b"0000000000000000_0000000000000000_0010010000011100_0101101011010001"; -- 0.14105765914592383
	pesos_i(5346) := b"1111111111111111_1111111111111111_1110100110100011_1010000001001100"; -- -0.08734701283155687
	pesos_i(5347) := b"1111111111111111_1111111111111111_1111111101010000_1110000011101011"; -- -0.0026721407069910303
	pesos_i(5348) := b"0000000000000000_0000000000000000_0000101110110010_0111111001010100"; -- 0.04569234415045239
	pesos_i(5349) := b"0000000000000000_0000000000000000_0001000000000100_0001100110100111"; -- 0.06256256416278401
	pesos_i(5350) := b"0000000000000000_0000000000000000_0001010001011000_0010011000100010"; -- 0.07947004643284744
	pesos_i(5351) := b"1111111111111111_1111111111111111_1110010000111000_1100111011110001"; -- -0.10850817319594698
	pesos_i(5352) := b"1111111111111111_1111111111111111_1101001100010001_1110101000000110"; -- -0.1755079016218974
	pesos_i(5353) := b"0000000000000000_0000000000000000_0001001010110010_1111110101111101"; -- 0.07304367364184482
	pesos_i(5354) := b"0000000000000000_0000000000000000_0000011110101011_1001001001110100"; -- 0.029961732310938335
	pesos_i(5355) := b"1111111111111111_1111111111111111_1111100011010100_0100111111110111"; -- -0.028010370554376187
	pesos_i(5356) := b"0000000000000000_0000000000000000_0001000001110011_1010101010100111"; -- 0.06426493238665891
	pesos_i(5357) := b"1111111111111111_1111111111111111_1111101010110111_1100111001011000"; -- -0.02063284246146615
	pesos_i(5358) := b"0000000000000000_0000000000000000_0000100111111011_0110000111011010"; -- 0.038992038563629844
	pesos_i(5359) := b"0000000000000000_0000000000000000_0001111101000001_1110100111101110"; -- 0.12209951454580031
	pesos_i(5360) := b"0000000000000000_0000000000000000_0001110100011100_0100101001100111"; -- 0.11371293073734254
	pesos_i(5361) := b"0000000000000000_0000000000000000_0010001111011100_0100011101011011"; -- 0.14007993669079927
	pesos_i(5362) := b"0000000000000000_0000000000000000_0000000100000000_1110110100111010"; -- 0.003920389813088862
	pesos_i(5363) := b"0000000000000000_0000000000000000_0001000011011100_0110011101110000"; -- 0.06586309895127991
	pesos_i(5364) := b"0000000000000000_0000000000000000_0000000100001101_0011010101100000"; -- 0.004107795639315381
	pesos_i(5365) := b"1111111111111111_1111111111111111_1111000010010101_0011000011011000"; -- -0.06022352910397215
	pesos_i(5366) := b"0000000000000000_0000000000000000_0010010001101000_0011101011011110"; -- 0.14221542288832986
	pesos_i(5367) := b"1111111111111111_1111111111111111_1110110000111010_1110011111010101"; -- -0.07722617190483717
	pesos_i(5368) := b"1111111111111111_1111111111111111_1110010101011101_0101100111010100"; -- -0.1040443284322669
	pesos_i(5369) := b"1111111111111111_1111111111111111_1110011100110001_0011000101001001"; -- -0.0969056317693725
	pesos_i(5370) := b"0000000000000000_0000000000000000_0000101100011111_1010000110010001"; -- 0.04345140250316637
	pesos_i(5371) := b"1111111111111111_1111111111111111_1101101100100001_1101001101001100"; -- -0.14401511578790357
	pesos_i(5372) := b"1111111111111111_1111111111111111_1111100010001001_0100111101000100"; -- -0.029154821327566634
	pesos_i(5373) := b"0000000000000000_0000000000000000_0000011100101010_0100101000001101"; -- 0.027989032975271683
	pesos_i(5374) := b"0000000000000000_0000000000000000_0001010010000111_0101000001101101"; -- 0.08018973027332184
	pesos_i(5375) := b"0000000000000000_0000000000000000_0000110101000011_0110100000101111"; -- 0.05180979872051179
	pesos_i(5376) := b"1111111111111111_1111111111111111_1111000110001110_0011010100010111"; -- -0.05642383763469311
	pesos_i(5377) := b"0000000000000000_0000000000000000_0000000110111001_1100011011010001"; -- 0.006740976399041833
	pesos_i(5378) := b"0000000000000000_0000000000000000_0000101100001100_1100011010011010"; -- 0.04316369302424475
	pesos_i(5379) := b"0000000000000000_0000000000000000_0001100101110110_0101001101010010"; -- 0.09946175337253799
	pesos_i(5380) := b"0000000000000000_0000000000000000_0001001000110000_1000010011001111"; -- 0.07105283791058868
	pesos_i(5381) := b"0000000000000000_0000000000000000_0010101111000111_1111110110011101"; -- 0.17102036564403567
	pesos_i(5382) := b"1111111111111111_1111111111111111_1110011111100000_0011010011001001"; -- -0.09423513511383172
	pesos_i(5383) := b"0000000000000000_0000000000000000_0000001010001001_0000111110111010"; -- 0.009903891504245865
	pesos_i(5384) := b"1111111111111111_1111111111111111_1100110001110011_1101111000000001"; -- -0.20135700688882366
	pesos_i(5385) := b"1111111111111111_1111111111111111_1110101001011011_1110000000010000"; -- -0.0845355950783715
	pesos_i(5386) := b"0000000000000000_0000000000000000_0001101101110110_1110101001111101"; -- 0.1072832637920722
	pesos_i(5387) := b"1111111111111111_1111111111111111_1111111011110001_0011001110010001"; -- -0.004132058228020094
	pesos_i(5388) := b"1111111111111111_1111111111111111_1111010110000110_0010111100010100"; -- -0.040921266144767224
	pesos_i(5389) := b"0000000000000000_0000000000000000_0010100001010001_1101100011000000"; -- 0.15749888111083105
	pesos_i(5390) := b"0000000000000000_0000000000000000_0000101110111100_1000100100110110"; -- 0.04584558070778883
	pesos_i(5391) := b"0000000000000000_0000000000000000_0000000011111111_1111011110111011"; -- 0.003905757195198952
	pesos_i(5392) := b"0000000000000000_0000000000000000_0001110011101000_0000101100001101"; -- 0.11291569782221358
	pesos_i(5393) := b"1111111111111111_1111111111111111_1110100000111100_1010100000110110"; -- -0.09282444645455147
	pesos_i(5394) := b"1111111111111111_1111111111111111_1110101100110111_0111000110100100"; -- -0.0811852430131491
	pesos_i(5395) := b"0000000000000000_0000000000000000_0000001001100010_0010011111010000"; -- 0.009310234329842041
	pesos_i(5396) := b"0000000000000000_0000000000000000_0001100111011011_0100100110111010"; -- 0.10100231915347417
	pesos_i(5397) := b"0000000000000000_0000000000000000_0000011001011011_1001011001000110"; -- 0.024835006835641233
	pesos_i(5398) := b"1111111111111111_1111111111111111_1110110011000111_1011011101110100"; -- -0.07507756631141643
	pesos_i(5399) := b"1111111111111111_1111111111111111_1111010111101001_0100110000011101"; -- -0.03940891538863932
	pesos_i(5400) := b"1111111111111111_1111111111111111_1101011111010101_1100000111111111"; -- -0.15689456476237804
	pesos_i(5401) := b"1111111111111111_1111111111111111_1111111010000000_1010010000111100"; -- -0.0058495857938047685
	pesos_i(5402) := b"1111111111111111_1111111111111111_1101111100001110_1010100101010011"; -- -0.12868253444924949
	pesos_i(5403) := b"0000000000000000_0000000000000000_0001111010110110_1111001100001110"; -- 0.11997908676898096
	pesos_i(5404) := b"1111111111111111_1111111111111111_1111001010111011_0100010010010110"; -- -0.05183001844527445
	pesos_i(5405) := b"0000000000000000_0000000000000000_0000110111000010_0001000110010000"; -- 0.053742501956323886
	pesos_i(5406) := b"0000000000000000_0000000000000000_0001111010001011_1101100011010101"; -- 0.11932139594847128
	pesos_i(5407) := b"1111111111111111_1111111111111111_1101111111001001_1101111110100101"; -- -0.12582590313355907
	pesos_i(5408) := b"1111111111111111_1111111111111111_1111011110010010_1100010100101111"; -- -0.03291671365517912
	pesos_i(5409) := b"1111111111111111_1111111111111111_1101011001110110_1000010111011010"; -- -0.1622539847878263
	pesos_i(5410) := b"0000000000000000_0000000000000000_0000011100101010_0100011011110010"; -- 0.027988847731843677
	pesos_i(5411) := b"0000000000000000_0000000000000000_0010000101110001_0001100001101110"; -- 0.1306319492164674
	pesos_i(5412) := b"1111111111111111_1111111111111111_1101001011000100_1000011100001101"; -- -0.17668872773985222
	pesos_i(5413) := b"0000000000000000_0000000000000000_0000011010011010_0110100011010011"; -- 0.02579360164144923
	pesos_i(5414) := b"0000000000000000_0000000000000000_0000000011001001_1110110110000110"; -- 0.003081174194834323
	pesos_i(5415) := b"1111111111111111_1111111111111111_1101101101101110_1111010010100101"; -- -0.1428382011451609
	pesos_i(5416) := b"1111111111111111_1111111111111111_1110000000010100_0000110011001011"; -- -0.12469406179201725
	pesos_i(5417) := b"1111111111111111_1111111111111111_1110100010011110_1110110000100100"; -- -0.09132503622198251
	pesos_i(5418) := b"0000000000000000_0000000000000000_0001011010001111_0011001001100111"; -- 0.08812251110678299
	pesos_i(5419) := b"1111111111111111_1111111111111111_1110001111000000_1101010001000110"; -- -0.11033891005349435
	pesos_i(5420) := b"0000000000000000_0000000000000000_0010100100101000_1110010011110101"; -- 0.16078024840562422
	pesos_i(5421) := b"0000000000000000_0000000000000000_0010101101111000_0000001001100101"; -- 0.16979994729886946
	pesos_i(5422) := b"1111111111111111_1111111111111111_1111111011011001_0111110110011110"; -- -0.004493855304400353
	pesos_i(5423) := b"0000000000000000_0000000000000000_0001111101100110_0111110000001000"; -- 0.12265753925587783
	pesos_i(5424) := b"1111111111111111_1111111111111111_1110001101001001_1110100100111001"; -- -0.11215345723560215
	pesos_i(5425) := b"0000000000000000_0000000000000000_0001100100111011_1101011111000100"; -- 0.09856937922371593
	pesos_i(5426) := b"0000000000000000_0000000000000000_0010001001101100_0010110101110001"; -- 0.13446315771134973
	pesos_i(5427) := b"0000000000000000_0000000000000000_0000011110101001_0011101000111110"; -- 0.029925956824133123
	pesos_i(5428) := b"1111111111111111_1111111111111111_1101010100110001_1011011101111000"; -- -0.16721013374932525
	pesos_i(5429) := b"1111111111111111_1111111111111111_1110101011110000_0011110000010010"; -- -0.08227181005820616
	pesos_i(5430) := b"0000000000000000_0000000000000000_0001101001000100_0001111100010001"; -- 0.10260194940431905
	pesos_i(5431) := b"1111111111111111_1111111111111111_1111110111110001_1100100101010111"; -- -0.008029381098244479
	pesos_i(5432) := b"1111111111111111_1111111111111111_1101110001000110_1111111011100111"; -- -0.13954169133645206
	pesos_i(5433) := b"1111111111111111_1111111111111111_1111000101111010_0111111111001001"; -- -0.05672456110912221
	pesos_i(5434) := b"0000000000000000_0000000000000000_0001100100100001_0111110101011100"; -- 0.09816726212888287
	pesos_i(5435) := b"0000000000000000_0000000000000000_0001110101110001_0111000001010111"; -- 0.11501218915100896
	pesos_i(5436) := b"1111111111111111_1111111111111111_1111111011001111_0011110010101100"; -- -0.00465031441912887
	pesos_i(5437) := b"0000000000000000_0000000000000000_0010101111010010_0110100100010101"; -- 0.17117935904744683
	pesos_i(5438) := b"1111111111111111_1111111111111111_1101000110110011_1010110000000001"; -- -0.1808521744750385
	pesos_i(5439) := b"0000000000000000_0000000000000000_0010010111111000_1011001000011110"; -- 0.1483260463955351
	pesos_i(5440) := b"0000000000000000_0000000000000000_0010000010100101_1101100010010000"; -- 0.12753060828249732
	pesos_i(5441) := b"1111111111111111_1111111111111111_1110100010010101_1100011100001010"; -- -0.09146457688337407
	pesos_i(5442) := b"1111111111111111_1111111111111111_1101101100000110_0101111011101110"; -- -0.14443403897447812
	pesos_i(5443) := b"0000000000000000_0000000000000000_0001010000100000_0100000100001111"; -- 0.07861715893225599
	pesos_i(5444) := b"0000000000000000_0000000000000000_0000100011000111_1110000100101100"; -- 0.034299920386990895
	pesos_i(5445) := b"0000000000000000_0000000000000000_0010010101100100_0101010010001000"; -- 0.14606216741488903
	pesos_i(5446) := b"0000000000000000_0000000000000000_0001100011000101_1011100011000100"; -- 0.09676699442251054
	pesos_i(5447) := b"1111111111111111_1111111111111111_1111101110110101_0100101011001110"; -- -0.016764950493529145
	pesos_i(5448) := b"1111111111111111_1111111111111111_1111101110110110_0001001010010110"; -- -0.016753042524020743
	pesos_i(5449) := b"0000000000000000_0000000000000000_0000011100110000_0100000000111101"; -- 0.028080000747128325
	pesos_i(5450) := b"0000000000000000_0000000000000000_0000111110111110_0011010101000001"; -- 0.06149609415934458
	pesos_i(5451) := b"0000000000000000_0000000000000000_0000010010001010_1111111000110000"; -- 0.017745863744223888
	pesos_i(5452) := b"1111111111111111_1111111111111111_1111011001010001_0100111111110000"; -- -0.03782177352930925
	pesos_i(5453) := b"1111111111111111_1111111111111111_1111001010010111_0100111011000111"; -- -0.052378727450328864
	pesos_i(5454) := b"1111111111111111_1111111111111111_1101010010101011_0010110001011100"; -- -0.16926310312946743
	pesos_i(5455) := b"1111111111111111_1111111111111111_1101110010101110_0001110111000001"; -- -0.13796819711817984
	pesos_i(5456) := b"0000000000000000_0000000000000000_0001110011011111_0011000101111110"; -- 0.11278065986032534
	pesos_i(5457) := b"0000000000000000_0000000000000000_0001011011011011_1010111100010001"; -- 0.08928960966106206
	pesos_i(5458) := b"0000000000000000_0000000000000000_0001001011001100_1000000011110101"; -- 0.07343297930203567
	pesos_i(5459) := b"1111111111111111_1111111111111111_1111101110101111_1001101001111000"; -- -0.01685175488230435
	pesos_i(5460) := b"0000000000000000_0000000000000000_0000100111000000_0100001100010101"; -- 0.0380899359715092
	pesos_i(5461) := b"1111111111111111_1111111111111111_1111111111110110_0011011100010111"; -- -0.0001493042538499265
	pesos_i(5462) := b"0000000000000000_0000000000000000_0001110101010111_1000001011101100"; -- 0.11461656817363264
	pesos_i(5463) := b"1111111111111111_1111111111111111_1111100110000110_1110101110101000"; -- -0.025285026026842523
	pesos_i(5464) := b"1111111111111111_1111111111111111_1111110011000111_1110010010010110"; -- -0.012574876116710819
	pesos_i(5465) := b"1111111111111111_1111111111111111_1111101111101010_0111010101110010"; -- -0.015953693037454586
	pesos_i(5466) := b"0000000000000000_0000000000000000_0010110001010110_1101101001110000"; -- 0.17320027568758703
	pesos_i(5467) := b"1111111111111111_1111111111111111_1101011111101110_0111001011001100"; -- -0.15651781583093174
	pesos_i(5468) := b"0000000000000000_0000000000000000_0000100011011110_0001001101101110"; -- 0.034638609304150476
	pesos_i(5469) := b"1111111111111111_1111111111111111_1111010001010011_1111111000001001"; -- -0.04559337879569027
	pesos_i(5470) := b"1111111111111111_1111111111111111_1111111000101111_1111000101111001"; -- -0.007080943945978081
	pesos_i(5471) := b"1111111111111111_1111111111111111_1101010110111010_1111111011000001"; -- -0.16511543060973335
	pesos_i(5472) := b"1111111111111111_1111111111111111_1101100010100001_1010010111110001"; -- -0.15378344415298373
	pesos_i(5473) := b"1111111111111111_1111111111111111_1110001010111010_1011000110010000"; -- -0.11433878173282175
	pesos_i(5474) := b"1111111111111111_1111111111111111_1110110101101001_0000100001110100"; -- -0.07261607341427687
	pesos_i(5475) := b"0000000000000000_0000000000000000_0000010111101101_1000111110001000"; -- 0.023156138121902325
	pesos_i(5476) := b"0000000000000000_0000000000000000_0010000001101110_1011001110101111"; -- 0.12668917679168878
	pesos_i(5477) := b"1111111111111111_1111111111111111_1110001001000010_1010110100110000"; -- -0.11617009709915073
	pesos_i(5478) := b"0000000000000000_0000000000000000_0001100011000000_0001110100111100"; -- 0.09668143008831416
	pesos_i(5479) := b"0000000000000000_0000000000000000_0001011000011000_1100000010101101"; -- 0.08631519530849138
	pesos_i(5480) := b"0000000000000000_0000000000000000_0000110011000100_1101101110011000"; -- 0.049878811432262915
	pesos_i(5481) := b"1111111111111111_1111111111111111_1111001111101000_0110010110100001"; -- -0.047235153320252354
	pesos_i(5482) := b"1111111111111111_1111111111111111_1111111000000001_0111010000100101"; -- -0.007790318536319732
	pesos_i(5483) := b"0000000000000000_0000000000000000_0000001101011000_0101110010000010"; -- 0.013067037249819877
	pesos_i(5484) := b"0000000000000000_0000000000000000_0010011100111100_1100001010001000"; -- 0.1532708722933576
	pesos_i(5485) := b"0000000000000000_0000000000000000_0000101101001111_1100111111010100"; -- 0.04418658186361686
	pesos_i(5486) := b"1111111111111111_1111111111111111_1101110110100011_0001111011111110"; -- -0.13422972017405094
	pesos_i(5487) := b"0000000000000000_0000000000000000_0010011101111111_0010001000101110"; -- 0.15428365348079864
	pesos_i(5488) := b"0000000000000000_0000000000000000_0001010111101101_1011000001100101"; -- 0.08565809693059859
	pesos_i(5489) := b"1111111111111111_1111111111111111_1111000001110100_0111010100110000"; -- -0.06072299563685985
	pesos_i(5490) := b"1111111111111111_1111111111111111_1111010000010001_0000001010010000"; -- -0.04661544783546118
	pesos_i(5491) := b"1111111111111111_1111111111111111_1111100101110100_1100010111111100"; -- -0.025561929739818662
	pesos_i(5492) := b"1111111111111111_1111111111111111_1111010000000100_0110000111011011"; -- -0.04680813227759691
	pesos_i(5493) := b"1111111111111111_1111111111111111_1101101101000110_1100101100101010"; -- -0.1434510251577776
	pesos_i(5494) := b"1111111111111111_1111111111111111_1111100100100010_1001000111111011"; -- -0.02681624997681027
	pesos_i(5495) := b"1111111111111111_1111111111111111_1111100100011010_1000001010000100"; -- -0.026939242116153308
	pesos_i(5496) := b"0000000000000000_0000000000000000_0010101111000111_0101111110110101"; -- 0.1710109535107762
	pesos_i(5497) := b"1111111111111111_1111111111111111_1110001100111111_1111100010010110"; -- -0.11230512929658402
	pesos_i(5498) := b"1111111111111111_1111111111111111_1101011100001101_1101110101011000"; -- -0.15994469259790695
	pesos_i(5499) := b"0000000000000000_0000000000000000_0001010100001110_0010101000001100"; -- 0.0822473792899075
	pesos_i(5500) := b"1111111111111111_1111111111111111_1101101001100100_1111111110011100"; -- -0.1468963855465185
	pesos_i(5501) := b"0000000000000000_0000000000000000_0010011001011011_1000110010010100"; -- 0.1498344288210802
	pesos_i(5502) := b"1111111111111111_1111111111111111_1110111010011101_0110111001011101"; -- -0.06791029194765105
	pesos_i(5503) := b"0000000000000000_0000000000000000_0001010110111001_1101111110010000"; -- 0.08486745137248076
	pesos_i(5504) := b"0000000000000000_0000000000000000_0010100000111111_0001101010101000"; -- 0.1572128925817213
	pesos_i(5505) := b"1111111111111111_1111111111111111_1110010100000000_1000110001001001"; -- -0.10546038825615851
	pesos_i(5506) := b"1111111111111111_1111111111111111_1110001100010100_0101110101000001"; -- -0.11297051586860865
	pesos_i(5507) := b"1111111111111111_1111111111111111_1101110101000111_1010010111101101"; -- -0.13562548614209938
	pesos_i(5508) := b"1111111111111111_1111111111111111_1101111101010000_0011101001011000"; -- -0.1276820693077145
	pesos_i(5509) := b"1111111111111111_1111111111111111_1111000011110011_1000110111100111"; -- -0.058783656202688814
	pesos_i(5510) := b"0000000000000000_0000000000000000_0001010000011010_1110110011011001"; -- 0.0785358456979956
	pesos_i(5511) := b"0000000000000000_0000000000000000_0001101000101000_1011011101110110"; -- 0.10218378657165765
	pesos_i(5512) := b"0000000000000000_0000000000000000_0010011111011110_0110001100011101"; -- 0.15573710879257535
	pesos_i(5513) := b"0000000000000000_0000000000000000_0010100000010110_1111001010001100"; -- 0.15660015022572513
	pesos_i(5514) := b"1111111111111111_1111111111111111_1110100010111101_0010100101010010"; -- -0.09086362606250056
	pesos_i(5515) := b"1111111111111111_1111111111111111_1101111101100111_1100000110110101"; -- -0.12732304886284618
	pesos_i(5516) := b"1111111111111111_1111111111111111_1110100011110110_1001111110011010"; -- -0.08998682485993612
	pesos_i(5517) := b"1111111111111111_1111111111111111_1111101110110011_1101001110101100"; -- -0.016787310118984846
	pesos_i(5518) := b"0000000000000000_0000000000000000_0001111011100101_0111100111011011"; -- 0.12068902587197886
	pesos_i(5519) := b"1111111111111111_1111111111111111_1111101010110101_0100100011100111"; -- -0.020671313815202444
	pesos_i(5520) := b"1111111111111111_1111111111111111_1110101100010011_1100110011110111"; -- -0.08172911626350715
	pesos_i(5521) := b"0000000000000000_0000000000000000_0001101010011101_0111111101010001"; -- 0.10396571863152694
	pesos_i(5522) := b"0000000000000000_0000000000000000_0000100000001001_0010111011011111"; -- 0.031390122943314676
	pesos_i(5523) := b"0000000000000000_0000000000000000_0000001101010010_1010110001100001"; -- 0.012980245291528426
	pesos_i(5524) := b"1111111111111111_1111111111111111_1110100100011110_0111011101110001"; -- -0.08937886704100122
	pesos_i(5525) := b"0000000000000000_0000000000000000_0001111001101001_1010001110001010"; -- 0.11879942057857446
	pesos_i(5526) := b"0000000000000000_0000000000000000_0001011011111110_1011001110011000"; -- 0.0898239370280217
	pesos_i(5527) := b"0000000000000000_0000000000000000_0001110111111010_0110010101011000"; -- 0.11710198788240189
	pesos_i(5528) := b"0000000000000000_0000000000000000_0000101100110001_1000101000000011"; -- 0.04372465670963379
	pesos_i(5529) := b"0000000000000000_0000000000000000_0000110101100010_1101111100111101"; -- 0.05228991727736439
	pesos_i(5530) := b"0000000000000000_0000000000000000_0001011000101000_1100110000010000"; -- 0.0865600146643554
	pesos_i(5531) := b"1111111111111111_1111111111111111_1110001101010110_1010110001100000"; -- -0.11195871968852451
	pesos_i(5532) := b"1111111111111111_1111111111111111_1101111010001010_1101011001010110"; -- -0.1306940117565195
	pesos_i(5533) := b"1111111111111111_1111111111111111_1110001110001010_1111110110100011"; -- -0.11116041922939729
	pesos_i(5534) := b"0000000000000000_0000000000000000_0000001101011110_0001000101100010"; -- 0.013154112270999356
	pesos_i(5535) := b"0000000000000000_0000000000000000_0000011111111100_0010101010011110"; -- 0.031191504940866394
	pesos_i(5536) := b"0000000000000000_0000000000000000_0000111101110001_1011010110100001"; -- 0.06032881916286156
	pesos_i(5537) := b"0000000000000000_0000000000000000_0000001101101111_0010001001001101"; -- 0.013414520136489975
	pesos_i(5538) := b"1111111111111111_1111111111111111_1110010101011111_1101111110100011"; -- -0.10400583522446624
	pesos_i(5539) := b"0000000000000000_0000000000000000_0010000010101010_0001011111001000"; -- 0.12759541167968885
	pesos_i(5540) := b"0000000000000000_0000000000000000_0001101011101100_0000011100101111"; -- 0.10516400246225314
	pesos_i(5541) := b"1111111111111111_1111111111111111_1110001011000010_1001111101011110"; -- -0.11421779600007527
	pesos_i(5542) := b"0000000000000000_0000000000000000_0010100001111100_1111010000111111"; -- 0.15815664813258065
	pesos_i(5543) := b"0000000000000000_0000000000000000_0001101000011100_1110111100100001"; -- 0.10200399927166168
	pesos_i(5544) := b"1111111111111111_1111111111111111_1101011110010000_1101000011000101"; -- -0.15794654077639592
	pesos_i(5545) := b"1111111111111111_1111111111111111_1101010001010101_0011110001100100"; -- -0.17057440330356835
	pesos_i(5546) := b"0000000000000000_0000000000000000_0001111111011101_1011001100100000"; -- 0.12447661909732854
	pesos_i(5547) := b"1111111111111111_1111111111111111_1110101010001111_0011000100010011"; -- -0.08375256803265166
	pesos_i(5548) := b"0000000000000000_0000000000000000_0010110101110111_0001101101101011"; -- 0.177598680145113
	pesos_i(5549) := b"1111111111111111_1111111111111111_1111010011111101_1110011001000111"; -- -0.04300080073597158
	pesos_i(5550) := b"1111111111111111_1111111111111111_1101101000101000_0111110110001000"; -- -0.14781966618755277
	pesos_i(5551) := b"1111111111111111_1111111111111111_1100110001100000_0100000100010101"; -- -0.20165627700585315
	pesos_i(5552) := b"0000000000000000_0000000000000000_0001101100100110_1101111001100011"; -- 0.10606183928574867
	pesos_i(5553) := b"1111111111111111_1111111111111111_1110101011011110_1110100111000100"; -- -0.08253611524174637
	pesos_i(5554) := b"1111111111111111_1111111111111111_1101000100010010_1110000001101010"; -- -0.18330571557243522
	pesos_i(5555) := b"1111111111111111_1111111111111111_1101111010000100_1110011100010110"; -- -0.13078456601266536
	pesos_i(5556) := b"1111111111111111_1111111111111111_1101101110111110_1000101111110110"; -- -0.14162373776572337
	pesos_i(5557) := b"0000000000000000_0000000000000000_0001101111001100_1000000101010000"; -- 0.10858925064987991
	pesos_i(5558) := b"1111111111111111_1111111111111111_1101011110100101_0101010101101001"; -- -0.1576334589702993
	pesos_i(5559) := b"0000000000000000_0000000000000000_0001010100011000_1110000110101000"; -- 0.08241091120479295
	pesos_i(5560) := b"1111111111111111_1111111111111111_1111111000110000_1011111001011000"; -- -0.007068732792123278
	pesos_i(5561) := b"1111111111111111_1111111111111111_1101101001111010_1010110101101111"; -- -0.1465655902614607
	pesos_i(5562) := b"1111111111111111_1111111111111111_1111101100111010_1111011101011010"; -- -0.018631496872230972
	pesos_i(5563) := b"1111111111111111_1111111111111111_1111100000101000_0000100001100100"; -- -0.030639148301376942
	pesos_i(5564) := b"1111111111111111_1111111111111111_1110110000010111_1001000111111110"; -- -0.07776534599480445
	pesos_i(5565) := b"0000000000000000_0000000000000000_0010100001010100_1111100001011111"; -- 0.15754654234021015
	pesos_i(5566) := b"0000000000000000_0000000000000000_0001011000000110_1111101101111111"; -- 0.08604404305031318
	pesos_i(5567) := b"0000000000000000_0000000000000000_0001101111101010_0000110000001110"; -- 0.10904002504816887
	pesos_i(5568) := b"1111111111111111_1111111111111111_1111101110100000_1100000100010111"; -- -0.017078334648885612
	pesos_i(5569) := b"0000000000000000_0000000000000000_0010001100111101_1000100011101010"; -- 0.13765769691208368
	pesos_i(5570) := b"1111111111111111_1111111111111111_1111110111011100_1101100110000011"; -- -0.00834885164710608
	pesos_i(5571) := b"0000000000000000_0000000000000000_0001011011111011_1100111011011111"; -- 0.08977978661849303
	pesos_i(5572) := b"1111111111111111_1111111111111111_1110010101000000_1000101100111001"; -- -0.1044838891416545
	pesos_i(5573) := b"1111111111111111_1111111111111111_1110011110000001_0100000010100001"; -- -0.09568401410596374
	pesos_i(5574) := b"1111111111111111_1111111111111111_1111111110001111_0010010101010011"; -- -0.001722018574157723
	pesos_i(5575) := b"0000000000000000_0000000000000000_0001001111000000_0001011111011100"; -- 0.07714985955472621
	pesos_i(5576) := b"1111111111111111_1111111111111111_1110110110111011_0011101111001010"; -- -0.07136179262309464
	pesos_i(5577) := b"1111111111111111_1111111111111111_1110011110010000_0010000010010011"; -- -0.09545704270099972
	pesos_i(5578) := b"1111111111111111_1111111111111111_1111011101111001_1100101101111011"; -- -0.03329780803416957
	pesos_i(5579) := b"0000000000000000_0000000000000000_0000001000111111_0010010011100111"; -- 0.008776003204718125
	pesos_i(5580) := b"0000000000000000_0000000000000000_0001110111001001_1100111100000101"; -- 0.11636060591745961
	pesos_i(5581) := b"0000000000000000_0000000000000000_0001100001111110_0000101111001011"; -- 0.09567331022419732
	pesos_i(5582) := b"0000000000000000_0000000000000000_0001111110001010_1010100000110110"; -- 0.12320948895179637
	pesos_i(5583) := b"0000000000000000_0000000000000000_0001011111001001_0011001000001100"; -- 0.09291374963635357
	pesos_i(5584) := b"1111111111111111_1111111111111111_1111011001110111_0010010010001000"; -- -0.03724452656089636
	pesos_i(5585) := b"1111111111111111_1111111111111111_1110000110100110_0110101101100100"; -- -0.11855439013857375
	pesos_i(5586) := b"1111111111111111_1111111111111111_1111110011000111_0110101000111011"; -- -0.012582169124083727
	pesos_i(5587) := b"1111111111111111_1111111111111111_1111010100111011_1110111110000111"; -- -0.042054204549938946
	pesos_i(5588) := b"0000000000000000_0000000000000000_0010001101001111_1100000110110101"; -- 0.1379357400625214
	pesos_i(5589) := b"0000000000000000_0000000000000000_0001110000100011_0101010010010110"; -- 0.10991409940450535
	pesos_i(5590) := b"0000000000000000_0000000000000000_0010000110001000_1000111011100011"; -- 0.13098996200235538
	pesos_i(5591) := b"1111111111111111_1111111111111111_1101001001001101_0101010110101001"; -- -0.17850746740973908
	pesos_i(5592) := b"1111111111111111_1111111111111111_1100101000011101_0001111110100110"; -- -0.21049310874999447
	pesos_i(5593) := b"1111111111111111_1111111111111111_1101100111100011_1011111101110010"; -- -0.14886859375382339
	pesos_i(5594) := b"1111111111111111_1111111111111111_1111001110110111_0010010001000111"; -- -0.04798672930388655
	pesos_i(5595) := b"1111111111111111_1111111111111111_1111001110011100_1111011011011001"; -- -0.048386165699732676
	pesos_i(5596) := b"0000000000000000_0000000000000000_0000000100011111_1000110100010000"; -- 0.004387680332004481
	pesos_i(5597) := b"0000000000000000_0000000000000000_0001101110000111_1101001100010110"; -- 0.10754126820031976
	pesos_i(5598) := b"1111111111111111_1111111111111111_1101111011111111_1001100100011101"; -- -0.12891238253142429
	pesos_i(5599) := b"1111111111111111_1111111111111111_1110010001101011_1011001011010101"; -- -0.10773165031317623
	pesos_i(5600) := b"1111111111111111_1111111111111111_1111010011110001_1011010000010100"; -- -0.04318689844830639
	pesos_i(5601) := b"0000000000000000_0000000000000000_0000100101100101_0001101000001111"; -- 0.036698940970456714
	pesos_i(5602) := b"0000000000000000_0000000000000000_0001101011101101_1111111111011001"; -- 0.10519408271331791
	pesos_i(5603) := b"0000000000000000_0000000000000000_0001010011000001_1011010111111101"; -- 0.0810807935365466
	pesos_i(5604) := b"1111111111111111_1111111111111111_1111111000101011_0111111010010001"; -- -0.007148828164091335
	pesos_i(5605) := b"0000000000000000_0000000000000000_0001010001000001_1100111101010001"; -- 0.07912917841694699
	pesos_i(5606) := b"1111111111111111_1111111111111111_1110010110001111_0011111001011010"; -- -0.10328302664938055
	pesos_i(5607) := b"1111111111111111_1111111111111111_1110000111000110_1010101101100000"; -- -0.11806229502142296
	pesos_i(5608) := b"1111111111111111_1111111111111111_1110111011001101_0110000101111000"; -- -0.06717863867074227
	pesos_i(5609) := b"1111111111111111_1111111111111111_1110101001011010_0001000100001011"; -- -0.08456319315881523
	pesos_i(5610) := b"0000000000000000_0000000000000000_0010001100010001_1011010011001111"; -- 0.1369889264623837
	pesos_i(5611) := b"1111111111111111_1111111111111111_1110000111100010_0110101001100111"; -- -0.11763892152410921
	pesos_i(5612) := b"0000000000000000_0000000000000000_0001000001101010_0011010110100011"; -- 0.06412062860659892
	pesos_i(5613) := b"0000000000000000_0000000000000000_0000111011100001_0111011010011000"; -- 0.05812779637978541
	pesos_i(5614) := b"0000000000000000_0000000000000000_0010011011111011_1100111100100001"; -- 0.15227980190770712
	pesos_i(5615) := b"1111111111111111_1111111111111111_1110111000010111_1101010111000111"; -- -0.06994880578900556
	pesos_i(5616) := b"0000000000000000_0000000000000000_0001101011011001_0011010111001110"; -- 0.10487686421746537
	pesos_i(5617) := b"1111111111111111_1111111111111111_1111100100110111_1100111011000111"; -- -0.02649219160500405
	pesos_i(5618) := b"1111111111111111_1111111111111111_1101111010011010_1110100011010001"; -- -0.13044876944785988
	pesos_i(5619) := b"1111111111111111_1111111111111111_1111110001011111_1111001101001001"; -- -0.014160914105126583
	pesos_i(5620) := b"1111111111111111_1111111111111111_1101100101001011_1000000000000100"; -- -0.1511917105817652
	pesos_i(5621) := b"1111111111111111_1111111111111111_1101110001000011_0101100101100011"; -- -0.13959733337378763
	pesos_i(5622) := b"0000000000000000_0000000000000000_0001110111011101_1111111010001100"; -- 0.11666861449365862
	pesos_i(5623) := b"1111111111111111_1111111111111111_1111011110001001_0010011010111010"; -- -0.033063487589447264
	pesos_i(5624) := b"0000000000000000_0000000000000000_0001010011101111_0100001001100001"; -- 0.08177580715852814
	pesos_i(5625) := b"1111111111111111_1111111111111111_1110010111101001_0001101100010001"; -- -0.10191183876887404
	pesos_i(5626) := b"1111111111111111_1111111111111111_1101110001011011_0011101111000101"; -- -0.1392328875985052
	pesos_i(5627) := b"1111111111111111_1111111111111111_1110001011001011_0000010111010000"; -- -0.11408961928942572
	pesos_i(5628) := b"1111111111111111_1111111111111111_1101011101100110_0111110100100010"; -- -0.1585923949091457
	pesos_i(5629) := b"0000000000000000_0000000000000000_0001011001001010_0000000101001010"; -- 0.08706672715857947
	pesos_i(5630) := b"1111111111111111_1111111111111111_1101100011100010_0000011000001100"; -- -0.15280115316776618
	pesos_i(5631) := b"1111111111111111_1111111111111111_1111111101001110_0011000011011101"; -- -0.002713152077379365
	pesos_i(5632) := b"1111111111111111_1111111111111111_1111011110110010_1011000011010011"; -- -0.03242964604910739
	pesos_i(5633) := b"1111111111111111_1111111111111111_1111100101110111_1101011101010100"; -- -0.025515119514024798
	pesos_i(5634) := b"0000000000000000_0000000000000000_0001100010001111_1010110101111100"; -- 0.09594234733373402
	pesos_i(5635) := b"1111111111111111_1111111111111111_1111100010000001_0101011010001100"; -- -0.029276457720278672
	pesos_i(5636) := b"1111111111111111_1111111111111111_1110101100101101_1111101000111011"; -- -0.08132968966244021
	pesos_i(5637) := b"1111111111111111_1111111111111111_1111001000100111_0001000101011010"; -- -0.05409137308139478
	pesos_i(5638) := b"0000000000000000_0000000000000000_0000101010001100_0111000110101100"; -- 0.04120550589772493
	pesos_i(5639) := b"1111111111111111_1111111111111111_1111101011001010_1100000101100000"; -- -0.020343698457823262
	pesos_i(5640) := b"1111111111111111_1111111111111111_1110111010110000_1101011001000000"; -- -0.06761418281501044
	pesos_i(5641) := b"0000000000000000_0000000000000000_0000001001110000_0110101100111101"; -- 0.009527876290227921
	pesos_i(5642) := b"0000000000000000_0000000000000000_0001111010110010_1110101101101101"; -- 0.11991759689390652
	pesos_i(5643) := b"1111111111111111_1111111111111111_1111011110100000_1111011100001000"; -- -0.03270011956093629
	pesos_i(5644) := b"1111111111111111_1111111111111111_1110100110100000_1000011111110100"; -- -0.08739424040254401
	pesos_i(5645) := b"0000000000000000_0000000000000000_0010011001100111_1111010101011010"; -- 0.1500237794824288
	pesos_i(5646) := b"0000000000000000_0000000000000000_0010001101010000_0100000000010110"; -- 0.13794327300189196
	pesos_i(5647) := b"0000000000000000_0000000000000000_0010011100001011_1011111010111010"; -- 0.1525229649033828
	pesos_i(5648) := b"0000000000000000_0000000000000000_0001101010011101_0100011101100001"; -- 0.10396238429128976
	pesos_i(5649) := b"1111111111111111_1111111111111111_1111000000001111_1111110000100111"; -- -0.0622560886378903
	pesos_i(5650) := b"1111111111111111_1111111111111111_1111010010010000_0100010011010000"; -- -0.04467363275261421
	pesos_i(5651) := b"1111111111111111_1111111111111111_1110000000100001_1110101011100000"; -- -0.12448246036027134
	pesos_i(5652) := b"1111111111111111_1111111111111111_1111111111000110_1001001011100101"; -- -0.0008762541907404826
	pesos_i(5653) := b"0000000000000000_0000000000000000_0000101111100111_0101100101110111"; -- 0.04649886287951082
	pesos_i(5654) := b"0000000000000000_0000000000000000_0001011111111001_1011100000010111"; -- 0.09365416109298223
	pesos_i(5655) := b"0000000000000000_0000000000000000_0000010001100100_1010111001001001"; -- 0.017161267048319804
	pesos_i(5656) := b"1111111111111111_1111111111111111_1110000101000000_1110010111000100"; -- -0.12010349231708731
	pesos_i(5657) := b"1111111111111111_1111111111111111_1111111100000101_0110111100000111"; -- -0.00382333822584348
	pesos_i(5658) := b"0000000000000000_0000000000000000_0000110101000010_1010100011100010"; -- 0.05179839631444783
	pesos_i(5659) := b"0000000000000000_0000000000000000_0001101110000001_1110100101000100"; -- 0.10745103751964466
	pesos_i(5660) := b"1111111111111111_1111111111111111_1110100001000001_1010110011101100"; -- -0.09274787174620673
	pesos_i(5661) := b"0000000000000000_0000000000000000_0000011011100100_0011111100101101"; -- 0.026920269499808108
	pesos_i(5662) := b"1111111111111111_1111111111111111_1110111110111110_0101100011100111"; -- -0.0635017811129952
	pesos_i(5663) := b"1111111111111111_1111111111111111_1110001011011010_1001100110100010"; -- -0.11385192679670146
	pesos_i(5664) := b"1111111111111111_1111111111111111_1111111001000011_1000000100100011"; -- -0.006782463973882991
	pesos_i(5665) := b"0000000000000000_0000000000000000_0000000000011001_0100001100101011"; -- 0.0003854732161306904
	pesos_i(5666) := b"1111111111111111_1111111111111111_1111101010001110_0000101100111000"; -- -0.02127008318949898
	pesos_i(5667) := b"0000000000000000_0000000000000000_0001100000111101_0110111110101001"; -- 0.09468744148285792
	pesos_i(5668) := b"1111111111111111_1111111111111111_1110010110100111_1011111101001001"; -- -0.10290913068453231
	pesos_i(5669) := b"1111111111111111_1111111111111111_1101100101110111_0100110010010000"; -- -0.15052339052644578
	pesos_i(5670) := b"1111111111111111_1111111111111111_1111001010100000_1001110110001100"; -- -0.05223670318540517
	pesos_i(5671) := b"1111111111111111_1111111111111111_1110001110110001_1111110001001010"; -- -0.11056540685168377
	pesos_i(5672) := b"0000000000000000_0000000000000000_0010101010001100_0001110100010101"; -- 0.16620046381842665
	pesos_i(5673) := b"1111111111111111_1111111111111111_1111010111010000_1110010100111010"; -- -0.039781258927419516
	pesos_i(5674) := b"0000000000000000_0000000000000000_0000111110111101_1101001010101111"; -- 0.06149021877115958
	pesos_i(5675) := b"0000000000000000_0000000000000000_0001101110010001_0111111100010000"; -- 0.10768884794499566
	pesos_i(5676) := b"0000000000000000_0000000000000000_0001101100010111_0100100001110110"; -- 0.10582402124140752
	pesos_i(5677) := b"0000000000000000_0000000000000000_0000000000100011_0001001100011010"; -- 0.0005351961978555914
	pesos_i(5678) := b"1111111111111111_1111111111111111_1111111001111110_1100000110111111"; -- -0.005878344495609203
	pesos_i(5679) := b"0000000000000000_0000000000000000_0001110100010100_1000011101010110"; -- 0.11359449233951248
	pesos_i(5680) := b"0000000000000000_0000000000000000_0000101110010111_0010110110000110"; -- 0.04527554055365629
	pesos_i(5681) := b"0000000000000000_0000000000000000_0001101100110110_1010111100100000"; -- 0.10630316282989569
	pesos_i(5682) := b"1111111111111111_1111111111111111_1111011001011000_1001001000000110"; -- -0.037711022897809476
	pesos_i(5683) := b"0000000000000000_0000000000000000_0001111011110010_1101000110111000"; -- 0.12089262727017108
	pesos_i(5684) := b"0000000000000000_0000000000000000_0001110101010110_0100011101000001"; -- 0.11459775300629609
	pesos_i(5685) := b"0000000000000000_0000000000000000_0001011100101100_1011101101001011"; -- 0.09052630020167869
	pesos_i(5686) := b"1111111111111111_1111111111111111_1111000000001111_1111111111100001"; -- -0.06225586654608499
	pesos_i(5687) := b"1111111111111111_1111111111111111_1110111010110010_1101001001101010"; -- -0.06758389397562374
	pesos_i(5688) := b"1111111111111111_1111111111111111_1111100010110100_0000101011010001"; -- -0.028502773174902574
	pesos_i(5689) := b"0000000000000000_0000000000000000_0001000110100011_0100111101001101"; -- 0.06889815922053201
	pesos_i(5690) := b"0000000000000000_0000000000000000_0000001110101001_1011101111001010"; -- 0.014308678460021818
	pesos_i(5691) := b"0000000000000000_0000000000000000_0010010100010110_1001111100011010"; -- 0.1448764265509947
	pesos_i(5692) := b"1111111111111111_1111111111111111_1110111000011010_1010000100011111"; -- -0.06990616789904901
	pesos_i(5693) := b"1111111111111111_1111111111111111_1111011011000101_0111101001011011"; -- -0.036049225621972984
	pesos_i(5694) := b"0000000000000000_0000000000000000_0010011011011100_1110111011011010"; -- 0.15180867030434947
	pesos_i(5695) := b"1111111111111111_1111111111111111_1111100010111111_1001110010101101"; -- -0.028326232754934105
	pesos_i(5696) := b"0000000000000000_0000000000000000_0001001011000100_0011000000110100"; -- 0.07330609585081863
	pesos_i(5697) := b"0000000000000000_0000000000000000_0001101010101010_0011001100111001"; -- 0.1041595471725809
	pesos_i(5698) := b"1111111111111111_1111111111111111_1101011001110011_0011101011110001"; -- -0.16230422615725168
	pesos_i(5699) := b"1111111111111111_1111111111111111_1110111001100111_0111111110100110"; -- -0.0687332362195909
	pesos_i(5700) := b"0000000000000000_0000000000000000_0001000100110001_0011101100000000"; -- 0.06715744729255549
	pesos_i(5701) := b"0000000000000000_0000000000000000_0010010101001110_1100110000001111"; -- 0.1457335984619493
	pesos_i(5702) := b"0000000000000000_0000000000000000_0010001010110011_0101010011000011"; -- 0.13554887545820235
	pesos_i(5703) := b"0000000000000000_0000000000000000_0001010001010111_0101011111010010"; -- 0.07945774914882016
	pesos_i(5704) := b"1111111111111111_1111111111111111_1110000010001100_0100000000110110"; -- -0.12285994235195283
	pesos_i(5705) := b"1111111111111111_1111111111111111_1101011111111101_1000010111110011"; -- -0.1562877922800504
	pesos_i(5706) := b"1111111111111111_1111111111111111_1111010100111100_0001000001010011"; -- -0.04205224974006531
	pesos_i(5707) := b"0000000000000000_0000000000000000_0000011010011011_0010110110000011"; -- 0.025805324996688462
	pesos_i(5708) := b"1111111111111111_1111111111111111_1110011111110011_1110100111110010"; -- -0.09393442010139119
	pesos_i(5709) := b"0000000000000000_0000000000000000_0000001111100001_1001010000000010"; -- 0.015160799483863367
	pesos_i(5710) := b"0000000000000000_0000000000000000_0000111110101001_1100101000110001"; -- 0.061184537009584004
	pesos_i(5711) := b"0000000000000000_0000000000000000_0001000100011000_1001011011100011"; -- 0.06678145437870986
	pesos_i(5712) := b"1111111111111111_1111111111111111_1110000110000101_1110100111100100"; -- -0.11905039012027815
	pesos_i(5713) := b"0000000000000000_0000000000000000_0001110101000001_0101011111001011"; -- 0.1142783041306139
	pesos_i(5714) := b"0000000000000000_0000000000000000_0000011111010001_0101010011101111"; -- 0.03053789925543407
	pesos_i(5715) := b"0000000000000000_0000000000000000_0001011001101101_0000000010000101"; -- 0.08760073904243415
	pesos_i(5716) := b"0000000000000000_0000000000000000_0001110101000011_0000101010100001"; -- 0.11430422238974175
	pesos_i(5717) := b"0000000000000000_0000000000000000_0000100010010110_1010101101111111"; -- 0.03354904036669926
	pesos_i(5718) := b"1111111111111111_1111111111111111_1101100101110100_1010010101110010"; -- -0.15056386925143353
	pesos_i(5719) := b"0000000000000000_0000000000000000_0001100001010011_1110110001001110"; -- 0.09503056432540176
	pesos_i(5720) := b"0000000000000000_0000000000000000_0010001110010001_0011001100011000"; -- 0.1389343198250971
	pesos_i(5721) := b"0000000000000000_0000000000000000_0010001001101001_1100011011111010"; -- 0.13442653279855848
	pesos_i(5722) := b"0000000000000000_0000000000000000_0000000100101110_0111111011111010"; -- 0.004615722633102105
	pesos_i(5723) := b"1111111111111111_1111111111111111_1101110100101001_1010000010011110"; -- -0.13608356602725402
	pesos_i(5724) := b"1111111111111111_1111111111111111_1111001011000010_0010111010110111"; -- -0.051724510476763914
	pesos_i(5725) := b"1111111111111111_1111111111111111_1111100100000000_1111100101110001"; -- -0.027328882030043942
	pesos_i(5726) := b"1111111111111111_1111111111111111_1111110100000100_0111101010110111"; -- -0.011650400553525167
	pesos_i(5727) := b"0000000000000000_0000000000000000_0001110100111110_1001100011111100"; -- 0.11423641349267763
	pesos_i(5728) := b"0000000000000000_0000000000000000_0001111010001001_0100110010010110"; -- 0.11928251888911104
	pesos_i(5729) := b"1111111111111111_1111111111111111_1101110000001100_0000110001011001"; -- -0.14044115853244146
	pesos_i(5730) := b"0000000000000000_0000000000000000_0001100110010001_1011100101011101"; -- 0.09987982295617057
	pesos_i(5731) := b"0000000000000000_0000000000000000_0000101001111001_1000101011011101"; -- 0.040917090486827026
	pesos_i(5732) := b"0000000000000000_0000000000000000_0010010011010011_1011001100000001"; -- 0.1438552740271792
	pesos_i(5733) := b"1111111111111111_1111111111111111_1110000000011110_1100100110010110"; -- -0.12453022088842867
	pesos_i(5734) := b"1111111111111111_1111111111111111_1110000011010101_0011010011011111"; -- -0.12174672667812193
	pesos_i(5735) := b"0000000000000000_0000000000000000_0001011010100010_1010111000010100"; -- 0.08841979968165622
	pesos_i(5736) := b"1111111111111111_1111111111111111_1110101101111101_1010011011100000"; -- -0.080113954739148
	pesos_i(5737) := b"1111111111111111_1111111111111111_1110110000100111_0001001100110100"; -- -0.07752876257656297
	pesos_i(5738) := b"1111111111111111_1111111111111111_1110001111010011_1111111111101000"; -- -0.11004639237666919
	pesos_i(5739) := b"0000000000000000_0000000000000000_0010010111111101_1111000101100001"; -- 0.14840611088085678
	pesos_i(5740) := b"1111111111111111_1111111111111111_1111011111000111_0101011010100101"; -- -0.03211458648554142
	pesos_i(5741) := b"0000000000000000_0000000000000000_0001001111010010_1111010100010100"; -- 0.07743770345564042
	pesos_i(5742) := b"0000000000000000_0000000000000000_0001010000001000_0100000101000011"; -- 0.07825096013830346
	pesos_i(5743) := b"1111111111111111_1111111111111111_1111000001000001_1101111000110110"; -- -0.06149493394773845
	pesos_i(5744) := b"1111111111111111_1111111111111111_1101101000111011_0111100110000000"; -- -0.14752998954077462
	pesos_i(5745) := b"0000000000000000_0000000000000000_0001000000010001_0010101100101110"; -- 0.06276197320705172
	pesos_i(5746) := b"0000000000000000_0000000000000000_0000110110001110_0010100111000000"; -- 0.05295048657574728
	pesos_i(5747) := b"1111111111111111_1111111111111111_1110111100100100_0001111111110011"; -- -0.0658550292587509
	pesos_i(5748) := b"1111111111111111_1111111111111111_1111101111011101_0001010001101000"; -- -0.016157841244655833
	pesos_i(5749) := b"1111111111111111_1111111111111111_1111001001100110_0101111111000111"; -- -0.053125394747531716
	pesos_i(5750) := b"1111111111111111_1111111111111111_1110010011111111_0101101101011000"; -- -0.10547856428943873
	pesos_i(5751) := b"1111111111111111_1111111111111111_1111100000001101_0101100110110010"; -- -0.03104628953856341
	pesos_i(5752) := b"1111111111111111_1111111111111111_1110000001111110_1000111110100010"; -- -0.1230688314088382
	pesos_i(5753) := b"1111111111111111_1111111111111111_1110001010011101_1101001011101010"; -- -0.11477929861816247
	pesos_i(5754) := b"0000000000000000_0000000000000000_0001001111000000_1001111000100101"; -- 0.07715786358073737
	pesos_i(5755) := b"0000000000000000_0000000000000000_0001001000111000_0010011110000000"; -- 0.07116934653717409
	pesos_i(5756) := b"1111111111111111_1111111111111111_1101101000000000_0011011000001001"; -- -0.1484342791733257
	pesos_i(5757) := b"1111111111111111_1111111111111111_1110100000001110_0101010111011000"; -- -0.09353126036771582
	pesos_i(5758) := b"0000000000000000_0000000000000000_0000011001100110_0001110000100000"; -- 0.024995572863616488
	pesos_i(5759) := b"0000000000000000_0000000000000000_0010000010001000_1001010110010010"; -- 0.12708411028321798
	pesos_i(5760) := b"0000000000000000_0000000000000000_0000001100011000_0101001010101101"; -- 0.012089888777094854
	pesos_i(5761) := b"0000000000000000_0000000000000000_0001000011000101_0001101001101010"; -- 0.06550755573981297
	pesos_i(5762) := b"0000000000000000_0000000000000000_0010010111001100_1010000111000110"; -- 0.14765368546298346
	pesos_i(5763) := b"0000000000000000_0000000000000000_0010100100100111_0100111000110111"; -- 0.16075600469548026
	pesos_i(5764) := b"1111111111111111_1111111111111111_1111000011100111_1101100100011011"; -- -0.058962279214516466
	pesos_i(5765) := b"0000000000000000_0000000000000000_0010000100000110_0111010001011111"; -- 0.12900473900359946
	pesos_i(5766) := b"1111111111111111_1111111111111111_1111010111101100_0100100011001010"; -- -0.039363337207347006
	pesos_i(5767) := b"1111111111111111_1111111111111111_1111111110111000_1110001100110000"; -- -0.0010850913073726794
	pesos_i(5768) := b"1111111111111111_1111111111111111_1101001111101111_1011011011101100"; -- -0.17212349632746737
	pesos_i(5769) := b"1111111111111111_1111111111111111_1101110110100000_1011100001101110"; -- -0.13426635093267408
	pesos_i(5770) := b"0000000000000000_0000000000000000_0001011001101010_0101111100011100"; -- 0.08756060067490752
	pesos_i(5771) := b"0000000000000000_0000000000000000_0001111110100101_0100010101101001"; -- 0.12361558743662698
	pesos_i(5772) := b"1111111111111111_1111111111111111_1111000100110111_0110111110111110"; -- -0.05774785613748852
	pesos_i(5773) := b"0000000000000000_0000000000000000_0000111010110100_1110100111100001"; -- 0.057448022335387275
	pesos_i(5774) := b"1111111111111111_1111111111111111_1101100011110111_1100111000010000"; -- -0.1524687967873667
	pesos_i(5775) := b"0000000000000000_0000000000000000_0001101011010011_1111101010101001"; -- 0.10479704493684851
	pesos_i(5776) := b"1111111111111111_1111111111111111_1110100101001001_0100011100011011"; -- -0.08872562024036273
	pesos_i(5777) := b"0000000000000000_0000000000000000_0001110011101001_1111001001110100"; -- 0.1129447490930602
	pesos_i(5778) := b"0000000000000000_0000000000000000_0001011010101001_0111100011010011"; -- 0.0885234370283148
	pesos_i(5779) := b"1111111111111111_1111111111111111_1111000110100101_0010011010100111"; -- -0.05607374584652096
	pesos_i(5780) := b"1111111111111111_1111111111111111_1110101110101110_0010100011011010"; -- -0.07937378578699437
	pesos_i(5781) := b"0000000000000000_0000000000000000_0000010000111100_0101101010011011"; -- 0.016545927872091432
	pesos_i(5782) := b"0000000000000000_0000000000000000_0001110010101001_0100000100101010"; -- 0.11195761954521
	pesos_i(5783) := b"0000000000000000_0000000000000000_0010011000010111_0101001011111000"; -- 0.14879339736954084
	pesos_i(5784) := b"1111111111111111_1111111111111111_1110110111111110_1000101000101100"; -- -0.07033478186017278
	pesos_i(5785) := b"0000000000000000_0000000000000000_0001001010010001_1010010110001010"; -- 0.07253489134199614
	pesos_i(5786) := b"1111111111111111_1111111111111111_1111000011110010_0010101011111100"; -- -0.058804810927624455
	pesos_i(5787) := b"1111111111111111_1111111111111111_1110000101110111_1101100111101011"; -- -0.11926496517076968
	pesos_i(5788) := b"1111111111111111_1111111111111111_1110111101000101_1010000110101011"; -- -0.06534375743116048
	pesos_i(5789) := b"1111111111111111_1111111111111111_1101010000011111_0000111001011111"; -- -0.17140112095450738
	pesos_i(5790) := b"1111111111111111_1111111111111111_1110110001010000_1010101101011010"; -- -0.0768940834539354
	pesos_i(5791) := b"1111111111111111_1111111111111111_1111101100111110_1111001111100111"; -- -0.018570667300231297
	pesos_i(5792) := b"0000000000000000_0000000000000000_0000011110110101_1110110110110000"; -- 0.03011975814720297
	pesos_i(5793) := b"0000000000000000_0000000000000000_0001101101100100_0110101110101010"; -- 0.10700104609294446
	pesos_i(5794) := b"1111111111111111_1111111111111111_1110001100110110_1111010110000011"; -- -0.11244264175917949
	pesos_i(5795) := b"1111111111111111_1111111111111111_1101011000010000_0010111100010110"; -- -0.1638155527719158
	pesos_i(5796) := b"0000000000000000_0000000000000000_0000010101011111_0010100011111100"; -- 0.020983277728771576
	pesos_i(5797) := b"0000000000000000_0000000000000000_0000100110101101_1100111001110101"; -- 0.037808326413958974
	pesos_i(5798) := b"1111111111111111_1111111111111111_1111110011110100_0001011011101010"; -- -0.011900489699552114
	pesos_i(5799) := b"0000000000000000_0000000000000000_0000111101010011_1110010010010010"; -- 0.059873853301005836
	pesos_i(5800) := b"0000000000000000_0000000000000000_0001010110100100_1100010111001000"; -- 0.08454548016826705
	pesos_i(5801) := b"0000000000000000_0000000000000000_0001001011101110_1111111111000010"; -- 0.07395933625521543
	pesos_i(5802) := b"1111111111111111_1111111111111111_1111011111100101_0001011100111010"; -- -0.03166060284515098
	pesos_i(5803) := b"0000000000000000_0000000000000000_0001001001001000_1110001001011001"; -- 0.0714246242228899
	pesos_i(5804) := b"0000000000000000_0000000000000000_0001000011101000_0110111101010100"; -- 0.06604667468483767
	pesos_i(5805) := b"1111111111111111_1111111111111111_1101110110011001_1111001011100011"; -- -0.134369678018483
	pesos_i(5806) := b"0000000000000000_0000000000000000_0010011101001100_0010100011110110"; -- 0.15350585943911532
	pesos_i(5807) := b"0000000000000000_0000000000000000_0000001100111110_1110000010101101"; -- 0.012678186593998499
	pesos_i(5808) := b"1111111111111111_1111111111111111_1101101000101110_1011010100100111"; -- -0.14772479807233752
	pesos_i(5809) := b"1111111111111111_1111111111111111_1101110111001110_0011101100100010"; -- -0.1335719149375707
	pesos_i(5810) := b"0000000000000000_0000000000000000_0010010010111100_1001100011100000"; -- 0.1435027643269885
	pesos_i(5811) := b"0000000000000000_0000000000000000_0010101011101101_1111001100100110"; -- 0.16769332585921043
	pesos_i(5812) := b"0000000000000000_0000000000000000_0000011000001000_1111010001111011"; -- 0.02357414237379492
	pesos_i(5813) := b"0000000000000000_0000000000000000_0010011010010110_0110111000110001"; -- 0.15073288637846086
	pesos_i(5814) := b"1111111111111111_1111111111111111_1110110011000100_1011110110000111"; -- -0.07512298066928852
	pesos_i(5815) := b"0000000000000000_0000000000000000_0000111000011011_0000011011000001"; -- 0.055099889753487355
	pesos_i(5816) := b"0000000000000000_0000000000000000_0001000001110000_1010001110101100"; -- 0.06421873999865915
	pesos_i(5817) := b"1111111111111111_1111111111111111_1111001000110000_0111001001110000"; -- -0.053948257154257745
	pesos_i(5818) := b"1111111111111111_1111111111111111_1111101010011000_1111001010011010"; -- -0.0211037038204572
	pesos_i(5819) := b"1111111111111111_1111111111111111_1101111000110100_0010010111111011"; -- -0.13201677919133986
	pesos_i(5820) := b"1111111111111111_1111111111111111_1111101011010000_1010011010000100"; -- -0.020253746869452815
	pesos_i(5821) := b"1111111111111111_1111111111111111_1111101110001101_1011000100100011"; -- -0.017369202680780915
	pesos_i(5822) := b"1111111111111111_1111111111111111_1111001101001110_1111011110111110"; -- -0.04957629790504837
	pesos_i(5823) := b"0000000000000000_0000000000000000_0001011011111101_1011101100111111"; -- 0.08980913427074957
	pesos_i(5824) := b"1111111111111111_1111111111111111_1110011110100011_1110100011100111"; -- -0.09515518542176965
	pesos_i(5825) := b"0000000000000000_0000000000000000_0001110110110011_1011110110100000"; -- 0.11602387568306516
	pesos_i(5826) := b"0000000000000000_0000000000000000_0000100010100011_0101011100101000"; -- 0.03374237752411195
	pesos_i(5827) := b"0000000000000000_0000000000000000_0000101110110110_0010101010110110"; -- 0.04574839531618019
	pesos_i(5828) := b"1111111111111111_1111111111111111_1101110110101110_0100101111001010"; -- -0.1340592032779819
	pesos_i(5829) := b"1111111111111111_1111111111111111_1101111101000110_1011010100111111"; -- -0.12782733169308907
	pesos_i(5830) := b"1111111111111111_1111111111111111_1101011010110000_0000011001010101"; -- -0.16137657566728617
	pesos_i(5831) := b"0000000000000000_0000000000000000_0001011010011110_0011100110000110"; -- 0.08835181739474253
	pesos_i(5832) := b"1111111111111111_1111111111111111_1110100000110111_0011111101011011"; -- -0.0929069902206394
	pesos_i(5833) := b"1111111111111111_1111111111111111_1110111100010101_1000011111111010"; -- -0.06607771056854739
	pesos_i(5834) := b"1111111111111111_1111111111111111_1110101001010001_1100101110110011"; -- -0.0846893967618187
	pesos_i(5835) := b"1111111111111111_1111111111111111_1110001010110011_1011110001111011"; -- -0.11444494252539601
	pesos_i(5836) := b"0000000000000000_0000000000000000_0010111100010100_0010111000100011"; -- 0.1839016757039866
	pesos_i(5837) := b"1111111111111111_1111111111111111_1111111000100011_1110100110100001"; -- -0.007264516937704028
	pesos_i(5838) := b"1111111111111111_1111111111111111_1110011111101010_1110100110110101"; -- -0.09407176337374781
	pesos_i(5839) := b"0000000000000000_0000000000000000_0010100110000110_1111011000011000"; -- 0.16221559606301852
	pesos_i(5840) := b"0000000000000000_0000000000000000_0010000101000001_0101010001010000"; -- 0.12990309677143788
	pesos_i(5841) := b"0000000000000000_0000000000000000_0010101010111100_1000111101001010"; -- 0.16693969303238743
	pesos_i(5842) := b"1111111111111111_1111111111111111_1110101001101000_1111011110001011"; -- -0.08433583127463816
	pesos_i(5843) := b"0000000000000000_0000000000000000_0000100101000011_0111010100001110"; -- 0.03618556575704429
	pesos_i(5844) := b"1111111111111111_1111111111111111_1111100000011011_1111001011010111"; -- -0.03082353823694533
	pesos_i(5845) := b"1111111111111111_1111111111111111_1111111011000111_0010001101101100"; -- -0.004773889600082521
	pesos_i(5846) := b"0000000000000000_0000000000000000_0001011111110100_0101000001101111"; -- 0.0935716887854344
	pesos_i(5847) := b"0000000000000000_0000000000000000_0000100101001011_1100010010010111"; -- 0.03631237678215726
	pesos_i(5848) := b"0000000000000000_0000000000000000_0000111100100011_0111010000111011"; -- 0.05913473538396671
	pesos_i(5849) := b"0000000000000000_0000000000000000_0000010101100111_0000010010111010"; -- 0.021103187107628762
	pesos_i(5850) := b"0000000000000000_0000000000000000_0001001010011011_1000110101001001"; -- 0.07268603353957417
	pesos_i(5851) := b"1111111111111111_1111111111111111_1111111101100010_1001110100101010"; -- -0.0024015209396175026
	pesos_i(5852) := b"1111111111111111_1111111111111111_1101000001100101_1111110001000000"; -- -0.1859438271090963
	pesos_i(5853) := b"0000000000000000_0000000000000000_0001010000010010_1001010101101110"; -- 0.07840856491101103
	pesos_i(5854) := b"0000000000000000_0000000000000000_0000011011000001_0011011000110010"; -- 0.02638567657048816
	pesos_i(5855) := b"1111111111111111_1111111111111111_1110111010100101_1110000001101100"; -- -0.06778142326975514
	pesos_i(5856) := b"0000000000000000_0000000000000000_0010110010100111_1000100010000101"; -- 0.17443135501979376
	pesos_i(5857) := b"0000000000000000_0000000000000000_0010101011001101_0000111010000101"; -- 0.1671914170738037
	pesos_i(5858) := b"0000000000000000_0000000000000000_0001101100001110_1111000101110011"; -- 0.1056967644614513
	pesos_i(5859) := b"0000000000000000_0000000000000000_0001001010111111_0001100100010001"; -- 0.07322842283478531
	pesos_i(5860) := b"1111111111111111_1111111111111111_1110101110001001_0000000100010110"; -- -0.07994073118496307
	pesos_i(5861) := b"0000000000000000_0000000000000000_0010111001110001_1110100111010011"; -- 0.18142568013457688
	pesos_i(5862) := b"0000000000000000_0000000000000000_0001111011010101_0010001011100001"; -- 0.12043970092613909
	pesos_i(5863) := b"0000000000000000_0000000000000000_0000010011111111_0000110110111011"; -- 0.019516809601533347
	pesos_i(5864) := b"0000000000000000_0000000000000000_0010011111110111_0110001111101100"; -- 0.15611862669817486
	pesos_i(5865) := b"0000000000000000_0000000000000000_0001011011011101_0010101000010010"; -- 0.08931219992321965
	pesos_i(5866) := b"1111111111111111_1111111111111111_1111000111101101_0000110000011011"; -- -0.05497669544310625
	pesos_i(5867) := b"0000000000000000_0000000000000000_0000011001011101_1111000011011001"; -- 0.024870922926077222
	pesos_i(5868) := b"0000000000000000_0000000000000000_0000101111011100_1000001000100101"; -- 0.046333440791464287
	pesos_i(5869) := b"0000000000000000_0000000000000000_0000111101000000_0110011111000101"; -- 0.05957649760333472
	pesos_i(5870) := b"0000000000000000_0000000000000000_0000011111000011_0010111000001001"; -- 0.03032195767386234
	pesos_i(5871) := b"0000000000000000_0000000000000000_0011010010101010_0000001001010101"; -- 0.2057191331258061
	pesos_i(5872) := b"0000000000000000_0000000000000000_0001111100101111_0000110010011001"; -- 0.12181166398666007
	pesos_i(5873) := b"1111111111111111_1111111111111111_1111100100110011_0011011101010011"; -- -0.026562254155543204
	pesos_i(5874) := b"1111111111111111_1111111111111111_1110001100100011_0111000011010010"; -- -0.11274046788194513
	pesos_i(5875) := b"1111111111111111_1111111111111111_1111111100101100_0001010111001010"; -- -0.0032335645860942833
	pesos_i(5876) := b"1111111111111111_1111111111111111_1110110110111001_0000110000001011"; -- -0.07139515624048941
	pesos_i(5877) := b"0000000000000000_0000000000000000_0000001110011010_0010101001001110"; -- 0.014071124982920099
	pesos_i(5878) := b"1111111111111111_1111111111111111_1110010000101001_1101000100010100"; -- -0.1087369276613489
	pesos_i(5879) := b"0000000000000000_0000000000000000_0010110111010010_1011101111010101"; -- 0.17899679132872004
	pesos_i(5880) := b"1111111111111111_1111111111111111_1101101100000101_1010100001100000"; -- -0.14444492012203008
	pesos_i(5881) := b"1111111111111111_1111111111111111_1111010011001111_1010001111100111"; -- -0.04370666134125518
	pesos_i(5882) := b"0000000000000000_0000000000000000_0000111001101100_1101011001110000"; -- 0.05634823073863213
	pesos_i(5883) := b"0000000000000000_0000000000000000_0001011010001001_0000111110110100"; -- 0.0880288901737334
	pesos_i(5884) := b"0000000000000000_0000000000000000_0000010001011010_1110111000111100"; -- 0.017012490992042367
	pesos_i(5885) := b"1111111111111111_1111111111111111_1110001001010110_1001111010110101"; -- -0.11586578446592981
	pesos_i(5886) := b"1111111111111111_1111111111111111_1101011111010110_1101101001111010"; -- -0.15687784695720966
	pesos_i(5887) := b"1111111111111111_1111111111111111_1101101000111010_0001110001010000"; -- -0.14755080269756182
	pesos_i(5888) := b"0000000000000000_0000000000000000_0000001100110010_1101110110110010"; -- 0.012494903413970526
	pesos_i(5889) := b"0000000000000000_0000000000000000_0001101110100110_0000101001111011"; -- 0.10800233360320993
	pesos_i(5890) := b"1111111111111111_1111111111111111_1110101101001110_0100101110110001"; -- -0.08083655280757947
	pesos_i(5891) := b"0000000000000000_0000000000000000_0000110101010010_0000100010000010"; -- 0.052032977696641974
	pesos_i(5892) := b"1111111111111111_1111111111111111_1111110011110000_0011111010110101"; -- -0.011959153110116411
	pesos_i(5893) := b"1111111111111111_1111111111111111_1101110100110000_0000010010001110"; -- -0.13598605672868705
	pesos_i(5894) := b"0000000000000000_0000000000000000_0001100000001001_1000001101011000"; -- 0.09389515772853987
	pesos_i(5895) := b"1111111111111111_1111111111111111_1101111010011010_0011101010011000"; -- -0.1304591541012383
	pesos_i(5896) := b"0000000000000000_0000000000000000_0000011110111100_0111000010011001"; -- 0.030219113570869857
	pesos_i(5897) := b"0000000000000000_0000000000000000_0001111101010110_0011111000011010"; -- 0.12240970735750631
	pesos_i(5898) := b"1111111111111111_1111111111111111_1101010110001000_1010110001101011"; -- -0.16588327768342748
	pesos_i(5899) := b"1111111111111111_1111111111111111_1111101011011011_1000110011010101"; -- -0.020087430884820217
	pesos_i(5900) := b"0000000000000000_0000000000000000_0000000110100011_1011000111000111"; -- 0.006404028913254279
	pesos_i(5901) := b"0000000000000000_0000000000000000_0010011010001011_0010111001011111"; -- 0.15056123572681332
	pesos_i(5902) := b"0000000000000000_0000000000000000_0010100001101100_1011011001100000"; -- 0.15790881964956166
	pesos_i(5903) := b"0000000000000000_0000000000000000_0010010100000100_1110001101101001"; -- 0.14460583981348937
	pesos_i(5904) := b"1111111111111111_1111111111111111_1110110000100001_0001100010010000"; -- -0.07761999599115249
	pesos_i(5905) := b"1111111111111111_1111111111111111_1110010010110111_1111001011000010"; -- -0.1065681720805166
	pesos_i(5906) := b"0000000000000000_0000000000000000_0000100110000110_0000100010001110"; -- 0.03720143772542753
	pesos_i(5907) := b"0000000000000000_0000000000000000_0000010110001100_1111101011011101"; -- 0.02168243319519141
	pesos_i(5908) := b"1111111111111111_1111111111111111_1110010111001111_0011110101000100"; -- -0.10230652899866376
	pesos_i(5909) := b"1111111111111111_1111111111111111_1101011100010010_0001101001100010"; -- -0.15988001924457876
	pesos_i(5910) := b"1111111111111111_1111111111111111_1110010100111010_0101010110010010"; -- -0.10457863988541728
	pesos_i(5911) := b"1111111111111111_1111111111111111_1111010000001001_1000110010001000"; -- -0.046729294573828066
	pesos_i(5912) := b"0000000000000000_0000000000000000_0000100011100000_0010100010010101"; -- 0.03467038762429743
	pesos_i(5913) := b"0000000000000000_0000000000000000_0000010000100111_0001101110001110"; -- 0.01622173513857524
	pesos_i(5914) := b"1111111111111111_1111111111111111_1101011111111111_1000101100011001"; -- -0.1562569678803622
	pesos_i(5915) := b"1111111111111111_1111111111111111_1101010010111100_1111000101101100"; -- -0.16899195785993576
	pesos_i(5916) := b"1111111111111111_1111111111111111_1110111111011000_0100100001111111"; -- -0.0631060305683049
	pesos_i(5917) := b"1111111111111111_1111111111111111_1111111110100001_0001001101101101"; -- -0.0014484270810693953
	pesos_i(5918) := b"1111111111111111_1111111111111111_1110010001111011_1001111010111011"; -- -0.1074887079854306
	pesos_i(5919) := b"0000000000000000_0000000000000000_0000000000010101_0000110110001101"; -- 0.0003212421664343934
	pesos_i(5920) := b"1111111111111111_1111111111111111_1110101101001000_1111000111010100"; -- -0.08091820305397755
	pesos_i(5921) := b"0000000000000000_0000000000000000_0001000110110001_0001101110100011"; -- 0.06910870293530536
	pesos_i(5922) := b"1111111111111111_1111111111111111_1101010001001110_0111000000101110"; -- -0.17067812792646425
	pesos_i(5923) := b"1111111111111111_1111111111111111_1101110001000111_0101000000001111"; -- -0.13953685422089274
	pesos_i(5924) := b"0000000000000000_0000000000000000_0001001000110100_0110100100111100"; -- 0.0711122295318002
	pesos_i(5925) := b"1111111111111111_1111111111111111_1111110010101111_0011001001111001"; -- -0.01295170342656442
	pesos_i(5926) := b"1111111111111111_1111111111111111_1101110000111010_0011110101110110"; -- -0.13973632690882185
	pesos_i(5927) := b"0000000000000000_0000000000000000_0001000011111101_1000100000010110"; -- 0.06636858488196248
	pesos_i(5928) := b"1111111111111111_1111111111111111_1110011011100011_1011110100000010"; -- -0.09808748906241399
	pesos_i(5929) := b"0000000000000000_0000000000000000_0010011101011010_0110101100110000"; -- 0.15372342996329721
	pesos_i(5930) := b"1111111111111111_1111111111111111_1111011010011000_1110101111000101"; -- -0.03672911121773073
	pesos_i(5931) := b"1111111111111111_1111111111111111_1111111100110000_0001011110000010"; -- -0.003172426897433604
	pesos_i(5932) := b"0000000000000000_0000000000000000_0001010100001000_0010101001111110"; -- 0.08215585306049161
	pesos_i(5933) := b"1111111111111111_1111111111111111_1101101100000000_1100100111011010"; -- -0.1445192186937091
	pesos_i(5934) := b"0000000000000000_0000000000000000_0000001011000000_1101010110110011"; -- 0.010754924906474799
	pesos_i(5935) := b"0000000000000000_0000000000000000_0001111011011101_0101001011000100"; -- 0.12056462571227711
	pesos_i(5936) := b"1111111111111111_1111111111111111_1111001010101100_1101000001101101"; -- -0.05205056511399017
	pesos_i(5937) := b"1111111111111111_1111111111111111_1110000111111001_1100010110111010"; -- -0.11728252603881763
	pesos_i(5938) := b"1111111111111111_1111111111111111_1110011101001111_1010010100111011"; -- -0.09644095719721128
	pesos_i(5939) := b"1111111111111111_1111111111111111_1110110100111000_1101101010000010"; -- -0.07335123384070888
	pesos_i(5940) := b"0000000000000000_0000000000000000_0001000110010101_1001000100110101"; -- 0.068688464572574
	pesos_i(5941) := b"1111111111111111_1111111111111111_1101101111000110_1110101100100010"; -- -0.14149599477620933
	pesos_i(5942) := b"1111111111111111_1111111111111111_1110011111000000_0010010010001001"; -- -0.09472438472504045
	pesos_i(5943) := b"0000000000000000_0000000000000000_0001010000000100_0111011100011111"; -- 0.07819313531559509
	pesos_i(5944) := b"0000000000000000_0000000000000000_0001100101100100_1101001110011001"; -- 0.09919474115550406
	pesos_i(5945) := b"1111111111111111_1111111111111111_1110000000101010_1101101010010001"; -- -0.12434610334447234
	pesos_i(5946) := b"1111111111111111_1111111111111111_1111010000111010_0101011111001001"; -- -0.045984757898890526
	pesos_i(5947) := b"1111111111111111_1111111111111111_1101010000000111_1000010001110011"; -- -0.17176029390189115
	pesos_i(5948) := b"0000000000000000_0000000000000000_0000000000010100_1110010100110100"; -- 0.0003188374263029848
	pesos_i(5949) := b"0000000000000000_0000000000000000_0010010110000101_0100001000000010"; -- 0.1465646033837495
	pesos_i(5950) := b"0000000000000000_0000000000000000_0001111101100101_1000000010101011"; -- 0.12264255690857395
	pesos_i(5951) := b"1111111111111111_1111111111111111_1101101101010000_1111100000000011"; -- -0.14329576417159476
	pesos_i(5952) := b"1111111111111111_1111111111111111_1101100011111111_0001101011100111"; -- -0.15235740530161535
	pesos_i(5953) := b"0000000000000000_0000000000000000_0000100011010011_0001111010010001"; -- 0.03447142650068126
	pesos_i(5954) := b"1111111111111111_1111111111111111_1111000101001001_0001000011011011"; -- -0.05747885362080043
	pesos_i(5955) := b"0000000000000000_0000000000000000_0000101101100110_1100111010000010"; -- 0.044537455392020524
	pesos_i(5956) := b"0000000000000000_0000000000000000_0001011001000111_1110111110001001"; -- 0.08703515153151202
	pesos_i(5957) := b"1111111111111111_1111111111111111_1110000011110111_1001110110001000"; -- -0.12122168947394217
	pesos_i(5958) := b"1111111111111111_1111111111111111_1111000001110100_1000000001110101"; -- -0.06072232383278469
	pesos_i(5959) := b"1111111111111111_1111111111111111_1111101101011101_1010000100111011"; -- -0.018102572426938024
	pesos_i(5960) := b"1111111111111111_1111111111111111_1100000001100011_1110011001100010"; -- -0.24847564788436124
	pesos_i(5961) := b"1111111111111111_1111111111111111_1101111110101001_1101100111001011"; -- -0.1263145330734745
	pesos_i(5962) := b"0000000000000000_0000000000000000_0001001000111101_0111000100111001"; -- 0.07125003475110558
	pesos_i(5963) := b"0000000000000000_0000000000000000_0010010111101110_1011100011001010"; -- 0.1481738561540176
	pesos_i(5964) := b"0000000000000000_0000000000000000_0010000100111001_1101110110101001"; -- 0.12978921283860276
	pesos_i(5965) := b"1111111111111111_1111111111111111_1110011101010010_1001000011100101"; -- -0.09639639282354943
	pesos_i(5966) := b"0000000000000000_0000000000000000_0001111100001101_0000010001010001"; -- 0.1212923715559717
	pesos_i(5967) := b"0000000000000000_0000000000000000_0001100000110111_0011010010011100"; -- 0.09459236909517568
	pesos_i(5968) := b"1111111111111111_1111111111111111_1101111011001100_0010011111000110"; -- -0.1296973363363597
	pesos_i(5969) := b"1111111111111111_1111111111111111_1111111100010000_0000011110011101"; -- -0.003661655525673041
	pesos_i(5970) := b"0000000000000000_0000000000000000_0001101100111111_1110011101100111"; -- 0.10644384646536771
	pesos_i(5971) := b"1111111111111111_1111111111111111_1110000010101001_0100100111001001"; -- -0.12241686673226196
	pesos_i(5972) := b"1111111111111111_1111111111111111_1101001000100111_1001011011110100"; -- -0.17908340980605558
	pesos_i(5973) := b"0000000000000000_0000000000000000_0001011010110111_1110111011000110"; -- 0.08874409033896709
	pesos_i(5974) := b"0000000000000000_0000000000000000_0010011010111101_0100010000001100"; -- 0.15132546695349594
	pesos_i(5975) := b"1111111111111111_1111111111111111_1101001101001001_0000010101100001"; -- -0.17466703789044638
	pesos_i(5976) := b"1111111111111111_1111111111111111_1111110001001001_0100000110101100"; -- -0.01450719395799233
	pesos_i(5977) := b"0000000000000000_0000000000000000_0000111001110000_0101101000101101"; -- 0.056401859174799174
	pesos_i(5978) := b"1111111111111111_1111111111111111_1110001110011110_0001111110001110"; -- -0.11086848048362571
	pesos_i(5979) := b"0000000000000000_0000000000000000_0001011001011001_0010101000100110"; -- 0.08729804441584484
	pesos_i(5980) := b"0000000000000000_0000000000000000_0000001011111100_0101111001001101"; -- 0.011663335495923943
	pesos_i(5981) := b"0000000000000000_0000000000000000_0010111100100101_0111001110101110"; -- 0.18416522022048362
	pesos_i(5982) := b"1111111111111111_1111111111111111_1101011110100100_0100011110011110"; -- -0.15764953989350283
	pesos_i(5983) := b"0000000000000000_0000000000000000_0000011010101000_0010101001001101"; -- 0.026003497769587464
	pesos_i(5984) := b"1111111111111111_1111111111111111_1101011010011011_1110010010000011"; -- -0.16168376735618714
	pesos_i(5985) := b"1111111111111111_1111111111111111_1101111011101001_1111000010000110"; -- -0.12924286588347514
	pesos_i(5986) := b"1111111111111111_1111111111111111_1111010010010110_0110100101110011"; -- -0.044579896327330955
	pesos_i(5987) := b"1111111111111111_1111111111111111_1111010010010010_1000100101111001"; -- -0.04463902281346436
	pesos_i(5988) := b"1111111111111111_1111111111111111_1111011111100001_1001001110011001"; -- -0.03171422507024262
	pesos_i(5989) := b"0000000000000000_0000000000000000_0001000101110100_0010001111011001"; -- 0.0681784061686881
	pesos_i(5990) := b"1111111111111111_1111111111111111_1111011010101110_0101110101011101"; -- -0.036401905811407294
	pesos_i(5991) := b"1111111111111111_1111111111111111_1101011111000001_1110110110010100"; -- -0.15719714298996512
	pesos_i(5992) := b"0000000000000000_0000000000000000_0001111001111101_0010111001100011"; -- 0.11909761353004636
	pesos_i(5993) := b"1111111111111111_1111111111111111_1111000010001001_0011001001011011"; -- -0.0604065445905922
	pesos_i(5994) := b"0000000000000000_0000000000000000_0001100000011101_0000110100111010"; -- 0.09419329321073144
	pesos_i(5995) := b"1111111111111111_1111111111111111_1101100111000001_1000100101101111"; -- -0.14939061211947482
	pesos_i(5996) := b"1111111111111111_1111111111111111_1111001010110011_1110011111101110"; -- -0.051942352730126366
	pesos_i(5997) := b"1111111111111111_1111111111111111_1111111000000101_1011100101001110"; -- -0.007725161122909311
	pesos_i(5998) := b"1111111111111111_1111111111111111_1110100101101001_1001100010100111"; -- -0.08823247836403746
	pesos_i(5999) := b"0000000000000000_0000000000000000_0010001100000110_0100001101010101"; -- 0.13681431609071792
	pesos_i(6000) := b"1111111111111111_1111111111111111_1111101011101100_0110100010110000"; -- -0.019830185885973545
	pesos_i(6001) := b"1111111111111111_1111111111111111_1111011110111101_1001111101110001"; -- -0.032262835341764294
	pesos_i(6002) := b"1111111111111111_1111111111111111_1101101110110010_1101100100110110"; -- -0.1418022388451401
	pesos_i(6003) := b"0000000000000000_0000000000000000_0000101101100010_1010001101011001"; -- 0.0444738475841143
	pesos_i(6004) := b"0000000000000000_0000000000000000_0000110001010111_1001001001010100"; -- 0.04821123652774348
	pesos_i(6005) := b"1111111111111111_1111111111111111_1111010010110110_1100001000100100"; -- -0.04408632859789073
	pesos_i(6006) := b"0000000000000000_0000000000000000_0000000110111011_1001011101111110"; -- 0.00676867324247877
	pesos_i(6007) := b"1111111111111111_1111111111111111_1110000111010001_0101011110011001"; -- -0.11789944196204151
	pesos_i(6008) := b"0000000000000000_0000000000000000_0010101000111111_1001101010001010"; -- 0.16503301492692848
	pesos_i(6009) := b"1111111111111111_1111111111111111_1110110101110010_1111010000011001"; -- -0.07246469879173265
	pesos_i(6010) := b"0000000000000000_0000000000000000_0001111111001100_1010100111011010"; -- 0.12421666700440809
	pesos_i(6011) := b"1111111111111111_1111111111111111_1101111110010111_1110011000010111"; -- -0.12658845847507144
	pesos_i(6012) := b"1111111111111111_1111111111111111_1101110100101111_1000000101101010"; -- -0.13599387321645398
	pesos_i(6013) := b"0000000000000000_0000000000000000_0000101100111100_0110110110110011"; -- 0.04389081604213929
	pesos_i(6014) := b"0000000000000000_0000000000000000_0001100111010101_0000101100001000"; -- 0.10090702956311604
	pesos_i(6015) := b"1111111111111111_1111111111111111_1110101100110011_1101110000001010"; -- -0.08123993636488874
	pesos_i(6016) := b"1111111111111111_1111111111111111_1110000101100000_0011110110001011"; -- -0.11962523802869347
	pesos_i(6017) := b"1111111111111111_1111111111111111_1111100111011001_0110010110100100"; -- -0.024026534475333424
	pesos_i(6018) := b"0000000000000000_0000000000000000_0000101101110011_1110101011001110"; -- 0.04473750627021783
	pesos_i(6019) := b"1111111111111111_1111111111111111_1111000100010100_0111011101010000"; -- -0.058281462660719825
	pesos_i(6020) := b"1111111111111111_1111111111111111_1111011100110001_0010001101110010"; -- -0.03440645673528983
	pesos_i(6021) := b"1111111111111111_1111111111111111_1100111100111111_0011000001011100"; -- -0.19044206388166812
	pesos_i(6022) := b"0000000000000000_0000000000000000_0000001010110100_0111011011010101"; -- 0.010566164955638653
	pesos_i(6023) := b"0000000000000000_0000000000000000_0001110001000000_1000101001111110"; -- 0.1103598173526288
	pesos_i(6024) := b"0000000000000000_0000000000000000_0000100110111001_1011110010001010"; -- 0.03799036387078166
	pesos_i(6025) := b"1111111111111111_1111111111111111_1110011001101001_1111011100101001"; -- -0.09994559532533255
	pesos_i(6026) := b"0000000000000000_0000000000000000_0001010111000111_0101010000100000"; -- 0.08507276326699352
	pesos_i(6027) := b"1111111111111111_1111111111111111_1110100111011000_1000101000101100"; -- -0.0865396158023464
	pesos_i(6028) := b"0000000000000000_0000000000000000_0000010011101111_0110000101111110"; -- 0.019277661521927166
	pesos_i(6029) := b"0000000000000000_0000000000000000_0010101000000100_0001011000100011"; -- 0.16412485449224423
	pesos_i(6030) := b"0000000000000000_0000000000000000_0001001010000111_0011000010010110"; -- 0.07237533255892417
	pesos_i(6031) := b"0000000000000000_0000000000000000_0010011110010001_1111101000001000"; -- 0.15457117737037782
	pesos_i(6032) := b"0000000000000000_0000000000000000_0001100000100011_0001100001000000"; -- 0.09428550299944874
	pesos_i(6033) := b"1111111111111111_1111111111111111_1110101101100010_0100000000111100"; -- -0.08053205993247184
	pesos_i(6034) := b"1111111111111111_1111111111111111_1111110100111000_1010001111011110"; -- -0.010854490609231743
	pesos_i(6035) := b"0000000000000000_0000000000000000_0000001101110000_1001100010100111"; -- 0.013436833087432265
	pesos_i(6036) := b"0000000000000000_0000000000000000_0000101101110000_1111101101111101"; -- 0.04469272426784462
	pesos_i(6037) := b"1111111111111111_1111111111111111_1101110011111101_0101111111101111"; -- -0.1367588081886365
	pesos_i(6038) := b"0000000000000000_0000000000000000_0000100100101110_0001001011111011"; -- 0.03585928551349761
	pesos_i(6039) := b"1111111111111111_1111111111111111_1101011110110110_1101011011101000"; -- -0.15736634108272068
	pesos_i(6040) := b"0000000000000000_0000000000000000_0000001010001111_0000111010110000"; -- 0.009995382251905726
	pesos_i(6041) := b"1111111111111111_1111111111111111_1110000111011000_1101000101001110"; -- -0.11778537598266685
	pesos_i(6042) := b"0000000000000000_0000000000000000_0001001001010101_0000101101000001"; -- 0.0716101678010545
	pesos_i(6043) := b"1111111111111111_1111111111111111_1111110110101011_0000011100110001"; -- -0.009109068436369355
	pesos_i(6044) := b"1111111111111111_1111111111111111_1111001000001101_0110100101011011"; -- -0.054482856136800255
	pesos_i(6045) := b"0000000000000000_0000000000000000_0000111111001010_1101011000000000"; -- 0.06168878088152279
	pesos_i(6046) := b"0000000000000000_0000000000000000_0000111101001010_1000000101111110"; -- 0.05973061871395378
	pesos_i(6047) := b"1111111111111111_1111111111111111_1110001001010000_1000000111011011"; -- -0.11595905691225905
	pesos_i(6048) := b"1111111111111111_1111111111111111_1111010001101101_1110001110111111"; -- -0.04519821715871997
	pesos_i(6049) := b"1111111111111111_1111111111111111_1111000000001110_1000100001101011"; -- -0.06227824590401752
	pesos_i(6050) := b"1111111111111111_1111111111111111_1110000110011101_0001101110100101"; -- -0.11869647231101611
	pesos_i(6051) := b"0000000000000000_0000000000000000_0001100000000111_1010000101101110"; -- 0.0938664333691717
	pesos_i(6052) := b"1111111111111111_1111111111111111_1101100011111111_1110010110111000"; -- -0.15234531649498895
	pesos_i(6053) := b"0000000000000000_0000000000000000_0000101111001100_0100000011011111"; -- 0.04608540955286364
	pesos_i(6054) := b"0000000000000000_0000000000000000_0001000111010100_0001001101001000"; -- 0.06964226260873574
	pesos_i(6055) := b"1111111111111111_1111111111111111_1111000100110110_0110100011000001"; -- -0.057763531526290865
	pesos_i(6056) := b"0000000000000000_0000000000000000_0000011110100000_1111101100000110"; -- 0.02980011848101899
	pesos_i(6057) := b"0000000000000000_0000000000000000_0000000101111011_0111011001101011"; -- 0.005790139210106026
	pesos_i(6058) := b"1111111111111111_1111111111111111_1101010011110010_0101110110000010"; -- -0.16817679955674067
	pesos_i(6059) := b"0000000000000000_0000000000000000_0001010100110100_1011000000000101"; -- 0.08283519864524495
	pesos_i(6060) := b"1111111111111111_1111111111111111_1111000011110010_0101010010001011"; -- -0.05880233394323801
	pesos_i(6061) := b"1111111111111111_1111111111111111_1101000111010110_0110000000110010"; -- -0.18032263546066357
	pesos_i(6062) := b"0000000000000000_0000000000000000_0000100111100001_1110010010001011"; -- 0.03860309980147915
	pesos_i(6063) := b"1111111111111111_1111111111111111_1101111110001000_1111010010010101"; -- -0.12681647636900187
	pesos_i(6064) := b"1111111111111111_1111111111111111_1101001101011001_1100110001010000"; -- -0.17441103991027068
	pesos_i(6065) := b"0000000000000000_0000000000000000_0010010100011101_0111000101000011"; -- 0.14498050579010754
	pesos_i(6066) := b"0000000000000000_0000000000000000_0000111011111111_1011011110011111"; -- 0.058589435914632705
	pesos_i(6067) := b"0000000000000000_0000000000000000_0000011000011011_1001110010001000"; -- 0.023858817370382975
	pesos_i(6068) := b"1111111111111111_1111111111111111_1111110001000100_0001111010011110"; -- -0.014585577489577499
	pesos_i(6069) := b"0000000000000000_0000000000000000_0000101001100101_1111010010101101"; -- 0.04061822142162243
	pesos_i(6070) := b"0000000000000000_0000000000000000_0001110101010111_0111100010111100"; -- 0.11461596101871241
	pesos_i(6071) := b"0000000000000000_0000000000000000_0010011110101010_1101011110001111"; -- 0.15495059252266707
	pesos_i(6072) := b"1111111111111111_1111111111111111_1110111110011111_1101100110001110"; -- -0.06396713517374822
	pesos_i(6073) := b"1111111111111111_1111111111111111_1111110111010100_1001011110100111"; -- -0.008474847527232633
	pesos_i(6074) := b"0000000000000000_0000000000000000_0000101100100101_0100001101100100"; -- 0.04353734210153342
	pesos_i(6075) := b"0000000000000000_0000000000000000_0010001110000010_0111100010000101"; -- 0.13870957599032804
	pesos_i(6076) := b"0000000000000000_0000000000000000_0001110010111110_0000111111011000"; -- 0.11227511419615621
	pesos_i(6077) := b"0000000000000000_0000000000000000_0000111011010110_0001010100100110"; -- 0.057954141368011004
	pesos_i(6078) := b"0000000000000000_0000000000000000_0010100100110111_0110101011100001"; -- 0.16100185385440122
	pesos_i(6079) := b"0000000000000000_0000000000000000_0001110101011011_0100001000110100"; -- 0.1146737458201739
	pesos_i(6080) := b"0000000000000000_0000000000000000_0000010000001100_1100101101010100"; -- 0.01582022475588113
	pesos_i(6081) := b"0000000000000000_0000000000000000_0010001010100000_1110110101100000"; -- 0.1352680549727663
	pesos_i(6082) := b"1111111111111111_1111111111111111_1110011001100000_1001100011010010"; -- -0.10008854739897521
	pesos_i(6083) := b"0000000000000000_0000000000000000_0000000000000100_1110000100011100"; -- 7.44527304618723e-05
	pesos_i(6084) := b"0000000000000000_0000000000000000_0000111111111001_0101110111000110"; -- 0.062398777725294285
	pesos_i(6085) := b"1111111111111111_1111111111111111_1110100111010100_0111101001100100"; -- -0.08660159161821179
	pesos_i(6086) := b"0000000000000000_0000000000000000_0000110010011011_0010100111101110"; -- 0.04924261155850365
	pesos_i(6087) := b"0000000000000000_0000000000000000_0000101111100101_0100111011111100"; -- 0.046467720420680265
	pesos_i(6088) := b"1111111111111111_1111111111111111_1110001100100010_0001100010101001"; -- -0.11276098138999678
	pesos_i(6089) := b"0000000000000000_0000000000000000_0010011000100010_1010011000000111"; -- 0.1489661949096767
	pesos_i(6090) := b"0000000000000000_0000000000000000_0010000101011000_0101001100110101"; -- 0.13025398297644866
	pesos_i(6091) := b"1111111111111111_1111111111111111_1111000111111100_1111000100111100"; -- -0.05473415640296534
	pesos_i(6092) := b"1111111111111111_1111111111111111_1110011011011100_1010100101010100"; -- -0.09819547367750535
	pesos_i(6093) := b"0000000000000000_0000000000000000_0010010110101000_1000111010001111"; -- 0.14710322368555986
	pesos_i(6094) := b"0000000000000000_0000000000000000_0001111100000001_1101111011010110"; -- 0.12112229095307496
	pesos_i(6095) := b"1111111111111111_1111111111111111_1110101100110010_0100000011001100"; -- -0.08126444830092037
	pesos_i(6096) := b"1111111111111111_1111111111111111_1101011100110111_0011000111111011"; -- -0.15931403753295928
	pesos_i(6097) := b"1111111111111111_1111111111111111_1111101111001100_1111000111011111"; -- -0.016404040463811484
	pesos_i(6098) := b"1111111111111111_1111111111111111_1111101011101001_1010111010110001"; -- -0.019871789754841045
	pesos_i(6099) := b"0000000000000000_0000000000000000_0000000010001110_0001110011111001"; -- 0.00216847505601617
	pesos_i(6100) := b"1111111111111111_1111111111111111_1101111011010010_0010001000000110"; -- -0.1296061264036348
	pesos_i(6101) := b"1111111111111111_1111111111111111_1110100110101111_1101110100000010"; -- -0.08716028885443938
	pesos_i(6102) := b"0000000000000000_0000000000000000_0010001101001010_0001010001011101"; -- 0.13784911405914774
	pesos_i(6103) := b"1111111111111111_1111111111111111_1110001111101110_1100010000110110"; -- -0.1096379631043102
	pesos_i(6104) := b"1111111111111111_1111111111111111_1111011110111001_1111000001111010"; -- -0.03231904049658839
	pesos_i(6105) := b"1111111111111111_1111111111111111_1110010010111110_1100000101011001"; -- -0.10646430567133126
	pesos_i(6106) := b"1111111111111111_1111111111111111_1101001101010011_0011011101101111"; -- -0.17451146650207408
	pesos_i(6107) := b"1111111111111111_1111111111111111_1110011101110010_1100011101101001"; -- -0.09590486227614843
	pesos_i(6108) := b"1111111111111111_1111111111111111_1101011010001111_0001100011000000"; -- -0.16187901805855964
	pesos_i(6109) := b"1111111111111111_1111111111111111_1111111111011011_1011010100111010"; -- -0.0005537732699124998
	pesos_i(6110) := b"1111111111111111_1111111111111111_1111000010010010_1010001011000111"; -- -0.06026251450384482
	pesos_i(6111) := b"1111111111111111_1111111111111111_1101110001111101_1100101111010101"; -- -0.13870550200969162
	pesos_i(6112) := b"0000000000000000_0000000000000000_0000011011100001_1110000000010110"; -- 0.02688408405081333
	pesos_i(6113) := b"0000000000000000_0000000000000000_0010110001100100_1101000111110001"; -- 0.17341339232043199
	pesos_i(6114) := b"0000000000000000_0000000000000000_0000100101010010_0111010001011100"; -- 0.03641440625398069
	pesos_i(6115) := b"1111111111111111_1111111111111111_1110111010100011_0010001100111011"; -- -0.06782321752840388
	pesos_i(6116) := b"1111111111111111_1111111111111111_1110110010001010_1110001100111000"; -- -0.07600574386969682
	pesos_i(6117) := b"1111111111111111_1111111111111111_1111101111101001_0001101110001101"; -- -0.015974310094510603
	pesos_i(6118) := b"1111111111111111_1111111111111111_1110010011110010_0011110110100001"; -- -0.10567869957647634
	pesos_i(6119) := b"1111111111111111_1111111111111111_1110000101010100_1111011110010000"; -- -0.11979725591681267
	pesos_i(6120) := b"1111111111111111_1111111111111111_1101011000100010_1101010110011111"; -- -0.16353096841461615
	pesos_i(6121) := b"0000000000000000_0000000000000000_0001100000111010_1000111100100110"; -- 0.0946435420774144
	pesos_i(6122) := b"0000000000000000_0000000000000000_0010101000100111_1010000101101101"; -- 0.16466721460297626
	pesos_i(6123) := b"1111111111111111_1111111111111111_1111001010110111_0110101100111110"; -- -0.05188874938888459
	pesos_i(6124) := b"0000000000000000_0000000000000000_0000011001101010_0001011100001100"; -- 0.025056305366963433
	pesos_i(6125) := b"0000000000000000_0000000000000000_0010001010011101_1111010111101011"; -- 0.13522278762230927
	pesos_i(6126) := b"1111111111111111_1111111111111111_1101011100000001_1001000000001100"; -- -0.16013240531078649
	pesos_i(6127) := b"1111111111111111_1111111111111111_1101101101010100_0110110001010110"; -- -0.1432430543205583
	pesos_i(6128) := b"1111111111111111_1111111111111111_1101011100011010_1010011111110011"; -- -0.15974951086492525
	pesos_i(6129) := b"0000000000000000_0000000000000000_0010011000001100_0111111101110010"; -- 0.1486282017143565
	pesos_i(6130) := b"1111111111111111_1111111111111111_1111100010011101_1011000111011000"; -- -0.02884376978163426
	pesos_i(6131) := b"1111111111111111_1111111111111111_1110100101111101_0101101000100100"; -- -0.08793102847950343
	pesos_i(6132) := b"0000000000000000_0000000000000000_0010100010101100_0011000000110001"; -- 0.15887738405195356
	pesos_i(6133) := b"0000000000000000_0000000000000000_0010010000000010_0011101100101110"; -- 0.1406590450703116
	pesos_i(6134) := b"0000000000000000_0000000000000000_0010001000000011_0001110111000100"; -- 0.1328600505422996
	pesos_i(6135) := b"0000000000000000_0000000000000000_0000100000101110_0001010011010110"; -- 0.031953146203962314
	pesos_i(6136) := b"0000000000000000_0000000000000000_0010001011011111_1101111101011100"; -- 0.13622852332305294
	pesos_i(6137) := b"1111111111111111_1111111111111111_1110110010111010_1101101110110000"; -- -0.075273770806697
	pesos_i(6138) := b"1111111111111111_1111111111111111_1111001101110100_1110101101101101"; -- -0.04899719799698533
	pesos_i(6139) := b"1111111111111111_1111111111111111_1101110001111011_1010001010001001"; -- -0.13873848117913995
	pesos_i(6140) := b"0000000000000000_0000000000000000_0001100110001110_1110011100011110"; -- 0.09983677373946996
	pesos_i(6141) := b"0000000000000000_0000000000000000_0001000001100111_0000100100001011"; -- 0.06407219421397323
	pesos_i(6142) := b"0000000000000000_0000000000000000_0001110000001010_0000000101110110"; -- 0.10952767502167356
	pesos_i(6143) := b"1111111111111111_1111111111111111_1111010110001101_1011111001001000"; -- -0.04080591902182392
	pesos_i(6144) := b"0000000000000000_0000000000000000_0001010001111100_1010010101000000"; -- 0.08002693945165792
	pesos_i(6145) := b"1111111111111111_1111111111111111_1101011101110101_1011001010110110"; -- -0.15836031958165941
	pesos_i(6146) := b"0000000000000000_0000000000000000_0000101000001111_1000101000001000"; -- 0.03929960911445355
	pesos_i(6147) := b"1111111111111111_1111111111111111_1110100011100010_0000000101010110"; -- -0.09030143400735233
	pesos_i(6148) := b"0000000000000000_0000000000000000_0001010010110111_1011110110110001"; -- 0.08092866481719654
	pesos_i(6149) := b"0000000000000000_0000000000000000_0001100100111101_1011111101100000"; -- 0.0985984428704223
	pesos_i(6150) := b"0000000000000000_0000000000000000_0000100010001000_0101111010100111"; -- 0.03333083698356092
	pesos_i(6151) := b"1111111111111111_1111111111111111_1101011111100001_1010010011010000"; -- -0.15671319878011783
	pesos_i(6152) := b"1111111111111111_1111111111111111_1100010010000010_0110001100010000"; -- -0.23238545280570677
	pesos_i(6153) := b"1111111111111111_1111111111111111_1111010000110001_1010011101111000"; -- -0.04611733746166701
	pesos_i(6154) := b"0000000000000000_0000000000000000_0000000110100100_0101111100101100"; -- 0.006414364102369825
	pesos_i(6155) := b"1111111111111111_1111111111111111_1110100011101111_0111000011100011"; -- -0.0900964208393601
	pesos_i(6156) := b"0000000000000000_0000000000000000_0010100011101011_1001011011100101"; -- 0.1598448094115621
	pesos_i(6157) := b"1111111111111111_1111111111111111_1101110000000111_1001010100110100"; -- -0.1405092953634838
	pesos_i(6158) := b"1111111111111111_1111111111111111_1111010101010101_1111011111111110"; -- -0.04165697133777322
	pesos_i(6159) := b"1111111111111111_1111111111111111_1110010111111000_1101111011010100"; -- -0.1016712886120228
	pesos_i(6160) := b"1111111111111111_1111111111111111_1110011100000111_1100100110001111"; -- -0.09753742458958674
	pesos_i(6161) := b"1111111111111111_1111111111111111_1110011110010000_0001101011010010"; -- -0.09545738570303282
	pesos_i(6162) := b"1111111111111111_1111111111111111_1101111111111001_1100111000000010"; -- -0.12509453240074989
	pesos_i(6163) := b"0000000000000000_0000000000000000_0000001011011001_1100000001111101"; -- 0.011135130424397144
	pesos_i(6164) := b"1111111111111111_1111111111111111_1111010101111011_0010001100000111"; -- -0.041089831060551266
	pesos_i(6165) := b"0000000000000000_0000000000000000_0001001011001000_1001110110000010"; -- 0.07337364595113621
	pesos_i(6166) := b"1111111111111111_1111111111111111_1110001100110111_0111111101111100"; -- -0.11243441794114632
	pesos_i(6167) := b"1111111111111111_1111111111111111_1101110011000010_0001111110001100"; -- -0.1376629145247982
	pesos_i(6168) := b"1111111111111111_1111111111111111_1110011101010111_0011101100110100"; -- -0.09632520663406118
	pesos_i(6169) := b"0000000000000000_0000000000000000_0000011111011111_0011100111101011"; -- 0.030749912060640684
	pesos_i(6170) := b"1111111111111111_1111111111111111_1110100010011110_1000011011100101"; -- -0.09133107098968636
	pesos_i(6171) := b"0000000000000000_0000000000000000_0010010111111101_0111001010001010"; -- 0.14839855070385527
	pesos_i(6172) := b"1111111111111111_1111111111111111_1111101010001101_1000101001010010"; -- -0.02127776631011374
	pesos_i(6173) := b"0000000000000000_0000000000000000_0000011011101001_1000100011010101"; -- 0.027000953675592607
	pesos_i(6174) := b"0000000000000000_0000000000000000_0001100001101000_1001011110111111"; -- 0.0953459588617889
	pesos_i(6175) := b"1111111111111111_1111111111111111_1111110111101011_1111000110001100"; -- -0.008118537294625056
	pesos_i(6176) := b"0000000000000000_0000000000000000_0001101011101111_1010000100001100"; -- 0.10521894981390997
	pesos_i(6177) := b"0000000000000000_0000000000000000_0010010001001110_0001001110101000"; -- 0.14181635725635358
	pesos_i(6178) := b"0000000000000000_0000000000000000_0000000000100010_1011100010000010"; -- 0.000529796313066585
	pesos_i(6179) := b"0000000000000000_0000000000000000_0000000011000000_0001100010101010"; -- 0.0029311576719666848
	pesos_i(6180) := b"0000000000000000_0000000000000000_0001001101000000_0001101011001001"; -- 0.07519690891618512
	pesos_i(6181) := b"1111111111111111_1111111111111111_1110010100111110_1101010001010010"; -- -0.1045100497128279
	pesos_i(6182) := b"1111111111111111_1111111111111111_1110011011101100_0011111111011000"; -- -0.09795762050766696
	pesos_i(6183) := b"1111111111111111_1111111111111111_1110011010100100_0100000001111100"; -- -0.09905621510011565
	pesos_i(6184) := b"1111111111111111_1111111111111111_1111100010100111_0010011010111101"; -- -0.028699473341338266
	pesos_i(6185) := b"0000000000000000_0000000000000000_0000110110000001_1011101001101011"; -- 0.05276074509098706
	pesos_i(6186) := b"0000000000000000_0000000000000000_0000100000111100_0000110011001011"; -- 0.03216628988757278
	pesos_i(6187) := b"1111111111111111_1111111111111111_1111011101111101_1000111111010101"; -- -0.03324032832632118
	pesos_i(6188) := b"1111111111111111_1111111111111111_1111010100101011_0010010101101001"; -- -0.042310392343865716
	pesos_i(6189) := b"0000000000000000_0000000000000000_0010001111111111_1101100111001111"; -- 0.1406227235030493
	pesos_i(6190) := b"1111111111111111_1111111111111111_1110001111101110_1100100101110101"; -- -0.10963765046326127
	pesos_i(6191) := b"0000000000000000_0000000000000000_0000011100011111_1010110101101101"; -- 0.027827109501944378
	pesos_i(6192) := b"0000000000000000_0000000000000000_0000111100101101_0100111100000001"; -- 0.05928510443858129
	pesos_i(6193) := b"0000000000000000_0000000000000000_0001000000110101_0111100001110111"; -- 0.0633158961838802
	pesos_i(6194) := b"1111111111111111_1111111111111111_1110001010110111_0110011010111110"; -- -0.11438901778728947
	pesos_i(6195) := b"0000000000000000_0000000000000000_0001010101010000_0111011101101010"; -- 0.08325907078339147
	pesos_i(6196) := b"1111111111111111_1111111111111111_1111000100010010_0011001101010100"; -- -0.05831603236153268
	pesos_i(6197) := b"1111111111111111_1111111111111111_1111100001111100_0010110110011010"; -- -0.02935519215639861
	pesos_i(6198) := b"0000000000000000_0000000000000000_0000110011101110_0111010001000101"; -- 0.05051352202444077
	pesos_i(6199) := b"0000000000000000_0000000000000000_0010011110101100_0100001000110000"; -- 0.1549722067536025
	pesos_i(6200) := b"1111111111111111_1111111111111111_1101010011000001_0110000101011101"; -- -0.16892425037189446
	pesos_i(6201) := b"0000000000000000_0000000000000000_0000000100111100_1101100110011000"; -- 0.004834746899814866
	pesos_i(6202) := b"0000000000000000_0000000000000000_0010101001011101_0100010000011010"; -- 0.16548562649529294
	pesos_i(6203) := b"0000000000000000_0000000000000000_0000110100010000_1010000111100110"; -- 0.05103504057520696
	pesos_i(6204) := b"1111111111111111_1111111111111111_1101100100111100_1100001100010010"; -- -0.15141659551128764
	pesos_i(6205) := b"1111111111111111_1111111111111111_1110010001101000_0110100111000101"; -- -0.10778178167362278
	pesos_i(6206) := b"0000000000000000_0000000000000000_0001000000000010_1111011000110101"; -- 0.06254519277525715
	pesos_i(6207) := b"1111111111111111_1111111111111111_1101101100100100_0010100010011011"; -- -0.143979513340045
	pesos_i(6208) := b"1111111111111111_1111111111111111_1110101000101010_1001100110011010"; -- -0.08528747543736291
	pesos_i(6209) := b"1111111111111111_1111111111111111_1101011000110101_0100100010011110"; -- -0.16324945592999043
	pesos_i(6210) := b"0000000000000000_0000000000000000_0010000100110111_0011001011111011"; -- 0.1297485221334166
	pesos_i(6211) := b"1111111111111111_1111111111111111_1101010111000111_0110010100110110"; -- -0.16492621838618926
	pesos_i(6212) := b"0000000000000000_0000000000000000_0010000011011011_1000010110110000"; -- 0.12834964313242703
	pesos_i(6213) := b"0000000000000000_0000000000000000_0010101111010011_0110010011000000"; -- 0.17119435955012033
	pesos_i(6214) := b"0000000000000000_0000000000000000_0001100000111010_0110111010101110"; -- 0.09464160679272136
	pesos_i(6215) := b"1111111111111111_1111111111111111_1111001000011110_1110001011111111"; -- -0.05421620633468169
	pesos_i(6216) := b"1111111111111111_1111111111111111_1110011000000100_0110101110001001"; -- -0.10149505535533691
	pesos_i(6217) := b"1111111111111111_1111111111111111_1110101101101000_1001100011010001"; -- -0.08043522728488794
	pesos_i(6218) := b"0000000000000000_0000000000000000_0010010111001011_1110110010011100"; -- 0.1476428871726254
	pesos_i(6219) := b"0000000000000000_0000000000000000_0000110101110110_0101100100101001"; -- 0.05258710157528786
	pesos_i(6220) := b"1111111111111111_1111111111111111_1101101011110011_1011100011010011"; -- -0.14471859776766186
	pesos_i(6221) := b"0000000000000000_0000000000000000_0000111011010110_1101101011001010"; -- 0.05796592165046316
	pesos_i(6222) := b"0000000000000000_0000000000000000_0000010101111010_1000011101100001"; -- 0.02140089147277636
	pesos_i(6223) := b"0000000000000000_0000000000000000_0001100001111110_1100001101000000"; -- 0.09568424518510038
	pesos_i(6224) := b"0000000000000000_0000000000000000_0010110000001100_0000111101011111"; -- 0.1720590215762741
	pesos_i(6225) := b"1111111111111111_1111111111111111_1110100000001001_0111010010011101"; -- -0.0936057200990251
	pesos_i(6226) := b"1111111111111111_1111111111111111_1101011111011110_1111100011011000"; -- -0.15675396653016346
	pesos_i(6227) := b"1111111111111111_1111111111111111_1101111001101010_1110101110010101"; -- -0.13118102650475133
	pesos_i(6228) := b"0000000000000000_0000000000000000_0010110010101111_1110000111011100"; -- 0.1745587502417765
	pesos_i(6229) := b"0000000000000000_0000000000000000_0001010101011110_1110111011010101"; -- 0.0834798117699156
	pesos_i(6230) := b"1111111111111111_1111111111111111_1110101011100100_1011100101111111"; -- -0.08244743970677251
	pesos_i(6231) := b"0000000000000000_0000000000000000_0011010010000110_0100110100100011"; -- 0.20517427550280168
	pesos_i(6232) := b"1111111111111111_1111111111111111_1101100011011001_0011110100111101"; -- -0.15293519259381427
	pesos_i(6233) := b"0000000000000000_0000000000000000_0000011111010111_0001011001000001"; -- 0.030625716011555337
	pesos_i(6234) := b"1111111111111111_1111111111111111_1110010110001100_1000101101001001"; -- -0.10332421741981697
	pesos_i(6235) := b"0000000000000000_0000000000000000_0001110010011100_1100111011110100"; -- 0.11176770637863315
	pesos_i(6236) := b"1111111111111111_1111111111111111_1111011010110100_0001111010010000"; -- -0.03631409630655598
	pesos_i(6237) := b"1111111111111111_1111111111111111_1101110111100110_0111111000110100"; -- -0.13320170631573558
	pesos_i(6238) := b"1111111111111111_1111111111111111_1110001100001111_0011111000010101"; -- -0.11304866778859923
	pesos_i(6239) := b"0000000000000000_0000000000000000_0000110001101100_1011001111010010"; -- 0.04853366733726888
	pesos_i(6240) := b"1111111111111111_1111111111111111_1101100001011110_1110010000000101"; -- -0.15480208270500503
	pesos_i(6241) := b"0000000000000000_0000000000000000_0001000101110111_0101000101100111"; -- 0.0682268979136637
	pesos_i(6242) := b"1111111111111111_1111111111111111_1110010011100110_1001001010000001"; -- -0.10585674611236864
	pesos_i(6243) := b"1111111111111111_1111111111111111_1111111110001100_1001000011011011"; -- -0.0017613855605989842
	pesos_i(6244) := b"0000000000000000_0000000000000000_0001001100111100_1111101101001110"; -- 0.07514925616783323
	pesos_i(6245) := b"0000000000000000_0000000000000000_0010110000100011_1110010011100011"; -- 0.1724227002448544
	pesos_i(6246) := b"1111111111111111_1111111111111111_1110000100011101_0111111000001011"; -- -0.12064373229109916
	pesos_i(6247) := b"0000000000000000_0000000000000000_0001011010101001_1011111011001011"; -- 0.08852760760959608
	pesos_i(6248) := b"0000000000000000_0000000000000000_0000110111000010_0111000100100000"; -- 0.05374819783318033
	pesos_i(6249) := b"1111111111111111_1111111111111111_1111011010010111_1001101100111000"; -- -0.03674917102287035
	pesos_i(6250) := b"0000000000000000_0000000000000000_0000000111110000_0000111100110100"; -- 0.007569265608372765
	pesos_i(6251) := b"0000000000000000_0000000000000000_0001100111000100_1001010001111000"; -- 0.10065582209650584
	pesos_i(6252) := b"1111111111111111_1111111111111111_1111111100011011_0000101011111111"; -- -0.0034936073453753456
	pesos_i(6253) := b"1111111111111111_1111111111111111_1110000111110000_1101000011010001"; -- -0.11741919430059677
	pesos_i(6254) := b"0000000000000000_0000000000000000_0000010101011100_1011101010000011"; -- 0.020946175655307882
	pesos_i(6255) := b"0000000000000000_0000000000000000_0000111110110101_0101100010000010"; -- 0.06136086640939596
	pesos_i(6256) := b"0000000000000000_0000000000000000_0000100110011010_0001101111111111"; -- 0.037507772266392514
	pesos_i(6257) := b"0000000000000000_0000000000000000_0000001000101111_0001111010111000"; -- 0.0085314941542389
	pesos_i(6258) := b"0000000000000000_0000000000000000_0001111010110001_1010111001000010"; -- 0.11989869213298618
	pesos_i(6259) := b"0000000000000000_0000000000000000_0001100101100111_0000111000110010"; -- 0.09922875127068144
	pesos_i(6260) := b"0000000000000000_0000000000000000_0010100011011100_0001100101000001"; -- 0.1596084389016593
	pesos_i(6261) := b"1111111111111111_1111111111111111_1111110001111001_1111010001101101"; -- -0.013764117525299113
	pesos_i(6262) := b"1111111111111111_1111111111111111_1110001101101111_0010010000010011"; -- -0.11158537421215654
	pesos_i(6263) := b"1111111111111111_1111111111111111_1111010011001101_1100101100010101"; -- -0.04373484356106249
	pesos_i(6264) := b"1111111111111111_1111111111111111_1110000111100101_1111011101000011"; -- -0.11758474936200544
	pesos_i(6265) := b"1111111111111111_1111111111111111_1101011001101101_1001000011100111"; -- -0.1623906551554861
	pesos_i(6266) := b"0000000000000000_0000000000000000_0001010011011100_1010000101101000"; -- 0.08149155425440423
	pesos_i(6267) := b"1111111111111111_1111111111111111_1111100011000011_0101011101010010"; -- -0.0282693313591264
	pesos_i(6268) := b"1111111111111111_1111111111111111_1111101011100001_0001100110111010"; -- -0.020002738948761704
	pesos_i(6269) := b"1111111111111111_1111111111111111_1110001110000100_0111000011011010"; -- -0.11126036337352356
	pesos_i(6270) := b"1111111111111111_1111111111111111_1110010101100101_1100001101000001"; -- -0.10391597429433162
	pesos_i(6271) := b"1111111111111111_1111111111111111_1111111000011101_0101001111011011"; -- -0.007364996915053151
	pesos_i(6272) := b"1111111111111111_1111111111111111_1110100111100111_0000011000100111"; -- -0.08631860312036037
	pesos_i(6273) := b"0000000000000000_0000000000000000_0000101011100110_1011011000100000"; -- 0.042582877033023464
	pesos_i(6274) := b"1111111111111111_1111111111111111_1101101010000001_1110010101000001"; -- -0.14645545166157645
	pesos_i(6275) := b"1111111111111111_1111111111111111_1110010011001100_0101001110011010"; -- -0.1062572240156103
	pesos_i(6276) := b"0000000000000000_0000000000000000_0000000011100010_1110000101001100"; -- 0.0034619151295790817
	pesos_i(6277) := b"0000000000000000_0000000000000000_0001110000110011_0000100000100100"; -- 0.11015368335809517
	pesos_i(6278) := b"1111111111111111_1111111111111111_1101111100011111_1110110000110011"; -- -0.12841914891210454
	pesos_i(6279) := b"0000000000000000_0000000000000000_0000101100000101_1110101010111101"; -- 0.043059035440543555
	pesos_i(6280) := b"1111111111111111_1111111111111111_1110100001010010_1111111000000100"; -- -0.09248363879960152
	pesos_i(6281) := b"0000000000000000_0000000000000000_0000010001101011_0111110000010100"; -- 0.017265086063643555
	pesos_i(6282) := b"1111111111111111_1111111111111111_1101011100001101_1010010110101011"; -- -0.1599480110716869
	pesos_i(6283) := b"0000000000000000_0000000000000000_0000000001110110_0010100100110101"; -- 0.0018029931689397833
	pesos_i(6284) := b"1111111111111111_1111111111111111_1101110100111110_1011000001010110"; -- -0.13576219469444745
	pesos_i(6285) := b"0000000000000000_0000000000000000_0000001100101001_1110111110001101"; -- 0.012358638761397946
	pesos_i(6286) := b"1111111111111111_1111111111111111_1111000101100101_1111111011110011"; -- -0.05703741621092084
	pesos_i(6287) := b"0000000000000000_0000000000000000_0010100011001110_0111010001101011"; -- 0.15940024954554508
	pesos_i(6288) := b"1111111111111111_1111111111111111_1111001101001011_0011111000010010"; -- -0.049633141247006796
	pesos_i(6289) := b"0000000000000000_0000000000000000_0010001011110010_1001100011011111"; -- 0.136514238845861
	pesos_i(6290) := b"0000000000000000_0000000000000000_0000001011101110_1011101000110111"; -- 0.0114551911764659
	pesos_i(6291) := b"1111111111111111_1111111111111111_1110011101111011_0001011011000100"; -- -0.09577806209067867
	pesos_i(6292) := b"1111111111111111_1111111111111111_1111111110001100_0110001001000011"; -- -0.0017641626726191096
	pesos_i(6293) := b"1111111111111111_1111111111111111_1101100111101110_1001101111101111"; -- -0.14870286387847467
	pesos_i(6294) := b"1111111111111111_1111111111111111_1111111000011100_1101111010000111"; -- -0.007371990265767319
	pesos_i(6295) := b"1111111111111111_1111111111111111_1110001000000010_0100100011101011"; -- -0.11715263614960525
	pesos_i(6296) := b"0000000000000000_0000000000000000_0011010110111100_0010100100001000"; -- 0.20990234796941692
	pesos_i(6297) := b"1111111111111111_1111111111111111_1101110001001110_0110001101111001"; -- -0.139428885480714
	pesos_i(6298) := b"0000000000000000_0000000000000000_0000110111111001_0101100001000110"; -- 0.054585950066795313
	pesos_i(6299) := b"1111111111111111_1111111111111111_1101101000011101_1001010100111101"; -- -0.1479860998577301
	pesos_i(6300) := b"0000000000000000_0000000000000000_0000110111011010_0011101110100011"; -- 0.05411122061015085
	pesos_i(6301) := b"1111111111111111_1111111111111111_1110001011001001_0011000110110111"; -- -0.11411752019980416
	pesos_i(6302) := b"1111111111111111_1111111111111111_1111000110011110_0010010001110000"; -- -0.05618068943891775
	pesos_i(6303) := b"1111111111111111_1111111111111111_1101111000100000_1010110110001001"; -- -0.13231387514799853
	pesos_i(6304) := b"1111111111111111_1111111111111111_1111110010110000_0010011110110001"; -- -0.01293708729648968
	pesos_i(6305) := b"0000000000000000_0000000000000000_0001001000101111_1100000000000010"; -- 0.07104110767223137
	pesos_i(6306) := b"1111111111111111_1111111111111111_1110110111010010_1001010011111010"; -- -0.07100552464677413
	pesos_i(6307) := b"1111111111111111_1111111111111111_1111110111000110_1010000010100001"; -- -0.008687935622150342
	pesos_i(6308) := b"0000000000000000_0000000000000000_0000111010110100_1001001100100100"; -- 0.057442852261544226
	pesos_i(6309) := b"1111111111111111_1111111111111111_1101011110110000_1001001010111100"; -- -0.15746195709073268
	pesos_i(6310) := b"1111111111111111_1111111111111111_1111110010000101_1010001100100001"; -- -0.013585857835756993
	pesos_i(6311) := b"0000000000000000_0000000000000000_0010010011100010_0101110100100101"; -- 0.14407903822548304
	pesos_i(6312) := b"1111111111111111_1111111111111111_1110100111100100_0110110010011000"; -- -0.0863582735045668
	pesos_i(6313) := b"0000000000000000_0000000000000000_0000100101011001_1011010111001000"; -- 0.0365251171542428
	pesos_i(6314) := b"1111111111111111_1111111111111111_1101100000000001_0101010000011101"; -- -0.1562297276483748
	pesos_i(6315) := b"1111111111111111_1111111111111111_1111010000011011_0000110101001100"; -- -0.046462220248619596
	pesos_i(6316) := b"0000000000000000_0000000000000000_0010000011011000_0010111001001000"; -- 0.12829865695715095
	pesos_i(6317) := b"1111111111111111_1111111111111111_1110011111111011_0111110110010101"; -- -0.09381880872551944
	pesos_i(6318) := b"0000000000000000_0000000000000000_0000000110001111_0111101001111001"; -- 0.006095556834066099
	pesos_i(6319) := b"0000000000000000_0000000000000000_0001110000010110_0101011011111001"; -- 0.10971587741323505
	pesos_i(6320) := b"0000000000000000_0000000000000000_0000100011100101_0111010001000111"; -- 0.034751193262015756
	pesos_i(6321) := b"0000000000000000_0000000000000000_0001010000000010_0010110101100000"; -- 0.07815822210867815
	pesos_i(6322) := b"0000000000000000_0000000000000000_0001110001110011_1100010100100000"; -- 0.11114151031820496
	pesos_i(6323) := b"1111111111111111_1111111111111111_1101011010111111_1110110111101101"; -- -0.16113388983573865
	pesos_i(6324) := b"0000000000000000_0000000000000000_0010000101110101_0110001111000010"; -- 0.13069747432398107
	pesos_i(6325) := b"0000000000000000_0000000000000000_0010011111001100_0111001111010101"; -- 0.15546344720045752
	pesos_i(6326) := b"1111111111111111_1111111111111111_1111011100000000_1010000011011111"; -- -0.03514666139420655
	pesos_i(6327) := b"0000000000000000_0000000000000000_0000100100000001_0010111101001101"; -- 0.0351743280242939
	pesos_i(6328) := b"1111111111111111_1111111111111111_1110001111111110_0101111111110110"; -- -0.1093997977637583
	pesos_i(6329) := b"1111111111111111_1111111111111111_1101100011001100_0110001011111010"; -- -0.1531313076062993
	pesos_i(6330) := b"0000000000000000_0000000000000000_0001110001101010_0100100101001110"; -- 0.1109968010117725
	pesos_i(6331) := b"0000000000000000_0000000000000000_0010001011101000_0100111011000111"; -- 0.13635723454538046
	pesos_i(6332) := b"0000000000000000_0000000000000000_0001001100001010_1010101111111000"; -- 0.07438158799308088
	pesos_i(6333) := b"1111111111111111_1111111111111111_1101101001000101_1011001000110001"; -- -0.14737402248414558
	pesos_i(6334) := b"0000000000000000_0000000000000000_0000100101100110_0001110101000001"; -- 0.03671439006482427
	pesos_i(6335) := b"1111111111111111_1111111111111111_1110100100001111_0110000010010000"; -- -0.0896091125302681
	pesos_i(6336) := b"1111111111111111_1111111111111111_1110010101101110_0111010010001001"; -- -0.10378333711847727
	pesos_i(6337) := b"0000000000000000_0000000000000000_0001011100010001_1010100011010100"; -- 0.09011321227127836
	pesos_i(6338) := b"0000000000000000_0000000000000000_0001010110010101_1111100010011010"; -- 0.08431962736987555
	pesos_i(6339) := b"1111111111111111_1111111111111111_1111111101100111_0000111001001111"; -- -0.002333741766043319
	pesos_i(6340) := b"0000000000000000_0000000000000000_0010010101110111_0000100100100011"; -- 0.14634759058200286
	pesos_i(6341) := b"1111111111111111_1111111111111111_1110100010110000_0111011000011011"; -- -0.09105741341533467
	pesos_i(6342) := b"0000000000000000_0000000000000000_0000000100000100_0100111110000110"; -- 0.003972025107138759
	pesos_i(6343) := b"1111111111111111_1111111111111111_1110000000001011_1100000010111111"; -- -0.12482066471417369
	pesos_i(6344) := b"1111111111111111_1111111111111111_1110000001010001_1110111111011100"; -- -0.12374974125390509
	pesos_i(6345) := b"0000000000000000_0000000000000000_0000000001100000_0011101001010110"; -- 0.0014683208165722338
	pesos_i(6346) := b"1111111111111111_1111111111111111_1101111111100001_0011000000010110"; -- -0.12547015641224327
	pesos_i(6347) := b"1111111111111111_1111111111111111_1101010110100000_0010101000000100"; -- -0.16552483948609417
	pesos_i(6348) := b"0000000000000000_0000000000000000_0001101001010001_1000111000001001"; -- 0.1028069278944807
	pesos_i(6349) := b"1111111111111111_1111111111111111_1110100111101110_1100110010100110"; -- -0.08619996018471143
	pesos_i(6350) := b"0000000000000000_0000000000000000_0010111011000011_0101101000100001"; -- 0.1826683358811816
	pesos_i(6351) := b"0000000000000000_0000000000000000_0000000101110000_1011110101001010"; -- 0.005626516807557082
	pesos_i(6352) := b"1111111111111111_1111111111111111_1110000111010110_0111100111011100"; -- -0.1178211057340493
	pesos_i(6353) := b"0000000000000000_0000000000000000_0010010011111000_1100110111011010"; -- 0.14442144932578904
	pesos_i(6354) := b"0000000000000000_0000000000000000_0000110100110101_0110010101011111"; -- 0.051596008084508635
	pesos_i(6355) := b"1111111111111111_1111111111111111_1110111100010000_1100100000011101"; -- -0.0661501816743951
	pesos_i(6356) := b"1111111111111111_1111111111111111_1110101011000100_0011001000100011"; -- -0.08294378891651873
	pesos_i(6357) := b"0000000000000000_0000000000000000_0001100100000011_0011111011100001"; -- 0.09770577432896609
	pesos_i(6358) := b"1111111111111111_1111111111111111_1101111110110011_0101100001011111"; -- -0.12616965952558318
	pesos_i(6359) := b"0000000000000000_0000000000000000_0000110111000111_0010010011001001"; -- 0.053819941554615336
	pesos_i(6360) := b"0000000000000000_0000000000000000_0001101101111000_0111111010110001"; -- 0.10730735610289412
	pesos_i(6361) := b"0000000000000000_0000000000000000_0000001010011101_1110110100011010"; -- 0.010222262331843531
	pesos_i(6362) := b"1111111111111111_1111111111111111_1101101111010110_1111100100110010"; -- -0.14125101604897491
	pesos_i(6363) := b"1111111111111111_1111111111111111_1110011011110011_1001001101111110"; -- -0.09784582294069115
	pesos_i(6364) := b"1111111111111111_1111111111111111_1111010010111001_0011010000100111"; -- -0.04404901544147804
	pesos_i(6365) := b"0000000000000000_0000000000000000_0001101110000100_1100001100110000"; -- 0.10749454415916412
	pesos_i(6366) := b"1111111111111111_1111111111111111_1101111110110100_1010100101010101"; -- -0.12614957496256532
	pesos_i(6367) := b"0000000000000000_0000000000000000_0001110011110001_0000110100011001"; -- 0.11305314891017973
	pesos_i(6368) := b"0000000000000000_0000000000000000_0001000100001001_0111000001100000"; -- 0.06655027728327931
	pesos_i(6369) := b"0000000000000000_0000000000000000_0000100000000011_0010100111010001"; -- 0.031298268746527795
	pesos_i(6370) := b"1111111111111111_1111111111111111_1101010101010010_0011010101111100"; -- -0.166714341355732
	pesos_i(6371) := b"1111111111111111_1111111111111111_1111100110010010_1010011111010110"; -- -0.0251059630818877
	pesos_i(6372) := b"1111111111111111_1111111111111111_1101111011101001_0000000010001111"; -- -0.12925716884983535
	pesos_i(6373) := b"1111111111111111_1111111111111111_1110101110110111_0001110110100010"; -- -0.07923712523822653
	pesos_i(6374) := b"0000000000000000_0000000000000000_0000000100110001_0011011100010011"; -- 0.004657213322886193
	pesos_i(6375) := b"1111111111111111_1111111111111111_1110100101011010_1011100000001001"; -- -0.08845948959137526
	pesos_i(6376) := b"0000000000000000_0000000000000000_0000011010000100_1010010000000101"; -- 0.025461436494922052
	pesos_i(6377) := b"1111111111111111_1111111111111111_1111111001001000_1110100100111011"; -- -0.006699965621537735
	pesos_i(6378) := b"0000000000000000_0000000000000000_0000000110111111_1110100101010100"; -- 0.006834586214758826
	pesos_i(6379) := b"0000000000000000_0000000000000000_0010101000010001_1110000010011010"; -- 0.1643352867919864
	pesos_i(6380) := b"1111111111111111_1111111111111111_1110110100011111_1010111111011101"; -- -0.07373524531361253
	pesos_i(6381) := b"0000000000000000_0000000000000000_0000100010000001_0100101101100111"; -- 0.03322287803228365
	pesos_i(6382) := b"0000000000000000_0000000000000000_0001000101001011_1010000011101101"; -- 0.06756025121088438
	pesos_i(6383) := b"1111111111111111_1111111111111111_1110111100111001_1010101001110001"; -- -0.06552633987816761
	pesos_i(6384) := b"0000000000000000_0000000000000000_0010110001011010_1111100000111000"; -- 0.17326308596270615
	pesos_i(6385) := b"1111111111111111_1111111111111111_1111110001101101_1111001001011011"; -- -0.013947346553856781
	pesos_i(6386) := b"0000000000000000_0000000000000000_0000100011000100_1100000001001101"; -- 0.034252184565601286
	pesos_i(6387) := b"1111111111111111_1111111111111111_1111101111111000_0010101000110101"; -- -0.015744554617158457
	pesos_i(6388) := b"1111111111111111_1111111111111111_1110000101000111_0111100110100000"; -- -0.12000312648096578
	pesos_i(6389) := b"1111111111111111_1111111111111111_1101111001010101_0000110001101000"; -- -0.13151476341081225
	pesos_i(6390) := b"1111111111111111_1111111111111111_1110110101111110_1101111001010100"; -- -0.07228289087807901
	pesos_i(6391) := b"0000000000000000_0000000000000000_0010000100011101_1111000011011010"; -- 0.1293631107901359
	pesos_i(6392) := b"1111111111111111_1111111111111111_1110001000111010_0011001101100111"; -- -0.11629942641960661
	pesos_i(6393) := b"0000000000000000_0000000000000000_0001011101010011_1110110010110001"; -- 0.09112433745051125
	pesos_i(6394) := b"1111111111111111_1111111111111111_1111011100000001_0111101001000011"; -- -0.03513370384825379
	pesos_i(6395) := b"1111111111111111_1111111111111111_1111010110001110_1000101000010110"; -- -0.04079377146248589
	pesos_i(6396) := b"0000000000000000_0000000000000000_0000101111100111_1001101010111111"; -- 0.04650275380414276
	pesos_i(6397) := b"0000000000000000_0000000000000000_0010100100000011_0111011000001111"; -- 0.16020906310746486
	pesos_i(6398) := b"0000000000000000_0000000000000000_0010001011110000_0111111001001110"; -- 0.13648213774601559
	pesos_i(6399) := b"0000000000000000_0000000000000000_0000010011101000_0011110110100101"; -- 0.019168713292586955
	pesos_i(6400) := b"0000000000000000_0000000000000000_0000010011001001_0100010010000111"; -- 0.01869610122720003
	pesos_i(6401) := b"0000000000000000_0000000000000000_0000111001101101_1110010100100101"; -- 0.056364366072867815
	pesos_i(6402) := b"0000000000000000_0000000000000000_0010010100000000_1011100100110000"; -- 0.1445422879817493
	pesos_i(6403) := b"0000000000000000_0000000000000000_0000010011010010_1011001111011000"; -- 0.018840065118153233
	pesos_i(6404) := b"1111111111111111_1111111111111111_1110111100111001_0101011100100000"; -- -0.06553130599946985
	pesos_i(6405) := b"0000000000000000_0000000000000000_0001110000001001_1101110100011001"; -- 0.10952550744284485
	pesos_i(6406) := b"1111111111111111_1111111111111111_1110011111111100_1011010011000010"; -- -0.09380026124692595
	pesos_i(6407) := b"1111111111111111_1111111111111111_1111111101011101_1110101000011011"; -- -0.00247322883280678
	pesos_i(6408) := b"1111111111111111_1111111111111111_1101011000110011_0011100011110110"; -- -0.1632809065645486
	pesos_i(6409) := b"1111111111111111_1111111111111111_1111000101110001_1100110000011000"; -- -0.05685734179554027
	pesos_i(6410) := b"0000000000000000_0000000000000000_0000001100111001_1001010111101000"; -- 0.012597436006248837
	pesos_i(6411) := b"1111111111111111_1111111111111111_1111101101001101_1101010011111111"; -- -0.01834362767887544
	pesos_i(6412) := b"1111111111111111_1111111111111111_1111001111100111_0011010000010010"; -- -0.04725336613942914
	pesos_i(6413) := b"0000000000000000_0000000000000000_0010000000000111_1010010110110011"; -- 0.12511668792021968
	pesos_i(6414) := b"1111111111111111_1111111111111111_1101011001001101_0011001000001110"; -- -0.1628845897542444
	pesos_i(6415) := b"1111111111111111_1111111111111111_1101110100010001_1001010110100001"; -- -0.1364504320722391
	pesos_i(6416) := b"0000000000000000_0000000000000000_0001111111011111_1100001001100101"; -- 0.12450804671194979
	pesos_i(6417) := b"0000000000000000_0000000000000000_0010110111111001_0001101110000001"; -- 0.17958232779644015
	pesos_i(6418) := b"0000000000000000_0000000000000000_0001100100110011_1111011101000000"; -- 0.0984491853933478
	pesos_i(6419) := b"0000000000000000_0000000000000000_0010011101100000_1001110101011000"; -- 0.15381797206376627
	pesos_i(6420) := b"0000000000000000_0000000000000000_0001101011101000_0111000001100010"; -- 0.10510923749822107
	pesos_i(6421) := b"1111111111111111_1111111111111111_1111100110101110_1000011111111000"; -- -0.024680616356766938
	pesos_i(6422) := b"1111111111111111_1111111111111111_1110001110111110_0101100000001000"; -- -0.11037683304886646
	pesos_i(6423) := b"1111111111111111_1111111111111111_1111111010101011_0111011001101011"; -- -0.005196188880017929
	pesos_i(6424) := b"0000000000000000_0000000000000000_0001000000001100_0011111101011000"; -- 0.0626868811330989
	pesos_i(6425) := b"1111111111111111_1111111111111111_1110011010100100_1000110000101001"; -- -0.09905170431235165
	pesos_i(6426) := b"0000000000000000_0000000000000000_0000110000000100_1000010001000111"; -- 0.046943919463166305
	pesos_i(6427) := b"0000000000000000_0000000000000000_0000101011001000_1010001010101000"; -- 0.04212395286795204
	pesos_i(6428) := b"1111111111111111_1111111111111111_1101100000100100_1010110000100100"; -- -0.15569042316354587
	pesos_i(6429) := b"0000000000000000_0000000000000000_0010001000011010_1011000110000110"; -- 0.1332198097171248
	pesos_i(6430) := b"0000000000000000_0000000000000000_0001101001001111_1100111010101100"; -- 0.10278026297585334
	pesos_i(6431) := b"1111111111111111_1111111111111111_1111010111000110_1001011101010001"; -- -0.0399384905993187
	pesos_i(6432) := b"0000000000000000_0000000000000000_0001101100110010_1100010111101110"; -- 0.10624348694383404
	pesos_i(6433) := b"0000000000000000_0000000000000000_0001011000001011_1101111001001110"; -- 0.08611859696801477
	pesos_i(6434) := b"0000000000000000_0000000000000000_0010010010100111_1011011011100001"; -- 0.14318411828462999
	pesos_i(6435) := b"0000000000000000_0000000000000000_0001011101101100_0101010101000111"; -- 0.09149678216963285
	pesos_i(6436) := b"0000000000000000_0000000000000000_0000111101010100_0110011001101000"; -- 0.05988159207529001
	pesos_i(6437) := b"0000000000000000_0000000000000000_0001001011001110_0111001001001011"; -- 0.0734626229657223
	pesos_i(6438) := b"1111111111111111_1111111111111111_1111010000111101_1100010101001100"; -- -0.04593245408935103
	pesos_i(6439) := b"0000000000000000_0000000000000000_0000101001000010_0111010001100010"; -- 0.04007651703360057
	pesos_i(6440) := b"0000000000000000_0000000000000000_0010100000001001_1110100100101000"; -- 0.15640122625484568
	pesos_i(6441) := b"0000000000000000_0000000000000000_0000010100110100_1001100101110011"; -- 0.020333853216977706
	pesos_i(6442) := b"1111111111111111_1111111111111111_1101110000000011_1100001011010101"; -- -0.14056761083726274
	pesos_i(6443) := b"1111111111111111_1111111111111111_1101010010000100_0010111000110000"; -- -0.16985808691454848
	pesos_i(6444) := b"0000000000000000_0000000000000000_0010101000100010_1100111010101110"; -- 0.16459361797162486
	pesos_i(6445) := b"1111111111111111_1111111111111111_1111101111111010_1101111011110000"; -- -0.015703264552632743
	pesos_i(6446) := b"0000000000000000_0000000000000000_0000100000000011_0101111000010100"; -- 0.031301383880224555
	pesos_i(6447) := b"0000000000000000_0000000000000000_0010001110111011_1110010111001100"; -- 0.1395858406024005
	pesos_i(6448) := b"1111111111111111_1111111111111111_1111010110100010_1100110100001001"; -- -0.040484605048995564
	pesos_i(6449) := b"1111111111111111_1111111111111111_1111011010011101_0100000111100101"; -- -0.036662942533709005
	pesos_i(6450) := b"0000000000000000_0000000000000000_0010101101100001_0111010111010010"; -- 0.169455875186643
	pesos_i(6451) := b"0000000000000000_0000000000000000_0000001111001001_0000001101010100"; -- 0.014785964962593164
	pesos_i(6452) := b"0000000000000000_0000000000000000_0001000011011100_0100110111111100"; -- 0.06586158178180776
	pesos_i(6453) := b"1111111111111111_1111111111111111_1101101100110001_0001110011111001"; -- -0.1437818425424279
	pesos_i(6454) := b"0000000000000000_0000000000000000_0001100101110011_0101011001111010"; -- 0.09941616508364026
	pesos_i(6455) := b"1111111111111111_1111111111111111_1111001010110001_0101100111111111"; -- -0.05198133018390357
	pesos_i(6456) := b"0000000000000000_0000000000000000_0000100001000101_0001100000101110"; -- 0.03230429768079651
	pesos_i(6457) := b"0000000000000000_0000000000000000_0010010011101111_0110111010110111"; -- 0.14427844978175575
	pesos_i(6458) := b"1111111111111111_1111111111111111_1110000101011010_0101001000111011"; -- -0.11971555768549438
	pesos_i(6459) := b"1111111111111111_1111111111111111_1111110001001111_1000101011011000"; -- -0.014411279862951463
	pesos_i(6460) := b"0000000000000000_0000000000000000_0000000110111010_1011011100000101"; -- 0.006755293622802397
	pesos_i(6461) := b"1111111111111111_1111111111111111_1111100001010101_1011011010001010"; -- -0.029942122816394825
	pesos_i(6462) := b"1111111111111111_1111111111111111_1111010011101110_1001101001110100"; -- -0.043234201982873983
	pesos_i(6463) := b"1111111111111111_1111111111111111_1111011100111101_0111111110010110"; -- -0.03421785916305668
	pesos_i(6464) := b"1111111111111111_1111111111111111_1110000000111111_0011010111100010"; -- -0.12403548465729497
	pesos_i(6465) := b"0000000000000000_0000000000000000_0000011111111001_1110110101110001"; -- 0.03115734109695605
	pesos_i(6466) := b"1111111111111111_1111111111111111_1111110111000100_0110101000111100"; -- -0.008721695239099549
	pesos_i(6467) := b"1111111111111111_1111111111111111_1101011001101000_1011011001100001"; -- -0.1624647152264678
	pesos_i(6468) := b"0000000000000000_0000000000000000_0000110001011111_0101110010101010"; -- 0.04833010818890511
	pesos_i(6469) := b"0000000000000000_0000000000000000_0000000001100011_1110101100001011"; -- 0.0015246296642395611
	pesos_i(6470) := b"0000000000000000_0000000000000000_0000010011000101_1101101000011100"; -- 0.018643981893436364
	pesos_i(6471) := b"0000000000000000_0000000000000000_0001111010110001_1010011110111101"; -- 0.11989830364164679
	pesos_i(6472) := b"1111111111111111_1111111111111111_1111001101111101_0001000010100010"; -- -0.0488729100273449
	pesos_i(6473) := b"0000000000000000_0000000000000000_0000110100101110_0110111110001011"; -- 0.05148980277182623
	pesos_i(6474) := b"1111111111111111_1111111111111111_1110101001010101_1010111000110111"; -- -0.08463011880980054
	pesos_i(6475) := b"0000000000000000_0000000000000000_0001111010001010_1011100010110011"; -- 0.11930422173983184
	pesos_i(6476) := b"0000000000000000_0000000000000000_0000101000000101_0011010000000010"; -- 0.03914189382753897
	pesos_i(6477) := b"0000000000000000_0000000000000000_0001100110101100_1001101101100011"; -- 0.10029002357100024
	pesos_i(6478) := b"0000000000000000_0000000000000000_0001100110010011_0000001110010001"; -- 0.09989950447901316
	pesos_i(6479) := b"1111111111111111_1111111111111111_1101111001110010_0101101001000010"; -- -0.13106761816791448
	pesos_i(6480) := b"1111111111111111_1111111111111111_1101010010001101_0000011111011101"; -- -0.16972304198962634
	pesos_i(6481) := b"0000000000000000_0000000000000000_0010100111011101_0010001010011101"; -- 0.16353050555272222
	pesos_i(6482) := b"1111111111111111_1111111111111111_1111001001100110_1110110101011011"; -- -0.05311695608996839
	pesos_i(6483) := b"0000000000000000_0000000000000000_0010010001111111_1000111011111010"; -- 0.1425713883409873
	pesos_i(6484) := b"0000000000000000_0000000000000000_0010101110101010_1111111101110101"; -- 0.17057797050632476
	pesos_i(6485) := b"0000000000000000_0000000000000000_0010000001011001_1101011111110101"; -- 0.12637090433849357
	pesos_i(6486) := b"0000000000000000_0000000000000000_0000100001011110_0011100111011000"; -- 0.03268777396935976
	pesos_i(6487) := b"0000000000000000_0000000000000000_0000011000100010_1011110100011001"; -- 0.0239675699260818
	pesos_i(6488) := b"0000000000000000_0000000000000000_0001110101101111_1001011011000100"; -- 0.11498396198509069
	pesos_i(6489) := b"1111111111111111_1111111111111111_1111111110011000_1100001111110101"; -- -0.0015752340950660052
	pesos_i(6490) := b"0000000000000000_0000000000000000_0001101100110100_0110111011110010"; -- 0.10626881984915482
	pesos_i(6491) := b"1111111111111111_1111111111111111_1111001111010101_1000110010110011"; -- -0.04752274158343558
	pesos_i(6492) := b"0000000000000000_0000000000000000_0010010111011011_1011101011111110"; -- 0.14788407044855348
	pesos_i(6493) := b"1111111111111111_1111111111111111_1111001110110101_1100011010100111"; -- -0.04800756862753902
	pesos_i(6494) := b"0000000000000000_0000000000000000_0000001000011001_0000101100010011"; -- 0.008194629715196071
	pesos_i(6495) := b"0000000000000000_0000000000000000_0010101000001110_0111011001101111"; -- 0.1642831822822405
	pesos_i(6496) := b"1111111111111111_1111111111111111_1110010000110001_0011010010001100"; -- -0.10862418723435942
	pesos_i(6497) := b"1111111111111111_1111111111111111_1101110010000111_1001011100010101"; -- -0.13855605834210186
	pesos_i(6498) := b"1111111111111111_1111111111111111_1101100000111000_0111111011001001"; -- -0.155387950891111
	pesos_i(6499) := b"0000000000000000_0000000000000000_0000001110101010_1110101111111100"; -- 0.014326809817882556
	pesos_i(6500) := b"1111111111111111_1111111111111111_1111111100010111_0111100010110000"; -- -0.0035481043620193987
	pesos_i(6501) := b"1111111111111111_1111111111111111_1111100110100011_1000100001111000"; -- -0.02484843326288925
	pesos_i(6502) := b"1111111111111111_1111111111111111_1110001111001001_1010000010110011"; -- -0.1102046550364088
	pesos_i(6503) := b"0000000000000000_0000000000000000_0000111011001100_1000111011101100"; -- 0.057808811685022
	pesos_i(6504) := b"0000000000000000_0000000000000000_0010001111010111_1011000100000110"; -- 0.14000994098616784
	pesos_i(6505) := b"0000000000000000_0000000000000000_0010000110111010_1011110011000011"; -- 0.13175563580177943
	pesos_i(6506) := b"0000000000000000_0000000000000000_0000000011010011_0011100000100001"; -- 0.0032229500321174368
	pesos_i(6507) := b"0000000000000000_0000000000000000_0001100001101111_0000111011001011"; -- 0.09544460736022399
	pesos_i(6508) := b"1111111111111111_1111111111111111_1110110100111111_1100110110001100"; -- -0.07324519482849894
	pesos_i(6509) := b"1111111111111111_1111111111111111_1111000010111100_1011101010110000"; -- -0.0596202201377545
	pesos_i(6510) := b"0000000000000000_0000000000000000_0000111100111001_1110101010010100"; -- 0.059477482989754686
	pesos_i(6511) := b"1111111111111111_1111111111111111_1101111010111100_1010011101101011"; -- -0.129933868655606
	pesos_i(6512) := b"0000000000000000_0000000000000000_0000000111101000_1010100110101101"; -- 0.007456402622649488
	pesos_i(6513) := b"1111111111111111_1111111111111111_1111101111010101_0111011010101110"; -- -0.016274054062033666
	pesos_i(6514) := b"1111111111111111_1111111111111111_1101100000111001_0110111000100000"; -- -0.15537368507809124
	pesos_i(6515) := b"0000000000000000_0000000000000000_0001001000110011_0000110001000110"; -- 0.07109142982863226
	pesos_i(6516) := b"1111111111111111_1111111111111111_1101110011001111_1000100110010100"; -- -0.13745823025361797
	pesos_i(6517) := b"0000000000000000_0000000000000000_0001011111001100_1000001011101000"; -- 0.09296434566214795
	pesos_i(6518) := b"0000000000000000_0000000000000000_0001110011101100_1010111100001001"; -- 0.11298650704329301
	pesos_i(6519) := b"0000000000000000_0000000000000000_0010110101001101_0010101011111000"; -- 0.17695873778896037
	pesos_i(6520) := b"1111111111111111_1111111111111111_1110001100001011_1111110100101100"; -- -0.11309831305457393
	pesos_i(6521) := b"0000000000000000_0000000000000000_0001001011011110_0001000100001001"; -- 0.07370096659759086
	pesos_i(6522) := b"0000000000000000_0000000000000000_0000100010011100_0100110011011000"; -- 0.033634951366049166
	pesos_i(6523) := b"1111111111111111_1111111111111111_1110110001001001_0100000000101000"; -- -0.07700728434672273
	pesos_i(6524) := b"0000000000000000_0000000000000000_0000100000111110_1010101000010011"; -- 0.03220618206551225
	pesos_i(6525) := b"0000000000000000_0000000000000000_0010101000011000_1100010101001100"; -- 0.16444047077890978
	pesos_i(6526) := b"1111111111111111_1111111111111111_1111111001011000_1001001011001110"; -- -0.006460976356471511
	pesos_i(6527) := b"0000000000000000_0000000000000000_0001000010010010_1111010101111100"; -- 0.06474241528707919
	pesos_i(6528) := b"1111111111111111_1111111111111111_1110100110111101_0101001010011101"; -- -0.08695491472272582
	pesos_i(6529) := b"0000000000000000_0000000000000000_0011000110011110_1010101000100110"; -- 0.1938272802538662
	pesos_i(6530) := b"0000000000000000_0000000000000000_0000011111011111_1110010011011101"; -- 0.03076010119549945
	pesos_i(6531) := b"1111111111111111_1111111111111111_1110010110110110_1010110001101001"; -- -0.10268137396582157
	pesos_i(6532) := b"0000000000000000_0000000000000000_0000001011100001_0010110011011000"; -- 0.01124840052098825
	pesos_i(6533) := b"0000000000000000_0000000000000000_0001100011010011_1101100111100101"; -- 0.09698259207903188
	pesos_i(6534) := b"0000000000000000_0000000000000000_0001101001111101_0110011010100010"; -- 0.10347596606466736
	pesos_i(6535) := b"1111111111111111_1111111111111111_1111110110100111_0001011111000011"; -- -0.009169115819356548
	pesos_i(6536) := b"1111111111111111_1111111111111111_1100010011010001_1110101000111011"; -- -0.2311719519639876
	pesos_i(6537) := b"1111111111111111_1111111111111111_1110001000110010_1000100011101010"; -- -0.11641639990466866
	pesos_i(6538) := b"1111111111111111_1111111111111111_1110011000101101_0100100000010000"; -- -0.10087155923768162
	pesos_i(6539) := b"0000000000000000_0000000000000000_0000111000011001_0101100000110111"; -- 0.05507422773737498
	pesos_i(6540) := b"1111111111111111_1111111111111111_1110110101110100_1000110111011011"; -- -0.07244027530191002
	pesos_i(6541) := b"1111111111111111_1111111111111111_1110011000100100_1000000001000101"; -- -0.10100553821387877
	pesos_i(6542) := b"0000000000000000_0000000000000000_0001110010110110_0011111000101000"; -- 0.11215580442160246
	pesos_i(6543) := b"1111111111111111_1111111111111111_1110100110101000_1011100010100010"; -- -0.08726926850613163
	pesos_i(6544) := b"1111111111111111_1111111111111111_1111110110001000_1001100001011111"; -- -0.009634472601652788
	pesos_i(6545) := b"0000000000000000_0000000000000000_0001110000010111_1101100100001100"; -- 0.10973888911375657
	pesos_i(6546) := b"0000000000000000_0000000000000000_0001111011010101_1111001111000100"; -- 0.12045215172770486
	pesos_i(6547) := b"1111111111111111_1111111111111111_1111011000011101_1101010110110101"; -- -0.03860725714279164
	pesos_i(6548) := b"1111111111111111_1111111111111111_1110011100101111_0110010111111001"; -- -0.09693300885915575
	pesos_i(6549) := b"0000000000000000_0000000000000000_0001110111011010_1010100000010111"; -- 0.11661768485181578
	pesos_i(6550) := b"0000000000000000_0000000000000000_0010101001010111_0100010100011110"; -- 0.1653941343861296
	pesos_i(6551) := b"0000000000000000_0000000000000000_0010000000011000_0100100011001100"; -- 0.12537054998410319
	pesos_i(6552) := b"0000000000000000_0000000000000000_0010100001001110_1001000001100001"; -- 0.15744879110878698
	pesos_i(6553) := b"1111111111111111_1111111111111111_1111110010100011_0101110011101011"; -- -0.013132278961850824
	pesos_i(6554) := b"1111111111111111_1111111111111111_1101010101110101_1110011101110000"; -- -0.16616967704000618
	pesos_i(6555) := b"0000000000000000_0000000000000000_0000001010010101_0110100101100011"; -- 0.010092341119773699
	pesos_i(6556) := b"1111111111111111_1111111111111111_1101100100111001_1000001000010100"; -- -0.1514662457915765
	pesos_i(6557) := b"0000000000000000_0000000000000000_0000001000101011_0110110000100001"; -- 0.008475072798404835
	pesos_i(6558) := b"0000000000000000_0000000000000000_0001111110011100_1001110110010111"; -- 0.12348351419319212
	pesos_i(6559) := b"0000000000000000_0000000000000000_0000101010000101_0010110111101011"; -- 0.04109465591968578
	pesos_i(6560) := b"0000000000000000_0000000000000000_0000000100011111_0110001001011000"; -- 0.00438513415768696
	pesos_i(6561) := b"0000000000000000_0000000000000000_0000000100000100_0101110110001010"; -- 0.003972860593191726
	pesos_i(6562) := b"1111111111111111_1111111111111111_1110010111101000_0101101000011111"; -- -0.10192333940778495
	pesos_i(6563) := b"1111111111111111_1111111111111111_1101111110001010_0111001100011100"; -- -0.12679367599080682
	pesos_i(6564) := b"0000000000000000_0000000000000000_0010011001011010_1100101101010100"; -- 0.1498229104132771
	pesos_i(6565) := b"1111111111111111_1111111111111111_1110111110100111_1000001010000000"; -- -0.06385025390513903
	pesos_i(6566) := b"0000000000000000_0000000000000000_0010110100111010_1011100000010011"; -- 0.1766772314532375
	pesos_i(6567) := b"1111111111111111_1111111111111111_1101111010000001_0011000100001110"; -- -0.13084119226517654
	pesos_i(6568) := b"0000000000000000_0000000000000000_0001010100001100_1010110111011000"; -- 0.08222471739478829
	pesos_i(6569) := b"1111111111111111_1111111111111111_1110110101101001_1001110001010101"; -- -0.07260725895774386
	pesos_i(6570) := b"0000000000000000_0000000000000000_0010011001100011_0011111100001100"; -- 0.1499518779244767
	pesos_i(6571) := b"0000000000000000_0000000000000000_0000101100010001_1100111010011101"; -- 0.0432404645759097
	pesos_i(6572) := b"1111111111111111_1111111111111111_1111011110100000_1101001101101101"; -- -0.032702241842644725
	pesos_i(6573) := b"1111111111111111_1111111111111111_1111010100010011_1111000100101101"; -- -0.04266445781092166
	pesos_i(6574) := b"0000000000000000_0000000000000000_0000001000101111_0101110010110110"; -- 0.008535189113123839
	pesos_i(6575) := b"1111111111111111_1111111111111111_1111000111011110_1011000101001000"; -- -0.05519573207294735
	pesos_i(6576) := b"1111111111111111_1111111111111111_1110100000111111_1100001110101011"; -- -0.09277703350587892
	pesos_i(6577) := b"0000000000000000_0000000000000000_0010000100101000_0111000101011000"; -- 0.12952335747271806
	pesos_i(6578) := b"1111111111111111_1111111111111111_1111011101010110_0001111101001000"; -- -0.0338421297017068
	pesos_i(6579) := b"0000000000000000_0000000000000000_0001100110000110_1000010011100110"; -- 0.0997088491115502
	pesos_i(6580) := b"1111111111111111_1111111111111111_1111011011010001_0011100101100100"; -- -0.035869992263649134
	pesos_i(6581) := b"0000000000000000_0000000000000000_0011001101010101_1101001111001001"; -- 0.20052837053335273
	pesos_i(6582) := b"0000000000000000_0000000000000000_0000110001101100_1110011111000110"; -- 0.048536764031172484
	pesos_i(6583) := b"0000000000000000_0000000000000000_0001101111110101_0011010110101111"; -- 0.10921035302215691
	pesos_i(6584) := b"1111111111111111_1111111111111111_1101101100010010_1100101000110010"; -- -0.14424454008271986
	pesos_i(6585) := b"1111111111111111_1111111111111111_1110001101011000_1100101000110011"; -- -0.11192642461086759
	pesos_i(6586) := b"0000000000000000_0000000000000000_0000110100000011_0010111001010010"; -- 0.050829787165842924
	pesos_i(6587) := b"0000000000000000_0000000000000000_0010101000111000_0000010101101011"; -- 0.16491731507486398
	pesos_i(6588) := b"1111111111111111_1111111111111111_1110011110101001_1111010111101111"; -- -0.09506285584031865
	pesos_i(6589) := b"1111111111111111_1111111111111111_1111001110110001_1100101010101011"; -- -0.04806836429707261
	pesos_i(6590) := b"1111111111111111_1111111111111111_1101101100110101_1011011011110010"; -- -0.1437116297788041
	pesos_i(6591) := b"0000000000000000_0000000000000000_0010101010110010_0011001111010000"; -- 0.166781652807702
	pesos_i(6592) := b"1111111111111111_1111111111111111_1111101001000110_1111110111011010"; -- -0.02235425405006755
	pesos_i(6593) := b"1111111111111111_1111111111111111_1110011000011110_0100101010001111"; -- -0.10110029221613936
	pesos_i(6594) := b"1111111111111111_1111111111111111_1111111110010101_0100000110111011"; -- -0.0016287726356247444
	pesos_i(6595) := b"0000000000000000_0000000000000000_0000001110111010_0100011110101111"; -- 0.014561157436106077
	pesos_i(6596) := b"1111111111111111_1111111111111111_1111010010011100_0100111111011111"; -- -0.044489868129559636
	pesos_i(6597) := b"0000000000000000_0000000000000000_0001111101010101_0111100110000010"; -- 0.12239798951718626
	pesos_i(6598) := b"1111111111111111_1111111111111111_1111000110100011_1100000010100001"; -- -0.05609508591903946
	pesos_i(6599) := b"0000000000000000_0000000000000000_0000010000011111_1110101100000011"; -- 0.016112030190041936
	pesos_i(6600) := b"1111111111111111_1111111111111111_1110111010101011_1010010110001010"; -- -0.0676933801748579
	pesos_i(6601) := b"0000000000000000_0000000000000000_0001111110011101_1010110100000001"; -- 0.12349969166438719
	pesos_i(6602) := b"1111111111111111_1111111111111111_1111101111001101_0110011010001011"; -- -0.01639708622550295
	pesos_i(6603) := b"0000000000000000_0000000000000000_0001000110001111_0000010011011001"; -- 0.06858854581847428
	pesos_i(6604) := b"1111111111111111_1111111111111111_1101001111111000_1011000100000101"; -- -0.17198651918549313
	pesos_i(6605) := b"1111111111111111_1111111111111111_1101101110100111_1010011001110001"; -- -0.14197311153178332
	pesos_i(6606) := b"0000000000000000_0000000000000000_0001011011111111_1101010111010101"; -- 0.08984123661769743
	pesos_i(6607) := b"0000000000000000_0000000000000000_0000010011111001_0011000101101110"; -- 0.01942738478716145
	pesos_i(6608) := b"1111111111111111_1111111111111111_1101101010101001_1100100101001110"; -- -0.14584676592791904
	pesos_i(6609) := b"1111111111111111_1111111111111111_1101110011100100_1011010101010001"; -- -0.13713518869949873
	pesos_i(6610) := b"0000000000000000_0000000000000000_0001111100000000_0111000000010000"; -- 0.12110042936756944
	pesos_i(6611) := b"0000000000000000_0000000000000000_0001011001100110_0101011111000010"; -- 0.08749912715777787
	pesos_i(6612) := b"1111111111111111_1111111111111111_1111011110001010_1011111111001000"; -- -0.03303910605286467
	pesos_i(6613) := b"1111111111111111_1111111111111111_1111101101110001_1100000101010110"; -- -0.01779548312432311
	pesos_i(6614) := b"1111111111111111_1111111111111111_1110111110110011_0111010000000100"; -- -0.06366801169456768
	pesos_i(6615) := b"1111111111111111_1111111111111111_1111010100100001_0100110110000000"; -- -0.042460590577934165
	pesos_i(6616) := b"1111111111111111_1111111111111111_1111110011110011_0010101111101110"; -- -0.011914495915273889
	pesos_i(6617) := b"1111111111111111_1111111111111111_1110011111110110_0001100000101111"; -- -0.09390114643918736
	pesos_i(6618) := b"0000000000000000_0000000000000000_0010011011000111_0101001101011000"; -- 0.1514789667862237
	pesos_i(6619) := b"0000000000000000_0000000000000000_0001000110100100_0101010011101110"; -- 0.06891375353797506
	pesos_i(6620) := b"1111111111111111_1111111111111111_1101011001010100_1100000111010001"; -- -0.16276920937693115
	pesos_i(6621) := b"1111111111111111_1111111111111111_1110110010010001_0101110011111001"; -- -0.075906933962917
	pesos_i(6622) := b"0000000000000000_0000000000000000_0000100100110110_1011001000101010"; -- 0.03599084399465907
	pesos_i(6623) := b"1111111111111111_1111111111111111_1111000001011110_1000101011010100"; -- -0.06105739901227476
	pesos_i(6624) := b"0000000000000000_0000000000000000_0000010000001010_0111101100111010"; -- 0.01578493274804252
	pesos_i(6625) := b"1111111111111111_1111111111111111_1110001110101111_0010110111111011"; -- -0.11060822117969604
	pesos_i(6626) := b"0000000000000000_0000000000000000_0000110011001111_1100001010110110"; -- 0.05004517494339513
	pesos_i(6627) := b"0000000000000000_0000000000000000_0000010110101001_0011000111100001"; -- 0.02211295835547614
	pesos_i(6628) := b"0000000000000000_0000000000000000_0001110011101011_0010001010101011"; -- 0.11296288188153994
	pesos_i(6629) := b"0000000000000000_0000000000000000_0010100011001000_0001010010101101"; -- 0.1593029901598606
	pesos_i(6630) := b"0000000000000000_0000000000000000_0010000010110110_1010001010101101"; -- 0.1277867958299482
	pesos_i(6631) := b"1111111111111111_1111111111111111_1101100110100110_1000001000111010"; -- -0.14980302890406927
	pesos_i(6632) := b"1111111111111111_1111111111111111_1111100011000001_1100011111111011"; -- -0.02829313392584032
	pesos_i(6633) := b"0000000000000000_0000000000000000_0000101010111001_0010011110000100"; -- 0.04188773125292154
	pesos_i(6634) := b"1111111111111111_1111111111111111_1110100101000110_0101101100111101"; -- -0.08877019644758831
	pesos_i(6635) := b"0000000000000000_0000000000000000_0000011000110010_0110000001110100"; -- 0.02420618851546356
	pesos_i(6636) := b"1111111111111111_1111111111111111_1110011110111100_1010010101000010"; -- -0.094777747452165
	pesos_i(6637) := b"1111111111111111_1111111111111111_1111000011110111_1100100111001101"; -- -0.058719050945949605
	pesos_i(6638) := b"0000000000000000_0000000000000000_0001100000011010_0011100011110001"; -- 0.09415012252113081
	pesos_i(6639) := b"1111111111111111_1111111111111111_1101100111000011_1100010001011001"; -- -0.14935658283061004
	pesos_i(6640) := b"0000000000000000_0000000000000000_0000100111101100_1001000110011000"; -- 0.03876600239750491
	pesos_i(6641) := b"1111111111111111_1111111111111111_1100101100110010_1010011110010100"; -- -0.20625832221838422
	pesos_i(6642) := b"1111111111111111_1111111111111111_1101110110110001_0001101011101101"; -- -0.13401633937141244
	pesos_i(6643) := b"0000000000000000_0000000000000000_0010100010111000_0000101111111011"; -- 0.15905833118492346
	pesos_i(6644) := b"1111111111111111_1111111111111111_1110011000011101_1000110100010101"; -- -0.10111158597316415
	pesos_i(6645) := b"0000000000000000_0000000000000000_0001001111000111_0110111001011011"; -- 0.07726182661744632
	pesos_i(6646) := b"0000000000000000_0000000000000000_0010100011011010_0111101010111100"; -- 0.1595837314901221
	pesos_i(6647) := b"0000000000000000_0000000000000000_0000001010000111_0010001000000010"; -- 0.009874463623228509
	pesos_i(6648) := b"0000000000000000_0000000000000000_0000001000001110_0101110011111100"; -- 0.008031665314395309
	pesos_i(6649) := b"1111111111111111_1111111111111111_1111000100100111_0001010010100110"; -- -0.057997426532116654
	pesos_i(6650) := b"0000000000000000_0000000000000000_0001001110100001_0010100010000001"; -- 0.0766778293401718
	pesos_i(6651) := b"0000000000000000_0000000000000000_0001010010001001_0001111011001001"; -- 0.08021728911106904
	pesos_i(6652) := b"0000000000000000_0000000000000000_0000111100110011_1011011111001000"; -- 0.059382902459156374
	pesos_i(6653) := b"1111111111111111_1111111111111111_1111011001111000_1110100100001010"; -- -0.03721755499829078
	pesos_i(6654) := b"1111111111111111_1111111111111111_1101111101010111_1100110100010000"; -- -0.12756651258457094
	pesos_i(6655) := b"0000000000000000_0000000000000000_0001001101111001_1101111010110011"; -- 0.07607833739037329
	pesos_i(6656) := b"1111111111111111_1111111111111111_1101100100111111_0110010000100111"; -- -0.15137647668714133
	pesos_i(6657) := b"1111111111111111_1111111111111111_1111111000001110_0111001100101101"; -- -0.007592011892951164
	pesos_i(6658) := b"1111111111111111_1111111111111111_1110011110010100_0000000001110000"; -- -0.09539792321749191
	pesos_i(6659) := b"1111111111111111_1111111111111111_1110100001001110_1010000111110110"; -- -0.09255016073423325
	pesos_i(6660) := b"1111111111111111_1111111111111111_1111011011111011_1010100001000100"; -- -0.0352225144836761
	pesos_i(6661) := b"0000000000000000_0000000000000000_0000100000001100_1011111010011001"; -- 0.03144446602456237
	pesos_i(6662) := b"1111111111111111_1111111111111111_1111001100011111_1111001111000000"; -- -0.0502936988854327
	pesos_i(6663) := b"0000000000000000_0000000000000000_0001100011000111_0001100001000110"; -- 0.09678794584806923
	pesos_i(6664) := b"1111111111111111_1111111111111111_1110000111011011_1010010010111010"; -- -0.11774225678888726
	pesos_i(6665) := b"0000000000000000_0000000000000000_0001001101110001_0000111010011011"; -- 0.07594386362632419
	pesos_i(6666) := b"1111111111111111_1111111111111111_1110010100001101_1001000011100101"; -- -0.10526174936175976
	pesos_i(6667) := b"1111111111111111_1111111111111111_1101010110011010_1111000110010111"; -- -0.16560449652196058
	pesos_i(6668) := b"1111111111111111_1111111111111111_1111110110111101_1010111001111001"; -- -0.008824439516469409
	pesos_i(6669) := b"0000000000000000_0000000000000000_0001100111001010_0101001111000011"; -- 0.10074351793358073
	pesos_i(6670) := b"0000000000000000_0000000000000000_0000000011101010_1001111101100111"; -- 0.0035800578451646733
	pesos_i(6671) := b"1111111111111111_1111111111111111_1101110010010000_1011011000011000"; -- -0.13841688066163835
	pesos_i(6672) := b"1111111111111111_1111111111111111_1101001110101000_1101011111101000"; -- -0.17320490442091255
	pesos_i(6673) := b"1111111111111111_1111111111111111_1111111010101000_0111101000111111"; -- -0.005241737070052162
	pesos_i(6674) := b"1111111111111111_1111111111111111_1101110110010110_1010011011011101"; -- -0.13441998589159526
	pesos_i(6675) := b"1111111111111111_1111111111111111_1101110011010100_0110000011010100"; -- -0.1373843653980417
	pesos_i(6676) := b"0000000000000000_0000000000000000_0010011011110000_1000011100101001"; -- 0.15210766558823177
	pesos_i(6677) := b"0000000000000000_0000000000000000_0010100010101010_1101110000001000"; -- 0.15885710903837483
	pesos_i(6678) := b"0000000000000000_0000000000000000_0000101001001011_0011011110011000"; -- 0.04021022274405808
	pesos_i(6679) := b"0000000000000000_0000000000000000_0011000011100100_1100010111110000"; -- 0.19099080196779433
	pesos_i(6680) := b"0000000000000000_0000000000000000_0001010111001011_0110100111000010"; -- 0.08513508780027647
	pesos_i(6681) := b"0000000000000000_0000000000000000_0001110100100100_0001000010110010"; -- 0.11383156147223027
	pesos_i(6682) := b"1111111111111111_1111111111111111_1110010111010001_1011000010101011"; -- -0.10226913296935364
	pesos_i(6683) := b"1111111111111111_1111111111111111_1110100001111100_0110010000000010"; -- -0.09185194922786491
	pesos_i(6684) := b"0000000000000000_0000000000000000_0010101000111001_1110110000010010"; -- 0.16494632176587173
	pesos_i(6685) := b"0000000000000000_0000000000000000_0000001110110000_1111111110000011"; -- 0.014419526516484866
	pesos_i(6686) := b"1111111111111111_1111111111111111_1111000011101101_1010011100011111"; -- -0.05887370588864171
	pesos_i(6687) := b"1111111111111111_1111111111111111_1111001010000101_1101101110100110"; -- -0.05264498892231291
	pesos_i(6688) := b"1111111111111111_1111111111111111_1111000000101101_1100000111101010"; -- -0.06180179636058676
	pesos_i(6689) := b"1111111111111111_1111111111111111_1111001110111101_0100011110011000"; -- -0.047893071592724656
	pesos_i(6690) := b"1111111111111111_1111111111111111_1111110111101010_1001000110101101"; -- -0.008139510504615324
	pesos_i(6691) := b"1111111111111111_1111111111111111_1110001000011010_0101100001010111"; -- -0.11678550600250004
	pesos_i(6692) := b"1111111111111111_1111111111111111_1111100101110001_0110011001101100"; -- -0.02561340192537499
	pesos_i(6693) := b"1111111111111111_1111111111111111_1111111001010010_0101011100001101"; -- -0.006556090705308057
	pesos_i(6694) := b"1111111111111111_1111111111111111_1111000110010111_1101010110010110"; -- -0.05627694223629915
	pesos_i(6695) := b"1111111111111111_1111111111111111_1101101111111011_1010111000001011"; -- -0.14069092006445166
	pesos_i(6696) := b"1111111111111111_1111111111111111_1111111000000110_1011100101010010"; -- -0.007709901243639544
	pesos_i(6697) := b"0000000000000000_0000000000000000_0000101010111011_1001100011011100"; -- 0.04192500468700763
	pesos_i(6698) := b"0000000000000000_0000000000000000_0001110011100001_0000101001010110"; -- 0.11280884350411999
	pesos_i(6699) := b"0000000000000000_0000000000000000_0001101001000111_0101101001010010"; -- 0.10265125743288453
	pesos_i(6700) := b"1111111111111111_1111111111111111_1110010001110110_1001010110110000"; -- -0.10756554092292453
	pesos_i(6701) := b"0000000000000000_0000000000000000_0000101011111111_0110101111010000"; -- 0.04295991725849829
	pesos_i(6702) := b"0000000000000000_0000000000000000_0010010110011110_0101110100010001"; -- 0.1469476859682334
	pesos_i(6703) := b"0000000000000000_0000000000000000_0001101101000000_0110001001001001"; -- 0.10645117075498618
	pesos_i(6704) := b"0000000000000000_0000000000000000_0010110000101001_1011101111110101"; -- 0.17251181345017544
	pesos_i(6705) := b"0000000000000000_0000000000000000_0010010001101011_1100101100110110"; -- 0.14226980265212702
	pesos_i(6706) := b"0000000000000000_0000000000000000_0001100100011100_0110010111001111"; -- 0.09808956424490176
	pesos_i(6707) := b"1111111111111111_1111111111111111_1111110111100101_1001001010000100"; -- -0.008215754375654853
	pesos_i(6708) := b"1111111111111111_1111111111111111_1110111101100000_0100010001001011"; -- -0.0649373357418944
	pesos_i(6709) := b"0000000000000000_0000000000000000_0001011000001111_0100010010110101"; -- 0.0861704770470908
	pesos_i(6710) := b"1111111111111111_1111111111111111_1101101100010001_1011111111001000"; -- -0.14426041953692895
	pesos_i(6711) := b"0000000000000000_0000000000000000_0000110000111001_0111000001101000"; -- 0.04775145088143702
	pesos_i(6712) := b"1111111111111111_1111111111111111_1101101000011100_1001110111100010"; -- -0.1480008432466902
	pesos_i(6713) := b"1111111111111111_1111111111111111_1101011000010110_0010000110111100"; -- -0.16372479596153913
	pesos_i(6714) := b"1111111111111111_1111111111111111_1111111011010110_0000010110111001"; -- -0.004546778074912395
	pesos_i(6715) := b"0000000000000000_0000000000000000_0001000101100001_1001110111000111"; -- 0.06789575669877859
	pesos_i(6716) := b"1111111111111111_1111111111111111_1101100100011100_1011010100001111"; -- -0.15190571189000598
	pesos_i(6717) := b"0000000000000000_0000000000000000_0001100011000110_0010000011001010"; -- 0.09677319465234982
	pesos_i(6718) := b"0000000000000000_0000000000000000_0001001101001010_1001010001011101"; -- 0.07535674361233918
	pesos_i(6719) := b"1111111111111111_1111111111111111_1101110010000111_0011001011101001"; -- -0.13856202889587396
	pesos_i(6720) := b"1111111111111111_1111111111111111_1101111101110110_1110001000101001"; -- -0.12709223277158208
	pesos_i(6721) := b"1111111111111111_1111111111111111_1110000011000101_1100011001111110"; -- -0.12198218757917412
	pesos_i(6722) := b"0000000000000000_0000000000000000_0001010000000101_1101111111100111"; -- 0.07821463968063345
	pesos_i(6723) := b"0000000000000000_0000000000000000_0001110000111000_0011000101101010"; -- 0.11023243750083916
	pesos_i(6724) := b"1111111111111111_1111111111111111_1110011110100111_1111001010111111"; -- -0.09509356350141897
	pesos_i(6725) := b"1111111111111111_1111111111111111_1111011100011110_0001111010100010"; -- -0.034696660386404087
	pesos_i(6726) := b"0000000000000000_0000000000000000_0001011011101100_0101001110101011"; -- 0.08954356117558351
	pesos_i(6727) := b"1111111111111111_1111111111111111_1101111100001111_1111100000000001"; -- -0.12866258604667694
	pesos_i(6728) := b"1111111111111111_1111111111111111_1101100110110110_1111101101110000"; -- -0.14955166353164234
	pesos_i(6729) := b"0000000000000000_0000000000000000_0010101011001000_1111010100111010"; -- 0.16712887440020105
	pesos_i(6730) := b"1111111111111111_1111111111111111_1101101101001011_0100110101101101"; -- -0.14338222589322674
	pesos_i(6731) := b"1111111111111111_1111111111111111_1101011011000000_1001110010010100"; -- -0.16112347963721654
	pesos_i(6732) := b"0000000000000000_0000000000000000_0010001110110110_0100000111011100"; -- 0.13949977520785434
	pesos_i(6733) := b"1111111111111111_1111111111111111_1110011010010000_0110011111001001"; -- -0.09935904821004868
	pesos_i(6734) := b"0000000000000000_0000000000000000_0001101111111101_0101100100110010"; -- 0.10933453997618892
	pesos_i(6735) := b"1111111111111111_1111111111111111_1110111001111001_0010110110111010"; -- -0.06846346093984003
	pesos_i(6736) := b"1111111111111111_1111111111111111_1110000111110001_0101010011111001"; -- -0.11741131707764701
	pesos_i(6737) := b"0000000000000000_0000000000000000_0001000101010011_1000111000010010"; -- 0.06768119759063887
	pesos_i(6738) := b"0000000000000000_0000000000000000_0010011100000010_0100001010111001"; -- 0.15237824460678245
	pesos_i(6739) := b"0000000000000000_0000000000000000_0001000011001101_0000000110110011"; -- 0.06562815300624063
	pesos_i(6740) := b"1111111111111111_1111111111111111_1111100101110001_1011011010000100"; -- -0.025608628141764633
	pesos_i(6741) := b"0000000000000000_0000000000000000_0000000101100111_0101000110101111"; -- 0.005482773974058436
	pesos_i(6742) := b"1111111111111111_1111111111111111_1101100100111001_1000010001111111"; -- -0.15146610166585156
	pesos_i(6743) := b"0000000000000000_0000000000000000_0001000000100001_0111100011111110"; -- 0.06301075168614145
	pesos_i(6744) := b"0000000000000000_0000000000000000_0010111101001111_1111101001000100"; -- 0.18481411125556918
	pesos_i(6745) := b"0000000000000000_0000000000000000_0001100011101001_1101101110001101"; -- 0.09731838403982
	pesos_i(6746) := b"1111111111111111_1111111111111111_1110110111000010_0100010100111111"; -- -0.0712544176051487
	pesos_i(6747) := b"1111111111111111_1111111111111111_1101000100001001_1111001111001100"; -- -0.1834418895801796
	pesos_i(6748) := b"1111111111111111_1111111111111111_1110010010100101_1100101010011100"; -- -0.10684522326374002
	pesos_i(6749) := b"0000000000000000_0000000000000000_0000111111011001_1001001100101010"; -- 0.061913678827579546
	pesos_i(6750) := b"1111111111111111_1111111111111111_1110010110010010_0010100001110101"; -- -0.10323855538458815
	pesos_i(6751) := b"1111111111111111_1111111111111111_1110011011111001_1010110011001110"; -- -0.09775276145189207
	pesos_i(6752) := b"0000000000000000_0000000000000000_0001000110010011_0010011110101001"; -- 0.06865165580604263
	pesos_i(6753) := b"0000000000000000_0000000000000000_0010110011101011_0110111101010010"; -- 0.17546745058426322
	pesos_i(6754) := b"0000000000000000_0000000000000000_0001001110000000_1001101000000000"; -- 0.07618105422613207
	pesos_i(6755) := b"0000000000000000_0000000000000000_0000010011010100_1011001101111110"; -- 0.018870561763168738
	pesos_i(6756) := b"0000000000000000_0000000000000000_0001011010100001_1101111110111101"; -- 0.08840750080373581
	pesos_i(6757) := b"1111111111111111_1111111111111111_1101010101100001_0010101100110111"; -- -0.16648607169323845
	pesos_i(6758) := b"0000000000000000_0000000000000000_0010111010110110_0011100000011001"; -- 0.18246794329461336
	pesos_i(6759) := b"0000000000000000_0000000000000000_0010101101101101_1011100101101010"; -- 0.16964300952122777
	pesos_i(6760) := b"1111111111111111_1111111111111111_1111110111000110_0111100101000001"; -- -0.008690282396558308
	pesos_i(6761) := b"0000000000000000_0000000000000000_0000101000001001_0111010001000011"; -- 0.03920675875939902
	pesos_i(6762) := b"0000000000000000_0000000000000000_0000101011000011_0011001110010001"; -- 0.04204103740930891
	pesos_i(6763) := b"0000000000000000_0000000000000000_0010000100010110_1100100010101001"; -- 0.12925390369098755
	pesos_i(6764) := b"0000000000000000_0000000000000000_0000000110100111_1011011001001010"; -- 0.006465333084274026
	pesos_i(6765) := b"0000000000000000_0000000000000000_0000111000101000_0010001101111100"; -- 0.05529996667680931
	pesos_i(6766) := b"1111111111111111_1111111111111111_1110010000100000_0000010101011000"; -- -0.10888640013436388
	pesos_i(6767) := b"0000000000000000_0000000000000000_0010111000110010_0000110111110000"; -- 0.18045127010741452
	pesos_i(6768) := b"0000000000000000_0000000000000000_0000010010100000_0001100010000010"; -- 0.01806786702273297
	pesos_i(6769) := b"0000000000000000_0000000000000000_0000101100010111_0110111100101110"; -- 0.043326329000001926
	pesos_i(6770) := b"1111111111111111_1111111111111111_1110110011100111_1001110111111100"; -- -0.07459080322949635
	pesos_i(6771) := b"1111111111111111_1111111111111111_1111011000001100_1011000110000000"; -- -0.03886881478468016
	pesos_i(6772) := b"1111111111111111_1111111111111111_1101110011100110_1011001001101110"; -- -0.1371048433024575
	pesos_i(6773) := b"0000000000000000_0000000000000000_0001110101101001_0111110101001111"; -- 0.11489089174382308
	pesos_i(6774) := b"0000000000000000_0000000000000000_0000000110001110_1011011011101100"; -- 0.0060839010761475215
	pesos_i(6775) := b"1111111111111111_1111111111111111_1101111110111111_0010111000111111"; -- -0.12598906469144733
	pesos_i(6776) := b"0000000000000000_0000000000000000_0000100101000000_0011100110010101"; -- 0.03613624455874473
	pesos_i(6777) := b"0000000000000000_0000000000000000_0000000111101100_0111101001101100"; -- 0.007514621031605422
	pesos_i(6778) := b"1111111111111111_1111111111111111_1110011001100100_0010000110110011"; -- -0.10003461240022588
	pesos_i(6779) := b"0000000000000000_0000000000000000_0000010001001001_1000010111110111"; -- 0.016746876590213098
	pesos_i(6780) := b"0000000000000000_0000000000000000_0010100001010100_0001110000110001"; -- 0.15753341850774355
	pesos_i(6781) := b"1111111111111111_1111111111111111_1110111000110011_1100101010010011"; -- -0.0695222274713111
	pesos_i(6782) := b"1111111111111111_1111111111111111_1111111001100010_1010111010110110"; -- -0.006306725125646026
	pesos_i(6783) := b"0000000000000000_0000000000000000_0000001001000010_0101110111011000"; -- 0.008825173488242983
	pesos_i(6784) := b"1111111111111111_1111111111111111_1101110000111101_1000111010001110"; -- -0.13968571686050016
	pesos_i(6785) := b"1111111111111111_1111111111111111_1110001000001000_0001101101011010"; -- -0.11706379933578247
	pesos_i(6786) := b"0000000000000000_0000000000000000_0001111110001111_1000111110110100"; -- 0.12328432209954815
	pesos_i(6787) := b"0000000000000000_0000000000000000_0010100011110000_1010000010011101"; -- 0.15992168268241413
	pesos_i(6788) := b"1111111111111111_1111111111111111_1111101101111100_0101001110010101"; -- -0.017634178199923783
	pesos_i(6789) := b"0000000000000000_0000000000000000_0001111111010010_0100100110000001"; -- 0.12430247690100636
	pesos_i(6790) := b"0000000000000000_0000000000000000_0000010110000101_0111100000111011"; -- 0.021567835250325903
	pesos_i(6791) := b"1111111111111111_1111111111111111_1110111101011000_0000101101010110"; -- -0.06506280096467065
	pesos_i(6792) := b"1111111111111111_1111111111111111_1110100101011100_1101010011010100"; -- -0.08842725584578014
	pesos_i(6793) := b"0000000000000000_0000000000000000_0000111001101111_1110110000100001"; -- 0.056395299869759496
	pesos_i(6794) := b"1111111111111111_1111111111111111_1101110111011101_1101001000100111"; -- -0.13333403152266177
	pesos_i(6795) := b"0000000000000000_0000000000000000_0000111111000010_0010100000011101"; -- 0.06155634604686321
	pesos_i(6796) := b"0000000000000000_0000000000000000_0000010011111110_1100000100011000"; -- 0.01951224164248263
	pesos_i(6797) := b"1111111111111111_1111111111111111_1110100101110100_1011011010010111"; -- -0.0880628472434852
	pesos_i(6798) := b"1111111111111111_1111111111111111_1101110001101110_1010010011100001"; -- -0.1389367056196197
	pesos_i(6799) := b"1111111111111111_1111111111111111_1101111101011010_0010011000111111"; -- -0.12753067942772345
	pesos_i(6800) := b"1111111111111111_1111111111111111_1101110110110010_0010101011000010"; -- -0.13400013697468044
	pesos_i(6801) := b"0000000000000000_0000000000000000_0001000101101100_1101000010001000"; -- 0.06806662869430809
	pesos_i(6802) := b"0000000000000000_0000000000000000_0001100010001000_1101101110111100"; -- 0.09583829253242766
	pesos_i(6803) := b"1111111111111111_1111111111111111_1111010111001111_0010010011101100"; -- -0.039807979945373585
	pesos_i(6804) := b"1111111111111111_1111111111111111_1110010011110001_1101011100000001"; -- -0.10568481656005094
	pesos_i(6805) := b"0000000000000000_0000000000000000_0001111101100001_1100011010100100"; -- 0.12258569241051881
	pesos_i(6806) := b"0000000000000000_0000000000000000_0001001000000000_1000110101010110"; -- 0.07032092424522396
	pesos_i(6807) := b"0000000000000000_0000000000000000_0010011010001001_1100000011001011"; -- 0.15053944556978233
	pesos_i(6808) := b"1111111111111111_1111111111111111_1101111111101010_0111010001000001"; -- -0.1253287640891649
	pesos_i(6809) := b"0000000000000000_0000000000000000_0010011011101110_1001111011001010"; -- 0.15207855631438413
	pesos_i(6810) := b"1111111111111111_1111111111111111_1110011001001100_0111101001001111"; -- -0.10039554188659945
	pesos_i(6811) := b"1111111111111111_1111111111111111_1111101001010110_0000101000110101"; -- -0.02212463565228928
	pesos_i(6812) := b"1111111111111111_1111111111111111_1101100111111100_0011101010101100"; -- -0.14849503806448427
	pesos_i(6813) := b"1111111111111111_1111111111111111_1110001000011101_0011110101101100"; -- -0.11674133408439193
	pesos_i(6814) := b"0000000000000000_0000000000000000_0000010001001111_0110111000110001"; -- 0.01683701235841655
	pesos_i(6815) := b"1111111111111111_1111111111111111_1111111000111001_0100110110101011"; -- -0.006938119697731532
	pesos_i(6816) := b"0000000000000000_0000000000000000_0000000110010001_0100110111010100"; -- 0.006123413366740854
	pesos_i(6817) := b"0000000000000000_0000000000000000_0001000011010010_1000111111100000"; -- 0.06571292125072875
	pesos_i(6818) := b"0000000000000000_0000000000000000_0010101110010011_1101111110101101"; -- 0.17022512405468038
	pesos_i(6819) := b"1111111111111111_1111111111111111_1111100100011001_0000010100001101"; -- -0.026961979272758296
	pesos_i(6820) := b"0000000000000000_0000000000000000_0000011111010011_0101000111110101"; -- 0.03056823951182446
	pesos_i(6821) := b"0000000000000000_0000000000000000_0000001011001011_1111111110001001"; -- 0.010925265318196806
	pesos_i(6822) := b"0000000000000000_0000000000000000_0000000010010110_1000011110111000"; -- 0.002296907847382517
	pesos_i(6823) := b"0000000000000000_0000000000000000_0010000110010010_1000011010101101"; -- 0.13114206060256847
	pesos_i(6824) := b"0000000000000000_0000000000000000_0001010111100110_0000001010000011"; -- 0.08554092126241783
	pesos_i(6825) := b"1111111111111111_1111111111111111_1111101000011100_1010110111111011"; -- -0.022999883775736224
	pesos_i(6826) := b"1111111111111111_1111111111111111_1101010111000111_0111000111001011"; -- -0.1649254682967765
	pesos_i(6827) := b"1111111111111111_1111111111111111_1110001010010100_0001101110110000"; -- -0.1149275490138554
	pesos_i(6828) := b"1111111111111111_1111111111111111_1110111101101011_0111011000001000"; -- -0.06476652439606244
	pesos_i(6829) := b"0000000000000000_0000000000000000_0010001101011101_1010110101100101"; -- 0.13814815253777007
	pesos_i(6830) := b"0000000000000000_0000000000000000_0000011110110111_1110010010111101"; -- 0.030149742190950103
	pesos_i(6831) := b"0000000000000000_0000000000000000_0001101100111001_0011001011100001"; -- 0.10634153351669715
	pesos_i(6832) := b"0000000000000000_0000000000000000_0000000000001110_1001010100100110"; -- 0.00022251294645031505
	pesos_i(6833) := b"0000000000000000_0000000000000000_0010010111010000_1100100111010001"; -- 0.14771710733105994
	pesos_i(6834) := b"1111111111111111_1111111111111111_1101101100100100_0100000100110111"; -- -0.14397804641810982
	pesos_i(6835) := b"0000000000000000_0000000000000000_0010010101111100_0111111110000101"; -- 0.14643094063528578
	pesos_i(6836) := b"0000000000000000_0000000000000000_0001110110101000_0100010110001111"; -- 0.11584887259117255
	pesos_i(6837) := b"0000000000000000_0000000000000000_0010010100110101_0011010100010001"; -- 0.14534312876883582
	pesos_i(6838) := b"0000000000000000_0000000000000000_0001001000101100_0100000101010111"; -- 0.07098778118900084
	pesos_i(6839) := b"1111111111111111_1111111111111111_1101110001111001_1000001010100110"; -- -0.1387708992692967
	pesos_i(6840) := b"1111111111111111_1111111111111111_1110010010110110_1000100000111100"; -- -0.1065897801398084
	pesos_i(6841) := b"1111111111111111_1111111111111111_1110110100011100_0011011101000111"; -- -0.0737882091283254
	pesos_i(6842) := b"0000000000000000_0000000000000000_0001111011100000_0011001100010100"; -- 0.1206085133084835
	pesos_i(6843) := b"1111111111111111_1111111111111111_1101100001101100_1010111000011111"; -- -0.15459167231872395
	pesos_i(6844) := b"0000000000000000_0000000000000000_0000111010111001_1100011111001011"; -- 0.05752228466518758
	pesos_i(6845) := b"0000000000000000_0000000000000000_0001101100000100_0001100110100111"; -- 0.105531314176382
	pesos_i(6846) := b"1111111111111111_1111111111111111_1101110010100010_0001101100101100"; -- -0.1381514566228378
	pesos_i(6847) := b"1111111111111111_1111111111111111_1110001100011010_1111110001111101"; -- -0.11286947194763502
	pesos_i(6848) := b"0000000000000000_0000000000000000_0000101010011111_0111101001100000"; -- 0.04149594159267336
	pesos_i(6849) := b"1111111111111111_1111111111111111_1101110010001110_1100110000010110"; -- -0.13844608743097944
	pesos_i(6850) := b"0000000000000000_0000000000000000_0010010100010111_1101101001110111"; -- 0.14489522364183594
	pesos_i(6851) := b"0000000000000000_0000000000000000_0000000111001101_1010000000011111"; -- 0.007043845792144663
	pesos_i(6852) := b"0000000000000000_0000000000000000_0000100000110110_1011101111110001"; -- 0.03208517673786275
	pesos_i(6853) := b"1111111111111111_1111111111111111_1111001100111011_1000100010001000"; -- -0.04987284351338679
	pesos_i(6854) := b"1111111111111111_1111111111111111_1111110111000100_0101001010110100"; -- -0.00872309776277269
	pesos_i(6855) := b"1111111111111111_1111111111111111_1101001001111110_0010100100001111"; -- -0.1777624453341697
	pesos_i(6856) := b"1111111111111111_1111111111111111_1111011100011101_0110110101001011"; -- -0.034707230763527955
	pesos_i(6857) := b"1111111111111111_1111111111111111_1101111100010010_1001011100010001"; -- -0.12862258748768768
	pesos_i(6858) := b"0000000000000000_0000000000000000_0010000010001010_1110011101010110"; -- 0.1271195015395365
	pesos_i(6859) := b"1111111111111111_1111111111111111_1111101001110010_0110111100111101"; -- -0.02169136765963341
	pesos_i(6860) := b"0000000000000000_0000000000000000_0010000111110110_0011100101001000"; -- 0.13266332625535482
	pesos_i(6861) := b"1111111111111111_1111111111111111_1111101000111100_1001011001111011"; -- -0.022513003258901366
	pesos_i(6862) := b"1111111111111111_1111111111111111_1111000010000010_0010011111100100"; -- -0.060513979712010744
	pesos_i(6863) := b"0000000000000000_0000000000000000_0010010100111100_0111010100000111"; -- 0.14545375265132587
	pesos_i(6864) := b"1111111111111111_1111111111111111_1111110010000010_0001101010111010"; -- -0.013639764421660011
	pesos_i(6865) := b"1111111111111111_1111111111111111_1110110011000110_1111011010010111"; -- -0.07508906190153236
	pesos_i(6866) := b"1111111111111111_1111111111111111_1110111111010110_0111001000001111"; -- -0.06313407065192517
	pesos_i(6867) := b"0000000000000000_0000000000000000_0001000001111111_1010110010100100"; -- 0.06444815637533802
	pesos_i(6868) := b"0000000000000000_0000000000000000_0001101100000010_0111111100110110"; -- 0.10550684997738355
	pesos_i(6869) := b"0000000000000000_0000000000000000_0001101000010011_0000101111010010"; -- 0.10185312159370416
	pesos_i(6870) := b"0000000000000000_0000000000000000_0000101001110111_0001011000111111"; -- 0.04087962192924777
	pesos_i(6871) := b"0000000000000000_0000000000000000_0000011100001111_1011000110110100"; -- 0.02758322366639806
	pesos_i(6872) := b"0000000000000000_0000000000000000_0011001010000010_0110001111001111"; -- 0.19730209155306444
	pesos_i(6873) := b"0000000000000000_0000000000000000_0011001101111011_0111010110111111"; -- 0.20110259937115504
	pesos_i(6874) := b"1111111111111111_1111111111111111_1101011110100111_0011000011101101"; -- -0.1576051161158345
	pesos_i(6875) := b"1111111111111111_1111111111111111_1110000011000011_0011100111000100"; -- -0.12202109312690519
	pesos_i(6876) := b"1111111111111111_1111111111111111_1110001000110000_1011101111001111"; -- -0.11644388394478704
	pesos_i(6877) := b"1111111111111111_1111111111111111_1101011001111001_1101111000110100"; -- -0.16220294211160874
	pesos_i(6878) := b"1111111111111111_1111111111111111_1101011110111011_1110100010111101"; -- -0.15728898425553817
	pesos_i(6879) := b"1111111111111111_1111111111111111_1111101000110100_0100110010100000"; -- -0.02263947566766114
	pesos_i(6880) := b"1111111111111111_1111111111111111_1111001100010010_1100110001101100"; -- -0.050494407303905364
	pesos_i(6881) := b"1111111111111111_1111111111111111_1111000101011000_0001001101001010"; -- -0.057249826738400504
	pesos_i(6882) := b"0000000000000000_0000000000000000_0000100010101000_0011000011100100"; -- 0.03381639064450289
	pesos_i(6883) := b"1111111111111111_1111111111111111_1110010011100110_1111001100011011"; -- -0.1058509882905144
	pesos_i(6884) := b"0000000000000000_0000000000000000_0001110010111010_0100011100100100"; -- 0.11221737506134034
	pesos_i(6885) := b"1111111111111111_1111111111111111_1101001110010001_1101110010001111"; -- -0.17355557916029785
	pesos_i(6886) := b"1111111111111111_1111111111111111_1110101011000110_1001100010101001"; -- -0.08290716043389336
	pesos_i(6887) := b"0000000000000000_0000000000000000_0001010011010010_0011110110010100"; -- 0.08133301598476553
	pesos_i(6888) := b"1111111111111111_1111111111111111_1101001101101001_0010100011000100"; -- -0.1741766472620272
	pesos_i(6889) := b"0000000000000000_0000000000000000_0001100000110010_0001111011001000"; -- 0.09451477411402628
	pesos_i(6890) := b"0000000000000000_0000000000000000_0001110100101100_0111111011110000"; -- 0.11396020285039399
	pesos_i(6891) := b"1111111111111111_1111111111111111_1111100000111001_0111001100011011"; -- -0.03037338817880837
	pesos_i(6892) := b"1111111111111111_1111111111111111_1111010100011100_0010001001000010"; -- -0.042539461978915206
	pesos_i(6893) := b"0000000000000000_0000000000000000_0000010001110111_0101111110101110"; -- 0.017446498937589077
	pesos_i(6894) := b"1111111111111111_1111111111111111_1110000111100000_0100001111010110"; -- -0.11767173784786637
	pesos_i(6895) := b"0000000000000000_0000000000000000_0000000100100001_0011010011010011"; -- 0.0044129385270216094
	pesos_i(6896) := b"1111111111111111_1111111111111111_1101101001001111_1111011000100001"; -- -0.14721738527949266
	pesos_i(6897) := b"1111111111111111_1111111111111111_1110001111010110_1000111010100001"; -- -0.11000736787137794
	pesos_i(6898) := b"1111111111111111_1111111111111111_1101001010110100_0010101100100011"; -- -0.17693834674791561
	pesos_i(6899) := b"0000000000000000_0000000000000000_0001111100111000_0100001001100011"; -- 0.12195219923812024
	pesos_i(6900) := b"1111111111111111_1111111111111111_1111000100010001_1001010110111011"; -- -0.05832542596834642
	pesos_i(6901) := b"1111111111111111_1111111111111111_1111111001011100_0000000101110110"; -- -0.0064086042676482985
	pesos_i(6902) := b"1111111111111111_1111111111111111_1101101000010001_0111000011111000"; -- -0.14817136707913672
	pesos_i(6903) := b"1111111111111111_1111111111111111_1111101001110100_0011110101001101"; -- -0.021663826688115683
	pesos_i(6904) := b"1111111111111111_1111111111111111_1111111110110000_0010101111101110"; -- -0.0012180847378538695
	pesos_i(6905) := b"1111111111111111_1111111111111111_1111011010010011_0001000000011110"; -- -0.03681849731396086
	pesos_i(6906) := b"0000000000000000_0000000000000000_0010100110011000_0100100110011010"; -- 0.1624799730283027
	pesos_i(6907) := b"0000000000000000_0000000000000000_0010110000000100_1101101001000010"; -- 0.17194904445187387
	pesos_i(6908) := b"1111111111111111_1111111111111111_1111111011011001_1001010001000101"; -- -0.004492505263395423
	pesos_i(6909) := b"0000000000000000_0000000000000000_0001101110110010_0100001000010010"; -- 0.10818875254922987
	pesos_i(6910) := b"1111111111111111_1111111111111111_1110000010001111_0110001000111100"; -- -0.12281213782659363
	pesos_i(6911) := b"0000000000000000_0000000000000000_0000110101100101_0110000010101111"; -- 0.052328150585552985
	pesos_i(6912) := b"1111111111111111_1111111111111111_1101001111101100_1100100101100111"; -- -0.17216817118205346
	pesos_i(6913) := b"0000000000000000_0000000000000000_0001000001110110_1001100111000001"; -- 0.06430970158539137
	pesos_i(6914) := b"0000000000000000_0000000000000000_0000011011001100_0101111001111100"; -- 0.026555924762251916
	pesos_i(6915) := b"0000000000000000_0000000000000000_0001111101111011_1110101010111110"; -- 0.1229845728601074
	pesos_i(6916) := b"0000000000000000_0000000000000000_0010101101111001_0111010011011101"; -- 0.1698220291049052
	pesos_i(6917) := b"1111111111111111_1111111111111111_1101101010111010_1001110010100110"; -- -0.14559002822120654
	pesos_i(6918) := b"0000000000000000_0000000000000000_0001000111110011_1110100000111000"; -- 0.07012797699593885
	pesos_i(6919) := b"1111111111111111_1111111111111111_1101011010011011_0000110110101110"; -- -0.16169657237698856
	pesos_i(6920) := b"0000000000000000_0000000000000000_0000010010101110_0111011100111100"; -- 0.018287136227750172
	pesos_i(6921) := b"1111111111111111_1111111111111111_1110111010111001_1100101111100111"; -- -0.06747747051314809
	pesos_i(6922) := b"1111111111111111_1111111111111111_1111011010001011_0001011110101111"; -- -0.036940116669603056
	pesos_i(6923) := b"1111111111111111_1111111111111111_1101111001001010_1110001101000011"; -- -0.13166980378782742
	pesos_i(6924) := b"1111111111111111_1111111111111111_1110010000110000_0110001000010101"; -- -0.10863673189220444
	pesos_i(6925) := b"1111111111111111_1111111111111111_1111011111110001_1100000000000001"; -- -0.031467437574729196
	pesos_i(6926) := b"0000000000000000_0000000000000000_0000011101111110_0001001001001100"; -- 0.02926744788881113
	pesos_i(6927) := b"1111111111111111_1111111111111111_1111111101111111_1000001110000110"; -- -0.0019605443680432155
	pesos_i(6928) := b"1111111111111111_1111111111111111_1110101001100011_1101100011010011"; -- -0.08441395607674966
	pesos_i(6929) := b"1111111111111111_1111111111111111_1101000101101001_1011101011001001"; -- -0.18198044387987822
	pesos_i(6930) := b"0000000000000000_0000000000000000_0000011011011001_0111110101001110"; -- 0.02675612587497329
	pesos_i(6931) := b"0000000000000000_0000000000000000_0000011000001001_0011111011010110"; -- 0.023578574457250017
	pesos_i(6932) := b"1111111111111111_1111111111111111_1111010111001100_0000101111010001"; -- -0.039855252634149095
	pesos_i(6933) := b"1111111111111111_1111111111111111_1101100000001000_0001110011110011"; -- -0.15612620409207645
	pesos_i(6934) := b"0000000000000000_0000000000000000_0001101000111011_0011101000100001"; -- 0.10246623319759487
	pesos_i(6935) := b"1111111111111111_1111111111111111_1111010111000101_0001111011111011"; -- -0.03996092189219907
	pesos_i(6936) := b"1111111111111111_1111111111111111_1110100001011110_1010100000001100"; -- -0.09230565734515933
	pesos_i(6937) := b"0000000000000000_0000000000000000_0000001110111011_1101100100110001"; -- 0.014585089281625843
	pesos_i(6938) := b"1111111111111111_1111111111111111_1110001110010000_1111001110101000"; -- -0.11106946137253561
	pesos_i(6939) := b"0000000000000000_0000000000000000_0000011011100010_1110101110000001"; -- 0.026900023559140913
	pesos_i(6940) := b"0000000000000000_0000000000000000_0010001010111110_1100000110110001"; -- 0.1357232149311354
	pesos_i(6941) := b"1111111111111111_1111111111111111_1110111000111001_1110110001100011"; -- -0.06942865924884606
	pesos_i(6942) := b"0000000000000000_0000000000000000_0001000101110110_1110001001001001"; -- 0.06822027467557891
	pesos_i(6943) := b"0000000000000000_0000000000000000_0000001000111000_1101011001010110"; -- 0.00867976750938923
	pesos_i(6944) := b"1111111111111111_1111111111111111_1111110011011010_1100000101010110"; -- -0.012287060206423395
	pesos_i(6945) := b"1111111111111111_1111111111111111_1111110110111001_0011011110111011"; -- -0.008892552191299221
	pesos_i(6946) := b"0000000000000000_0000000000000000_0010100111101001_1101101000100101"; -- 0.1637245502567817
	pesos_i(6947) := b"0000000000000000_0000000000000000_0001011100011000_0011011100001101"; -- 0.09021324219656907
	pesos_i(6948) := b"0000000000000000_0000000000000000_0000011010110011_0010101101100000"; -- 0.026171408522347978
	pesos_i(6949) := b"1111111111111111_1111111111111111_1111000111011111_0000101101001011"; -- -0.05519036702634397
	pesos_i(6950) := b"0000000000000000_0000000000000000_0000000001100011_0101101100001101"; -- 0.0015160472592719908
	pesos_i(6951) := b"1111111111111111_1111111111111111_1101010001011111_1011010001011000"; -- -0.17041466569557145
	pesos_i(6952) := b"0000000000000000_0000000000000000_0010101110101011_0101011000111100"; -- 0.1705831429980523
	pesos_i(6953) := b"1111111111111111_1111111111111111_1111111110100110_0100011101101110"; -- -0.0013690334000880057
	pesos_i(6954) := b"1111111111111111_1111111111111111_1110110101001011_1000111100001000"; -- -0.07306581546360597
	pesos_i(6955) := b"1111111111111111_1111111111111111_1111111000110111_1001110101101101"; -- -0.0069638832106620795
	pesos_i(6956) := b"0000000000000000_0000000000000000_0010100010000010_1111001011101101"; -- 0.1582481219988148
	pesos_i(6957) := b"1111111111111111_1111111111111111_1101100110010100_0101100100110010"; -- -0.15008013268327755
	pesos_i(6958) := b"1111111111111111_1111111111111111_1110011100000111_0100010010011101"; -- -0.09754534890570347
	pesos_i(6959) := b"1111111111111111_1111111111111111_1110011001101011_1000010111111001"; -- -0.09992182426141592
	pesos_i(6960) := b"1111111111111111_1111111111111111_1111101110000001_1100011101101011"; -- -0.017550979910538667
	pesos_i(6961) := b"1111111111111111_1111111111111111_1101110101001001_0101011101100111"; -- -0.13559964875589356
	pesos_i(6962) := b"0000000000000000_0000000000000000_0001100111011010_1011101111111110"; -- 0.10099387114117675
	pesos_i(6963) := b"0000000000000000_0000000000000000_0010000011010110_1111101011001101"; -- 0.12828032985330726
	pesos_i(6964) := b"1111111111111111_1111111111111111_1110010101011010_0100001100010110"; -- -0.10409146039952599
	pesos_i(6965) := b"1111111111111111_1111111111111111_1110010110101011_1000011100001110"; -- -0.10285144712315322
	pesos_i(6966) := b"0000000000000000_0000000000000000_0000011100000000_0011110101110010"; -- 0.027347412319170327
	pesos_i(6967) := b"0000000000000000_0000000000000000_0001011011111110_0110100011001001"; -- 0.08981947803756878
	pesos_i(6968) := b"0000000000000000_0000000000000000_0001000110010100_1111000100101101"; -- 0.06867892607761406
	pesos_i(6969) := b"0000000000000000_0000000000000000_0001001001000110_1101101001100111"; -- 0.07139363292598894
	pesos_i(6970) := b"1111111111111111_1111111111111111_1111100111111011_0010011011100110"; -- -0.02351147535702015
	pesos_i(6971) := b"1111111111111111_1111111111111111_1110001011010110_1101001100000010"; -- -0.11390954210069826
	pesos_i(6972) := b"0000000000000000_0000000000000000_0000111001001001_0010000100010111"; -- 0.05580336383837045
	pesos_i(6973) := b"1111111111111111_1111111111111111_1111011001111011_1011110010001100"; -- -0.03717443059922012
	pesos_i(6974) := b"0000000000000000_0000000000000000_0000011101111101_0001010101010101"; -- 0.029252370108922038
	pesos_i(6975) := b"1111111111111111_1111111111111111_1110110101100000_0110110001001010"; -- -0.07274745162613547
	pesos_i(6976) := b"1111111111111111_1111111111111111_1101001110100001_1101111010110100"; -- -0.1733113107727897
	pesos_i(6977) := b"0000000000000000_0000000000000000_0001101111111011_1100101100110011"; -- 0.10931081766424897
	pesos_i(6978) := b"0000000000000000_0000000000000000_0000100110011101_1111111001100010"; -- 0.03756704232364398
	pesos_i(6979) := b"1111111111111111_1111111111111111_1110100000100100_1011001100101011"; -- -0.09319000439525908
	pesos_i(6980) := b"0000000000000000_0000000000000000_0000010010010101_0000100101011011"; -- 0.01789911710870278
	pesos_i(6981) := b"1111111111111111_1111111111111111_1111101100000010_0110101010010111"; -- -0.01949437910887652
	pesos_i(6982) := b"0000000000000000_0000000000000000_0001101111011001_0111110101001010"; -- 0.10878737510415885
	pesos_i(6983) := b"0000000000000000_0000000000000000_0010010110101111_1001000001111010"; -- 0.1472101495335526
	pesos_i(6984) := b"1111111111111111_1111111111111111_1111011100110010_1010000001101110"; -- -0.03438374821673182
	pesos_i(6985) := b"0000000000000000_0000000000000000_0001111110110100_0011111001000010"; -- 0.1238440429008401
	pesos_i(6986) := b"1111111111111111_1111111111111111_1101001001001100_0001000111100101"; -- -0.17852676551661897
	pesos_i(6987) := b"0000000000000000_0000000000000000_0001111101010101_1111110001010011"; -- 0.12240578669709123
	pesos_i(6988) := b"1111111111111111_1111111111111111_1111110010010111_1111010111111011"; -- -0.013306261354584296
	pesos_i(6989) := b"0000000000000000_0000000000000000_0000111011101111_1100011110111110"; -- 0.05834625615196261
	pesos_i(6990) := b"1111111111111111_1111111111111111_1111000000010010_1011100010010011"; -- -0.062214340386075054
	pesos_i(6991) := b"1111111111111111_1111111111111111_1111111010001100_1111101001010011"; -- -0.0056613490561392065
	pesos_i(6992) := b"1111111111111111_1111111111111111_1101001111110000_1101100001000001"; -- -0.17210625095011897
	pesos_i(6993) := b"0000000000000000_0000000000000000_0001010100000100_1000010011110100"; -- 0.08210020974059029
	pesos_i(6994) := b"1111111111111111_1111111111111111_1110000001011110_1011010000011001"; -- -0.12355493914121475
	pesos_i(6995) := b"1111111111111111_1111111111111111_1110100000000000_0111100100111100"; -- -0.09374277379532465
	pesos_i(6996) := b"1111111111111111_1111111111111111_1111110000001010_0001010110010111"; -- -0.01547112517344227
	pesos_i(6997) := b"1111111111111111_1111111111111111_1110101110111010_0011111100111110"; -- -0.07918934566766031
	pesos_i(6998) := b"0000000000000000_0000000000000000_0001001101001000_1110000110101010"; -- 0.07533083342865288
	pesos_i(6999) := b"1111111111111111_1111111111111111_1111101100110111_0001101010011101"; -- -0.018690430324061612
	pesos_i(7000) := b"0000000000000000_0000000000000000_0010010000110010_1101110111000010"; -- 0.14140115730792366
	pesos_i(7001) := b"1111111111111111_1111111111111111_1101110111111100_1001010100111010"; -- -0.13286464048797655
	pesos_i(7002) := b"0000000000000000_0000000000000000_0010011011111110_0001010000101100"; -- 0.15231443475333697
	pesos_i(7003) := b"0000000000000000_0000000000000000_0001100010111101_1000000110100101"; -- 0.09664163853422383
	pesos_i(7004) := b"0000000000000000_0000000000000000_0001111100000010_1010110010110000"; -- 0.12113456047654869
	pesos_i(7005) := b"0000000000000000_0000000000000000_0000100101001000_0100000100010100"; -- 0.03625876188705335
	pesos_i(7006) := b"0000000000000000_0000000000000000_0000011010101000_1100101001111110"; -- 0.026013046074437156
	pesos_i(7007) := b"1111111111111111_1111111111111111_1101011111101011_1111110001111010"; -- -0.15655538575580868
	pesos_i(7008) := b"0000000000000000_0000000000000000_0001010010001100_1100111100001101"; -- 0.08027357157547807
	pesos_i(7009) := b"0000000000000000_0000000000000000_0001110101000100_1111010000001110"; -- 0.11433339445418188
	pesos_i(7010) := b"1111111111111111_1111111111111111_1111111000010100_1000110010101100"; -- -0.007498939432678611
	pesos_i(7011) := b"1111111111111111_1111111111111111_1110111011011001_1000110111000001"; -- -0.06699289360242232
	pesos_i(7012) := b"0000000000000000_0000000000000000_0010001101000110_0001111001111110"; -- 0.13778868269981895
	pesos_i(7013) := b"1111111111111111_1111111111111111_1101111111011000_1011001101111111"; -- -0.1255996527206263
	pesos_i(7014) := b"0000000000000000_0000000000000000_0001101011000100_1000010000111111"; -- 0.1045611052242544
	pesos_i(7015) := b"1111111111111111_1111111111111111_1111100110010011_1101100110010110"; -- -0.025087738908403073
	pesos_i(7016) := b"0000000000000000_0000000000000000_0000011000011010_0111111111111100"; -- 0.023841856888866114
	pesos_i(7017) := b"0000000000000000_0000000000000000_0000101111000111_1110111101101110"; -- 0.04601952008466326
	pesos_i(7018) := b"1111111111111111_1111111111111111_1101101101010100_0010001111000100"; -- -0.14324737987637606
	pesos_i(7019) := b"1111111111111111_1111111111111111_1101010011111001_1000001011010101"; -- -0.16806776330287865
	pesos_i(7020) := b"0000000000000000_0000000000000000_0001111001111110_1101001100011001"; -- 0.11912268971703781
	pesos_i(7021) := b"1111111111111111_1111111111111111_1101110000100000_1001011011111101"; -- -0.14012771919849717
	pesos_i(7022) := b"1111111111111111_1111111111111111_1111100110011110_1010110101111010"; -- -0.024922521237068743
	pesos_i(7023) := b"1111111111111111_1111111111111111_1101011000110010_0110100011111101"; -- -0.16329330279153387
	pesos_i(7024) := b"0000000000000000_0000000000000000_0010001010011010_1001101100110111"; -- 0.13517160495129446
	pesos_i(7025) := b"1111111111111111_1111111111111111_1111111000011000_1011010000111111"; -- -0.0074355455170899976
	pesos_i(7026) := b"1111111111111111_1111111111111111_1111111100001101_1001101111000011"; -- -0.0036986015702073776
	pesos_i(7027) := b"1111111111111111_1111111111111111_1110000001011011_0011000111011110"; -- -0.12360847795322143
	pesos_i(7028) := b"0000000000000000_0000000000000000_0000101111001010_0000011000001101"; -- 0.04605138605876211
	pesos_i(7029) := b"0000000000000000_0000000000000000_0001011001101101_1100110101100001"; -- 0.08761294964074376
	pesos_i(7030) := b"1111111111111111_1111111111111111_1101100001010111_0001110011101001"; -- -0.1549207620993205
	pesos_i(7031) := b"0000000000000000_0000000000000000_0001111000010101_0000111101100001"; -- 0.11750885117883807
	pesos_i(7032) := b"1111111111111111_1111111111111111_1110101101010101_1010011010000101"; -- -0.0807243276172617
	pesos_i(7033) := b"1111111111111111_1111111111111111_1101000000011011_0000001001110011"; -- -0.18708786669262897
	pesos_i(7034) := b"0000000000000000_0000000000000000_0010001011101011_1100100001100000"; -- 0.13641025870071308
	pesos_i(7035) := b"0000000000000000_0000000000000000_0001000110001100_0010101110100010"; -- 0.06854508125872155
	pesos_i(7036) := b"0000000000000000_0000000000000000_0001010001110101_1101100011101111"; -- 0.0799232085582916
	pesos_i(7037) := b"0000000000000000_0000000000000000_0000001001100000_0100000110000111"; -- 0.009281249562141429
	pesos_i(7038) := b"1111111111111111_1111111111111111_1111011101010011_0000011001110011"; -- -0.03388938609201906
	pesos_i(7039) := b"1111111111111111_1111111111111111_1111001011110111_1011110000101001"; -- -0.05090736391972889
	pesos_i(7040) := b"1111111111111111_1111111111111111_1111111000000101_0110101000011101"; -- -0.007729881158737462
	pesos_i(7041) := b"0000000000000000_0000000000000000_0001101100110100_0010000100011101"; -- 0.10626418080871727
	pesos_i(7042) := b"1111111111111111_1111111111111111_1101111011100011_1111111101111000"; -- -0.1293335276497178
	pesos_i(7043) := b"0000000000000000_0000000000000000_0000111011001100_1000010101100010"; -- 0.05780824318850603
	pesos_i(7044) := b"0000000000000000_0000000000000000_0000011011011001_0011011111011011"; -- 0.026751986449215122
	pesos_i(7045) := b"0000000000000000_0000000000000000_0000001111101111_0011001100111101"; -- 0.015368654576329424
	pesos_i(7046) := b"0000000000000000_0000000000000000_0001010101100101_0000001111101110"; -- 0.08357262183012343
	pesos_i(7047) := b"1111111111111111_1111111111111111_1101100100000000_0010100001110010"; -- -0.15234133918553283
	pesos_i(7048) := b"0000000000000000_0000000000000000_0000111011101101_1111101010111110"; -- 0.05831877842784132
	pesos_i(7049) := b"0000000000000000_0000000000000000_0000000100101001_0110110111100010"; -- 0.004538409767930567
	pesos_i(7050) := b"0000000000000000_0000000000000000_0010111000110100_0110011110001010"; -- 0.1804871284883708
	pesos_i(7051) := b"0000000000000000_0000000000000000_0000000100100100_1110011000111001"; -- 0.004469288665830972
	pesos_i(7052) := b"1111111111111111_1111111111111111_1110110111000100_0101110100011010"; -- -0.07122247794674949
	pesos_i(7053) := b"0000000000000000_0000000000000000_0000101110001111_0001101101100001"; -- 0.04515238871695338
	pesos_i(7054) := b"1111111111111111_1111111111111111_1101010001000110_0101101101101001"; -- -0.17080143639128187
	pesos_i(7055) := b"0000000000000000_0000000000000000_0010100001010110_0101110100111010"; -- 0.15756781263482775
	pesos_i(7056) := b"1111111111111111_1111111111111111_1110110000110001_1100000001101101"; -- -0.0773658497847422
	pesos_i(7057) := b"0000000000000000_0000000000000000_0000000110111010_1100011100001111"; -- 0.006756249663595015
	pesos_i(7058) := b"1111111111111111_1111111111111111_1110011000111111_1100010101110010"; -- -0.10058942758036915
	pesos_i(7059) := b"0000000000000000_0000000000000000_0001110000011111_0011001101100101"; -- 0.10985108572566384
	pesos_i(7060) := b"0000000000000000_0000000000000000_0001010101010100_1110010011100001"; -- 0.08332663048550297
	pesos_i(7061) := b"1111111111111111_1111111111111111_1110100010001000_1001100101100101"; -- -0.09166566162129929
	pesos_i(7062) := b"1111111111111111_1111111111111111_1110011011100000_1111101100010001"; -- -0.0981295665130333
	pesos_i(7063) := b"1111111111111111_1111111111111111_1111101000101110_1100001001110000"; -- -0.02272400641470949
	pesos_i(7064) := b"1111111111111111_1111111111111111_1110111000100001_0010111111110111"; -- -0.0698061011014436
	pesos_i(7065) := b"0000000000000000_0000000000000000_0010000011110001_1101011000010101"; -- 0.12869012848651823
	pesos_i(7066) := b"1111111111111111_1111111111111111_1110010010000011_1100000101010101"; -- -0.10736457514948208
	pesos_i(7067) := b"1111111111111111_1111111111111111_1111101111010100_1010100011011110"; -- -0.016286321357230373
	pesos_i(7068) := b"0000000000000000_0000000000000000_0001101111011001_1010111110011110"; -- 0.10879037472699923
	pesos_i(7069) := b"1111111111111111_1111111111111111_1101100001110000_1101100011110001"; -- -0.15452808482211824
	pesos_i(7070) := b"1111111111111111_1111111111111111_1111101100000100_0110011011010101"; -- -0.019464085613002207
	pesos_i(7071) := b"1111111111111111_1111111111111111_1110100100100011_0100110111110000"; -- -0.0893050469283064
	pesos_i(7072) := b"0000000000000000_0000000000000000_0001010011100101_0000011110100010"; -- 0.08161971766937684
	pesos_i(7073) := b"1111111111111111_1111111111111111_1101110111010001_0001000010011110"; -- -0.1335286727013198
	pesos_i(7074) := b"0000000000000000_0000000000000000_0010011100011000_1010010001101000"; -- 0.15271976026878387
	pesos_i(7075) := b"0000000000000000_0000000000000000_0000110011111001_0001100011101001"; -- 0.05067592328609631
	pesos_i(7076) := b"0000000000000000_0000000000000000_0001110111011100_1000111010100111"; -- 0.11664668644017852
	pesos_i(7077) := b"0000000000000000_0000000000000000_0000110110101001_1010111001100011"; -- 0.053370379565537515
	pesos_i(7078) := b"1111111111111111_1111111111111111_1110111111100001_1001101010100110"; -- -0.06296380479626106
	pesos_i(7079) := b"1111111111111111_1111111111111111_1111011001011110_0111000110011100"; -- -0.03762140226350549
	pesos_i(7080) := b"0000000000000000_0000000000000000_0001010101011001_0011010110111111"; -- 0.08339248573237376
	pesos_i(7081) := b"1111111111111111_1111111111111111_1101110010011110_0101101010000001"; -- -0.13820871687998276
	pesos_i(7082) := b"1111111111111111_1111111111111111_1111011111010000_1111000100101011"; -- -0.031968047208413106
	pesos_i(7083) := b"1111111111111111_1111111111111111_1110011100101110_1011111001111010"; -- -0.09694299243502061
	pesos_i(7084) := b"1111111111111111_1111111111111111_1110100110010010_1100010000000100"; -- -0.08760428346591495
	pesos_i(7085) := b"1111111111111111_1111111111111111_1111000110101101_0100101110000111"; -- -0.05594947761033898
	pesos_i(7086) := b"1111111111111111_1111111111111111_1110010010011011_1111111011010000"; -- -0.10699469966256013
	pesos_i(7087) := b"1111111111111111_1111111111111111_1101111000100100_1011100110111010"; -- -0.13225211333854467
	pesos_i(7088) := b"0000000000000000_0000000000000000_0010110010011101_0100110000101011"; -- 0.17427516984085364
	pesos_i(7089) := b"0000000000000000_0000000000000000_0010011000011111_1101110110111000"; -- 0.14892373801989478
	pesos_i(7090) := b"0000000000000000_0000000000000000_0010100101111101_0011101001101110"; -- 0.16206708128405128
	pesos_i(7091) := b"1111111111111111_1111111111111111_1101010111111001_1110001000000001"; -- -0.1641558406356241
	pesos_i(7092) := b"0000000000000000_0000000000000000_0000011111010011_1101010011111110"; -- 0.030576049796509425
	pesos_i(7093) := b"0000000000000000_0000000000000000_0000011100010001_0101001001001000"; -- 0.02760805365727727
	pesos_i(7094) := b"1111111111111111_1111111111111111_1110010000011011_0101001000011110"; -- -0.10895811819057225
	pesos_i(7095) := b"1111111111111111_1111111111111111_1111011011111011_0101010011101100"; -- -0.0352274822448716
	pesos_i(7096) := b"0000000000000000_0000000000000000_0000010001001001_0010000000010010"; -- 0.01674080320051094
	pesos_i(7097) := b"0000000000000000_0000000000000000_0000100001010100_1010110001011000"; -- 0.03254201070340987
	pesos_i(7098) := b"0000000000000000_0000000000000000_0001010001110011_1110000001001001"; -- 0.07989312922438856
	pesos_i(7099) := b"1111111111111111_1111111111111111_1101010111100111_1101101100010100"; -- -0.16443091162066711
	pesos_i(7100) := b"1111111111111111_1111111111111111_1111000101011101_0001101011001011"; -- -0.05717308562801391
	pesos_i(7101) := b"0000000000000000_0000000000000000_0010100101001100_1110001100011100"; -- 0.16132945475103166
	pesos_i(7102) := b"1111111111111111_1111111111111111_1110010001011111_1010111010010100"; -- -0.10791500942496608
	pesos_i(7103) := b"0000000000000000_0000000000000000_0001111010000010_1111110000011000"; -- 0.11918616842705272
	pesos_i(7104) := b"0000000000000000_0000000000000000_0000000000010000_1001000101101111"; -- 0.0002528092562485429
	pesos_i(7105) := b"1111111111111111_1111111111111111_1101101110011101_1001100111101000"; -- -0.14212644662199644
	pesos_i(7106) := b"0000000000000000_0000000000000000_0000010100010110_1000111110001111"; -- 0.019875500067790215
	pesos_i(7107) := b"1111111111111111_1111111111111111_1110100001100011_0010011101011101"; -- -0.09223703363733937
	pesos_i(7108) := b"1111111111111111_1111111111111111_1110101100011001_1010100000111101"; -- -0.08163975244604603
	pesos_i(7109) := b"1111111111111111_1111111111111111_1111010000110111_0100010011101010"; -- -0.04603165906004337
	pesos_i(7110) := b"0000000000000000_0000000000000000_0001000011101000_0101000000100000"; -- 0.06604481480981766
	pesos_i(7111) := b"0000000000000000_0000000000000000_0010010110001100_0001110011100100"; -- 0.14666920246770548
	pesos_i(7112) := b"1111111111111111_1111111111111111_1110000000110011_0101101100100000"; -- -0.1242163701724046
	pesos_i(7113) := b"1111111111111111_1111111111111111_1110110110111111_0010111001011000"; -- -0.07130155895424112
	pesos_i(7114) := b"1111111111111111_1111111111111111_1111111001001001_0101101010011001"; -- -0.006693208254411622
	pesos_i(7115) := b"0000000000000000_0000000000000000_0010000010000110_0001110100000011"; -- 0.12704640686452132
	pesos_i(7116) := b"0000000000000000_0000000000000000_0001000111010110_0010010111111100"; -- 0.06967389497102683
	pesos_i(7117) := b"0000000000000000_0000000000000000_0010101001011111_0100100000101000"; -- 0.16551638588800777
	pesos_i(7118) := b"1111111111111111_1111111111111111_1101100001101110_1100011001000000"; -- -0.15455971650741068
	pesos_i(7119) := b"1111111111111111_1111111111111111_1101111110111100_1110110011010010"; -- -0.1260234821804908
	pesos_i(7120) := b"0000000000000000_0000000000000000_0001010011010011_1001000000111111"; -- 0.08135320220052797
	pesos_i(7121) := b"1111111111111111_1111111111111111_1110011101101011_0000000000110000"; -- -0.09602354835794612
	pesos_i(7122) := b"1111111111111111_1111111111111111_1101100110010000_1000101111101011"; -- -0.15013814468890674
	pesos_i(7123) := b"1111111111111111_1111111111111111_1110101000000010_1000101111111000"; -- -0.08589863952996286
	pesos_i(7124) := b"0000000000000000_0000000000000000_0001010101111001_0110011100110000"; -- 0.08388371389419795
	pesos_i(7125) := b"0000000000000000_0000000000000000_0000011011111000_1101110111101110"; -- 0.02723490774048036
	pesos_i(7126) := b"1111111111111111_1111111111111111_1110111110101100_0111011100011111"; -- -0.06377463806148273
	pesos_i(7127) := b"1111111111111111_1111111111111111_1111001100111101_0101111001011101"; -- -0.04984483932077419
	pesos_i(7128) := b"0000000000000000_0000000000000000_0010001111011001_1101011111110011"; -- 0.1400427788916417
	pesos_i(7129) := b"1111111111111111_1111111111111111_1111101011101101_0101011110001100"; -- -0.019815948836080562
	pesos_i(7130) := b"1111111111111111_1111111111111111_1110110110011010_0111001100010011"; -- -0.07186203758613895
	pesos_i(7131) := b"0000000000000000_0000000000000000_0001000010100100_0010011001100000"; -- 0.0650047287684026
	pesos_i(7132) := b"0000000000000000_0000000000000000_0001101101011001_1010110110100000"; -- 0.10683713116665437
	pesos_i(7133) := b"1111111111111111_1111111111111111_1110101010010100_1011010101101011"; -- -0.08366838581502058
	pesos_i(7134) := b"1111111111111111_1111111111111111_1110101111110010_1111010000011011"; -- -0.07832407313818794
	pesos_i(7135) := b"1111111111111111_1111111111111111_1111011011001001_0011100001101100"; -- -0.0359921204791992
	pesos_i(7136) := b"0000000000000000_0000000000000000_0010011101101001_1000110010000010"; -- 0.15395429788372164
	pesos_i(7137) := b"0000000000000000_0000000000000000_0001001110101010_1110111111101010"; -- 0.07682704421815835
	pesos_i(7138) := b"1111111111111111_1111111111111111_1101101100110111_1110111000101101"; -- -0.14367782015028585
	pesos_i(7139) := b"1111111111111111_1111111111111111_1101111001010011_1011010111011111"; -- -0.13153518014129126
	pesos_i(7140) := b"1111111111111111_1111111111111111_1110000000011011_0000000001011110"; -- -0.12458799077862787
	pesos_i(7141) := b"1111111111111111_1111111111111111_1110010111100000_0010000001010010"; -- -0.10204885485852624
	pesos_i(7142) := b"0000000000000000_0000000000000000_0010000101100111_1100011001101000"; -- 0.13048973127808974
	pesos_i(7143) := b"1111111111111111_1111111111111111_1111100001110101_1010010100000100"; -- -0.029454885992296703
	pesos_i(7144) := b"1111111111111111_1111111111111111_1101011110000000_1001110011001111"; -- -0.1581937784473829
	pesos_i(7145) := b"1111111111111111_1111111111111111_1110011111110100_0110010001100010"; -- -0.0939271222445451
	pesos_i(7146) := b"1111111111111111_1111111111111111_1101110001100111_1000011010011110"; -- -0.13904532096407854
	pesos_i(7147) := b"0000000000000000_0000000000000000_0000110111000111_0100000000110011"; -- 0.053821575621703456
	pesos_i(7148) := b"0000000000000000_0000000000000000_0001000011100001_0111011001010110"; -- 0.06594028099528139
	pesos_i(7149) := b"1111111111111111_1111111111111111_1101101010001001_1011011111000111"; -- -0.14633609194299846
	pesos_i(7150) := b"0000000000000000_0000000000000000_0001010100101011_1100001010101001"; -- 0.08269898064266326
	pesos_i(7151) := b"0000000000000000_0000000000000000_0000111010001010_1001010111000111"; -- 0.05680214034560446
	pesos_i(7152) := b"1111111111111111_1111111111111111_1110011000000011_1101101011000010"; -- -0.10150368468305915
	pesos_i(7153) := b"0000000000000000_0000000000000000_0010011100101000_0001001001011001"; -- 0.1529551951445497
	pesos_i(7154) := b"1111111111111111_1111111111111111_1101101101011010_0110101101111001"; -- -0.1431515531613535
	pesos_i(7155) := b"1111111111111111_1111111111111111_1110010010110111_0001111101001101"; -- -0.10658077598280576
	pesos_i(7156) := b"1111111111111111_1111111111111111_1111000110011101_1100011100111110"; -- -0.05618624424895765
	pesos_i(7157) := b"0000000000000000_0000000000000000_0001000001000000_1101000001111111"; -- 0.06348898992779017
	pesos_i(7158) := b"1111111111111111_1111111111111111_1111011010001011_1110011000101101"; -- -0.03692780875212593
	pesos_i(7159) := b"0000000000000000_0000000000000000_0000111101110100_0111100111000010"; -- 0.060371026857558255
	pesos_i(7160) := b"0000000000000000_0000000000000000_0001001000100110_0010110101110111"; -- 0.07089504394470056
	pesos_i(7161) := b"0000000000000000_0000000000000000_0010110010000000_1001111110011010"; -- 0.1738376380772797
	pesos_i(7162) := b"0000000000000000_0000000000000000_0010110011000011_1111110001010110"; -- 0.1748655042610581
	pesos_i(7163) := b"0000000000000000_0000000000000000_0010101010110000_1010100001110011"; -- 0.166758087164002
	pesos_i(7164) := b"0000000000000000_0000000000000000_0000001110101111_1011001110100110"; -- 0.014399745916486588
	pesos_i(7165) := b"1111111111111111_1111111111111111_1110101101100011_0111000101100011"; -- -0.0805138714561491
	pesos_i(7166) := b"0000000000000000_0000000000000000_0001001110111111_1101110110010000"; -- 0.07714638498007005
	pesos_i(7167) := b"0000000000000000_0000000000000000_0001000010100110_1111001111100110"; -- 0.06504749657522142
	pesos_i(7168) := b"1111111111111111_1111111111111111_1101111011011010_0101101010000110"; -- -0.12948068840373217
	pesos_i(7169) := b"0000000000000000_0000000000000000_0000000011111101_0000000011101001"; -- 0.003860527983445585
	pesos_i(7170) := b"1111111111111111_1111111111111111_1110110110110110_0111100000100111"; -- -0.07143448885121784
	pesos_i(7171) := b"0000000000000000_0000000000000000_0001011010111000_0011000000011010"; -- 0.088747984256875
	pesos_i(7172) := b"0000000000000000_0000000000000000_0001100110001111_0001110010101010"; -- 0.09983996528692517
	pesos_i(7173) := b"1111111111111111_1111111111111111_1101001001100001_1011100011110110"; -- -0.17819637282174308
	pesos_i(7174) := b"1111111111111111_1111111111111111_1101110000011000_1111001101010000"; -- -0.14024428659282628
	pesos_i(7175) := b"0000000000000000_0000000000000000_0001000011001100_1010010000000111"; -- 0.06562256985197693
	pesos_i(7176) := b"1111111111111111_1111111111111111_1110100110101000_1011111010011100"; -- -0.08726891216599675
	pesos_i(7177) := b"1111111111111111_1111111111111111_1111111011111100_0111011010111011"; -- -0.003960208307290821
	pesos_i(7178) := b"1111111111111111_1111111111111111_1101100110000110_1000110100111110"; -- -0.1502906536158642
	pesos_i(7179) := b"1111111111111111_1111111111111111_1110100100110111_1011110111000011"; -- -0.08899320582081993
	pesos_i(7180) := b"0000000000000000_0000000000000000_0000010100000010_1110011010011010"; -- 0.01957551252780794
	pesos_i(7181) := b"0000000000000000_0000000000000000_0010011010110010_0010100101000101"; -- 0.15115602429391375
	pesos_i(7182) := b"1111111111111111_1111111111111111_1101111001011001_0010101001000011"; -- -0.13145194881853195
	pesos_i(7183) := b"0000000000000000_0000000000000000_0010001000110101_0110010110000001"; -- 0.1336272659973311
	pesos_i(7184) := b"0000000000000000_0000000000000000_0000111000100111_0111011011011010"; -- 0.05528967678190094
	pesos_i(7185) := b"0000000000000000_0000000000000000_0010100111100010_0011011010110101"; -- 0.16360799723156466
	pesos_i(7186) := b"1111111111111111_1111111111111111_1101100010100111_0101101000001001"; -- -0.1536964157142472
	pesos_i(7187) := b"1111111111111111_1111111111111111_1111101011011101_1011101011001101"; -- -0.020054173308365213
	pesos_i(7188) := b"0000000000000000_0000000000000000_0010000111110011_1111011101111110"; -- 0.13262888745569254
	pesos_i(7189) := b"0000000000000000_0000000000000000_0000111101100110_0110010101100001"; -- 0.06015618917237109
	pesos_i(7190) := b"0000000000000000_0000000000000000_0001111010000100_1001000001001011"; -- 0.11921026063112816
	pesos_i(7191) := b"0000000000000000_0000000000000000_0011010010011001_1110010111110110"; -- 0.20547330146436524
	pesos_i(7192) := b"0000000000000000_0000000000000000_0010100111010010_0110101101110110"; -- 0.1633670008825381
	pesos_i(7193) := b"0000000000000000_0000000000000000_0000101001000100_0111110001101110"; -- 0.040107514211061804
	pesos_i(7194) := b"0000000000000000_0000000000000000_0010101100001111_0100100000100100"; -- 0.1682019317921008
	pesos_i(7195) := b"1111111111111111_1111111111111111_1111010111110101_1110000011000101"; -- -0.03921694940550275
	pesos_i(7196) := b"0000000000000000_0000000000000000_0001000000100000_0111111101011111"; -- 0.06299587316830198
	pesos_i(7197) := b"1111111111111111_1111111111111111_1101011111110101_0111010111001010"; -- -0.15641082592190939
	pesos_i(7198) := b"0000000000000000_0000000000000000_0000110111110000_1011000100111101"; -- 0.05445392370659694
	pesos_i(7199) := b"1111111111111111_1111111111111111_1111011111001111_0010111111101101"; -- -0.03199482397266831
	pesos_i(7200) := b"0000000000000000_0000000000000000_0010110100100000_0011001101011101"; -- 0.1762725927538997
	pesos_i(7201) := b"1111111111111111_1111111111111111_1101001100000011_0100101100000110"; -- -0.17573100187952487
	pesos_i(7202) := b"0000000000000000_0000000000000000_0001001111111111_1000100011011011"; -- 0.07811789848618758
	pesos_i(7203) := b"1111111111111111_1111111111111111_1111010000000110_0101001000001111"; -- -0.0467785561387559
	pesos_i(7204) := b"0000000000000000_0000000000000000_0001111011100111_1011000101011011"; -- 0.1207228514392898
	pesos_i(7205) := b"0000000000000000_0000000000000000_0010011010011010_1001101100011011"; -- 0.15079659841443696
	pesos_i(7206) := b"0000000000000000_0000000000000000_0010001000000010_0111000001101001"; -- 0.13284971775246565
	pesos_i(7207) := b"0000000000000000_0000000000000000_0010100001010111_0000010100010101"; -- 0.15757781745467217
	pesos_i(7208) := b"0000000000000000_0000000000000000_0001000001001110_0011010010001010"; -- 0.06369331718205432
	pesos_i(7209) := b"0000000000000000_0000000000000000_0010101001101010_0100000110010111"; -- 0.16568384100051362
	pesos_i(7210) := b"0000000000000000_0000000000000000_0000100010111101_1111100000111110"; -- 0.034148707500876584
	pesos_i(7211) := b"1111111111111111_1111111111111111_1111101010011010_1101110000100001"; -- -0.021074525663031723
	pesos_i(7212) := b"1111111111111111_1111111111111111_1111010000000010_1011011111110011"; -- -0.04683351818409468
	pesos_i(7213) := b"0000000000000000_0000000000000000_0000101100001001_1011111101010010"; -- 0.04311748268903534
	pesos_i(7214) := b"0000000000000000_0000000000000000_0000011101001000_0011001101110001"; -- 0.02844544898602131
	pesos_i(7215) := b"0000000000000000_0000000000000000_0000011111100010_0111010001010000"; -- 0.030799169106851265
	pesos_i(7216) := b"0000000000000000_0000000000000000_0000101010101101_1001110011011100"; -- 0.04171161996514702
	pesos_i(7217) := b"1111111111111111_1111111111111111_1110010111101001_0010011110110101"; -- -0.1019110853961524
	pesos_i(7218) := b"0000000000000000_0000000000000000_0010010010110100_1010100000101101"; -- 0.14338160614157244
	pesos_i(7219) := b"0000000000000000_0000000000000000_0010010111100010_0111001110011010"; -- 0.1479866266683992
	pesos_i(7220) := b"0000000000000000_0000000000000000_0000100110011000_1001000000010000"; -- 0.03748417267689044
	pesos_i(7221) := b"1111111111111111_1111111111111111_1111101100100111_1111011111101001"; -- -0.01892138072203075
	pesos_i(7222) := b"1111111111111111_1111111111111111_1110100101000001_0001111001110111"; -- -0.08885011289112411
	pesos_i(7223) := b"0000000000000000_0000000000000000_0000101111001000_1101000111110111"; -- 0.04603302258249409
	pesos_i(7224) := b"1111111111111111_1111111111111111_1111000111011101_1100011000110011"; -- -0.05520974396256634
	pesos_i(7225) := b"1111111111111111_1111111111111111_1111100101110101_1110000110010101"; -- -0.025545025858621326
	pesos_i(7226) := b"1111111111111111_1111111111111111_1110000110101100_0011101111100001"; -- -0.11846566918155765
	pesos_i(7227) := b"1111111111111111_1111111111111111_1101101000000111_1000110110100010"; -- -0.1483222464479125
	pesos_i(7228) := b"1111111111111111_1111111111111111_1101010011010011_0011000010001101"; -- -0.16865250169169493
	pesos_i(7229) := b"1111111111111111_1111111111111111_1110000100100011_0010110111100100"; -- -0.12055695706307805
	pesos_i(7230) := b"1111111111111111_1111111111111111_1101111000001000_1111000110011010"; -- -0.13267602904767745
	pesos_i(7231) := b"0000000000000000_0000000000000000_0001011110000110_0101000011111111"; -- 0.0918932555211921
	pesos_i(7232) := b"0000000000000000_0000000000000000_0000101101000010_1100101010101110"; -- 0.04398791066530419
	pesos_i(7233) := b"0000000000000000_0000000000000000_0010000101111001_0110110110010000"; -- 0.1307590938304116
	pesos_i(7234) := b"0000000000000000_0000000000000000_0001110110011010_0101100110000111"; -- 0.11563643986539686
	pesos_i(7235) := b"1111111111111111_1111111111111111_1101100101010001_0101111110011100"; -- -0.15110208928657437
	pesos_i(7236) := b"0000000000000000_0000000000000000_0010010111001100_1111100010101110"; -- 0.14765886538426773
	pesos_i(7237) := b"0000000000000000_0000000000000000_0001010110110010_0111000001111100"; -- 0.08475401894151617
	pesos_i(7238) := b"0000000000000000_0000000000000000_0011001110000111_1101101111001000"; -- 0.20129178647930795
	pesos_i(7239) := b"1111111111111111_1111111111111111_1101101010111101_1101110000100101"; -- -0.14554046732855744
	pesos_i(7240) := b"1111111111111111_1111111111111111_1101011100100110_1100110100101110"; -- -0.15956418639824196
	pesos_i(7241) := b"1111111111111111_1111111111111111_1111101110010111_1001101110011110"; -- -0.017217897438130965
	pesos_i(7242) := b"0000000000000000_0000000000000000_0000001011010000_1000111010010011"; -- 0.010994826146293683
	pesos_i(7243) := b"0000000000000000_0000000000000000_0000010101001101_1010010100001101"; -- 0.020716014500880085
	pesos_i(7244) := b"1111111111111111_1111111111111111_1111000000101011_1011011100111101"; -- -0.06183295025434903
	pesos_i(7245) := b"0000000000000000_0000000000000000_0000000001011011_0111011001110101"; -- 0.0013956104203510953
	pesos_i(7246) := b"0000000000000000_0000000000000000_0010000010110001_0110111111011001"; -- 0.12770747236159313
	pesos_i(7247) := b"0000000000000000_0000000000000000_0010000100010110_0011111011101101"; -- 0.12924569395743715
	pesos_i(7248) := b"1111111111111111_1111111111111111_1111000011101101_1110011010100110"; -- -0.05886991930895459
	pesos_i(7249) := b"0000000000000000_0000000000000000_0001010001101111_0110010000011000"; -- 0.07982469158955181
	pesos_i(7250) := b"1111111111111111_1111111111111111_1111001111011001_0010010001100010"; -- -0.047467924190616476
	pesos_i(7251) := b"0000000000000000_0000000000000000_0000000010011110_0100000101110101"; -- 0.002414790318889311
	pesos_i(7252) := b"1111111111111111_1111111111111111_1101010001111001_0100101110101010"; -- -0.1700241766851528
	pesos_i(7253) := b"1111111111111111_1111111111111111_1110010100001100_0001001100000001"; -- -0.10528451184737754
	pesos_i(7254) := b"0000000000000000_0000000000000000_0000000101001010_1110010001011001"; -- 0.0050490110043048125
	pesos_i(7255) := b"0000000000000000_0000000000000000_0001110111110001_0000000011011110"; -- 0.11695866993503416
	pesos_i(7256) := b"0000000000000000_0000000000000000_0010011100011111_0101001111011000"; -- 0.15282176982307635
	pesos_i(7257) := b"1111111111111111_1111111111111111_1111000001011100_1111110101000001"; -- -0.06108109627598746
	pesos_i(7258) := b"0000000000000000_0000000000000000_0001101010011100_1010111010110000"; -- 0.10395328328313044
	pesos_i(7259) := b"1111111111111111_1111111111111111_1110001000111111_0000001101001101"; -- -0.11622599959315966
	pesos_i(7260) := b"0000000000000000_0000000000000000_0010001011101011_0111010100010111"; -- 0.13640529449363167
	pesos_i(7261) := b"1111111111111111_1111111111111111_1111001000100010_0010010110110101"; -- -0.054166453596229756
	pesos_i(7262) := b"0000000000000000_0000000000000000_0001001000010110_0001101101010010"; -- 0.07064982167188233
	pesos_i(7263) := b"1111111111111111_1111111111111111_1111010010111000_0001000110000101"; -- -0.04406633866700771
	pesos_i(7264) := b"1111111111111111_1111111111111111_1111100001111100_1100111000011101"; -- -0.029345624805521553
	pesos_i(7265) := b"0000000000000000_0000000000000000_0001111111000100_1001010101101001"; -- 0.12409337827296386
	pesos_i(7266) := b"0000000000000000_0000000000000000_0001011101111011_1010111011010100"; -- 0.09173100166345831
	pesos_i(7267) := b"0000000000000000_0000000000000000_0010100110110100_1001011001111011"; -- 0.1629118013880833
	pesos_i(7268) := b"0000000000000000_0000000000000000_0010100110001101_0001011011100110"; -- 0.162309104096172
	pesos_i(7269) := b"0000000000000000_0000000000000000_0010011000011011_1001001011001101"; -- 0.1488582373037219
	pesos_i(7270) := b"0000000000000000_0000000000000000_0000011010111111_1001001110000101"; -- 0.026360721554949385
	pesos_i(7271) := b"1111111111111111_1111111111111111_1110111110100100_1010011101001100"; -- -0.06389383703567186
	pesos_i(7272) := b"0000000000000000_0000000000000000_0010001011111111_0011001100101111"; -- 0.13670654196158924
	pesos_i(7273) := b"0000000000000000_0000000000000000_0000001010100111_0011101101101001"; -- 0.010364258825616724
	pesos_i(7274) := b"1111111111111111_1111111111111111_1110111110110011_0010011110100011"; -- -0.0636725641845808
	pesos_i(7275) := b"0000000000000000_0000000000000000_0001110000111000_0111011010010011"; -- 0.11023655971850346
	pesos_i(7276) := b"1111111111111111_1111111111111111_1101110110100010_0111100101011100"; -- -0.13423959264695687
	pesos_i(7277) := b"0000000000000000_0000000000000000_0000110100000010_1110101100101111"; -- 0.050825785590043415
	pesos_i(7278) := b"0000000000000000_0000000000000000_0000110001011011_1111101010010010"; -- 0.048278485004031764
	pesos_i(7279) := b"1111111111111111_1111111111111111_1110010101001011_1100000000101001"; -- -0.10431288722278183
	pesos_i(7280) := b"1111111111111111_1111111111111111_1110011111100010_0111011010100101"; -- -0.09420069179994944
	pesos_i(7281) := b"1111111111111111_1111111111111111_1111110111101101_1011111011101100"; -- -0.008091037111698939
	pesos_i(7282) := b"1111111111111111_1111111111111111_1101110100000010_0110100000001011"; -- -0.13668203100574827
	pesos_i(7283) := b"0000000000000000_0000000000000000_0001010110010110_0101110010000101"; -- 0.08432558292297354
	pesos_i(7284) := b"0000000000000000_0000000000000000_0000011101011011_0011111110000001"; -- 0.028736084870997488
	pesos_i(7285) := b"0000000000000000_0000000000000000_0000000101110110_0111111101110001"; -- 0.00571438321991035
	pesos_i(7286) := b"0000000000000000_0000000000000000_0000000111111110_0001001000000010"; -- 0.007783055715749417
	pesos_i(7287) := b"0000000000000000_0000000000000000_0000001111001110_0011011000101010"; -- 0.014865288961930229
	pesos_i(7288) := b"0000000000000000_0000000000000000_0010010000100101_0101100100000010"; -- 0.14119488049220133
	pesos_i(7289) := b"1111111111111111_1111111111111111_1100111110010011_0110110000000101"; -- -0.1891567695453878
	pesos_i(7290) := b"1111111111111111_1111111111111111_1110010100000101_1100101001011011"; -- -0.10538039463979515
	pesos_i(7291) := b"1111111111111111_1111111111111111_1111100010010110_0001010011011100"; -- -0.028959938336322984
	pesos_i(7292) := b"1111111111111111_1111111111111111_1111100101000100_0000111101101000"; -- -0.02630523402418115
	pesos_i(7293) := b"1111111111111111_1111111111111111_1111101011001100_1011111001100101"; -- -0.020313358681648803
	pesos_i(7294) := b"0000000000000000_0000000000000000_0001110100101111_0110011000100011"; -- 0.11400450083841816
	pesos_i(7295) := b"1111111111111111_1111111111111111_1111000100111100_0111101000001110"; -- -0.05767094765387264
	pesos_i(7296) := b"1111111111111111_1111111111111111_1110111110101011_1111100001010000"; -- -0.06378219656416184
	pesos_i(7297) := b"1111111111111111_1111111111111111_1110010010110010_1000101011001100"; -- -0.10665066249397623
	pesos_i(7298) := b"0000000000000000_0000000000000000_0001111011011010_1111001011111010"; -- 0.120528398498891
	pesos_i(7299) := b"0000000000000000_0000000000000000_0001101011010110_0000111010011001"; -- 0.10482875090814228
	pesos_i(7300) := b"1111111111111111_1111111111111111_1111100101100011_1001011101110000"; -- -0.025824103596151407
	pesos_i(7301) := b"1111111111111111_1111111111111111_1111101111110010_0100111100100100"; -- -0.01583390593200419
	pesos_i(7302) := b"0000000000000000_0000000000000000_0001000010010000_0101111000000000"; -- 0.06470286840980106
	pesos_i(7303) := b"0000000000000000_0000000000000000_0001111110011100_1000001111001000"; -- 0.12348197587745613
	pesos_i(7304) := b"1111111111111111_1111111111111111_1101111010011010_1111100111010110"; -- -0.13044775503933895
	pesos_i(7305) := b"1111111111111111_1111111111111111_1111000101101011_0110000010001010"; -- -0.05695530547210873
	pesos_i(7306) := b"0000000000000000_0000000000000000_0001100000001011_0100110011011100"; -- 0.09392242777176754
	pesos_i(7307) := b"1111111111111111_1111111111111111_1110101000010111_1101011010100100"; -- -0.08557375418952197
	pesos_i(7308) := b"0000000000000000_0000000000000000_0000011000111011_0000000001101001"; -- 0.02433779308640638
	pesos_i(7309) := b"1111111111111111_1111111111111111_1110101111100000_0001011110010110"; -- -0.07861187535949768
	pesos_i(7310) := b"1111111111111111_1111111111111111_1110011100101001_0001010010100000"; -- -0.09702941029762129
	pesos_i(7311) := b"0000000000000000_0000000000000000_0001001101010010_1000011100110101"; -- 0.0754780296048396
	pesos_i(7312) := b"0000000000000000_0000000000000000_0010010000100000_0110010101111110"; -- 0.14111933074381175
	pesos_i(7313) := b"1111111111111111_1111111111111111_1111111110011100_0010111010110010"; -- -0.0015230957281736767
	pesos_i(7314) := b"0000000000000000_0000000000000000_0001011000110110_1111001010101000"; -- 0.08677593806191831
	pesos_i(7315) := b"1111111111111111_1111111111111111_1111101110101101_0000100111111000"; -- -0.016890885406570102
	pesos_i(7316) := b"0000000000000000_0000000000000000_0010001000111111_1011101101101011"; -- 0.13378497467357264
	pesos_i(7317) := b"1111111111111111_1111111111111111_1111100010100010_1100011110101100"; -- -0.028766174768024483
	pesos_i(7318) := b"1111111111111111_1111111111111111_1111011101110101_0011011101010011"; -- -0.03336767409774988
	pesos_i(7319) := b"0000000000000000_0000000000000000_0000111110011101_1001010011010001"; -- 0.06099824994289261
	pesos_i(7320) := b"1111111111111111_1111111111111111_1111101100100010_1011010111011011"; -- -0.01900161168402757
	pesos_i(7321) := b"1111111111111111_1111111111111111_1111011110010100_1101010010111110"; -- -0.03288526874984763
	pesos_i(7322) := b"1111111111111111_1111111111111111_1110100011111011_1010000111110110"; -- -0.08991039026942693
	pesos_i(7323) := b"1111111111111111_1111111111111111_1110100111111001_1011110001110011"; -- -0.0860330791486634
	pesos_i(7324) := b"0000000000000000_0000000000000000_0001101011110011_1000111101110010"; -- 0.10527893569829892
	pesos_i(7325) := b"0000000000000000_0000000000000000_0000101000000110_1100011010001100"; -- 0.039165886968131745
	pesos_i(7326) := b"0000000000000000_0000000000000000_0001000010010001_0000010000111101"; -- 0.06471277702437199
	pesos_i(7327) := b"1111111111111111_1111111111111111_1111000000010011_1101100001000011"; -- -0.06219719284042036
	pesos_i(7328) := b"1111111111111111_1111111111111111_1101101110100010_1111010011000100"; -- -0.1420447370435723
	pesos_i(7329) := b"0000000000000000_0000000000000000_0010010000101011_0000100001101110"; -- 0.14128163035239577
	pesos_i(7330) := b"0000000000000000_0000000000000000_0001010111100001_1001101000100001"; -- 0.08547366441192746
	pesos_i(7331) := b"1111111111111111_1111111111111111_1110100010000010_0011101011101110"; -- -0.09176284493251197
	pesos_i(7332) := b"1111111111111111_1111111111111111_1110110110000001_0011100010001001"; -- -0.07224699653486315
	pesos_i(7333) := b"0000000000000000_0000000000000000_0001000000111001_0001001110111011"; -- 0.06337092705806267
	pesos_i(7334) := b"0000000000000000_0000000000000000_0001110000011100_0111100111101111"; -- 0.10980951399488882
	pesos_i(7335) := b"0000000000000000_0000000000000000_0001101000101100_0011010110110100"; -- 0.1022370876075139
	pesos_i(7336) := b"0000000000000000_0000000000000000_0010100001101111_0111101101100110"; -- 0.15795108062301125
	pesos_i(7337) := b"0000000000000000_0000000000000000_0000101001110111_1000110011000001"; -- 0.04088668546031597
	pesos_i(7338) := b"0000000000000000_0000000000000000_0001011110101000_0111000001101111"; -- 0.09241392812156161
	pesos_i(7339) := b"1111111111111111_1111111111111111_1110010111110011_0110101100111111"; -- -0.10175447189889263
	pesos_i(7340) := b"1111111111111111_1111111111111111_1110011100010010_1000011000010111"; -- -0.09737359950814742
	pesos_i(7341) := b"1111111111111111_1111111111111111_1110001110101011_1001111101001101"; -- -0.11066250203842322
	pesos_i(7342) := b"0000000000000000_0000000000000000_0001111010110000_0001010111101010"; -- 0.11987435315063276
	pesos_i(7343) := b"0000000000000000_0000000000000000_0000111010011101_1101010101011010"; -- 0.05709584652782315
	pesos_i(7344) := b"1111111111111111_1111111111111111_1101101011110000_1000100011100101"; -- -0.14476723108457148
	pesos_i(7345) := b"0000000000000000_0000000000000000_0001100010101000_1100011000101001"; -- 0.09632528777288499
	pesos_i(7346) := b"1111111111111111_1111111111111111_1111100100101011_0000001001111100"; -- -0.026687474026696346
	pesos_i(7347) := b"1111111111111111_1111111111111111_1110111001100111_0100011110011010"; -- -0.06873657692839671
	pesos_i(7348) := b"0000000000000000_0000000000000000_0001010000010101_1101000110111011"; -- 0.0784579355852406
	pesos_i(7349) := b"1111111111111111_1111111111111111_1101010110110011_1001111101011101"; -- -0.1652279279748317
	pesos_i(7350) := b"0000000000000000_0000000000000000_0001001111100100_0101011011100001"; -- 0.0777029322588602
	pesos_i(7351) := b"0000000000000000_0000000000000000_0001110011100011_1101001000001100"; -- 0.11285126490178927
	pesos_i(7352) := b"0000000000000000_0000000000000000_0001000111101111_0101111011000111"; -- 0.07005874973784784
	pesos_i(7353) := b"0000000000000000_0000000000000000_0010001010011000_0110111010011101"; -- 0.13513842895549863
	pesos_i(7354) := b"0000000000000000_0000000000000000_0000110011101110_1001110011110111"; -- 0.05051594765220398
	pesos_i(7355) := b"0000000000000000_0000000000000000_0000000101010001_1100111000111100"; -- 0.005154504493041189
	pesos_i(7356) := b"0000000000000000_0000000000000000_0000011001001110_1010101110110110"; -- 0.024637920251846673
	pesos_i(7357) := b"0000000000000000_0000000000000000_0000100100100001_0001100100000001"; -- 0.03566128040619037
	pesos_i(7358) := b"0000000000000000_0000000000000000_0001100010101110_0011000111101001"; -- 0.09640800422711515
	pesos_i(7359) := b"1111111111111111_1111111111111111_1110101101111101_1011100111000100"; -- -0.08011282898863857
	pesos_i(7360) := b"1111111111111111_1111111111111111_1101110110000101_0100010011011111"; -- -0.1346852261214645
	pesos_i(7361) := b"0000000000000000_0000000000000000_0001111100000101_1110001011110100"; -- 0.12118357151708024
	pesos_i(7362) := b"0000000000000000_0000000000000000_0000010110011010_0011000101001000"; -- 0.02188404081787644
	pesos_i(7363) := b"0000000000000000_0000000000000000_0001111000011100_1000011101110001"; -- 0.11762281894473635
	pesos_i(7364) := b"1111111111111111_1111111111111111_1110111000000101_1100000010100000"; -- -0.07022472475397533
	pesos_i(7365) := b"0000000000000000_0000000000000000_0000111101011010_0011111011011100"; -- 0.05997078773384232
	pesos_i(7366) := b"0000000000000000_0000000000000000_0001000110100100_0001000110000101"; -- 0.06890973574138619
	pesos_i(7367) := b"1111111111111111_1111111111111111_1111111010000100_1010001100011010"; -- -0.005788618306825282
	pesos_i(7368) := b"0000000000000000_0000000000000000_0001010000101100_0101011111100101"; -- 0.07880162564207714
	pesos_i(7369) := b"0000000000000000_0000000000000000_0001000111010010_1010010011010010"; -- 0.06962041985114002
	pesos_i(7370) := b"0000000000000000_0000000000000000_0010001100001111_1011101110011001"; -- 0.1369588135560204
	pesos_i(7371) := b"0000000000000000_0000000000000000_0001001011110110_0011110010111111"; -- 0.0740697828425672
	pesos_i(7372) := b"0000000000000000_0000000000000000_0001111011110001_1000011110101000"; -- 0.12087295382793367
	pesos_i(7373) := b"1111111111111111_1111111111111111_1101111010100100_1000001001101011"; -- -0.1303022851715113
	pesos_i(7374) := b"1111111111111111_1111111111111111_1110001011010100_1011111011001010"; -- -0.11394126473492432
	pesos_i(7375) := b"1111111111111111_1111111111111111_1110101001100101_0111101100011101"; -- -0.08438902415390372
	pesos_i(7376) := b"1111111111111111_1111111111111111_1101010101101101_0110010010101010"; -- -0.16629954201357186
	pesos_i(7377) := b"1111111111111111_1111111111111111_1111001011011011_0010100000000100"; -- -0.051343440093094085
	pesos_i(7378) := b"0000000000000000_0000000000000000_0000110110111100_0001010001111001"; -- 0.053651122721702936
	pesos_i(7379) := b"0000000000000000_0000000000000000_0010001001001010_1100001011011110"; -- 0.1339532654120023
	pesos_i(7380) := b"1111111111111111_1111111111111111_1111101110101110_1011111001111100"; -- -0.016864866879792374
	pesos_i(7381) := b"0000000000000000_0000000000000000_0001010001111110_0100101010001011"; -- 0.08005205050308209
	pesos_i(7382) := b"0000000000000000_0000000000000000_0010000000011010_1010111100100001"; -- 0.12540716708594915
	pesos_i(7383) := b"0000000000000000_0000000000000000_0000111110000101_0010101110011100"; -- 0.06062576829107501
	pesos_i(7384) := b"1111111111111111_1111111111111111_1110000110001110_0011110011001100"; -- -0.11892337817715891
	pesos_i(7385) := b"1111111111111111_1111111111111111_1110011010110001_0001011100000110"; -- -0.09886032206093899
	pesos_i(7386) := b"1111111111111111_1111111111111111_1110101110011101_0110111100010010"; -- -0.07962899970988295
	pesos_i(7387) := b"0000000000000000_0000000000000000_0000011101101110_1101000100010010"; -- 0.02903467840444547
	pesos_i(7388) := b"1111111111111111_1111111111111111_1111110000001001_1001001100010000"; -- -0.015478905373227861
	pesos_i(7389) := b"1111111111111111_1111111111111111_1111000011011001_1010101100101110"; -- -0.0591786397471876
	pesos_i(7390) := b"1111111111111111_1111111111111111_1101111011111101_0010011110110110"; -- -0.1289496593246549
	pesos_i(7391) := b"0000000000000000_0000000000000000_0000001100100001_0010010011010011"; -- 0.012224484853150558
	pesos_i(7392) := b"1111111111111111_1111111111111111_1101011101010001_0010111111000000"; -- -0.15891744195132185
	pesos_i(7393) := b"1111111111111111_1111111111111111_1111001001101111_1011001101010010"; -- -0.05298308600305023
	pesos_i(7394) := b"1111111111111111_1111111111111111_1101111010111110_0011100110110100"; -- -0.12990989080384663
	pesos_i(7395) := b"0000000000000000_0000000000000000_0010011000101101_1100100000110101"; -- 0.1491360787082578
	pesos_i(7396) := b"1111111111111111_1111111111111111_1111110101111101_1010011001101111"; -- -0.00980148123721692
	pesos_i(7397) := b"1111111111111111_1111111111111111_1101011001110101_1010101110110001"; -- -0.162266987970736
	pesos_i(7398) := b"0000000000000000_0000000000000000_0001010110001010_0111001001100110"; -- 0.08414378150438773
	pesos_i(7399) := b"1111111111111111_1111111111111111_1111011000101110_0100100001001000"; -- -0.03835628741481345
	pesos_i(7400) := b"1111111111111111_1111111111111111_1101101000001011_0111101000011011"; -- -0.1482623752297816
	pesos_i(7401) := b"1111111111111111_1111111111111111_1111111100000000_1000110100100100"; -- -0.003897837358317453
	pesos_i(7402) := b"1111111111111111_1111111111111111_1111101010010001_0010000101101000"; -- -0.02122298443251383
	pesos_i(7403) := b"1111111111111111_1111111111111111_1101110101101000_0100101010010110"; -- -0.13512739026730358
	pesos_i(7404) := b"1111111111111111_1111111111111111_1110110010110110_1101110100010011"; -- -0.07533472324773773
	pesos_i(7405) := b"0000000000000000_0000000000000000_0001111100011100_0000110000111100"; -- 0.12152172526592336
	pesos_i(7406) := b"0000000000000000_0000000000000000_0001111010000001_0001001011010010"; -- 0.11915700549759253
	pesos_i(7407) := b"1111111111111111_1111111111111111_1101111111001001_1100110101111110"; -- -0.1258269850483644
	pesos_i(7408) := b"0000000000000000_0000000000000000_0001110110111100_1101001101110101"; -- 0.11616250625195204
	pesos_i(7409) := b"0000000000000000_0000000000000000_0001100111000010_0101110100010101"; -- 0.10062200308923751
	pesos_i(7410) := b"0000000000000000_0000000000000000_0001110000101011_1110101101010011"; -- 0.1100451542758665
	pesos_i(7411) := b"1111111111111111_1111111111111111_1110101111001010_1110010110011000"; -- -0.07893528983178194
	pesos_i(7412) := b"0000000000000000_0000000000000000_0000010101000000_1010011101101011"; -- 0.020517791399489282
	pesos_i(7413) := b"1111111111111111_1111111111111111_1111100010101111_1111001111000011"; -- -0.02856518265271989
	pesos_i(7414) := b"0000000000000000_0000000000000000_0010001110100100_1110101011010000"; -- 0.1392351873282496
	pesos_i(7415) := b"1111111111111111_1111111111111111_1111110110010010_0011110101001111"; -- -0.009487312452660077
	pesos_i(7416) := b"0000000000000000_0000000000000000_0000001001110011_1100100101111010"; -- 0.009579269768737214
	pesos_i(7417) := b"1111111111111111_1111111111111111_1110101001001101_1000010101111010"; -- -0.08475461738145297
	pesos_i(7418) := b"0000000000000000_0000000000000000_0000000000110111_0000010110100110"; -- 0.0008395700496999315
	pesos_i(7419) := b"0000000000000000_0000000000000000_0010010010110100_0101011111101100"; -- 0.14337682265757853
	pesos_i(7420) := b"1111111111111111_1111111111111111_1110010001000000_0100011111011011"; -- -0.10839415459422212
	pesos_i(7421) := b"0000000000000000_0000000000000000_0010011011101011_0100000000001001"; -- 0.1520271322889576
	pesos_i(7422) := b"1111111111111111_1111111111111111_1111011101100010_0000100001011111"; -- -0.03366038982915174
	pesos_i(7423) := b"0000000000000000_0000000000000000_0000010011011000_0000000011111101"; -- 0.018920957286766026
	pesos_i(7424) := b"1111111111111111_1111111111111111_1110110011010110_1110011000010011"; -- -0.07484590557596074
	pesos_i(7425) := b"1111111111111111_1111111111111111_1110100101000000_0011101010011000"; -- -0.08886369502858707
	pesos_i(7426) := b"0000000000000000_0000000000000000_0000110000011111_1111000110000010"; -- 0.047362417398090495
	pesos_i(7427) := b"0000000000000000_0000000000000000_0010001001101110_1111111000101001"; -- 0.1345061159631393
	pesos_i(7428) := b"1111111111111111_1111111111111111_1101011000010111_1111000101000111"; -- -0.1636971665342841
	pesos_i(7429) := b"0000000000000000_0000000000000000_0000100010101100_0001011000101111"; -- 0.03387583406447341
	pesos_i(7430) := b"0000000000000000_0000000000000000_0000010101111001_0110101101011000"; -- 0.02138396157644314
	pesos_i(7431) := b"1111111111111111_1111111111111111_1111000010100000_1101001010100011"; -- -0.0600460387554415
	pesos_i(7432) := b"0000000000000000_0000000000000000_0000000011100101_1001101110110110"; -- 0.0035035437319517306
	pesos_i(7433) := b"0000000000000000_0000000000000000_0001001111101110_1110010001111001"; -- 0.07786395973277398
	pesos_i(7434) := b"1111111111111111_1111111111111111_1101010011100111_1111001110100010"; -- -0.16833569798968767
	pesos_i(7435) := b"1111111111111111_1111111111111111_1110100100010000_1111000001001011"; -- -0.08958528673658958
	pesos_i(7436) := b"0000000000000000_0000000000000000_0010010000000100_1011100010100001"; -- 0.1406970398970811
	pesos_i(7437) := b"1111111111111111_1111111111111111_1101101010010100_1000110011000100"; -- -0.1461708089746254
	pesos_i(7438) := b"0000000000000000_0000000000000000_0000000001111001_0000000100101111"; -- 0.0018463840806712865
	pesos_i(7439) := b"0000000000000000_0000000000000000_0010000011110001_1100111001100111"; -- 0.12868967077277424
	pesos_i(7440) := b"1111111111111111_1111111111111111_1101011000111100_0100000000100110"; -- -0.16314314900185103
	pesos_i(7441) := b"0000000000000000_0000000000000000_0010110010000010_1111101000111100"; -- 0.1738735578095431
	pesos_i(7442) := b"0000000000000000_0000000000000000_0010011111111010_1000110110111011"; -- 0.1561668949631914
	pesos_i(7443) := b"0000000000000000_0000000000000000_0001011111110001_1101110101110011"; -- 0.09353431747666968
	pesos_i(7444) := b"1111111111111111_1111111111111111_1111100001110110_0101011010111011"; -- -0.029444293419514673
	pesos_i(7445) := b"1111111111111111_1111111111111111_1101110100101001_0110111000100001"; -- -0.1360865755195647
	pesos_i(7446) := b"0000000000000000_0000000000000000_0010011001000011_1100010100011011"; -- 0.14947158725050042
	pesos_i(7447) := b"0000000000000000_0000000000000000_0000001010111110_0100100000011101"; -- 0.01071596831824476
	pesos_i(7448) := b"1111111111111111_1111111111111111_1100011100001111_1111111001001100"; -- -0.22241221089714977
	pesos_i(7449) := b"1111111111111111_1111111111111111_1101111110110011_0111010101100010"; -- -0.12616793025272316
	pesos_i(7450) := b"1111111111111111_1111111111111111_1101110101001011_1110111001001110"; -- -0.13556013678712264
	pesos_i(7451) := b"0000000000000000_0000000000000000_0000000110010000_1001010001000111"; -- 0.006112353698398569
	pesos_i(7452) := b"1111111111111111_1111111111111111_1110010101100111_1010001000010001"; -- -0.10388743475454165
	pesos_i(7453) := b"0000000000000000_0000000000000000_0001001110101100_1010100000111001"; -- 0.07685328850748531
	pesos_i(7454) := b"1111111111111111_1111111111111111_1111010110011011_1000111100001111"; -- -0.04059511072599095
	pesos_i(7455) := b"0000000000000000_0000000000000000_0001000011001000_1010000011110100"; -- 0.0655613514221158
	pesos_i(7456) := b"0000000000000000_0000000000000000_0001110101101010_0111000110111010"; -- 0.11490546020010914
	pesos_i(7457) := b"0000000000000000_0000000000000000_0000001001100101_0000010000000111"; -- 0.009353877752621259
	pesos_i(7458) := b"0000000000000000_0000000000000000_0001101100110111_0101101011110010"; -- 0.10631340413900006
	pesos_i(7459) := b"0000000000000000_0000000000000000_0001110101011001_1011011101011100"; -- 0.11465021129296868
	pesos_i(7460) := b"0000000000000000_0000000000000000_0001000000010011_0010001011000001"; -- 0.06279198859276496
	pesos_i(7461) := b"1111111111111111_1111111111111111_1110111101101110_0000011001110111"; -- -0.06472739796546399
	pesos_i(7462) := b"0000000000000000_0000000000000000_0010001110011110_0000001101000010"; -- 0.13912983274727955
	pesos_i(7463) := b"0000000000000000_0000000000000000_0001010000100001_0010000101101011"; -- 0.07863053191256272
	pesos_i(7464) := b"1111111111111111_1111111111111111_1101100010010011_0010100100010100"; -- -0.15400450959234457
	pesos_i(7465) := b"0000000000000000_0000000000000000_0001000010101111_0001001011100011"; -- 0.06517141380927371
	pesos_i(7466) := b"1111111111111111_1111111111111111_1101001110100001_0000000001010100"; -- -0.17332456549248096
	pesos_i(7467) := b"0000000000000000_0000000000000000_0000101011010101_1111011111001000"; -- 0.042327391055470974
	pesos_i(7468) := b"0000000000000000_0000000000000000_0000111001110001_1110001011110010"; -- 0.056425270260279034
	pesos_i(7469) := b"1111111111111111_1111111111111111_1101101000001100_1100001110110000"; -- -0.14824273067266772
	pesos_i(7470) := b"1111111111111111_1111111111111111_1111011001011011_0001111101111100"; -- -0.03767207359227226
	pesos_i(7471) := b"1111111111111111_1111111111111111_1111110100110100_0001100100110001"; -- -0.010923791500675085
	pesos_i(7472) := b"0000000000000000_0000000000000000_0000100111110001_1101101001111001"; -- 0.03884664009570102
	pesos_i(7473) := b"1111111111111111_1111111111111111_1111110001110000_0101111001000000"; -- -0.013910397921416727
	pesos_i(7474) := b"0000000000000000_0000000000000000_0001001000011001_1000111011111101"; -- 0.07070249258568906
	pesos_i(7475) := b"0000000000000000_0000000000000000_0000000100101111_0100101001100000"; -- 0.004627846220319306
	pesos_i(7476) := b"0000000000000000_0000000000000000_0001110111100001_0100110110101111"; -- 0.11671910782399285
	pesos_i(7477) := b"0000000000000000_0000000000000000_0010101111001111_0111011101011000"; -- 0.17113443266978923
	pesos_i(7478) := b"0000000000000000_0000000000000000_0000111111011000_0000100011110111"; -- 0.06189018279399651
	pesos_i(7479) := b"0000000000000000_0000000000000000_0001100001000101_1001000011111100"; -- 0.09481149814641164
	pesos_i(7480) := b"0000000000000000_0000000000000000_0000000111000011_0110001000111110"; -- 0.006887569642320235
	pesos_i(7481) := b"1111111111111111_1111111111111111_1110111001000000_0001001110111000"; -- -0.06933476228296191
	pesos_i(7482) := b"0000000000000000_0000000000000000_0000011000111010_0000011001000101"; -- 0.024322883361032204
	pesos_i(7483) := b"1111111111111111_1111111111111111_1111110100011101_0000001000000110"; -- -0.011276124465307805
	pesos_i(7484) := b"0000000000000000_0000000000000000_0010010100000010_1100111100000110"; -- 0.1445741071501736
	pesos_i(7485) := b"1111111111111111_1111111111111111_1110101000011011_1001101100110110"; -- -0.0855162614997072
	pesos_i(7486) := b"1111111111111111_1111111111111111_1110000011111111_0101110110011011"; -- -0.12110342948313994
	pesos_i(7487) := b"0000000000000000_0000000000000000_0001110110100010_0101110010011011"; -- 0.1157586936022581
	pesos_i(7488) := b"1111111111111111_1111111111111111_1111100110001110_0111110110011110"; -- -0.025169514474327637
	pesos_i(7489) := b"1111111111111111_1111111111111111_1110000100000111_1111100010000011"; -- -0.12097212607510695
	pesos_i(7490) := b"0000000000000000_0000000000000000_0000111011001110_1101111100001011"; -- 0.05784410492584053
	pesos_i(7491) := b"0000000000000000_0000000000000000_0010101011100100_0101111101110101"; -- 0.16754719350850814
	pesos_i(7492) := b"1111111111111111_1111111111111111_1111000111101100_1011001100000110"; -- -0.054982005228957756
	pesos_i(7493) := b"1111111111111111_1111111111111111_1110101101111001_1110011011111001"; -- -0.08017116950593188
	pesos_i(7494) := b"1111111111111111_1111111111111111_1101111010010010_1011111110010110"; -- -0.13057329746319174
	pesos_i(7495) := b"0000000000000000_0000000000000000_0010000011100010_1010010011001011"; -- 0.12845830883646325
	pesos_i(7496) := b"0000000000000000_0000000000000000_0000111101101101_0010010110101010"; -- 0.060259203038055216
	pesos_i(7497) := b"0000000000000000_0000000000000000_0001101000110001_1111100101110111"; -- 0.10232504988040796
	pesos_i(7498) := b"1111111111111111_1111111111111111_1101011110010011_0101000001011001"; -- -0.1579084189989091
	pesos_i(7499) := b"1111111111111111_1111111111111111_1110000000100110_0101101110001101"; -- -0.12441470917836257
	pesos_i(7500) := b"1111111111111111_1111111111111111_1111011001110111_1011101100010101"; -- -0.037235553189784776
	pesos_i(7501) := b"1111111111111111_1111111111111111_1110101000010000_1110101111010111"; -- -0.08567930231471406
	pesos_i(7502) := b"0000000000000000_0000000000000000_0010100010100110_0111001110100110"; -- 0.15878985212013544
	pesos_i(7503) := b"0000000000000000_0000000000000000_0001010001011111_1111011110111000"; -- 0.07958935009392172
	pesos_i(7504) := b"1111111111111111_1111111111111111_1101011100010000_0110001000010000"; -- -0.15990626429935054
	pesos_i(7505) := b"0000000000000000_0000000000000000_0010110010010011_1000001101010101"; -- 0.17412586989019105
	pesos_i(7506) := b"0000000000000000_0000000000000000_0001111101101011_1011000101001010"; -- 0.12273700776441739
	pesos_i(7507) := b"1111111111111111_1111111111111111_1111111011011001_1110100110100101"; -- -0.004487416552674266
	pesos_i(7508) := b"0000000000000000_0000000000000000_0001000010101010_0100010110100110"; -- 0.0650981456216405
	pesos_i(7509) := b"0000000000000000_0000000000000000_0010000001111010_0011001111000001"; -- 0.12686465697630492
	pesos_i(7510) := b"0000000000000000_0000000000000000_0010000000000101_0101111110001000"; -- 0.12508198816485994
	pesos_i(7511) := b"0000000000000000_0000000000000000_0001101010001001_0001000001000011"; -- 0.10365392342846672
	pesos_i(7512) := b"1111111111111111_1111111111111111_1111100000101111_1101000000110100"; -- -0.030520426938700194
	pesos_i(7513) := b"1111111111111111_1111111111111111_1111000101000000_1011111001110000"; -- -0.05760583652490617
	pesos_i(7514) := b"1111111111111111_1111111111111111_1111101001010101_1000110010101000"; -- -0.022132119214937584
	pesos_i(7515) := b"1111111111111111_1111111111111111_1110100011010100_1111100100111010"; -- -0.09050028169402048
	pesos_i(7516) := b"0000000000000000_0000000000000000_0001010011011101_1011101100001010"; -- 0.08150834072289109
	pesos_i(7517) := b"1111111111111111_1111111111111111_1111011101001111_0001100100010111"; -- -0.033949310303759354
	pesos_i(7518) := b"1111111111111111_1111111111111111_1111100001000111_0100100100010011"; -- -0.03016227043130454
	pesos_i(7519) := b"1111111111111111_1111111111111111_1111110101110010_0010111111011001"; -- -0.009976396162323264
	pesos_i(7520) := b"1111111111111111_1111111111111111_1110110001011011_0101101010101110"; -- -0.07673104524741854
	pesos_i(7521) := b"0000000000000000_0000000000000000_0001011010001111_0011011000011100"; -- 0.0881227320701413
	pesos_i(7522) := b"0000000000000000_0000000000000000_0000011110111100_1011111010010111"; -- 0.030223762272230958
	pesos_i(7523) := b"1111111111111111_1111111111111111_1101101000110111_0000101010110111"; -- -0.14759762783940986
	pesos_i(7524) := b"0000000000000000_0000000000000000_0010100001000001_1101010111110001"; -- 0.1572545731761371
	pesos_i(7525) := b"1111111111111111_1111111111111111_1101011100001110_0001101101110110"; -- -0.15994099013610072
	pesos_i(7526) := b"0000000000000000_0000000000000000_0001011101001100_0111000111000011"; -- 0.09101019878980353
	pesos_i(7527) := b"1111111111111111_1111111111111111_1111101101001110_0010011110111110"; -- -0.018338695542104766
	pesos_i(7528) := b"1111111111111111_1111111111111111_1110101000110101_1111001110000010"; -- -0.08511427009185113
	pesos_i(7529) := b"1111111111111111_1111111111111111_1101110010011011_0100001000110100"; -- -0.13825594175189232
	pesos_i(7530) := b"1111111111111111_1111111111111111_1111111111010001_0111111011010010"; -- -0.0007096040639022437
	pesos_i(7531) := b"0000000000000000_0000000000000000_0010010001000111_0010111011010100"; -- 0.1417111651857448
	pesos_i(7532) := b"1111111111111111_1111111111111111_1111101001011110_0110011000111010"; -- -0.021997080612177783
	pesos_i(7533) := b"1111111111111111_1111111111111111_1110111100000100_0100100000111011"; -- -0.06634090950443089
	pesos_i(7534) := b"0000000000000000_0000000000000000_0000100011001010_1010000101010010"; -- 0.03434189093694014
	pesos_i(7535) := b"0000000000000000_0000000000000000_0001001110010001_1100000000100100"; -- 0.0764427269040011
	pesos_i(7536) := b"0000000000000000_0000000000000000_0010001011001110_0100111011010010"; -- 0.1359605085681321
	pesos_i(7537) := b"1111111111111111_1111111111111111_1110000111100100_1010110000100101"; -- -0.11760448537271538
	pesos_i(7538) := b"1111111111111111_1111111111111111_1111000010000001_0100011110111101"; -- -0.06052734020608327
	pesos_i(7539) := b"1111111111111111_1111111111111111_1111111000010100_0100000001010010"; -- -0.007503490438964498
	pesos_i(7540) := b"1111111111111111_1111111111111111_1111100110001111_0101010001110101"; -- -0.02515670915570692
	pesos_i(7541) := b"1111111111111111_1111111111111111_1110001010000010_0000001000010111"; -- -0.11520373275225719
	pesos_i(7542) := b"1111111111111111_1111111111111111_1111111000101011_0000100000010001"; -- -0.007155891295813142
	pesos_i(7543) := b"1111111111111111_1111111111111111_1101100011010010_0010000110100000"; -- -0.1530436501515382
	pesos_i(7544) := b"1111111111111111_1111111111111111_1101101111111000_1011110010011011"; -- -0.1407358284819447
	pesos_i(7545) := b"0000000000000000_0000000000000000_0001010100001110_1110100111100110"; -- 0.0822588145827655
	pesos_i(7546) := b"1111111111111111_1111111111111111_1101110010000011_0100010010000100"; -- -0.13862201484172448
	pesos_i(7547) := b"1111111111111111_1111111111111111_1111101010011011_1110001100010001"; -- -0.021058853558164108
	pesos_i(7548) := b"1111111111111111_1111111111111111_1111101011111010_0010000011000111"; -- -0.01962084899417478
	pesos_i(7549) := b"1111111111111111_1111111111111111_1110011111011010_1101010111010010"; -- -0.09431708928992474
	pesos_i(7550) := b"1111111111111111_1111111111111111_1111111010000110_0110010100111101"; -- -0.005761787905969135
	pesos_i(7551) := b"1111111111111111_1111111111111111_1111011111000010_0011101011010010"; -- -0.03219253905132679
	pesos_i(7552) := b"0000000000000000_0000000000000000_0001101011000110_1011111010010001"; -- 0.10459509886655141
	pesos_i(7553) := b"1111111111111111_1111111111111111_1101011110001000_1010111000100111"; -- -0.15807067439627884
	pesos_i(7554) := b"1111111111111111_1111111111111111_1111010111000000_1001000011011100"; -- -0.04003042829671764
	pesos_i(7555) := b"0000000000000000_0000000000000000_0000000110110011_1011001100110001"; -- 0.0066482539259704815
	pesos_i(7556) := b"0000000000000000_0000000000000000_0001111000100100_0000110110101110"; -- 0.11773763176890176
	pesos_i(7557) := b"1111111111111111_1111111111111111_1111111010001001_1101001001010110"; -- -0.005709508924611822
	pesos_i(7558) := b"0000000000000000_0000000000000000_0000000000110100_0010111001101011"; -- 0.0007962238405817853
	pesos_i(7559) := b"1111111111111111_1111111111111111_1110011000100000_0100101000011110"; -- -0.101069801049544
	pesos_i(7560) := b"1111111111111111_1111111111111111_1101101000000000_1101100001110000"; -- -0.14842459937957195
	pesos_i(7561) := b"1111111111111111_1111111111111111_1101100000100010_1111110111100100"; -- -0.15571606806363023
	pesos_i(7562) := b"1111111111111111_1111111111111111_1110110010111110_0001111111101001"; -- -0.0752239281024284
	pesos_i(7563) := b"0000000000000000_0000000000000000_0000000001101011_0000110111010000"; -- 0.0016335138183357922
	pesos_i(7564) := b"1111111111111111_1111111111111111_1110010010011010_1101000100010011"; -- -0.10701268467550425
	pesos_i(7565) := b"0000000000000000_0000000000000000_0001010001111011_0001001010001011"; -- 0.08000293635725826
	pesos_i(7566) := b"1111111111111111_1111111111111111_1110111010001111_0000111000111111"; -- -0.06812964393079741
	pesos_i(7567) := b"0000000000000000_0000000000000000_0001111000011001_1110100111010110"; -- 0.11758290737551756
	pesos_i(7568) := b"0000000000000000_0000000000000000_0010010111101100_1000101001010000"; -- 0.1481405682492354
	pesos_i(7569) := b"0000000000000000_0000000000000000_0010010101101111_1111000111001000"; -- 0.14623938695609712
	pesos_i(7570) := b"0000000000000000_0000000000000000_0000001010101010_0011110011101010"; -- 0.0104101248734515
	pesos_i(7571) := b"0000000000000000_0000000000000000_0010010111010011_0111100000100000"; -- 0.14775801442186537
	pesos_i(7572) := b"0000000000000000_0000000000000000_0001011000010111_1011010100000010"; -- 0.08629924112742127
	pesos_i(7573) := b"0000000000000000_0000000000000000_0010100011111001_1011000111101010"; -- 0.16006004301655619
	pesos_i(7574) := b"0000000000000000_0000000000000000_0010010001110110_1101001011010111"; -- 0.14243810410906446
	pesos_i(7575) := b"0000000000000000_0000000000000000_0000001010111001_0010001110011011"; -- 0.010637498141200477
	pesos_i(7576) := b"0000000000000000_0000000000000000_0010101010110101_0010010100001000"; -- 0.16682654796360283
	pesos_i(7577) := b"0000000000000000_0000000000000000_0001110001101101_0101110001011111"; -- 0.11104371370288521
	pesos_i(7578) := b"0000000000000000_0000000000000000_0001110110110111_0111001001001000"; -- 0.11608042019962048
	pesos_i(7579) := b"1111111111111111_1111111111111111_1111100010001101_1000111010001111"; -- -0.029090013573969637
	pesos_i(7580) := b"0000000000000000_0000000000000000_0010001001110111_1101011100010000"; -- 0.1346411145579428
	pesos_i(7581) := b"1111111111111111_1111111111111111_1111101011110010_0100011010111010"; -- -0.019740657438863645
	pesos_i(7582) := b"0000000000000000_0000000000000000_0001001000111001_1111110100101011"; -- 0.07119734103159571
	pesos_i(7583) := b"1111111111111111_1111111111111111_1111100001111000_0000010001001000"; -- -0.029418690171383294
	pesos_i(7584) := b"0000000000000000_0000000000000000_0010101001000011_1100010011010100"; -- 0.16509657065484565
	pesos_i(7585) := b"0000000000000000_0000000000000000_0000101101100110_0111000111110100"; -- 0.044531938681446115
	pesos_i(7586) := b"1111111111111111_1111111111111111_1101111010000011_0011110000111010"; -- -0.13081000876664173
	pesos_i(7587) := b"1111111111111111_1111111111111111_1110001011010001_0111110011010011"; -- -0.11399097298107187
	pesos_i(7588) := b"1111111111111111_1111111111111111_1111010010010100_1000011100100001"; -- -0.0446086450171803
	pesos_i(7589) := b"1111111111111111_1111111111111111_1110000010000001_1000010111101010"; -- -0.12302363433644369
	pesos_i(7590) := b"0000000000000000_0000000000000000_0000000101100100_1011001001001001"; -- 0.005442755539410509
	pesos_i(7591) := b"0000000000000000_0000000000000000_0000100001001001_1011100010110110"; -- 0.03237490113542851
	pesos_i(7592) := b"1111111111111111_1111111111111111_1110101011110001_1110101001000001"; -- -0.08224616926928463
	pesos_i(7593) := b"0000000000000000_0000000000000000_0000110110101101_0100100101001110"; -- 0.05342538986731552
	pesos_i(7594) := b"0000000000000000_0000000000000000_0000110000110001_1100111110010010"; -- 0.04763505272848889
	pesos_i(7595) := b"0000000000000000_0000000000000000_0000010010101011_0010111111011100"; -- 0.018237105471345706
	pesos_i(7596) := b"0000000000000000_0000000000000000_0010001011011010_1101101001011101"; -- 0.13615193144331703
	pesos_i(7597) := b"0000000000000000_0000000000000000_0001100100000110_0110100100000010"; -- 0.09775406159790181
	pesos_i(7598) := b"1111111111111111_1111111111111111_1111101100010100_1001000111111110"; -- -0.019217372481284793
	pesos_i(7599) := b"1111111111111111_1111111111111111_1110000111000011_0100111011011101"; -- -0.11811358540730614
	pesos_i(7600) := b"0000000000000000_0000000000000000_0000111010000001_0000001100000111"; -- 0.05665606415684574
	pesos_i(7601) := b"1111111111111111_1111111111111111_1110110010110111_0010110111011110"; -- -0.07532990770720019
	pesos_i(7602) := b"0000000000000000_0000000000000000_0010000101000010_1001100110101000"; -- 0.12992248874703613
	pesos_i(7603) := b"1111111111111111_1111111111111111_1111011000100000_0011111011001011"; -- -0.03857047608849233
	pesos_i(7604) := b"0000000000000000_0000000000000000_0001111001100110_1011010001110011"; -- 0.11875465219811623
	pesos_i(7605) := b"1111111111111111_1111111111111111_1111100111001101_1000100011100010"; -- -0.024207539330734367
	pesos_i(7606) := b"1111111111111111_1111111111111111_1101001001111100_1010001100001110"; -- -0.17778569135625652
	pesos_i(7607) := b"1111111111111111_1111111111111111_1110110100000000_1101011101011100"; -- -0.07420591358647909
	pesos_i(7608) := b"0000000000000000_0000000000000000_0000100101101000_1000010000100100"; -- 0.03675104023573478
	pesos_i(7609) := b"1111111111111111_1111111111111111_1110001000011100_1110011001111000"; -- -0.11674651681345673
	pesos_i(7610) := b"0000000000000000_0000000000000000_0001110010110110_1011100110000001"; -- 0.11216315657050446
	pesos_i(7611) := b"1111111111111111_1111111111111111_1110110101010000_0100111101001011"; -- -0.07299332070255822
	pesos_i(7612) := b"1111111111111111_1111111111111111_1111001111101111_1010100000100101"; -- -0.04712437718870929
	pesos_i(7613) := b"0000000000000000_0000000000000000_0000100010110010_0000100011000001"; -- 0.0339665863062356
	pesos_i(7614) := b"0000000000000000_0000000000000000_0000000101001001_0111111100000111"; -- 0.0050277129974657655
	pesos_i(7615) := b"0000000000000000_0000000000000000_0001000100101010_0110100000011100"; -- 0.06705332460868803
	pesos_i(7616) := b"0000000000000000_0000000000000000_0001011101111011_0111010001011011"; -- 0.09172751630054285
	pesos_i(7617) := b"1111111111111111_1111111111111111_1101001001111000_0011000111001011"; -- -0.17785347734932275
	pesos_i(7618) := b"1111111111111111_1111111111111111_1101010101111101_0000110000100111"; -- -0.1660606770034902
	pesos_i(7619) := b"0000000000000000_0000000000000000_0000100101111101_0000111001001001"; -- 0.03706445019925724
	pesos_i(7620) := b"0000000000000000_0000000000000000_0001100100011101_1011010000010111"; -- 0.09810948895928773
	pesos_i(7621) := b"0000000000000000_0000000000000000_0000101111111010_0110000100100111"; -- 0.046789237994321116
	pesos_i(7622) := b"0000000000000000_0000000000000000_0000101011101000_0100010011000001"; -- 0.04260663710194132
	pesos_i(7623) := b"1111111111111111_1111111111111111_1111101000101111_1111001010001110"; -- -0.022705879431327566
	pesos_i(7624) := b"0000000000000000_0000000000000000_0000111110100111_1010011101001111"; -- 0.06115194022242903
	pesos_i(7625) := b"0000000000000000_0000000000000000_0000010000100101_1100000001111011"; -- 0.0162010478793095
	pesos_i(7626) := b"0000000000000000_0000000000000000_0000110011110110_1100110001011011"; -- 0.05064084257159845
	pesos_i(7627) := b"1111111111111111_1111111111111111_1101010101010111_1111001100000111"; -- -0.16662674982045148
	pesos_i(7628) := b"1111111111111111_1111111111111111_1110101011010110_1100000011011101"; -- -0.08266062348257298
	pesos_i(7629) := b"1111111111111111_1111111111111111_1111000000011100_1111000110000100"; -- -0.06205835847798882
	pesos_i(7630) := b"0000000000000000_0000000000000000_0000000001111000_0111011010111101"; -- 0.0018381321478135957
	pesos_i(7631) := b"0000000000000000_0000000000000000_0010000001000100_0001101100010000"; -- 0.12603921076482652
	pesos_i(7632) := b"0000000000000000_0000000000000000_0000001111001101_0011111111101101"; -- 0.014850611936999825
	pesos_i(7633) := b"1111111111111111_1111111111111111_1101110100001110_1100100111110110"; -- -0.13649308904667537
	pesos_i(7634) := b"1111111111111111_1111111111111111_1111001110010110_1000011001000101"; -- -0.048484428493538824
	pesos_i(7635) := b"1111111111111111_1111111111111111_1110001110010100_1001011001101101"; -- -0.11101398323528847
	pesos_i(7636) := b"0000000000000000_0000000000000000_0000111000111101_1000000001000011"; -- 0.055625931067124504
	pesos_i(7637) := b"0000000000000000_0000000000000000_0010011100100111_1101001110111111"; -- 0.15295146391536685
	pesos_i(7638) := b"0000000000000000_0000000000000000_0000001011011001_0011011100111011"; -- 0.011126949184449543
	pesos_i(7639) := b"1111111111111111_1111111111111111_1110101110000110_1100101100111111"; -- -0.07997445787242866
	pesos_i(7640) := b"1111111111111111_1111111111111111_1100111110001001_0101001010001101"; -- -0.1893108754919276
	pesos_i(7641) := b"1111111111111111_1111111111111111_1110010011100000_0000100100110110"; -- -0.10595648219067809
	pesos_i(7642) := b"1111111111111111_1111111111111111_1111011011100011_0011111111011100"; -- -0.03559494846608529
	pesos_i(7643) := b"1111111111111111_1111111111111111_1111010100101011_1101100010100110"; -- -0.04229970889538112
	pesos_i(7644) := b"0000000000000000_0000000000000000_0001110000010110_0111100101010010"; -- 0.10971792454285612
	pesos_i(7645) := b"1111111111111111_1111111111111111_1110001010110001_0011010101001011"; -- -0.11448351793426322
	pesos_i(7646) := b"0000000000000000_0000000000000000_0001011010100101_1011000111101101"; -- 0.08846580549590471
	pesos_i(7647) := b"1111111111111111_1111111111111111_1111100111000110_0011001100101100"; -- -0.024319459570805113
	pesos_i(7648) := b"0000000000000000_0000000000000000_0010101110111010_0011110101000010"; -- 0.17081053611585031
	pesos_i(7649) := b"0000000000000000_0000000000000000_0000111001101000_1011010011110000"; -- 0.056285198874220045
	pesos_i(7650) := b"1111111111111111_1111111111111111_1111001010000111_1000010011100111"; -- -0.0526196419051458
	pesos_i(7651) := b"0000000000000000_0000000000000000_0001000001010011_1000010111110010"; -- 0.0637744632359685
	pesos_i(7652) := b"0000000000000000_0000000000000000_0010000000110100_0100101010001101"; -- 0.12579790049367093
	pesos_i(7653) := b"0000000000000000_0000000000000000_0001111011101010_0111010101000111"; -- 0.12076504681881485
	pesos_i(7654) := b"1111111111111111_1111111111111111_1101111101010011_0111001001001101"; -- -0.12763295758106546
	pesos_i(7655) := b"1111111111111111_1111111111111111_1110001100000011_1100110000011000"; -- -0.11322330875364883
	pesos_i(7656) := b"1111111111111111_1111111111111111_1111110010100111_0001000110010110"; -- -0.013075733932436717
	pesos_i(7657) := b"0000000000000000_0000000000000000_0010001000100110_1101110000010000"; -- 0.1334054507478129
	pesos_i(7658) := b"0000000000000000_0000000000000000_0010000001111100_0111011110010010"; -- 0.12689921677956995
	pesos_i(7659) := b"1111111111111111_1111111111111111_1111101101001100_1001011000111011"; -- -0.018362627492206966
	pesos_i(7660) := b"0000000000000000_0000000000000000_0001110001011000_1011110100100111"; -- 0.11072904774191066
	pesos_i(7661) := b"1111111111111111_1111111111111111_1110010010110011_0000011101100000"; -- -0.10664323717959985
	pesos_i(7662) := b"1111111111111111_1111111111111111_1110101011111010_1101000101001101"; -- -0.08211032748637347
	pesos_i(7663) := b"1111111111111111_1111111111111111_1111011011001101_0001001011001100"; -- -0.035933327758306356
	pesos_i(7664) := b"1111111111111111_1111111111111111_1111111011110010_1000010011010101"; -- -0.0041119556934643975
	pesos_i(7665) := b"0000000000000000_0000000000000000_0010001111000110_1110111100111001"; -- 0.1397542489071277
	pesos_i(7666) := b"1111111111111111_1111111111111111_1101111110001111_0101001011001010"; -- -0.12671930850651617
	pesos_i(7667) := b"0000000000000000_0000000000000000_0001100101011000_1001001111010001"; -- 0.09900783402122541
	pesos_i(7668) := b"1111111111111111_1111111111111111_1110111110100110_0011110101100100"; -- -0.06386963182182288
	pesos_i(7669) := b"0000000000000000_0000000000000000_0000111110000000_1110111011100101"; -- 0.06056111414498419
	pesos_i(7670) := b"1111111111111111_1111111111111111_1111110101111101_0110001011001111"; -- -0.009805511955738469
	pesos_i(7671) := b"1111111111111111_1111111111111111_1110001111101111_1011111110010101"; -- -0.10962298026543647
	pesos_i(7672) := b"1111111111111111_1111111111111111_1101010101101010_0000010101100100"; -- -0.16635099707377213
	pesos_i(7673) := b"1111111111111111_1111111111111111_1101111100011111_1010101101000000"; -- -0.12842302029844097
	pesos_i(7674) := b"0000000000000000_0000000000000000_0001101110110001_1111110101001001"; -- 0.10818465270475539
	pesos_i(7675) := b"1111111111111111_1111111111111111_1111011001011100_0111111111110110"; -- -0.037651064456087326
	pesos_i(7676) := b"0000000000000000_0000000000000000_0010000110011000_0111011110011101"; -- 0.13123271546672433
	pesos_i(7677) := b"1111111111111111_1111111111111111_1110110000100010_0011101010100100"; -- -0.07760270592332352
	pesos_i(7678) := b"1111111111111111_1111111111111111_1110011101110101_1111000111100000"; -- -0.09585655490191683
	pesos_i(7679) := b"0000000000000000_0000000000000000_0010001010010011_1110001001010110"; -- 0.13506903266231035
	pesos_i(7680) := b"0000000000000000_0000000000000000_0010110001010101_1010001100110001"; -- 0.17318172412324004
	pesos_i(7681) := b"1111111111111111_1111111111111111_1111100101000110_1001100100111010"; -- -0.02626650172899994
	pesos_i(7682) := b"0000000000000000_0000000000000000_0010100111000011_0001001101100111"; -- 0.16313287032898263
	pesos_i(7683) := b"0000000000000000_0000000000000000_0000101001110010_0000010101011000"; -- 0.040802320420766945
	pesos_i(7684) := b"1111111111111111_1111111111111111_1110011110001011_0001000000101000"; -- -0.09553431533113325
	pesos_i(7685) := b"0000000000000000_0000000000000000_0010101010011111_0100101101110000"; -- 0.16649314395538403
	pesos_i(7686) := b"1111111111111111_1111111111111111_1110110010011101_1011111000000010"; -- -0.07571804479644555
	pesos_i(7687) := b"1111111111111111_1111111111111111_1111011111100001_0111000110100010"; -- -0.03171624943897461
	pesos_i(7688) := b"0000000000000000_0000000000000000_0001000101110101_1011001010100011"; -- 0.06820217589245593
	pesos_i(7689) := b"0000000000000000_0000000000000000_0000101010111000_1110011100110101"; -- 0.04188389824908031
	pesos_i(7690) := b"0000000000000000_0000000000000000_0001110101110101_1111111001111101"; -- 0.11508169708440238
	pesos_i(7691) := b"0000000000000000_0000000000000000_0000001100110101_0100010001010100"; -- 0.012531538451207707
	pesos_i(7692) := b"0000000000000000_0000000000000000_0001111110001001_1000000000111000"; -- 0.12319184655517747
	pesos_i(7693) := b"1111111111111111_1111111111111111_1101010100001000_0111101010111111"; -- -0.16783936345597766
	pesos_i(7694) := b"0000000000000000_0000000000000000_0000010011001101_1000101100010011"; -- 0.01876134125273534
	pesos_i(7695) := b"0000000000000000_0000000000000000_0001000101110001_1100110000001000"; -- 0.0681426544483309
	pesos_i(7696) := b"0000000000000000_0000000000000000_0000011001110001_0101000010011110"; -- 0.02516654838927837
	pesos_i(7697) := b"1111111111111111_1111111111111111_1110000011001011_1011001010010110"; -- -0.12189182122133532
	pesos_i(7698) := b"1111111111111111_1111111111111111_1101101110010110_0010110101001001"; -- -0.1422397325332608
	pesos_i(7699) := b"1111111111111111_1111111111111111_1111010110010101_0111100101100110"; -- -0.040687954452830986
	pesos_i(7700) := b"1111111111111111_1111111111111111_1110111100001101_0000111010101100"; -- -0.06620701121849125
	pesos_i(7701) := b"1111111111111111_1111111111111111_1101011100111111_0100111000101011"; -- -0.15919028702347615
	pesos_i(7702) := b"0000000000000000_0000000000000000_0001111111000000_1111001000100001"; -- 0.1240378695223945
	pesos_i(7703) := b"0000000000000000_0000000000000000_0001111001100111_0000011010000110"; -- 0.11875954401105362
	pesos_i(7704) := b"0000000000000000_0000000000000000_0000111100110111_1111111110000001"; -- 0.059448212711825314
	pesos_i(7705) := b"1111111111111111_1111111111111111_1111010100110000_0100000110110110"; -- -0.04223241149857734
	pesos_i(7706) := b"1111111111111111_1111111111111111_1110010001111101_0000111010110011"; -- -0.10746677525845039
	pesos_i(7707) := b"1111111111111111_1111111111111111_1101010111011010_0101101101011011"; -- -0.16463688873351603
	pesos_i(7708) := b"0000000000000000_0000000000000000_0001101110011111_1110110100110110"; -- 0.107909036389859
	pesos_i(7709) := b"1111111111111111_1111111111111111_1110000110111110_1111110101001011"; -- -0.11817948255483447
	pesos_i(7710) := b"0000000000000000_0000000000000000_0000100111110000_0011110101010001"; -- 0.03882201401855239
	pesos_i(7711) := b"1111111111111111_1111111111111111_1110000100001001_1101101000001001"; -- -0.12094342504518914
	pesos_i(7712) := b"1111111111111111_1111111111111111_1101010100010100_1010100100010011"; -- -0.1676534965090695
	pesos_i(7713) := b"0000000000000000_0000000000000000_0000111100001011_0111010110111110"; -- 0.0587686147011229
	pesos_i(7714) := b"0000000000000000_0000000000000000_0010110011011000_0010110001000000"; -- 0.17517353603930605
	pesos_i(7715) := b"0000000000000000_0000000000000000_0000110000101100_0101011111101010"; -- 0.04755162675348572
	pesos_i(7716) := b"0000000000000000_0000000000000000_0000100000110111_0010100000011111"; -- 0.032091624886296057
	pesos_i(7717) := b"0000000000000000_0000000000000000_0000111010011011_0110101011111111"; -- 0.057058989702823304
	pesos_i(7718) := b"1111111111111111_1111111111111111_1111011010111110_0101001011000100"; -- -0.03615839686143729
	pesos_i(7719) := b"1111111111111111_1111111111111111_1111111101010110_0111111110010010"; -- -0.002586390406585065
	pesos_i(7720) := b"1111111111111111_1111111111111111_1101011110011011_1110111001111001"; -- -0.15777692361041587
	pesos_i(7721) := b"0000000000000000_0000000000000000_0001000000100000_1111011110001111"; -- 0.06300303680279444
	pesos_i(7722) := b"0000000000000000_0000000000000000_0010011001001001_0100001101111111"; -- 0.14955541479507614
	pesos_i(7723) := b"1111111111111111_1111111111111111_1111010000100011_1111010000000100"; -- -0.04632639800163332
	pesos_i(7724) := b"1111111111111111_1111111111111111_1110010101101110_1010100101110100"; -- -0.10378018294090785
	pesos_i(7725) := b"1111111111111111_1111111111111111_1111100110011111_1001000111000101"; -- -0.024908914033467334
	pesos_i(7726) := b"0000000000000000_0000000000000000_0001111110101111_0001010000011001"; -- 0.12376523602013567
	pesos_i(7727) := b"1111111111111111_1111111111111111_1111111100010011_0011011010101100"; -- -0.0036130743072050327
	pesos_i(7728) := b"0000000000000000_0000000000000000_0001011010110111_0110111100110111"; -- 0.08873648732134834
	pesos_i(7729) := b"0000000000000000_0000000000000000_0000000000011111_0001000100011000"; -- 0.00047404126780225327
	pesos_i(7730) := b"1111111111111111_1111111111111111_1110100010101010_1001011101010001"; -- -0.09114698681036132
	pesos_i(7731) := b"1111111111111111_1111111111111111_1111000110000111_1101011001101010"; -- -0.05652103341716461
	pesos_i(7732) := b"0000000000000000_0000000000000000_0010001010111100_1110100110011011"; -- 0.13569507632642597
	pesos_i(7733) := b"1111111111111111_1111111111111111_1101001011010110_1010010101111101"; -- -0.1764122553366308
	pesos_i(7734) := b"1111111111111111_1111111111111111_1111011100011010_0111100010011000"; -- -0.03475233363363175
	pesos_i(7735) := b"1111111111111111_1111111111111111_1111101001001110_0011001011000101"; -- -0.022244288342461206
	pesos_i(7736) := b"0000000000000000_0000000000000000_0010011101100000_1100001101101111"; -- 0.15382024241165707
	pesos_i(7737) := b"1111111111111111_1111111111111111_1101101111100001_0001001000110000"; -- -0.14109693849372829
	pesos_i(7738) := b"0000000000000000_0000000000000000_0000100011010001_0111111110100010"; -- 0.03444669442605618
	pesos_i(7739) := b"0000000000000000_0000000000000000_0000111011001101_0001111101100100"; -- 0.05781742269251853
	pesos_i(7740) := b"1111111111111111_1111111111111111_1110011100110101_0101010010011001"; -- -0.09684249188139721
	pesos_i(7741) := b"0000000000000000_0000000000000000_0010100101111110_1010001010110101"; -- 0.16208855553814752
	pesos_i(7742) := b"1111111111111111_1111111111111111_1110101101110001_0101010101100010"; -- -0.08030191765124657
	pesos_i(7743) := b"1111111111111111_1111111111111111_1111100001110001_0011001101110001"; -- -0.029522690690951828
	pesos_i(7744) := b"0000000000000000_0000000000000000_0000110000111001_1111101101000111"; -- 0.04775972822411245
	pesos_i(7745) := b"1111111111111111_1111111111111111_1101111101010011_0101000000010111"; -- -0.12763499671719894
	pesos_i(7746) := b"0000000000000000_0000000000000000_0001000000001111_1100010100101101"; -- 0.06274063435695887
	pesos_i(7747) := b"0000000000000000_0000000000000000_0010100000110100_1011010101111000"; -- 0.1570542734735634
	pesos_i(7748) := b"0000000000000000_0000000000000000_0001001110111001_1000011001110110"; -- 0.07704964044599218
	pesos_i(7749) := b"0000000000000000_0000000000000000_0010100110110000_0011110110010000"; -- 0.16284546636792463
	pesos_i(7750) := b"1111111111111111_1111111111111111_1111100111111000_1100011100001010"; -- -0.02354770669589271
	pesos_i(7751) := b"0000000000000000_0000000000000000_0001010000110111_1111000100010001"; -- 0.07897860195956158
	pesos_i(7752) := b"1111111111111111_1111111111111111_1111100100010011_0010000110100011"; -- -0.02705182800840903
	pesos_i(7753) := b"0000000000000000_0000000000000000_0001000101011111_1110100100110100"; -- 0.06786973486858178
	pesos_i(7754) := b"0000000000000000_0000000000000000_0001010001000011_1111111001001110"; -- 0.07916249670720538
	pesos_i(7755) := b"0000000000000000_0000000000000000_0010011110110101_1011010010000111"; -- 0.15511635106881505
	pesos_i(7756) := b"1111111111111111_1111111111111111_1101111111111110_1001101111110000"; -- -0.12502122289837653
	pesos_i(7757) := b"0000000000000000_0000000000000000_0001111010010000_0110010110111110"; -- 0.11939083004289422
	pesos_i(7758) := b"1111111111111111_1111111111111111_1111111110010011_1101011010000001"; -- -0.0016504226156221697
	pesos_i(7759) := b"1111111111111111_1111111111111111_1110011010000011_1011100001110111"; -- -0.09955260366422704
	pesos_i(7760) := b"1111111111111111_1111111111111111_1110111000100011_1111100111010000"; -- -0.06976355233741618
	pesos_i(7761) := b"0000000000000000_0000000000000000_0001000010110101_0111000010011101"; -- 0.06526855301613693
	pesos_i(7762) := b"1111111111111111_1111111111111111_1110101001101001_1111001011001011"; -- -0.08432085554475623
	pesos_i(7763) := b"0000000000000000_0000000000000000_0010011111011011_1010111010010111"; -- 0.1556958312718582
	pesos_i(7764) := b"1111111111111111_1111111111111111_1111111100110000_0100111100000101"; -- -0.003169118098088712
	pesos_i(7765) := b"0000000000000000_0000000000000000_0010010100111100_0011010001100110"; -- 0.14544990046108988
	pesos_i(7766) := b"0000000000000000_0000000000000000_0001010000110100_0011110010101010"; -- 0.07892207285582228
	pesos_i(7767) := b"1111111111111111_1111111111111111_1110001011010111_0101000001101101"; -- -0.11390206653507101
	pesos_i(7768) := b"0000000000000000_0000000000000000_0001100010010001_0000010011000011"; -- 0.09596280833911464
	pesos_i(7769) := b"1111111111111111_1111111111111111_1111011100000010_1110011001110101"; -- -0.03511199616195362
	pesos_i(7770) := b"0000000000000000_0000000000000000_0001101110110111_0011110100111000"; -- 0.10826475737420913
	pesos_i(7771) := b"1111111111111111_1111111111111111_1101100100010111_0010011110110001"; -- -0.1519904320730236
	pesos_i(7772) := b"1111111111111111_1111111111111111_1101010110000110_1100011100111110"; -- -0.16591219648111244
	pesos_i(7773) := b"0000000000000000_0000000000000000_0000110011110001_0011000011111100"; -- 0.05055528787694094
	pesos_i(7774) := b"0000000000000000_0000000000000000_0001100100010111_1001111011110011"; -- 0.09801667633942754
	pesos_i(7775) := b"1111111111111111_1111111111111111_1101101010010100_0110101110100001"; -- -0.14617278414466323
	pesos_i(7776) := b"0000000000000000_0000000000000000_0000011100011111_0101111001011010"; -- 0.027822396263414345
	pesos_i(7777) := b"1111111111111111_1111111111111111_1101101100001111_1111101111011100"; -- -0.14428735608147963
	pesos_i(7778) := b"0000000000000000_0000000000000000_0001100111110001_0011001111000011"; -- 0.10133670346218183
	pesos_i(7779) := b"0000000000000000_0000000000000000_0001011111001010_0001000111101110"; -- 0.09292709416436161
	pesos_i(7780) := b"0000000000000000_0000000000000000_0010100000000111_0101011101101001"; -- 0.15636202158588666
	pesos_i(7781) := b"1111111111111111_1111111111111111_1110111110101010_1001011010101111"; -- -0.0638032744424519
	pesos_i(7782) := b"0000000000000000_0000000000000000_0001101101000000_1000010001001001"; -- 0.10645319734166377
	pesos_i(7783) := b"1111111111111111_1111111111111111_1110011110001000_0110101001100000"; -- -0.09557471435254992
	pesos_i(7784) := b"1111111111111111_1111111111111111_1111110000000111_0001011000110010"; -- -0.015516865471471436
	pesos_i(7785) := b"1111111111111111_1111111111111111_1111111001100001_0100100010010101"; -- -0.006328071155779043
	pesos_i(7786) := b"1111111111111111_1111111111111111_1110111110001110_1101000101101000"; -- -0.06422702031929887
	pesos_i(7787) := b"0000000000000000_0000000000000000_0000100101000100_0010110011011010"; -- 0.036196520972060595
	pesos_i(7788) := b"0000000000000000_0000000000000000_0010011111110000_1000000010011101"; -- 0.15601352528379658
	pesos_i(7789) := b"0000000000000000_0000000000000000_0010100000110100_1100100110010110"; -- 0.15705547240950637
	pesos_i(7790) := b"1111111111111111_1111111111111111_1110100100011000_0100011110110100"; -- -0.08947326529628588
	pesos_i(7791) := b"1111111111111111_1111111111111111_1110101100010110_0000011001111000"; -- -0.08169517105799287
	pesos_i(7792) := b"1111111111111111_1111111111111111_1110001011110001_1111100010101100"; -- -0.11349530974161158
	pesos_i(7793) := b"0000000000000000_0000000000000000_0010011110101100_0011100101010110"; -- 0.15497167924945252
	pesos_i(7794) := b"1111111111111111_1111111111111111_1110100111011000_1101010111101100"; -- -0.08653510086625932
	pesos_i(7795) := b"0000000000000000_0000000000000000_0001110101101011_0010111010011101"; -- 0.11491671882280252
	pesos_i(7796) := b"0000000000000000_0000000000000000_0000010010001010_1001100100010110"; -- 0.0177398374870982
	pesos_i(7797) := b"1111111111111111_1111111111111111_1110100010110110_0100110010001111"; -- -0.09096833707474598
	pesos_i(7798) := b"1111111111111111_1111111111111111_1101011111001101_0110000011111001"; -- -0.1570224181594768
	pesos_i(7799) := b"0000000000000000_0000000000000000_0001100101110100_0001010101101011"; -- 0.0994275461355569
	pesos_i(7800) := b"1111111111111111_1111111111111111_1111000111011010_1010100011110100"; -- -0.05525726368508037
	pesos_i(7801) := b"1111111111111111_1111111111111111_1110110000011100_1010110011001100"; -- -0.07768745447428199
	pesos_i(7802) := b"0000000000000000_0000000000000000_0010000100011110_1111111111000100"; -- 0.1293792584681823
	pesos_i(7803) := b"1111111111111111_1111111111111111_1110111010011101_0001100001100000"; -- -0.06791541718917213
	pesos_i(7804) := b"0000000000000000_0000000000000000_0010001111000000_1011010011110000"; -- 0.13965922217382984
	pesos_i(7805) := b"1111111111111111_1111111111111111_1111110101010000_1101111011101111"; -- -0.010484758907272374
	pesos_i(7806) := b"1111111111111111_1111111111111111_1111111011000110_0110001011110011"; -- -0.004785361950186265
	pesos_i(7807) := b"0000000000000000_0000000000000000_0000111111110011_0100111110010001"; -- 0.06230637833256215
	pesos_i(7808) := b"1111111111111111_1111111111111111_1111010110110100_1001011001111011"; -- -0.04021319859483721
	pesos_i(7809) := b"0000000000000000_0000000000000000_0000001001001101_0101010100011110"; -- 0.008992500187068653
	pesos_i(7810) := b"0000000000000000_0000000000000000_0000100110101100_0010101100001101"; -- 0.03778332781923072
	pesos_i(7811) := b"1111111111111111_1111111111111111_1110000111100110_0011101000101101"; -- -0.11758076092816377
	pesos_i(7812) := b"0000000000000000_0000000000000000_0000001001000011_1110100010100001"; -- 0.008848704554984004
	pesos_i(7813) := b"1111111111111111_1111111111111111_1101111101011010_1111101000010101"; -- -0.1275180530398898
	pesos_i(7814) := b"1111111111111111_1111111111111111_1111000010010100_0011010011001111"; -- -0.06023855167943767
	pesos_i(7815) := b"0000000000000000_0000000000000000_0000100010011111_0100101010010111"; -- 0.033680593341469355
	pesos_i(7816) := b"0000000000000000_0000000000000000_0001010011000111_0010010011100001"; -- 0.08116369716613632
	pesos_i(7817) := b"0000000000000000_0000000000000000_0010110100110010_0010101101011110"; -- 0.1765467742679455
	pesos_i(7818) := b"1111111111111111_1111111111111111_1111001100000110_1010010111000000"; -- -0.05067981790015415
	pesos_i(7819) := b"1111111111111111_1111111111111111_1110011000001001_0110110001001001"; -- -0.10141871652541849
	pesos_i(7820) := b"1111111111111111_1111111111111111_1110100001110010_0010110100111101"; -- -0.09200780155560086
	pesos_i(7821) := b"0000000000000000_0000000000000000_0000011010000100_0000101110111110"; -- 0.025452360017393483
	pesos_i(7822) := b"1111111111111111_1111111111111111_1101011000101101_0001001100110111"; -- -0.16337470917779054
	pesos_i(7823) := b"0000000000000000_0000000000000000_0010001011100101_1000111001100000"; -- 0.13631524883176327
	pesos_i(7824) := b"0000000000000000_0000000000000000_0010001110001010_0101100100000110"; -- 0.13882976908556963
	pesos_i(7825) := b"1111111111111111_1111111111111111_1111110101011000_1111111110011011"; -- -0.01036074124865371
	pesos_i(7826) := b"0000000000000000_0000000000000000_0010001100001001_1101010110001000"; -- 0.13686880667223272
	pesos_i(7827) := b"1111111111111111_1111111111111111_1110111111110101_1001100010101010"; -- -0.06265874708045606
	pesos_i(7828) := b"1111111111111111_1111111111111111_1111110010100011_1100101111111010"; -- -0.01312565940681408
	pesos_i(7829) := b"1111111111111111_1111111111111111_1111111111000000_0101001000000001"; -- -0.0009716746194393062
	pesos_i(7830) := b"1111111111111111_1111111111111111_1111000001000101_0000010011001110"; -- -0.061446857247659845
	pesos_i(7831) := b"0000000000000000_0000000000000000_0001110000011111_1100101011011010"; -- 0.10986011337177591
	pesos_i(7832) := b"0000000000000000_0000000000000000_0001010000101100_0111110001110100"; -- 0.07880380468377562
	pesos_i(7833) := b"1111111111111111_1111111111111111_1101011011011000_0101011100001110"; -- -0.16076141278541012
	pesos_i(7834) := b"0000000000000000_0000000000000000_0001000101110101_1001001011111110"; -- 0.0682002896529437
	pesos_i(7835) := b"1111111111111111_1111111111111111_1110110101001100_1100110000000111"; -- -0.0730469209462034
	pesos_i(7836) := b"1111111111111111_1111111111111111_1110101110001000_0000100111010001"; -- -0.07995546965681259
	pesos_i(7837) := b"1111111111111111_1111111111111111_1111111101000001_0010001011010110"; -- -0.0029123523202265805
	pesos_i(7838) := b"1111111111111111_1111111111111111_1110010011011011_1000111000001100"; -- -0.10602485861603098
	pesos_i(7839) := b"1111111111111111_1111111111111111_1110111010101011_1100011111001100"; -- -0.06769133830474328
	pesos_i(7840) := b"1111111111111111_1111111111111111_1111000101010111_1010000010000001"; -- -0.05725666858528096
	pesos_i(7841) := b"1111111111111111_1111111111111111_1110011001001011_1101100011110111"; -- -0.10040515872764319
	pesos_i(7842) := b"0000000000000000_0000000000000000_0000110111111001_0101000001001100"; -- 0.05458547456474664
	pesos_i(7843) := b"0000000000000000_0000000000000000_0000001101000011_1000011111011000"; -- 0.012749185873754494
	pesos_i(7844) := b"0000000000000000_0000000000000000_0000001110001111_1101001011110101"; -- 0.0139133309442723
	pesos_i(7845) := b"1111111111111111_1111111111111111_1110001110001001_1101111111100010"; -- -0.1111774515057343
	pesos_i(7846) := b"1111111111111111_1111111111111111_1111101000010001_0011000111001011"; -- -0.023175132602772576
	pesos_i(7847) := b"0000000000000000_0000000000000000_0001000001000111_1110010110001000"; -- 0.06359705512664443
	pesos_i(7848) := b"0000000000000000_0000000000000000_0000111100100111_1111110100011101"; -- 0.05920392946623071
	pesos_i(7849) := b"0000000000000000_0000000000000000_0000000011001010_1001011111001110"; -- 0.003091323757080326
	pesos_i(7850) := b"0000000000000000_0000000000000000_0010000100101100_1111101100101100"; -- 0.12959260776400383
	pesos_i(7851) := b"0000000000000000_0000000000000000_0010111011000111_1100000000110111"; -- 0.1827354558407075
	pesos_i(7852) := b"1111111111111111_1111111111111111_1101010001101010_1000101101110000"; -- -0.17024925727654397
	pesos_i(7853) := b"0000000000000000_0000000000000000_0001111000001101_0101110110000101"; -- 0.11739143857145853
	pesos_i(7854) := b"0000000000000000_0000000000000000_0001011111001000_0000010000101100"; -- 0.09289575646297211
	pesos_i(7855) := b"1111111111111111_1111111111111111_1110100110011011_0000111110101111"; -- -0.08747770278591566
	pesos_i(7856) := b"0000000000000000_0000000000000000_0010011011010101_1011010011000001"; -- 0.15169839587479392
	pesos_i(7857) := b"0000000000000000_0000000000000000_0010011111111010_1001111010101000"; -- 0.1561679040296303
	pesos_i(7858) := b"1111111111111111_1111111111111111_1110111001000101_1000001101010101"; -- -0.06925181555336263
	pesos_i(7859) := b"1111111111111111_1111111111111111_1101010100000100_0001100111001000"; -- -0.16790617812592787
	pesos_i(7860) := b"1111111111111111_1111111111111111_1110101001010011_1010101100001011"; -- -0.08466082544572376
	pesos_i(7861) := b"1111111111111111_1111111111111111_1110101010010001_0000000011010011"; -- -0.08372492648568944
	pesos_i(7862) := b"1111111111111111_1111111111111111_1110110100011111_0010101010010000"; -- -0.07374319066864732
	pesos_i(7863) := b"1111111111111111_1111111111111111_1111111100010000_1110011000001010"; -- -0.0036483979141163137
	pesos_i(7864) := b"1111111111111111_1111111111111111_1110100101001110_1101010110000111"; -- -0.08864083733152266
	pesos_i(7865) := b"0000000000000000_0000000000000000_0000110000101001_0001110001100101"; -- 0.047502302859483744
	pesos_i(7866) := b"0000000000000000_0000000000000000_0000011101110001_1101010101010111"; -- 0.029080709252266395
	pesos_i(7867) := b"1111111111111111_1111111111111111_1110100000111100_0111011010011010"; -- -0.09282740347927804
	pesos_i(7868) := b"0000000000000000_0000000000000000_0000110110111100_0000011111100100"; -- 0.05365037262054407
	pesos_i(7869) := b"1111111111111111_1111111111111111_1101010000011000_0111000000100110"; -- -0.17150210449145084
	pesos_i(7870) := b"0000000000000000_0000000000000000_0001100011100001_1001000111011100"; -- 0.09719192143157587
	pesos_i(7871) := b"1111111111111111_1111111111111111_1111010100101000_1110010111010000"; -- -0.04234470052739987
	pesos_i(7872) := b"0000000000000000_0000000000000000_0010010000010101_0001011001111101"; -- 0.14094677503319294
	pesos_i(7873) := b"1111111111111111_1111111111111111_1111001000010000_0100001110011111"; -- -0.05443932884358832
	pesos_i(7874) := b"0000000000000000_0000000000000000_0001100011101100_1010010011100101"; -- 0.09736090263286923
	pesos_i(7875) := b"0000000000000000_0000000000000000_0001100101001010_1110011101000111"; -- 0.09879918550149049
	pesos_i(7876) := b"0000000000000000_0000000000000000_0001001001001101_0100010001011101"; -- 0.07149150153259187
	pesos_i(7877) := b"1111111111111111_1111111111111111_1111011111110111_1100001010000001"; -- -0.03137573573416025
	pesos_i(7878) := b"1111111111111111_1111111111111111_1111001011101011_1110000010111011"; -- -0.051088289655910314
	pesos_i(7879) := b"1111111111111111_1111111111111111_1111101100100010_1011111001110010"; -- -0.01900109971105707
	pesos_i(7880) := b"1111111111111111_1111111111111111_1111011000000001_1000001000001110"; -- -0.03903948938416825
	pesos_i(7881) := b"0000000000000000_0000000000000000_0010101100111000_0000011011101001"; -- 0.1688236541426683
	pesos_i(7882) := b"1111111111111111_1111111111111111_1101100111111001_1111100011010101"; -- -0.14852947993661791
	pesos_i(7883) := b"0000000000000000_0000000000000000_0010001000100000_0001110111100111"; -- 0.13330256360940215
	pesos_i(7884) := b"0000000000000000_0000000000000000_0001101000111101_0111011110010110"; -- 0.10250041411308805
	pesos_i(7885) := b"1111111111111111_1111111111111111_1101111010101100_1110010101001001"; -- -0.13017432185552588
	pesos_i(7886) := b"1111111111111111_1111111111111111_1111101101011101_1000001011100000"; -- -0.018104381910381925
	pesos_i(7887) := b"0000000000000000_0000000000000000_0000100000000111_1000011011110101"; -- 0.03136485557437525
	pesos_i(7888) := b"1111111111111111_1111111111111111_1111111100001111_1000100100001010"; -- -0.0036691999149156274
	pesos_i(7889) := b"1111111111111111_1111111111111111_1101101011111111_1011001010011001"; -- -0.1445358635945518
	pesos_i(7890) := b"1111111111111111_1111111111111111_1111011110111011_1001000111011111"; -- -0.032294161740982166
	pesos_i(7891) := b"1111111111111111_1111111111111111_1111010000001100_0001110001101111"; -- -0.04669019967154996
	pesos_i(7892) := b"1111111111111111_1111111111111111_1111011011100111_1001101011000010"; -- -0.035528495389609685
	pesos_i(7893) := b"1111111111111111_1111111111111111_1101011110010000_1010010011101100"; -- -0.15794915429687859
	pesos_i(7894) := b"1111111111111111_1111111111111111_1101101011100111_1110111000001101"; -- -0.14489853069781858
	pesos_i(7895) := b"0000000000000000_0000000000000000_0000111101000010_0110000010001000"; -- 0.05960658378458731
	pesos_i(7896) := b"1111111111111111_1111111111111111_1111110110011101_0000000001011001"; -- -0.009323099295311665
	pesos_i(7897) := b"1111111111111111_1111111111111111_1101110110111001_1111100100100000"; -- -0.13388102504557906
	pesos_i(7898) := b"1111111111111111_1111111111111111_1101111000001011_1001000100010100"; -- -0.13263600596899966
	pesos_i(7899) := b"0000000000000000_0000000000000000_0000011110101011_0111010111111100"; -- 0.029960035382654317
	pesos_i(7900) := b"1111111111111111_1111111111111111_1110100001000110_1001110101000110"; -- -0.09267251054904814
	pesos_i(7901) := b"0000000000000000_0000000000000000_0001110011011001_0111101010100111"; -- 0.1126934679538885
	pesos_i(7902) := b"1111111111111111_1111111111111111_1111011010000101_1001010111001010"; -- -0.03702415289909217
	pesos_i(7903) := b"1111111111111111_1111111111111111_1101010100110011_1101111001000100"; -- -0.167177303619273
	pesos_i(7904) := b"0000000000000000_0000000000000000_0010000011101100_1110000010111110"; -- 0.12861446978931787
	pesos_i(7905) := b"1111111111111111_1111111111111111_1101100101000111_1001110001000000"; -- -0.15125106265036697
	pesos_i(7906) := b"0000000000000000_0000000000000000_0010100110011011_0101111101110100"; -- 0.16252705185082938
	pesos_i(7907) := b"0000000000000000_0000000000000000_0001000101111001_0111011001100101"; -- 0.06825962032231797
	pesos_i(7908) := b"0000000000000000_0000000000000000_0010011001001111_0111111000100010"; -- 0.14965046243945374
	pesos_i(7909) := b"0000000000000000_0000000000000000_0010011010010110_1011000011000011"; -- 0.15073685410385615
	pesos_i(7910) := b"1111111111111111_1111111111111111_1111010001001100_1110100011010101"; -- -0.0457014542063221
	pesos_i(7911) := b"0000000000000000_0000000000000000_0000001000001110_1101101110011000"; -- 0.00803921175834954
	pesos_i(7912) := b"1111111111111111_1111111111111111_1101111001111001_0010010001011010"; -- -0.13096401989524112
	pesos_i(7913) := b"1111111111111111_1111111111111111_1101101110011000_1011110111001000"; -- -0.14220060233276358
	pesos_i(7914) := b"0000000000000000_0000000000000000_0001011101001101_1101101101100111"; -- 0.0910317540791874
	pesos_i(7915) := b"0000000000000000_0000000000000000_0000010001011001_1000100010100100"; -- 0.016991176752948218
	pesos_i(7916) := b"1111111111111111_1111111111111111_1111011100100111_1000001010010100"; -- -0.03455337422890199
	pesos_i(7917) := b"1111111111111111_1111111111111111_1110010001111001_1000101001010101"; -- -0.10752044139220729
	pesos_i(7918) := b"0000000000000000_0000000000000000_0010001101000011_1111000000011110"; -- 0.1377554008574485
	pesos_i(7919) := b"0000000000000000_0000000000000000_0000110011001000_1001101000110000"; -- 0.04993594817395777
	pesos_i(7920) := b"1111111111111111_1111111111111111_1111001011100110_1011111101000101"; -- -0.05116657796285798
	pesos_i(7921) := b"1111111111111111_1111111111111111_1101101000101100_1111110011101101"; -- -0.14775103763046296
	pesos_i(7922) := b"1111111111111111_1111111111111111_1111101000110111_0000101111010010"; -- -0.02259756198396685
	pesos_i(7923) := b"1111111111111111_1111111111111111_1110000001001000_1000000001010101"; -- -0.12389371807017407
	pesos_i(7924) := b"0000000000000000_0000000000000000_0010001001101010_1001110110000010"; -- 0.1344393198830335
	pesos_i(7925) := b"0000000000000000_0000000000000000_0001100001101111_1101001010010111"; -- 0.09545627779778387
	pesos_i(7926) := b"1111111111111111_1111111111111111_1110001000111001_1010101100010001"; -- -0.11630755259421076
	pesos_i(7927) := b"1111111111111111_1111111111111111_1111100011000000_1011001110000111"; -- -0.028309611763861143
	pesos_i(7928) := b"1111111111111111_1111111111111111_1101101010010111_1011001000000000"; -- -0.14612281321769197
	pesos_i(7929) := b"1111111111111111_1111111111111111_1110001101001100_1111011000110001"; -- -0.11210690779545761
	pesos_i(7930) := b"1111111111111111_1111111111111111_1111111101000110_1110001101100011"; -- -0.002824581453591201
	pesos_i(7931) := b"1111111111111111_1111111111111111_1110010011000100_0111001101111111"; -- -0.10637739313657639
	pesos_i(7932) := b"1111111111111111_1111111111111111_1110010111100011_0100011011110000"; -- -0.10200077656565133
	pesos_i(7933) := b"1111111111111111_1111111111111111_1101111001010011_0111110001001110"; -- -0.1315386113946572
	pesos_i(7934) := b"0000000000000000_0000000000000000_0010100011101110_1111110110110110"; -- 0.1598967141371629
	pesos_i(7935) := b"0000000000000000_0000000000000000_0010011001110100_1101001111110101"; -- 0.15022015325464055
	pesos_i(7936) := b"0000000000000000_0000000000000000_0001010001111001_1000110110001100"; -- 0.07997975035914437
	pesos_i(7937) := b"1111111111111111_1111111111111111_1101101111011100_1111011000000111"; -- -0.14115965196844754
	pesos_i(7938) := b"1111111111111111_1111111111111111_1111100100101010_1111010100000110"; -- -0.026688276318631275
	pesos_i(7939) := b"1111111111111111_1111111111111111_1110000101100000_0000111010111011"; -- -0.11962802825248188
	pesos_i(7940) := b"1111111111111111_1111111111111111_1110011001100011_1101010010101000"; -- -0.10003920451562573
	pesos_i(7941) := b"0000000000000000_0000000000000000_0000111111100010_0000001001100001"; -- 0.062042378228202605
	pesos_i(7942) := b"0000000000000000_0000000000000000_0000010100001000_0001100100010110"; -- 0.0196548155310556
	pesos_i(7943) := b"0000000000000000_0000000000000000_0000101100110011_1010110000011110"; -- 0.04375720733384009
	pesos_i(7944) := b"1111111111111111_1111111111111111_1111001110100001_0101101111010010"; -- -0.048319112046258904
	pesos_i(7945) := b"0000000000000000_0000000000000000_0001000010011110_1101101100010111"; -- 0.06492394740766595
	pesos_i(7946) := b"1111111111111111_1111111111111111_1110000100101011_1110110011000111"; -- -0.12042350907636983
	pesos_i(7947) := b"0000000000000000_0000000000000000_0010101001110011_1000011101110111"; -- 0.1658253349617387
	pesos_i(7948) := b"0000000000000000_0000000000000000_0000001010100100_0010011010011000"; -- 0.010317241793386054
	pesos_i(7949) := b"0000000000000000_0000000000000000_0010000111011000_1000110111010011"; -- 0.13221060183289698
	pesos_i(7950) := b"0000000000000000_0000000000000000_0000010111011000_1100010011101110"; -- 0.022838886347453242
	pesos_i(7951) := b"0000000000000000_0000000000000000_0001011000100001_0001000011011000"; -- 0.08644204405889212
	pesos_i(7952) := b"0000000000000000_0000000000000000_0010100001000001_0100000010101100"; -- 0.15724567604686465
	pesos_i(7953) := b"0000000000000000_0000000000000000_0010100111001011_1100000011110000"; -- 0.16326528404980808
	pesos_i(7954) := b"1111111111111111_1111111111111111_1110011111100101_1101100110000111"; -- -0.09414902155089712
	pesos_i(7955) := b"1111111111111111_1111111111111111_1110011001100111_0011110011001011"; -- -0.09998722129885296
	pesos_i(7956) := b"1111111111111111_1111111111111111_1111110111110001_0110001100110011"; -- -0.008035469174971147
	pesos_i(7957) := b"1111111111111111_1111111111111111_1101011101101101_1010011011101000"; -- -0.1584830936844727
	pesos_i(7958) := b"1111111111111111_1111111111111111_1111000000111001_1011011000011110"; -- -0.06161939392058285
	pesos_i(7959) := b"0000000000000000_0000000000000000_0010000110101001_0001001111110110"; -- 0.13148617502303211
	pesos_i(7960) := b"1111111111111111_1111111111111111_1111011011010000_0101111001110001"; -- -0.035883042612912905
	pesos_i(7961) := b"0000000000000000_0000000000000000_0000110100110010_0010101001001010"; -- 0.05154671009000292
	pesos_i(7962) := b"0000000000000000_0000000000000000_0000101101100100_1111001000110101"; -- 0.04450906561524323
	pesos_i(7963) := b"1111111111111111_1111111111111111_1101110011111001_0101010101110110"; -- -0.1368204677322957
	pesos_i(7964) := b"0000000000000000_0000000000000000_0010101100101000_0000110000100001"; -- 0.16857982449630607
	pesos_i(7965) := b"0000000000000000_0000000000000000_0001011010011101_1010011111101011"; -- 0.08834313848362113
	pesos_i(7966) := b"0000000000000000_0000000000000000_0010011100001100_0000100010001000"; -- 0.15252736401374803
	pesos_i(7967) := b"1111111111111111_1111111111111111_1110001000010001_1001000101001110"; -- -0.11691943985798267
	pesos_i(7968) := b"1111111111111111_1111111111111111_1101110111010010_1100100100101100"; -- -0.13350241352995373
	pesos_i(7969) := b"0000000000000000_0000000000000000_0010100011101101_1101101000100110"; -- 0.15987933569386406
	pesos_i(7970) := b"1111111111111111_1111111111111111_1110001001101001_1000111111101110"; -- -0.11557674815491728
	pesos_i(7971) := b"0000000000000000_0000000000000000_0010000001000010_1100101010110010"; -- 0.1260191615625538
	pesos_i(7972) := b"1111111111111111_1111111111111111_1111110011000111_0111001111000110"; -- -0.012581600363289216
	pesos_i(7973) := b"0000000000000000_0000000000000000_0010001011011011_0001010001101011"; -- 0.13615539170426283
	pesos_i(7974) := b"1111111111111111_1111111111111111_1111110111001001_0001001001111111"; -- -0.008650630861531207
	pesos_i(7975) := b"1111111111111111_1111111111111111_1110011001000100_0010011011101110"; -- -0.10052258191506568
	pesos_i(7976) := b"1111111111111111_1111111111111111_1110100111010011_0000011010010111"; -- -0.08662375276128037
	pesos_i(7977) := b"1111111111111111_1111111111111111_1111101010110100_1100111001010110"; -- -0.020678619484769248
	pesos_i(7978) := b"0000000000000000_0000000000000000_0010100001001100_0101001100110010"; -- 0.15741462677073234
	pesos_i(7979) := b"1111111111111111_1111111111111111_1110100010001110_0010100011101001"; -- -0.09158081344911904
	pesos_i(7980) := b"0000000000000000_0000000000000000_0001100000110110_1110011011110011"; -- 0.09458774014912455
	pesos_i(7981) := b"0000000000000000_0000000000000000_0010100011011010_0011100101010000"; -- 0.15957983208771834
	pesos_i(7982) := b"1111111111111111_1111111111111111_1111010110001011_0000000000010010"; -- -0.04084777418132084
	pesos_i(7983) := b"1111111111111111_1111111111111111_1101011101111111_0101100000110111"; -- -0.15821312576566443
	pesos_i(7984) := b"1111111111111111_1111111111111111_1110000001100101_1101111010101001"; -- -0.12344559069703867
	pesos_i(7985) := b"1111111111111111_1111111111111111_1101110110000010_1101110001010100"; -- -0.13472197473761965
	pesos_i(7986) := b"0000000000000000_0000000000000000_0010000010100000_0101111111110100"; -- 0.12744712551091708
	pesos_i(7987) := b"0000000000000000_0000000000000000_0010011101101000_1001101111100010"; -- 0.15393995542201977
	pesos_i(7988) := b"0000000000000000_0000000000000000_0000101111000001_1111110011000100"; -- 0.045928762365790236
	pesos_i(7989) := b"1111111111111111_1111111111111111_1111100011101010_0000010100010111"; -- -0.027679139970183435
	pesos_i(7990) := b"1111111111111111_1111111111111111_1110011100100011_1101000001011110"; -- -0.09710977268027973
	pesos_i(7991) := b"1111111111111111_1111111111111111_1111110000101011_0101010111001011"; -- -0.014963758521060107
	pesos_i(7992) := b"1111111111111111_1111111111111111_1111110010111001_0100010001010000"; -- -0.012798052172771829
	pesos_i(7993) := b"1111111111111111_1111111111111111_1101111010010010_0111010010111111"; -- -0.13057775808477817
	pesos_i(7994) := b"0000000000000000_0000000000000000_0000101101100011_0101101100100000"; -- 0.04448480150692091
	pesos_i(7995) := b"0000000000000000_0000000000000000_0001000101101010_0001000010000001"; -- 0.06802466539993147
	pesos_i(7996) := b"1111111111111111_1111111111111111_1111101010100011_1111101101011000"; -- -0.020935336099639282
	pesos_i(7997) := b"1111111111111111_1111111111111111_1101100010110011_1111011011101000"; -- -0.15350396000709204
	pesos_i(7998) := b"0000000000000000_0000000000000000_0001111011110000_0010111001010111"; -- 0.12085237150713332
	pesos_i(7999) := b"0000000000000000_0000000000000000_0001100000100010_1001001000011100"; -- 0.09427750764024788
	pesos_i(8000) := b"0000000000000000_0000000000000000_0000000111111010_0101010111101011"; -- 0.007726068408877351
	pesos_i(8001) := b"1111111111111111_1111111111111111_1110100110000010_0001110100001000"; -- -0.08785837692550197
	pesos_i(8002) := b"1111111111111111_1111111111111111_1110101001111000_1001011111011001"; -- -0.08409739438905381
	pesos_i(8003) := b"1111111111111111_1111111111111111_1111011110111010_0001011101001000"; -- -0.0323167275009009
	pesos_i(8004) := b"1111111111111111_1111111111111111_1101100011010000_1111110111111111"; -- -0.15306103244893327
	pesos_i(8005) := b"0000000000000000_0000000000000000_0001000000111011_1101011100111100"; -- 0.06341309744817293
	pesos_i(8006) := b"0000000000000000_0000000000000000_0000100010111010_0110111100000110"; -- 0.03409475237695802
	pesos_i(8007) := b"0000000000000000_0000000000000000_0000101100100010_1101111000001110"; -- 0.043500784247742265
	pesos_i(8008) := b"1111111111111111_1111111111111111_1111011111100011_1100010101111000"; -- -0.031680734717392016
	pesos_i(8009) := b"0000000000000000_0000000000000000_0001001100110011_1010010000000110"; -- 0.07500672484970622
	pesos_i(8010) := b"1111111111111111_1111111111111111_1110010000011000_0011010111100010"; -- -0.10900557740033816
	pesos_i(8011) := b"0000000000000000_0000000000000000_0010100010001011_1001111010001101"; -- 0.15838042213117268
	pesos_i(8012) := b"1111111111111111_1111111111111111_1110011100101100_0111111000100010"; -- -0.0969773450922045
	pesos_i(8013) := b"1111111111111111_1111111111111111_1111011001011100_1000000011011001"; -- -0.037651011470921474
	pesos_i(8014) := b"0000000000000000_0000000000000000_0010000100010111_0111011100011101"; -- 0.12926430176399015
	pesos_i(8015) := b"0000000000000000_0000000000000000_0001100110101111_1001101111011101"; -- 0.10033582829032016
	pesos_i(8016) := b"0000000000000000_0000000000000000_0001101000001110_1101000101111011"; -- 0.10178860895163236
	pesos_i(8017) := b"0000000000000000_0000000000000000_0010110001010110_1111110010100000"; -- 0.17320231338611383
	pesos_i(8018) := b"1111111111111111_1111111111111111_1111010100111001_1011000100111100"; -- -0.04208843510767673
	pesos_i(8019) := b"1111111111111111_1111111111111111_1101100100001011_1111100110100011"; -- -0.1521610238580701
	pesos_i(8020) := b"1111111111111111_1111111111111111_1110110011010101_0000001100000100"; -- -0.07487469808264127
	pesos_i(8021) := b"0000000000000000_0000000000000000_0010001011001010_0001101010001111"; -- 0.13589635831183375
	pesos_i(8022) := b"1111111111111111_1111111111111111_1111100011111111_0110100001010110"; -- -0.02735278980993437
	pesos_i(8023) := b"1111111111111111_1111111111111111_1101101000110100_0011111000111011"; -- -0.14764033368563495
	pesos_i(8024) := b"1111111111111111_1111111111111111_1111101111000101_0010101110001000"; -- -0.016522673795487074
	pesos_i(8025) := b"1111111111111111_1111111111111111_1101101010011110_0110010110000010"; -- -0.14602056097955382
	pesos_i(8026) := b"1111111111111111_1111111111111111_1101101101000001_0010100001001011"; -- -0.14353702697851764
	pesos_i(8027) := b"0000000000000000_0000000000000000_0001110000110010_0111100100011110"; -- 0.11014515859831177
	pesos_i(8028) := b"1111111111111111_1111111111111111_1101011111111101_1011000100100110"; -- -0.15628521749420102
	pesos_i(8029) := b"1111111111111111_1111111111111111_1101101000111001_1000010010100010"; -- -0.1475598436009519
	pesos_i(8030) := b"0000000000000000_0000000000000000_0001110001100100_1000110010101001"; -- 0.11090926293766859
	pesos_i(8031) := b"1111111111111111_1111111111111111_1111000001111101_1011011011100101"; -- -0.060581750056641445
	pesos_i(8032) := b"1111111111111111_1111111111111111_1101001011110111_0110101100010110"; -- -0.1759121963128056
	pesos_i(8033) := b"1111111111111111_1111111111111111_1111101001010111_1011110110011011"; -- -0.022098684030992837
	pesos_i(8034) := b"0000000000000000_0000000000000000_0000101100010011_0001001101010011"; -- 0.04325981875600717
	pesos_i(8035) := b"1111111111111111_1111111111111111_1110110101101000_1001001111010100"; -- -0.0726230247675656
	pesos_i(8036) := b"1111111111111111_1111111111111111_1101100010111110_1110110001110000"; -- -0.15333673737531658
	pesos_i(8037) := b"0000000000000000_0000000000000000_0010011100101001_0001100100100110"; -- 0.1529708592365327
	pesos_i(8038) := b"1111111111111111_1111111111111111_1110001001000111_1100100010100100"; -- -0.11609216681216991
	pesos_i(8039) := b"0000000000000000_0000000000000000_0000110111100000_1110001100100010"; -- 0.05421275687033461
	pesos_i(8040) := b"0000000000000000_0000000000000000_0001001010010010_0001111110001011"; -- 0.07254216323662169
	pesos_i(8041) := b"0000000000000000_0000000000000000_0010010100101101_1011100010000011"; -- 0.14522889336813563
	pesos_i(8042) := b"0000000000000000_0000000000000000_0001000011110010_1010011000111110"; -- 0.06620253567783736
	pesos_i(8043) := b"1111111111111111_1111111111111111_1110000010100111_0111001000010100"; -- -0.12244498258277615
	pesos_i(8044) := b"0000000000000000_0000000000000000_0001110011101010_0100110000110000"; -- 0.11295009768117623
	pesos_i(8045) := b"0000000000000000_0000000000000000_0010000000100110_0100000110100010"; -- 0.12558374597889288
	pesos_i(8046) := b"0000000000000000_0000000000000000_0010001101111000_1101001011010000"; -- 0.1385623700371695
	pesos_i(8047) := b"1111111111111111_1111111111111111_1110111100101011_1100111010110110"; -- -0.06573780108040063
	pesos_i(8048) := b"1111111111111111_1111111111111111_1110010011000000_0100111110100011"; -- -0.10644056587749003
	pesos_i(8049) := b"0000000000000000_0000000000000000_0000101010011101_0000010110001110"; -- 0.04145846095366136
	pesos_i(8050) := b"1111111111111111_1111111111111111_1111000100001010_1100010100010110"; -- -0.05842941478581139
	pesos_i(8051) := b"1111111111111111_1111111111111111_1101110010000101_0111101100010111"; -- -0.13858824433769162
	pesos_i(8052) := b"0000000000000000_0000000000000000_0000010011101010_1010111101101010"; -- 0.01920601211413879
	pesos_i(8053) := b"1111111111111111_1111111111111111_1111010010110100_0100110000000100"; -- -0.04412388718154537
	pesos_i(8054) := b"1111111111111111_1111111111111111_1110100011111101_1111110011101110"; -- -0.08987445063359892
	pesos_i(8055) := b"1111111111111111_1111111111111111_1110110001000010_1100101110111010"; -- -0.07710577695405661
	pesos_i(8056) := b"0000000000000000_0000000000000000_0010011111011010_1111101100010011"; -- 0.1556851313104037
	pesos_i(8057) := b"0000000000000000_0000000000000000_0010001101110001_0000111000000101"; -- 0.13844382873688774
	pesos_i(8058) := b"0000000000000000_0000000000000000_0001101011110011_0001111000001101"; -- 0.1052721770232586
	pesos_i(8059) := b"0000000000000000_0000000000000000_0000010100110011_1100111111000011"; -- 0.020321831881537175
	pesos_i(8060) := b"1111111111111111_1111111111111111_1111111001110101_1100010011111101"; -- -0.006015480157735129
	pesos_i(8061) := b"1111111111111111_1111111111111111_1110001101000111_1111111101000001"; -- -0.11218266174304718
	pesos_i(8062) := b"0000000000000000_0000000000000000_0001001010001011_1100101001100001"; -- 0.07244553430448811
	pesos_i(8063) := b"0000000000000000_0000000000000000_0001100101011011_1100010110110110"; -- 0.09905658431421176
	pesos_i(8064) := b"0000000000000000_0000000000000000_0000100001100010_0010111000010011"; -- 0.032748107609060106
	pesos_i(8065) := b"0000000000000000_0000000000000000_0001110011101101_0011000001110000"; -- 0.11299422022209805
	pesos_i(8066) := b"1111111111111111_1111111111111111_1111100111101010_1000101111001001"; -- -0.02376486160615383
	pesos_i(8067) := b"1111111111111111_1111111111111111_1101001001010110_0010101100010101"; -- -0.1783726763426941
	pesos_i(8068) := b"1111111111111111_1111111111111111_1111010110001001_1110111100100011"; -- -0.040864042289198384
	pesos_i(8069) := b"1111111111111111_1111111111111111_1101001110000100_1100010101000010"; -- -0.17375533237891497
	pesos_i(8070) := b"1111111111111111_1111111111111111_1110101001110100_1001000101100000"; -- -0.0841588154239745
	pesos_i(8071) := b"1111111111111111_1111111111111111_1111100010001001_0110011000011110"; -- -0.02915345932383567
	pesos_i(8072) := b"0000000000000000_0000000000000000_0000011111010010_1111010111110011"; -- 0.030562755444816334
	pesos_i(8073) := b"1111111111111111_1111111111111111_1111100000101110_1101110101010110"; -- -0.0305349031216602
	pesos_i(8074) := b"0000000000000000_0000000000000000_0001000011000010_1010100101110011"; -- 0.06547030500163285
	pesos_i(8075) := b"0000000000000000_0000000000000000_0010010111000001_0000001011101011"; -- 0.14747637017380366
	pesos_i(8076) := b"0000000000000000_0000000000000000_0001011011011000_1011101110100000"; -- 0.08924458183223052
	pesos_i(8077) := b"0000000000000000_0000000000000000_0001010011011101_0010000100101101"; -- 0.08149916990991368
	pesos_i(8078) := b"0000000000000000_0000000000000000_0000111001101111_0001101111111100"; -- 0.05638289349568808
	pesos_i(8079) := b"1111111111111111_1111111111111111_1101010010000000_0100001101011001"; -- -0.1699178608279473
	pesos_i(8080) := b"1111111111111111_1111111111111111_1110111011010011_1100010011101000"; -- -0.0670811588833386
	pesos_i(8081) := b"1111111111111111_1111111111111111_1101110100101001_0010010010110010"; -- -0.1360909525189619
	pesos_i(8082) := b"1111111111111111_1111111111111111_1110010001000000_0110010010011011"; -- -0.10839244083321802
	pesos_i(8083) := b"1111111111111111_1111111111111111_1111011001101101_0101111101101001"; -- -0.037393605149756245
	pesos_i(8084) := b"0000000000000000_0000000000000000_0010100011011001_1111110001000010"; -- 0.15957619285660207
	pesos_i(8085) := b"0000000000000000_0000000000000000_0000101000011010_1001010110100111"; -- 0.03946814845524193
	pesos_i(8086) := b"0000000000000000_0000000000000000_0010010100110001_1100101001101111"; -- 0.1452909967217804
	pesos_i(8087) := b"1111111111111111_1111111111111111_1111000011011010_1110111000001101"; -- -0.0591593951488776
	pesos_i(8088) := b"0000000000000000_0000000000000000_0000001001010001_0100110110011111"; -- 0.009053088400763479
	pesos_i(8089) := b"1111111111111111_1111111111111111_1111101110100000_1100011101101111"; -- -0.01707795661613892
	pesos_i(8090) := b"1111111111111111_1111111111111111_1101101100000111_1010010001000110"; -- -0.14441464700910622
	pesos_i(8091) := b"0000000000000000_0000000000000000_0000000001010011_0001000000000110"; -- 0.0012674346651258843
	pesos_i(8092) := b"0000000000000000_0000000000000000_0001010001111110_1110111100101011"; -- 0.08006186286154911
	pesos_i(8093) := b"1111111111111111_1111111111111111_1111101101000111_0110001100110111"; -- -0.018441962263800266
	pesos_i(8094) := b"0000000000000000_0000000000000000_0001010101011110_1111101101110001"; -- 0.08348056326536483
	pesos_i(8095) := b"1111111111111111_1111111111111111_1101100101110011_1101000000110000"; -- -0.1505765803942174
	pesos_i(8096) := b"0000000000000000_0000000000000000_0001100010111110_0010110010010110"; -- 0.09665182742777298
	pesos_i(8097) := b"1111111111111111_1111111111111111_1110000000010110_1001001010011101"; -- -0.12465556770226667
	pesos_i(8098) := b"1111111111111111_1111111111111111_1101010011010100_1110011111111110"; -- -0.16862630900432624
	pesos_i(8099) := b"1111111111111111_1111111111111111_1110101101110011_1101110110000010"; -- -0.08026328632148727
	pesos_i(8100) := b"0000000000000000_0000000000000000_0001100101000000_0011100100110110"; -- 0.09863622253366541
	pesos_i(8101) := b"1111111111111111_1111111111111111_1101010000110101_0010111110011110"; -- -0.17106344608260038
	pesos_i(8102) := b"0000000000000000_0000000000000000_0001001101011110_0100101111111111"; -- 0.07565760597985259
	pesos_i(8103) := b"0000000000000000_0000000000000000_0001111101001011_0000010101000110"; -- 0.12223847345742375
	pesos_i(8104) := b"1111111111111111_1111111111111111_1111010000100110_0101000110000111"; -- -0.046290306621673105
	pesos_i(8105) := b"0000000000000000_0000000000000000_0000100001100111_1011010101101010"; -- 0.03283246844072808
	pesos_i(8106) := b"1111111111111111_1111111111111111_1111010110000111_0110011110110011"; -- -0.04090263245455381
	pesos_i(8107) := b"1111111111111111_1111111111111111_1111100000101010_1110001110000111"; -- -0.030595569207633632
	pesos_i(8108) := b"1111111111111111_1111111111111111_1110011101101000_1111100101011110"; -- -0.09605447251520659
	pesos_i(8109) := b"0000000000000000_0000000000000000_0000110111001000_1100000001101101"; -- 0.05384447731216793
	pesos_i(8110) := b"0000000000000000_0000000000000000_0001100011111100_0011011000111100"; -- 0.09759844751210398
	pesos_i(8111) := b"1111111111111111_1111111111111111_1110110100100101_0111010100011111"; -- -0.0736471938026886
	pesos_i(8112) := b"1111111111111111_1111111111111111_1110101000000100_0011000000010010"; -- -0.08587359963276658
	pesos_i(8113) := b"0000000000000000_0000000000000000_0001001100001100_1011011010011010"; -- 0.07441273936840245
	pesos_i(8114) := b"1111111111111111_1111111111111111_1111001000000011_0110111000010010"; -- -0.054635162904636256
	pesos_i(8115) := b"1111111111111111_1111111111111111_1110111110011100_1000111100010100"; -- -0.06401735086941339
	pesos_i(8116) := b"1111111111111111_1111111111111111_1101101001000100_1100010011000010"; -- -0.1473881745940883
	pesos_i(8117) := b"1111111111111111_1111111111111111_1110010101010111_0001011000111001"; -- -0.10413991083634633
	pesos_i(8118) := b"0000000000000000_0000000000000000_0001001010101001_1001111101101111"; -- 0.07290073834303192
	pesos_i(8119) := b"1111111111111111_1111111111111111_1111011110100001_1110011110010110"; -- -0.032685781408008444
	pesos_i(8120) := b"1111111111111111_1111111111111111_1111000011000000_1101000010110010"; -- -0.05955787338435141
	pesos_i(8121) := b"0000000000000000_0000000000000000_0000110111111111_1100110011010110"; -- 0.05468445035480087
	pesos_i(8122) := b"0000000000000000_0000000000000000_0001101011111111_0100110100100111"; -- 0.1054580898125542
	pesos_i(8123) := b"0000000000000000_0000000000000000_0001110001100101_1010110011000100"; -- 0.11092643522250892
	pesos_i(8124) := b"1111111111111111_1111111111111111_1111111010010110_0001011100000101"; -- -0.005522309471564741
	pesos_i(8125) := b"1111111111111111_1111111111111111_1110101100101010_1001011110000111"; -- -0.08138134915434288
	pesos_i(8126) := b"1111111111111111_1111111111111111_1110010111000100_1000110111111001"; -- -0.10246956510179854
	pesos_i(8127) := b"0000000000000000_0000000000000000_0001100000000100_1001111100010110"; -- 0.0938205173811113
	pesos_i(8128) := b"0000000000000000_0000000000000000_0010000010001010_0101101001111000"; -- 0.12711110520066102
	pesos_i(8129) := b"0000000000000000_0000000000000000_0010010000101001_1110111011011011"; -- 0.14126484714371404
	pesos_i(8130) := b"1111111111111111_1111111111111111_1111100110111101_1001011111011110"; -- -0.02445078682546083
	pesos_i(8131) := b"1111111111111111_1111111111111111_1101100110101001_1111100011001101"; -- -0.14975018501707227
	pesos_i(8132) := b"1111111111111111_1111111111111111_1110110001000001_0101100011111011"; -- -0.07712787496410432
	pesos_i(8133) := b"1111111111111111_1111111111111111_1110111111100111_0111110011101010"; -- -0.0628740242289968
	pesos_i(8134) := b"1111111111111111_1111111111111111_1111010110111010_1110001111101001"; -- -0.04011703076230937
	pesos_i(8135) := b"0000000000000000_0000000000000000_0010100110101010_0111111111101100"; -- 0.16275786885583662
	pesos_i(8136) := b"0000000000000000_0000000000000000_0001100010001100_1000101000110001"; -- 0.09589446736499826
	pesos_i(8137) := b"0000000000000000_0000000000000000_0001000110011000_0100111001001100"; -- 0.06873025282825666
	pesos_i(8138) := b"1111111111111111_1111111111111111_1110101010101010_1010101010111010"; -- -0.08333332970188644
	pesos_i(8139) := b"0000000000000000_0000000000000000_0001100100001000_1110111010100000"; -- 0.0977925435542122
	pesos_i(8140) := b"0000000000000000_0000000000000000_0001011000111001_0101110100110001"; -- 0.0868128056958046
	pesos_i(8141) := b"0000000000000000_0000000000000000_0001110110001101_0010111001010001"; -- 0.11543550002742502
	pesos_i(8142) := b"0000000000000000_0000000000000000_0000100110000111_0010000000100001"; -- 0.03721810157906447
	pesos_i(8143) := b"1111111111111111_1111111111111111_1110111011011000_1001111011110000"; -- -0.06700712820074883
	pesos_i(8144) := b"1111111111111111_1111111111111111_1101011110110011_1010000111100110"; -- -0.1574152768529066
	pesos_i(8145) := b"0000000000000000_0000000000000000_0000111100111110_0010100100100000"; -- 0.059542246215349544
	pesos_i(8146) := b"1111111111111111_1111111111111111_1101111001010000_1100010101001001"; -- -0.13158003786469177
	pesos_i(8147) := b"0000000000000000_0000000000000000_0010011101110110_0111100101100001"; -- 0.15415152184964304
	pesos_i(8148) := b"0000000000000000_0000000000000000_0000010110000010_0011110100111100"; -- 0.021518542546217816
	pesos_i(8149) := b"1111111111111111_1111111111111111_1110101000100111_1011000111111011"; -- -0.08533179886089956
	pesos_i(8150) := b"0000000000000000_0000000000000000_0000101110000011_1111101110010010"; -- 0.044982646072210794
	pesos_i(8151) := b"1111111111111111_1111111111111111_1110101110100110_0101100100001110"; -- -0.07949298294221693
	pesos_i(8152) := b"0000000000000000_0000000000000000_0001111010011110_0110101010010001"; -- 0.1196047406196458
	pesos_i(8153) := b"1111111111111111_1111111111111111_1110100000111111_0100110111110110"; -- -0.09278404944943866
	pesos_i(8154) := b"0000000000000000_0000000000000000_0010110011001010_0000100011011010"; -- 0.17495780299371835
	pesos_i(8155) := b"1111111111111111_1111111111111111_1111010000110110_0000011111001011"; -- -0.046050560858520856
	pesos_i(8156) := b"1111111111111111_1111111111111111_1101110000111000_0010001010011001"; -- -0.13976844567553603
	pesos_i(8157) := b"0000000000000000_0000000000000000_0000100010110010_0001110110111100"; -- 0.033967836692282864
	pesos_i(8158) := b"1111111111111111_1111111111111111_1111101000111011_1001000000001010"; -- -0.02252864608465855
	pesos_i(8159) := b"1111111111111111_1111111111111111_1101111001111110_0100011111100111"; -- -0.13088560687917716
	pesos_i(8160) := b"0000000000000000_0000000000000000_0000000110000110_1101110100100000"; -- 0.005964107712839423
	pesos_i(8161) := b"0000000000000000_0000000000000000_0000010010001010_1101001101000100"; -- 0.017743305284409084
	pesos_i(8162) := b"1111111111111111_1111111111111111_1111111011100110_0100011100111010"; -- -0.004298733094321133
	pesos_i(8163) := b"1111111111111111_1111111111111111_1111000101111100_0001010100110111"; -- -0.056700395643184194
	pesos_i(8164) := b"0000000000000000_0000000000000000_0000101111010100_1110110100100111"; -- 0.046217748558335804
	pesos_i(8165) := b"0000000000000000_0000000000000000_0000101101110111_1100110110010111"; -- 0.04479679998222189
	pesos_i(8166) := b"0000000000000000_0000000000000000_0001111101110111_0011110001000011"; -- 0.12291313766347282
	pesos_i(8167) := b"0000000000000000_0000000000000000_0001110100001000_0111111010111111"; -- 0.11341087501373184
	pesos_i(8168) := b"1111111111111111_1111111111111111_1111011110000110_0110001010101111"; -- -0.03310569020817916
	pesos_i(8169) := b"1111111111111111_1111111111111111_1111101110100110_0001100101110111"; -- -0.016996773181084855
	pesos_i(8170) := b"0000000000000000_0000000000000000_0010011000110101_0110011101101111"; -- 0.14925238099477262
	pesos_i(8171) := b"1111111111111111_1111111111111111_1111000001100100_0001110011110110"; -- -0.060972394858640755
	pesos_i(8172) := b"0000000000000000_0000000000000000_0001001101110011_0111011101110101"; -- 0.07598063084446383
	pesos_i(8173) := b"0000000000000000_0000000000000000_0001110110111101_1000101000001100"; -- 0.11617338928631567
	pesos_i(8174) := b"1111111111111111_1111111111111111_1111110000000000_0101010010001110"; -- -0.015619960126442227
	pesos_i(8175) := b"1111111111111111_1111111111111111_1110111100100010_0011110011110101"; -- -0.06588381780600967
	pesos_i(8176) := b"0000000000000000_0000000000000000_0010010101010101_1011101110000010"; -- 0.14583942351332754
	pesos_i(8177) := b"1111111111111111_1111111111111111_1101101101010010_1101110111011100"; -- -0.14326680554134752
	pesos_i(8178) := b"1111111111111111_1111111111111111_1111010010010101_0000010101100100"; -- -0.04460111923322262
	pesos_i(8179) := b"1111111111111111_1111111111111111_1101001101101000_0111000100110111"; -- -0.17418758788940447
	pesos_i(8180) := b"0000000000000000_0000000000000000_0001011001111110_1010011111111101"; -- 0.08787012028686425
	pesos_i(8181) := b"0000000000000000_0000000000000000_0010010110101111_0000100100111011"; -- 0.14720208834002352
	pesos_i(8182) := b"0000000000000000_0000000000000000_0001101100011001_0000111110000100"; -- 0.10585114461608305
	pesos_i(8183) := b"0000000000000000_0000000000000000_0000111000111110_1111110100101000"; -- 0.05564863417630319
	pesos_i(8184) := b"1111111111111111_1111111111111111_1101100001000111_0101011011011011"; -- -0.15516144908963156
	pesos_i(8185) := b"0000000000000000_0000000000000000_0001101010111111_0100110111110100"; -- 0.10448157511508178
	pesos_i(8186) := b"1111111111111111_1111111111111111_1111101001011000_0010001011100110"; -- -0.022092646467763943
	pesos_i(8187) := b"0000000000000000_0000000000000000_0001110110110011_1111110001001000"; -- 0.11602761045340629
	pesos_i(8188) := b"1111111111111111_1111111111111111_1110100001001110_1000010101001001"; -- -0.09255186997484315
	pesos_i(8189) := b"1111111111111111_1111111111111111_1111011101100100_1110110100011011"; -- -0.03361623842099383
	pesos_i(8190) := b"0000000000000000_0000000000000000_0010101111101100_1100100110110101"; -- 0.17158184692714296
	pesos_i(8191) := b"0000000000000000_0000000000000000_0001000111010011_0011000010001001"; -- 0.06962874739101733
	pesos_i(8192) := b"1111111111111111_1111111111111111_1110000011111011_0011001110101110"; -- -0.12116696369704828
	pesos_i(8193) := b"1111111111111111_1111111111111111_1111110000101110_1111101011010111"; -- -0.014908144370054397
	pesos_i(8194) := b"1111111111111111_1111111111111111_1110110111111001_0100110000111110"; -- -0.0704147671769963
	pesos_i(8195) := b"0000000000000000_0000000000000000_0001001001011011_1011011010100010"; -- 0.07171193566245745
	pesos_i(8196) := b"0000000000000000_0000000000000000_0000111111101111_0011001000100011"; -- 0.06224358897012788
	pesos_i(8197) := b"1111111111111111_1111111111111111_1111101001100011_0011001011001000"; -- -0.021923853052800892
	pesos_i(8198) := b"0000000000000000_0000000000000000_0000001010011100_0111001101000110"; -- 0.010199741833003421
	pesos_i(8199) := b"1111111111111111_1111111111111111_1101101011010011_1100101011001011"; -- -0.14520580814599213
	pesos_i(8200) := b"1111111111111111_1111111111111111_1111010111100001_0101010001010101"; -- -0.03953049591506271
	pesos_i(8201) := b"1111111111111111_1111111111111111_1111010101110001_0100001001111001"; -- -0.04124054471274916
	pesos_i(8202) := b"0000000000000000_0000000000000000_0000010001011011_1010010000000001"; -- 0.017023325089029897
	pesos_i(8203) := b"0000000000000000_0000000000000000_0000110101000101_1111100101110110"; -- 0.05184897558104364
	pesos_i(8204) := b"0000000000000000_0000000000000000_0000010000110000_1111100011110011"; -- 0.016372260397841985
	pesos_i(8205) := b"0000000000000000_0000000000000000_0000100001100101_1101110010101011"; -- 0.03280429060483605
	pesos_i(8206) := b"0000000000000000_0000000000000000_0000011000111010_0000100001101011"; -- 0.024323011532009265
	pesos_i(8207) := b"0000000000000000_0000000000000000_0000000111101010_0110010011100011"; -- 0.007482820039348981
	pesos_i(8208) := b"1111111111111111_1111111111111111_1101101000100100_0101001111101011"; -- -0.14788318180536297
	pesos_i(8209) := b"0000000000000000_0000000000000000_0000000011011001_0010100011001110"; -- 0.0033135892976769695
	pesos_i(8210) := b"0000000000000000_0000000000000000_0000001100000100_0010000000001011"; -- 0.011781695125156658
	pesos_i(8211) := b"0000000000000000_0000000000000000_0000010100011100_0011010100011110"; -- 0.019961662057552888
	pesos_i(8212) := b"0000000000000000_0000000000000000_0001110010010101_1011111110001001"; -- 0.1116599759725442
	pesos_i(8213) := b"0000000000000000_0000000000000000_0000010010001100_0010001110010101"; -- 0.01776335140289306
	pesos_i(8214) := b"0000000000000000_0000000000000000_0001110101000100_1111111110111000"; -- 0.11433408956567533
	pesos_i(8215) := b"0000000000000000_0000000000000000_0001000000110111_0000100111001101"; -- 0.06333981755709556
	pesos_i(8216) := b"0000000000000000_0000000000000000_0000000101010101_0010100100001011"; -- 0.005205693510218446
	pesos_i(8217) := b"0000000000000000_0000000000000000_0001110011100011_1010100101001001"; -- 0.1128488352867532
	pesos_i(8218) := b"1111111111111111_1111111111111111_1111010100101100_0001111100010011"; -- -0.042295511025087974
	pesos_i(8219) := b"1111111111111111_1111111111111111_1110000000111100_1010011010011111"; -- -0.12407454115873251
	pesos_i(8220) := b"0000000000000000_0000000000000000_0001110111011000_1111111000110010"; -- 0.1165922997616667
	pesos_i(8221) := b"1111111111111111_1111111111111111_1101111010011000_1111111010011100"; -- -0.13047798815751702
	pesos_i(8222) := b"1111111111111111_1111111111111111_1111111111011000_1010001100111000"; -- -0.0006006229988983737
	pesos_i(8223) := b"0000000000000000_0000000000000000_0000111111110001_1010001000100000"; -- 0.06228078165540564
	pesos_i(8224) := b"0000000000000000_0000000000000000_0001010011000000_0100001011111101"; -- 0.08105868036190018
	pesos_i(8225) := b"1111111111111111_1111111111111111_1110110111100101_0110000011001111"; -- -0.07071871702632015
	pesos_i(8226) := b"0000000000000000_0000000000000000_0000011100000000_1011100010111010"; -- 0.02735476048014825
	pesos_i(8227) := b"1111111111111111_1111111111111111_1111010000111011_0101001110101111"; -- -0.04596974354229332
	pesos_i(8228) := b"1111111111111111_1111111111111111_1111000011010000_1110001110101000"; -- -0.0593126024476815
	pesos_i(8229) := b"0000000000000000_0000000000000000_0001110011001110_1111111111001011"; -- 0.11253355695796381
	pesos_i(8230) := b"0000000000000000_0000000000000000_0000010101110101_1101011010011100"; -- 0.02132932008746945
	pesos_i(8231) := b"0000000000000000_0000000000000000_0000111100000110_0000000001011001"; -- 0.0586853234003212
	pesos_i(8232) := b"0000000000000000_0000000000000000_0010100000111111_1001010111101001"; -- 0.157220239121795
	pesos_i(8233) := b"1111111111111111_1111111111111111_1110101111010101_0000101110000101"; -- -0.07878044127245233
	pesos_i(8234) := b"0000000000000000_0000000000000000_0001000110010010_1111000011001010"; -- 0.06864838531232463
	pesos_i(8235) := b"1111111111111111_1111111111111111_1101011111100111_0101111000101001"; -- -0.15662585732171863
	pesos_i(8236) := b"0000000000000000_0000000000000000_0001010011101111_0011011001001011"; -- 0.08177508666725823
	pesos_i(8237) := b"0000000000000000_0000000000000000_0000010111111100_1100110000100011"; -- 0.023388632450740177
	pesos_i(8238) := b"0000000000000000_0000000000000000_0000101010100000_1010011010100101"; -- 0.04151383909393852
	pesos_i(8239) := b"0000000000000000_0000000000000000_0001010101001010_1111011101001010"; -- 0.08317513987583912
	pesos_i(8240) := b"1111111111111111_1111111111111111_1110000100101101_1010011011100001"; -- -0.12039715768276572
	pesos_i(8241) := b"0000000000000000_0000000000000000_0010001101000110_1001001011010100"; -- 0.1377956167741362
	pesos_i(8242) := b"0000000000000000_0000000000000000_0001110100000001_0100000100111010"; -- 0.11330039657901891
	pesos_i(8243) := b"0000000000000000_0000000000000000_0000001110001111_1010111101101100"; -- 0.013911212857232172
	pesos_i(8244) := b"0000000000000000_0000000000000000_0001011000001101_1101001111001111"; -- 0.08614848899019567
	pesos_i(8245) := b"1111111111111111_1111111111111111_1111111100111110_1001100011101110"; -- -0.0029510897202629084
	pesos_i(8246) := b"1111111111111111_1111111111111111_1110000110011010_1101010100111110"; -- -0.11873118634267425
	pesos_i(8247) := b"1111111111111111_1111111111111111_1110110000011111_0001100110011010"; -- -0.0776504515468845
	pesos_i(8248) := b"1111111111111111_1111111111111111_1111100101101110_0101101100111101"; -- -0.025659844946069262
	pesos_i(8249) := b"0000000000000000_0000000000000000_0001000101101001_1101110110000110"; -- 0.0680216266999526
	pesos_i(8250) := b"1111111111111111_1111111111111111_1110110000100100_0010010010011010"; -- -0.07757350200604958
	pesos_i(8251) := b"0000000000000000_0000000000000000_0001110000000100_0001010001001010"; -- 0.10943724453823936
	pesos_i(8252) := b"0000000000000000_0000000000000000_0000000000101011_1011000001111011"; -- 0.0006666468868702463
	pesos_i(8253) := b"1111111111111111_1111111111111111_1111000111111110_0100011001111010"; -- -0.05471381685000536
	pesos_i(8254) := b"0000000000000000_0000000000000000_0001011110001001_1011000000101011"; -- 0.09194470457994007
	pesos_i(8255) := b"1111111111111111_1111111111111111_1111100100101110_1100111101011111"; -- -0.026629485476487115
	pesos_i(8256) := b"0000000000000000_0000000000000000_0000111011111011_0011010011010011"; -- 0.058520604537770915
	pesos_i(8257) := b"0000000000000000_0000000000000000_0001011000001000_0101001110010000"; -- 0.08606455094443072
	pesos_i(8258) := b"1111111111111111_1111111111111111_1101101011100010_1001101001111101"; -- -0.14497980554936638
	pesos_i(8259) := b"1111111111111111_1111111111111111_1111100100101000_1101001100010000"; -- -0.026720818233991396
	pesos_i(8260) := b"1111111111111111_1111111111111111_1111101000101000_1110000100100110"; -- -0.022813728508980287
	pesos_i(8261) := b"1111111111111111_1111111111111111_1110000101000000_1110010101010001"; -- -0.12010351914536545
	pesos_i(8262) := b"0000000000000000_0000000000000000_0001100101110100_1100110001011111"; -- 0.09943845088554085
	pesos_i(8263) := b"0000000000000000_0000000000000000_0000101000001011_0001011110111000"; -- 0.03923176053146882
	pesos_i(8264) := b"1111111111111111_1111111111111111_1111100101011001_0100010000110001"; -- -0.025981653207130362
	pesos_i(8265) := b"0000000000000000_0000000000000000_0000101101110110_1111010000100011"; -- 0.044783838736752936
	pesos_i(8266) := b"0000000000000000_0000000000000000_0010001110100011_1000011101101101"; -- 0.13921400470662412
	pesos_i(8267) := b"0000000000000000_0000000000000000_0000111100010000_1001011100001010"; -- 0.05884689327409383
	pesos_i(8268) := b"1111111111111111_1111111111111111_1111010110101011_1010111111011111"; -- -0.040349014282646437
	pesos_i(8269) := b"0000000000000000_0000000000000000_0000011101111000_0111100101011101"; -- 0.02918203855907261
	pesos_i(8270) := b"1111111111111111_1111111111111111_1101111000100110_1100110110010000"; -- -0.13222041351741745
	pesos_i(8271) := b"0000000000000000_0000000000000000_0000001000111101_1011011111111110"; -- 0.00875425296584279
	pesos_i(8272) := b"0000000000000000_0000000000000000_0000000000011111_1111001100001000"; -- 0.00048750829357580304
	pesos_i(8273) := b"0000000000000000_0000000000000000_0001100001001111_1110001010011000"; -- 0.09496895045198141
	pesos_i(8274) := b"0000000000000000_0000000000000000_0000011011011010_1110111101000010"; -- 0.026778176994500785
	pesos_i(8275) := b"0000000000000000_0000000000000000_0001010101000111_1100101101001101"; -- 0.08312674164904975
	pesos_i(8276) := b"0000000000000000_0000000000000000_0010000101010011_1100010100111111"; -- 0.13018448616206424
	pesos_i(8277) := b"1111111111111111_1111111111111111_1110010101000110_1110010101001000"; -- -0.10438696863277022
	pesos_i(8278) := b"1111111111111111_1111111111111111_1111110101101000_1011011111100111"; -- -0.010120874504959443
	pesos_i(8279) := b"1111111111111111_1111111111111111_1111110011010001_1111101110010100"; -- -0.012420917883121236
	pesos_i(8280) := b"0000000000000000_0000000000000000_0000001110011000_1111111011100101"; -- 0.01405327888961681
	pesos_i(8281) := b"0000000000000000_0000000000000000_0000000000101110_0110011011010100"; -- 0.0007080332998880462
	pesos_i(8282) := b"0000000000000000_0000000000000000_0001010101100111_0101000010010010"; -- 0.08360770768699176
	pesos_i(8283) := b"1111111111111111_1111111111111111_1101101111000010_0010000000101010"; -- -0.14156912790405748
	pesos_i(8284) := b"0000000000000000_0000000000000000_0010000100011110_1111011001111101"; -- 0.12937870562898576
	pesos_i(8285) := b"1111111111111111_1111111111111111_1111110101000010_1000001010010100"; -- -0.010703886925525848
	pesos_i(8286) := b"0000000000000000_0000000000000000_0000011001000100_1111100011111101"; -- 0.024489938605634986
	pesos_i(8287) := b"0000000000000000_0000000000000000_0000000001100111_0100111101101110"; -- 0.001576389755309708
	pesos_i(8288) := b"1111111111111111_1111111111111111_1111110100110001_1001100010100111"; -- -0.010961970536725643
	pesos_i(8289) := b"1111111111111111_1111111111111111_1101111000010001_1100101100011100"; -- -0.1325409942470623
	pesos_i(8290) := b"0000000000000000_0000000000000000_0001011001000001_1001100011000010"; -- 0.0869384262799171
	pesos_i(8291) := b"0000000000000000_0000000000000000_0001010001000110_1111111000101001"; -- 0.07920826434062954
	pesos_i(8292) := b"0000000000000000_0000000000000000_0001100011110000_1111010101100111"; -- 0.09742673654848164
	pesos_i(8293) := b"1111111111111111_1111111111111111_1110100101011111_1001100011010111"; -- -0.08838505496489274
	pesos_i(8294) := b"0000000000000000_0000000000000000_0001000110111011_1111101001100100"; -- 0.06927456794004563
	pesos_i(8295) := b"1111111111111111_1111111111111111_1111000111111010_0011011000000010"; -- -0.054775833565456074
	pesos_i(8296) := b"0000000000000000_0000000000000000_0001110011011110_0000111110010110"; -- 0.11276338022160948
	pesos_i(8297) := b"1111111111111111_1111111111111111_1111110001000101_1010000011011011"; -- -0.01456255585595431
	pesos_i(8298) := b"0000000000000000_0000000000000000_0000100110000000_0100111000000011"; -- 0.03711402479371814
	pesos_i(8299) := b"1111111111111111_1111111111111111_1111001110100111_0001110110011010"; -- -0.048231267818818854
	pesos_i(8300) := b"0000000000000000_0000000000000000_0000000010101010_1000100101110111"; -- 0.0026021875821781617
	pesos_i(8301) := b"0000000000000000_0000000000000000_0000110000001100_1011111100001110"; -- 0.047069493282955094
	pesos_i(8302) := b"0000000000000000_0000000000000000_0001101001000110_1011000010111110"; -- 0.10264114993228134
	pesos_i(8303) := b"1111111111111111_1111111111111111_1110011010001011_0100110000011100"; -- -0.09943699182882867
	pesos_i(8304) := b"0000000000000000_0000000000000000_0001101110111111_0101110000001001"; -- 0.10838866443301931
	pesos_i(8305) := b"1111111111111111_1111111111111111_1110101011101001_0110010110111000"; -- -0.08237613912663702
	pesos_i(8306) := b"0000000000000000_0000000000000000_0000010101010101_1100010111001100"; -- 0.020840036769931198
	pesos_i(8307) := b"0000000000000000_0000000000000000_0000011100111000_0000100000111110"; -- 0.028198733437896306
	pesos_i(8308) := b"0000000000000000_0000000000000000_0001110101010000_1000010000010110"; -- 0.11450982616190333
	pesos_i(8309) := b"1111111111111111_1111111111111111_1111001001000011_0011110110000011"; -- -0.05366149468420722
	pesos_i(8310) := b"0000000000000000_0000000000000000_0001010010101100_1100110110011100"; -- 0.08076176702896132
	pesos_i(8311) := b"0000000000000000_0000000000000000_0001001111111111_1010001011001100"; -- 0.07811944468959975
	pesos_i(8312) := b"1111111111111111_1111111111111111_1110111101001000_1101100010001001"; -- -0.06529471060857424
	pesos_i(8313) := b"0000000000000000_0000000000000000_0000001111000100_1101111110000101"; -- 0.014722795371631708
	pesos_i(8314) := b"0000000000000000_0000000000000000_0010010110000111_0001100000001010"; -- 0.14659261928805717
	pesos_i(8315) := b"1111111111111111_1111111111111111_1111101001010111_1011101011001010"; -- -0.022098851741498636
	pesos_i(8316) := b"0000000000000000_0000000000000000_0000111001001001_0100111001101010"; -- 0.05580606546038658
	pesos_i(8317) := b"0000000000000000_0000000000000000_0000000101111110_0111000111010100"; -- 0.005835642215357075
	pesos_i(8318) := b"1111111111111111_1111111111111111_1110010101111100_1011011111101010"; -- -0.10356569793532963
	pesos_i(8319) := b"0000000000000000_0000000000000000_0000100010111000_0100010001100000"; -- 0.03406169274143427
	pesos_i(8320) := b"1111111111111111_1111111111111111_1111100001011101_1001110111010001"; -- -0.029821526087237177
	pesos_i(8321) := b"1111111111111111_1111111111111111_1111110111110011_1101010001111100"; -- -0.007998199103179202
	pesos_i(8322) := b"0000000000000000_0000000000000000_0000101010011111_0000111010100011"; -- 0.04148951986416667
	pesos_i(8323) := b"1111111111111111_1111111111111111_1111001000101100_0010100010010001"; -- -0.054013695307370026
	pesos_i(8324) := b"0000000000000000_0000000000000000_0000011100111111_0100001010111110"; -- 0.028309031928362066
	pesos_i(8325) := b"0000000000000000_0000000000000000_0000000100111001_0001110010010000"; -- 0.004777703438984904
	pesos_i(8326) := b"1111111111111111_1111111111111111_1110100110011010_0011101111010101"; -- -0.08749033018831151
	pesos_i(8327) := b"0000000000000000_0000000000000000_0000111000111111_1111100110000001"; -- 0.05566367537887415
	pesos_i(8328) := b"1111111111111111_1111111111111111_1110000000010001_1000111100000101"; -- -0.12473207596987886
	pesos_i(8329) := b"1111111111111111_1111111111111111_1110111011101111_0110000000011011"; -- -0.06665992104898033
	pesos_i(8330) := b"1111111111111111_1111111111111111_1110110000111110_1101100110100001"; -- -0.07716598328565791
	pesos_i(8331) := b"0000000000000000_0000000000000000_0001001000000101_1010111100110000"; -- 0.07039923582906776
	pesos_i(8332) := b"1111111111111111_1111111111111111_1110111101101100_1000001100100110"; -- -0.06475048370672237
	pesos_i(8333) := b"1111111111111111_1111111111111111_1101111101111001_1101111011100011"; -- -0.12704665151168587
	pesos_i(8334) := b"0000000000000000_0000000000000000_0010100011100110_1111111011110000"; -- 0.15977471687710668
	pesos_i(8335) := b"1111111111111111_1111111111111111_1110011101000000_1111111001100000"; -- -0.09666452549835683
	pesos_i(8336) := b"0000000000000000_0000000000000000_0001010001001010_1000001111101011"; -- 0.07926201335346894
	pesos_i(8337) := b"1111111111111111_1111111111111111_1111111000101001_0100000011001100"; -- -0.007183027420306507
	pesos_i(8338) := b"0000000000000000_0000000000000000_0001100101010100_0000111110010001"; -- 0.09893891600850092
	pesos_i(8339) := b"1111111111111111_1111111111111111_1111000101010110_0000100111001011"; -- -0.05728091052877605
	pesos_i(8340) := b"1111111111111111_1111111111111111_1111010100100011_1100010011101001"; -- -0.042422955529224864
	pesos_i(8341) := b"1111111111111111_1111111111111111_1111010100110011_1110101110100011"; -- -0.04217650676719866
	pesos_i(8342) := b"0000000000000000_0000000000000000_0001101000101001_0010111101110101"; -- 0.10219093903370148
	pesos_i(8343) := b"1111111111111111_1111111111111111_1101011101111001_1110001100110000"; -- -0.1582963950309009
	pesos_i(8344) := b"1111111111111111_1111111111111111_1110100101101111_0110010100010100"; -- -0.0881439997989388
	pesos_i(8345) := b"1111111111111111_1111111111111111_1110110111001100_1011000010011101"; -- -0.0710954299851038
	pesos_i(8346) := b"1111111111111111_1111111111111111_1101110110000010_1001101111001000"; -- -0.13472582212574072
	pesos_i(8347) := b"0000000000000000_0000000000000000_0001111010011110_1100001011000010"; -- 0.11960999718887844
	pesos_i(8348) := b"0000000000000000_0000000000000000_0000111011011111_0100111010110111"; -- 0.05809490173487155
	pesos_i(8349) := b"0000000000000000_0000000000000000_0000010111010000_0011111110100111"; -- 0.022708872149688714
	pesos_i(8350) := b"1111111111111111_1111111111111111_1111001100110100_1010011101111100"; -- -0.04997781023769945
	pesos_i(8351) := b"0000000000000000_0000000000000000_0001100111100011_0110100100101000"; -- 0.10112626281114986
	pesos_i(8352) := b"0000000000000000_0000000000000000_0001100100011111_0100010001000001"; -- 0.09813334069010762
	pesos_i(8353) := b"1111111111111111_1111111111111111_1110011001000101_0000101010100001"; -- -0.10050900995302667
	pesos_i(8354) := b"0000000000000000_0000000000000000_0010100101010000_1000010000010101"; -- 0.16138482580488445
	pesos_i(8355) := b"0000000000000000_0000000000000000_0010001010011001_0001111001100111"; -- 0.13514890681755795
	pesos_i(8356) := b"1111111111111111_1111111111111111_1111000000101101_0101100101101111"; -- -0.061808023737674064
	pesos_i(8357) := b"1111111111111111_1111111111111111_1111110110011011_0110011101110111"; -- -0.009347470691870016
	pesos_i(8358) := b"1111111111111111_1111111111111111_1110001100110000_1000111101001001"; -- -0.11254028772206497
	pesos_i(8359) := b"0000000000000000_0000000000000000_0010001111010001_0101011100001110"; -- 0.1399130258475024
	pesos_i(8360) := b"1111111111111111_1111111111111111_1111101101000010_0100001001001010"; -- -0.018520218871932524
	pesos_i(8361) := b"0000000000000000_0000000000000000_0000001011011100_1000111110111110"; -- 0.011178001392066227
	pesos_i(8362) := b"1111111111111111_1111111111111111_1101101011011000_1011001101101101"; -- -0.14513090701573328
	pesos_i(8363) := b"1111111111111111_1111111111111111_1101011101010110_1000110011011011"; -- -0.15883559852718543
	pesos_i(8364) := b"1111111111111111_1111111111111111_1101100010101001_1111010100101000"; -- -0.1536566520906537
	pesos_i(8365) := b"0000000000000000_0000000000000000_0001110101001001_1010010001010011"; -- 0.11440493610882226
	pesos_i(8366) := b"0000000000000000_0000000000000000_0010000110001111_0110001000001010"; -- 0.13109410041050315
	pesos_i(8367) := b"0000000000000000_0000000000000000_0010000111001110_0110100011100101"; -- 0.1320558126483991
	pesos_i(8368) := b"1111111111111111_1111111111111111_1111101110110100_0000000010010110"; -- -0.016784633000334167
	pesos_i(8369) := b"0000000000000000_0000000000000000_0000010111100100_1011101010111010"; -- 0.023021383646599943
	pesos_i(8370) := b"1111111111111111_1111111111111111_1110101001111100_0110010111100001"; -- -0.08403933769199665
	pesos_i(8371) := b"1111111111111111_1111111111111111_1110100101110010_1001000110010011"; -- -0.08809557111016589
	pesos_i(8372) := b"0000000000000000_0000000000000000_0001010010000111_0000001101001011"; -- 0.08018513273945065
	pesos_i(8373) := b"1111111111111111_1111111111111111_1110001011011101_1111101001001111"; -- -0.11380038797920584
	pesos_i(8374) := b"0000000000000000_0000000000000000_0000110000011011_0011110010101011"; -- 0.04729060347170976
	pesos_i(8375) := b"0000000000000000_0000000000000000_0010001000001101_1111000100010100"; -- 0.13302523371239527
	pesos_i(8376) := b"1111111111111111_1111111111111111_1111010010110101_1010001010001000"; -- -0.044103471623653
	pesos_i(8377) := b"1111111111111111_1111111111111111_1111011011111100_0111101101110010"; -- -0.0352099272052801
	pesos_i(8378) := b"1111111111111111_1111111111111111_1110110010111001_1011101101101111"; -- -0.07529095212435981
	pesos_i(8379) := b"0000000000000000_0000000000000000_0001010110010001_0011000100011001"; -- 0.08424670096597908
	pesos_i(8380) := b"0000000000000000_0000000000000000_0000011101101101_0000001110010011"; -- 0.029007170960084133
	pesos_i(8381) := b"0000000000000000_0000000000000000_0000010101100101_1000000011100000"; -- 0.021080069249602602
	pesos_i(8382) := b"1111111111111111_1111111111111111_1110110110010111_1010111001001111"; -- -0.0719042833141604
	pesos_i(8383) := b"0000000000000000_0000000000000000_0000001111010110_0101111110110111"; -- 0.014989835889879555
	pesos_i(8384) := b"1111111111111111_1111111111111111_1101110100101001_1100100001100110"; -- -0.13608119489081408
	pesos_i(8385) := b"1111111111111111_1111111111111111_1111011101010110_0110110010011010"; -- -0.033837520964146384
	pesos_i(8386) := b"0000000000000000_0000000000000000_0000110011011000_0111000011111001"; -- 0.05017763213847548
	pesos_i(8387) := b"1111111111111111_1111111111111111_1111011111001000_1001000000110100"; -- -0.03209589711721361
	pesos_i(8388) := b"0000000000000000_0000000000000000_0000101110110100_1010101001011011"; -- 0.04572548605748224
	pesos_i(8389) := b"0000000000000000_0000000000000000_0001010010000011_1010011010110001"; -- 0.080133836894276
	pesos_i(8390) := b"1111111111111111_1111111111111111_1101111101010001_0000111010001000"; -- -0.12766942191667807
	pesos_i(8391) := b"0000000000000000_0000000000000000_0000111110110000_1101101000101011"; -- 0.06129230077540473
	pesos_i(8392) := b"0000000000000000_0000000000000000_0010000001000010_1110110000100111"; -- 0.12602115578777165
	pesos_i(8393) := b"0000000000000000_0000000000000000_0000111001010010_0100100001001010"; -- 0.05594302947931356
	pesos_i(8394) := b"0000000000000000_0000000000000000_0010001100010111_0001001000010100"; -- 0.1370707797744766
	pesos_i(8395) := b"0000000000000000_0000000000000000_0001001110000100_1110000111001110"; -- 0.07624636927356386
	pesos_i(8396) := b"0000000000000000_0000000000000000_0000101001011110_1011110111110010"; -- 0.040508147779627836
	pesos_i(8397) := b"0000000000000000_0000000000000000_0010010101110101_0000010110101000"; -- 0.14631686544075884
	pesos_i(8398) := b"0000000000000000_0000000000000000_0001001000001110_1001000011101010"; -- 0.07053476069743111
	pesos_i(8399) := b"0000000000000000_0000000000000000_0000011010110110_0010100110101111"; -- 0.026217084064255526
	pesos_i(8400) := b"0000000000000000_0000000000000000_0001100110110110_1101001110001000"; -- 0.10044595788979768
	pesos_i(8401) := b"1111111111111111_1111111111111111_1111000101001010_1111011000001101"; -- -0.057449933931628366
	pesos_i(8402) := b"0000000000000000_0000000000000000_0001111110011010_1101001100010000"; -- 0.12345618372799186
	pesos_i(8403) := b"1111111111111111_1111111111111111_1111000101001100_1000100001001000"; -- -0.05742595894438161
	pesos_i(8404) := b"1111111111111111_1111111111111111_1110010011001110_1000001000010001"; -- -0.10622393678302684
	pesos_i(8405) := b"0000000000000000_0000000000000000_0000000010111001_1001000110110110"; -- 0.0028315609810353544
	pesos_i(8406) := b"1111111111111111_1111111111111111_1110010101101101_0011010111001110"; -- -0.10380233500108473
	pesos_i(8407) := b"1111111111111111_1111111111111111_1101011011010101_0100110110011011"; -- -0.16080775232624092
	pesos_i(8408) := b"1111111111111111_1111111111111111_1110010100110000_1110001011110001"; -- -0.10472280135798775
	pesos_i(8409) := b"1111111111111111_1111111111111111_1111110010101010_1000000000000101"; -- -0.013023375256290307
	pesos_i(8410) := b"0000000000000000_0000000000000000_0001001110111011_1110100010000011"; -- 0.07708600228907012
	pesos_i(8411) := b"0000000000000000_0000000000000000_0000101110110001_1010010111100110"; -- 0.0456794440724962
	pesos_i(8412) := b"1111111111111111_1111111111111111_1111101000111111_1111010000100000"; -- -0.022461645395387368
	pesos_i(8413) := b"1111111111111111_1111111111111111_1101110111001110_0111010001101000"; -- -0.13356850103212814
	pesos_i(8414) := b"1111111111111111_1111111111111111_1110000110100001_1111101000010010"; -- -0.11862217959801839
	pesos_i(8415) := b"1111111111111111_1111111111111111_1111111110011010_1001101010000110"; -- -0.001547186108322081
	pesos_i(8416) := b"0000000000000000_0000000000000000_0000000000010011_0111000101010011"; -- 0.00029667161037519183
	pesos_i(8417) := b"0000000000000000_0000000000000000_0000001001100100_1110000000001111"; -- 0.009351733815907535
	pesos_i(8418) := b"1111111111111111_1111111111111111_1101110000011001_0010101011100001"; -- -0.1402409745432524
	pesos_i(8419) := b"1111111111111111_1111111111111111_1110101011101001_1011110011001000"; -- -0.0823709499470643
	pesos_i(8420) := b"0000000000000000_0000000000000000_0000100000101010_1110010011100010"; -- 0.03190451156321117
	pesos_i(8421) := b"1111111111111111_1111111111111111_1111110111000100_1100110100001000"; -- -0.008715806562013498
	pesos_i(8422) := b"0000000000000000_0000000000000000_0010010111100110_1111001110111001"; -- 0.14805529858460215
	pesos_i(8423) := b"1111111111111111_1111111111111111_1111011001101110_0010010001111011"; -- -0.03738185874085173
	pesos_i(8424) := b"1111111111111111_1111111111111111_1111000110110010_1011000110111110"; -- -0.055867091383848946
	pesos_i(8425) := b"0000000000000000_0000000000000000_0000111001110100_0110100001110000"; -- 0.056463744405204484
	pesos_i(8426) := b"0000000000000000_0000000000000000_0000101110100111_0100011011100111"; -- 0.045521193919464145
	pesos_i(8427) := b"1111111111111111_1111111111111111_1110101101100101_1110110001010101"; -- -0.08047602585790359
	pesos_i(8428) := b"1111111111111111_1111111111111111_1110100110100000_1100000011000000"; -- -0.08739085489392819
	pesos_i(8429) := b"1111111111111111_1111111111111111_1110111111101011_1100011010000100"; -- -0.06280860218663788
	pesos_i(8430) := b"1111111111111111_1111111111111111_1101100011001110_0101001001100111"; -- -0.1531017777932323
	pesos_i(8431) := b"0000000000000000_0000000000000000_0001011010101011_0100000001100111"; -- 0.08855059161376887
	pesos_i(8432) := b"1111111111111111_1111111111111111_1111000101010010_0011101100100111"; -- -0.05733900361285343
	pesos_i(8433) := b"1111111111111111_1111111111111111_1101110011010100_1111000000111001"; -- -0.13737581822900274
	pesos_i(8434) := b"1111111111111111_1111111111111111_1110011011101110_0000100111101100"; -- -0.0979303169274183
	pesos_i(8435) := b"0000000000000000_0000000000000000_0001110110011101_0000110010000001"; -- 0.11567762527126906
	pesos_i(8436) := b"0000000000000000_0000000000000000_0000111011100110_1001010010110011"; -- 0.05820588455131626
	pesos_i(8437) := b"0000000000000000_0000000000000000_0001000111101100_0001111111101010"; -- 0.0700092265256694
	pesos_i(8438) := b"1111111111111111_1111111111111111_1111100000000100_1000110011110001"; -- -0.031180564000244784
	pesos_i(8439) := b"1111111111111111_1111111111111111_1111111010100001_0110111000110001"; -- -0.005349267001675484
	pesos_i(8440) := b"0000000000000000_0000000000000000_0001101110001001_1101100110011010"; -- 0.10757217424695993
	pesos_i(8441) := b"1111111111111111_1111111111111111_1110010011011110_0100011101101001"; -- -0.10598329249017503
	pesos_i(8442) := b"1111111111111111_1111111111111111_1110000010110010_0000010101000000"; -- -0.12228362262826369
	pesos_i(8443) := b"0000000000000000_0000000000000000_0000101000001000_0100000101101101"; -- 0.039188469994811743
	pesos_i(8444) := b"0000000000000000_0000000000000000_0001010011101111_1101011010100100"; -- 0.08178464422495572
	pesos_i(8445) := b"0000000000000000_0000000000000000_0000011000110101_1010111101000001"; -- 0.024256661691755606
	pesos_i(8446) := b"0000000000000000_0000000000000000_0001101110001110_1100101000101100"; -- 0.10764754848960309
	pesos_i(8447) := b"1111111111111111_1111111111111111_1110110101010111_1000000100001101"; -- -0.07288354339525589
	pesos_i(8448) := b"0000000000000000_0000000000000000_0000101100111111_0110111100010011"; -- 0.0439366743401382
	pesos_i(8449) := b"1111111111111111_1111111111111111_1110001001011000_1011010101100110"; -- -0.11583391442516992
	pesos_i(8450) := b"0000000000000000_0000000000000000_0001000110101010_1101101111111011"; -- 0.06901335591714444
	pesos_i(8451) := b"1111111111111111_1111111111111111_1110111110011110_0111010000001111"; -- -0.06398844367348341
	pesos_i(8452) := b"1111111111111111_1111111111111111_1101100000100010_1011100001100110"; -- -0.1557202101183216
	pesos_i(8453) := b"0000000000000000_0000000000000000_0000000100100001_0010111110101100"; -- 0.00441263156013477
	pesos_i(8454) := b"0000000000000000_0000000000000000_0000011000110011_1001011100110111"; -- 0.02422471141540175
	pesos_i(8455) := b"0000000000000000_0000000000000000_0000000011001011_1001011100100011"; -- 0.003106542579480047
	pesos_i(8456) := b"0000000000000000_0000000000000000_0010001001110011_1010100000000011"; -- 0.1345772750659583
	pesos_i(8457) := b"0000000000000000_0000000000000000_0000011110111000_0101111000110011"; -- 0.030156981972328748
	pesos_i(8458) := b"0000000000000000_0000000000000000_0001010010011011_1000000100010011"; -- 0.08049780574080616
	pesos_i(8459) := b"0000000000000000_0000000000000000_0000101101011011_1111111011000100"; -- 0.044372485132233
	pesos_i(8460) := b"0000000000000000_0000000000000000_0001000001111111_1111011000110111"; -- 0.06445254173179217
	pesos_i(8461) := b"1111111111111111_1111111111111111_1110000100111110_0110010010111100"; -- -0.1201417008166458
	pesos_i(8462) := b"0000000000000000_0000000000000000_0000001110011001_1101010111000000"; -- 0.014066085223986185
	pesos_i(8463) := b"0000000000000000_0000000000000000_0000001000011011_1010010100001111"; -- 0.008234325566997873
	pesos_i(8464) := b"0000000000000000_0000000000000000_0001000111111011_1001011010011001"; -- 0.07024518239636449
	pesos_i(8465) := b"0000000000000000_0000000000000000_0000001011100000_1110000110101100"; -- 0.011243919726821762
	pesos_i(8466) := b"1111111111111111_1111111111111111_1110101011111101_1000100100001010"; -- -0.08206885818797034
	pesos_i(8467) := b"0000000000000000_0000000000000000_0000101011010101_0001001000101011"; -- 0.04231370505508246
	pesos_i(8468) := b"0000000000000000_0000000000000000_0010110110101101_1110000011110000"; -- 0.1784344279139567
	pesos_i(8469) := b"1111111111111111_1111111111111111_1111001111011011_0101010010100110"; -- -0.047434529701088114
	pesos_i(8470) := b"1111111111111111_1111111111111111_1111011101101010_0111100100110110"; -- -0.033531593738950316
	pesos_i(8471) := b"0000000000000000_0000000000000000_0001100101111010_1001010100110110"; -- 0.0995267158797069
	pesos_i(8472) := b"0000000000000000_0000000000000000_0000110100101011_0101110000010011"; -- 0.05144286601333527
	pesos_i(8473) := b"1111111111111111_1111111111111111_1110111001010010_1010010001101000"; -- -0.0690514799684162
	pesos_i(8474) := b"0000000000000000_0000000000000000_0001100010110101_0000110101110001"; -- 0.09651264204203444
	pesos_i(8475) := b"1111111111111111_1111111111111111_1111100100100110_1011010001111111"; -- -0.026753157618051047
	pesos_i(8476) := b"1111111111111111_1111111111111111_1111000000111010_0111001010111111"; -- -0.06160815079807923
	pesos_i(8477) := b"1111111111111111_1111111111111111_1111010110011011_1101011011100111"; -- -0.04059082861594338
	pesos_i(8478) := b"1111111111111111_1111111111111111_1110101101100101_0001111010000110"; -- -0.08048829303832417
	pesos_i(8479) := b"0000000000000000_0000000000000000_0001110000010111_0111011011000001"; -- 0.1097330305148305
	pesos_i(8480) := b"0000000000000000_0000000000000000_0001010101101100_0101000001100101"; -- 0.0836839911334392
	pesos_i(8481) := b"0000000000000000_0000000000000000_0001001100001011_1100010000110101"; -- 0.07439829149694026
	pesos_i(8482) := b"1111111111111111_1111111111111111_1111110010101100_1100111100100111"; -- -0.01298814104160187
	pesos_i(8483) := b"0000000000000000_0000000000000000_0001101110000010_0100000110100010"; -- 0.1074563045398002
	pesos_i(8484) := b"0000000000000000_0000000000000000_0001010111011100_1001000001101111"; -- 0.08539679256979064
	pesos_i(8485) := b"1111111111111111_1111111111111111_1111110000010010_0110010100011110"; -- -0.015344314712523325
	pesos_i(8486) := b"1111111111111111_1111111111111111_1110010011011101_0001000100011101"; -- -0.10600178754249337
	pesos_i(8487) := b"0000000000000000_0000000000000000_0000100000011011_1100000100111000"; -- 0.03167350407061622
	pesos_i(8488) := b"0000000000000000_0000000000000000_0000010101000111_1101101010011011"; -- 0.020627653854172128
	pesos_i(8489) := b"1111111111111111_1111111111111111_1101011110011101_0110111001001111"; -- -0.1577540451902287
	pesos_i(8490) := b"1111111111111111_1111111111111111_1111110111000101_0000010111101101"; -- -0.008712415436590699
	pesos_i(8491) := b"1111111111111111_1111111111111111_1111011000110000_1001100101101000"; -- -0.0383209343610914
	pesos_i(8492) := b"0000000000000000_0000000000000000_0000000100100001_0110000110110001"; -- 0.004415612861809508
	pesos_i(8493) := b"1111111111111111_1111111111111111_1110001101101100_0011001100100010"; -- -0.1116302530894504
	pesos_i(8494) := b"0000000000000000_0000000000000000_0010011011111101_0001100111010100"; -- 0.15229951307343267
	pesos_i(8495) := b"1111111111111111_1111111111111111_1111010010101110_0110010111011110"; -- -0.04421389901264241
	pesos_i(8496) := b"0000000000000000_0000000000000000_0010010101000100_0000101110000010"; -- 0.14556953359967578
	pesos_i(8497) := b"1111111111111111_1111111111111111_1111101101111000_0111101001001101"; -- -0.017692905528054276
	pesos_i(8498) := b"1111111111111111_1111111111111111_1111010111000010_0111001001101000"; -- -0.04000172579291724
	pesos_i(8499) := b"1111111111111111_1111111111111111_1111011000101101_1000100100001000"; -- -0.038367686712623035
	pesos_i(8500) := b"0000000000000000_0000000000000000_0000000000010100_0101100000011010"; -- 0.00031042711976760664
	pesos_i(8501) := b"0000000000000000_0000000000000000_0010100111110100_1111011011110111"; -- 0.16389411476829766
	pesos_i(8502) := b"1111111111111111_1111111111111111_1111110111010101_0111100101010011"; -- -0.008461396522644278
	pesos_i(8503) := b"1111111111111111_1111111111111111_1111111101111011_0110010100100101"; -- -0.002023390221074747
	pesos_i(8504) := b"1111111111111111_1111111111111111_1110000100000101_0111100111100110"; -- -0.12101019026946087
	pesos_i(8505) := b"0000000000000000_0000000000000000_0010010011100110_0110010010100000"; -- 0.1441405191301443
	pesos_i(8506) := b"1111111111111111_1111111111111111_1101111101101110_0101010010100001"; -- -0.12722273893044758
	pesos_i(8507) := b"1111111111111111_1111111111111111_1110000100110001_0001101110111100"; -- -0.12034441624122251
	pesos_i(8508) := b"1111111111111111_1111111111111111_1101101001001100_1000001010010101"; -- -0.14727004878877897
	pesos_i(8509) := b"0000000000000000_0000000000000000_0000111101100100_0011001100010100"; -- 0.06012267338883266
	pesos_i(8510) := b"1111111111111111_1111111111111111_1110111111000111_1110001000111001"; -- -0.0633562670178231
	pesos_i(8511) := b"1111111111111111_1111111111111111_1101101001001011_1011111000110111"; -- -0.14728175315634537
	pesos_i(8512) := b"1111111111111111_1111111111111111_1101111101111011_1100101000110011"; -- -0.1270173668869629
	pesos_i(8513) := b"0000000000000000_0000000000000000_0000101111110011_1111001100110001"; -- 0.046691131119009965
	pesos_i(8514) := b"1111111111111111_1111111111111111_1110010011001001_1111010001111100"; -- -0.10629341104210255
	pesos_i(8515) := b"1111111111111111_1111111111111111_1111110111010101_1101110110111111"; -- -0.00845541094229455
	pesos_i(8516) := b"1111111111111111_1111111111111111_1110101011010110_1011100110110010"; -- -0.08266105085479708
	pesos_i(8517) := b"0000000000000000_0000000000000000_0001101111100100_1010100111100010"; -- 0.10895787974614828
	pesos_i(8518) := b"1111111111111111_1111111111111111_1110110011101001_1100111101100111"; -- -0.07455734002997719
	pesos_i(8519) := b"0000000000000000_0000000000000000_0000100011110111_1011010000000110"; -- 0.035029651223554906
	pesos_i(8520) := b"1111111111111111_1111111111111111_1101101111111001_1101001010011011"; -- -0.14071925835156718
	pesos_i(8521) := b"0000000000000000_0000000000000000_0000101011010011_1001111111100100"; -- 0.04229163468266248
	pesos_i(8522) := b"0000000000000000_0000000000000000_0001101011010011_0101110100010001"; -- 0.10478765158701067
	pesos_i(8523) := b"0000000000000000_0000000000000000_0001011001011111_1010011010000111"; -- 0.08739701080902372
	pesos_i(8524) := b"0000000000000000_0000000000000000_0001010101011000_0001110111011100"; -- 0.08337580312136889
	pesos_i(8525) := b"1111111111111111_1111111111111111_1111110001111110_1001110110001001"; -- -0.013693002705650516
	pesos_i(8526) := b"0000000000000000_0000000000000000_0000110001100111_0010001011110111"; -- 0.04844873941945127
	pesos_i(8527) := b"0000000000000000_0000000000000000_0000101101110101_0101001100111000"; -- 0.04475898849826402
	pesos_i(8528) := b"1111111111111111_1111111111111111_1111101010001101_1111100001010110"; -- -0.021271208741932248
	pesos_i(8529) := b"0000000000000000_0000000000000000_0010000010010011_1101000100011101"; -- 0.12725550610976996
	pesos_i(8530) := b"0000000000000000_0000000000000000_0000100010110111_0011101011110111"; -- 0.03404587287303505
	pesos_i(8531) := b"0000000000000000_0000000000000000_0000011001011010_0110001000110100"; -- 0.02481664431251159
	pesos_i(8532) := b"1111111111111111_1111111111111111_1111011001011011_1011101110001010"; -- -0.037662771976797446
	pesos_i(8533) := b"0000000000000000_0000000000000000_0001111111110011_0110100110010101"; -- 0.12480792894877363
	pesos_i(8534) := b"1111111111111111_1111111111111111_1110000100000011_1010000000000101"; -- -0.12103843576315673
	pesos_i(8535) := b"0000000000000000_0000000000000000_0000001011010010_0001001100000110"; -- 0.0110179795962576
	pesos_i(8536) := b"1111111111111111_1111111111111111_1111011011000110_0000010000111100"; -- -0.0360410073872256
	pesos_i(8537) := b"1111111111111111_1111111111111111_1111110111011100_1001000011100001"; -- -0.008353180907225342
	pesos_i(8538) := b"0000000000000000_0000000000000000_0010010001010111_0000111010110000"; -- 0.14195339018954445
	pesos_i(8539) := b"0000000000000000_0000000000000000_0000100101111001_1100010100111101"; -- 0.037014319807329214
	pesos_i(8540) := b"1111111111111111_1111111111111111_1111000100000010_1001101110100011"; -- -0.05855395580922774
	pesos_i(8541) := b"1111111111111111_1111111111111111_1110010010011000_1000110001110110"; -- -0.10704729184966313
	pesos_i(8542) := b"1111111111111111_1111111111111111_1101010001110011_1110001001111111"; -- -0.17010673905890866
	pesos_i(8543) := b"1111111111111111_1111111111111111_1110010001001101_1001010110001000"; -- -0.10819116040322418
	pesos_i(8544) := b"1111111111111111_1111111111111111_1110000110001011_1010010011010011"; -- -0.11896295401516828
	pesos_i(8545) := b"0000000000000000_0000000000000000_0001101011000000_0010111111001111"; -- 0.1044950370078953
	pesos_i(8546) := b"0000000000000000_0000000000000000_0010000111001111_0101101111101110"; -- 0.13207029888537417
	pesos_i(8547) := b"1111111111111111_1111111111111111_1110000110100100_0000010101110111"; -- -0.11859098279311604
	pesos_i(8548) := b"1111111111111111_1111111111111111_1101110001011011_1010111111110110"; -- -0.1392259621982327
	pesos_i(8549) := b"0000000000000000_0000000000000000_0001100010111011_0010011000101111"; -- 0.09660566948398398
	pesos_i(8550) := b"0000000000000000_0000000000000000_0001100100101011_1000001110111001"; -- 0.09832022914287436
	pesos_i(8551) := b"0000000000000000_0000000000000000_0000000000100011_1000111101010011"; -- 0.0005426004786201409
	pesos_i(8552) := b"1111111111111111_1111111111111111_1111110100001101_1101011011100110"; -- -0.011507576830156373
	pesos_i(8553) := b"0000000000000000_0000000000000000_0001000011011000_1100011010110101"; -- 0.0658077422623154
	pesos_i(8554) := b"0000000000000000_0000000000000000_0000010001001010_1110010010011110"; -- 0.01676777712592217
	pesos_i(8555) := b"1111111111111111_1111111111111111_1111110111001010_1000011011101010"; -- -0.008628433131515824
	pesos_i(8556) := b"0000000000000000_0000000000000000_0010100010101010_1101110110100111"; -- 0.158857205755418
	pesos_i(8557) := b"1111111111111111_1111111111111111_1101101110000101_1011011010101111"; -- -0.142490942353738
	pesos_i(8558) := b"0000000000000000_0000000000000000_0001000010011101_1010111010001010"; -- 0.06490603318001209
	pesos_i(8559) := b"1111111111111111_1111111111111111_1111011010000111_0110100111001000"; -- -0.03699625842835012
	pesos_i(8560) := b"1111111111111111_1111111111111111_1110000011001111_1101011001111101"; -- -0.12182864612203852
	pesos_i(8561) := b"1111111111111111_1111111111111111_1110100111111011_1001111001110000"; -- -0.08600435022838251
	pesos_i(8562) := b"0000000000000000_0000000000000000_0000101000111011_1010011101010111"; -- 0.039972742724294484
	pesos_i(8563) := b"1111111111111111_1111111111111111_1110001000001110_1111010000110101"; -- -0.116959320984907
	pesos_i(8564) := b"1111111111111111_1111111111111111_1111000010101110_1010101101101011"; -- -0.05983475333447239
	pesos_i(8565) := b"0000000000000000_0000000000000000_0000011111101011_0111000101011011"; -- 0.030936321895256556
	pesos_i(8566) := b"0000000000000000_0000000000000000_0000111011110000_0111000001111011"; -- 0.05835631370958633
	pesos_i(8567) := b"1111111111111111_1111111111111111_1110110100010101_0101111000001011"; -- -0.07389271003795103
	pesos_i(8568) := b"1111111111111111_1111111111111111_1111000011111101_1011101101001010"; -- -0.05862836316459564
	pesos_i(8569) := b"0000000000000000_0000000000000000_0000100000010110_1010000110000100"; -- 0.03159532036428931
	pesos_i(8570) := b"0000000000000000_0000000000000000_0000001100110000_1001010001111111"; -- 0.012460022915312244
	pesos_i(8571) := b"0000000000000000_0000000000000000_0001001110011100_0010011110010101"; -- 0.07660148030040742
	pesos_i(8572) := b"1111111111111111_1111111111111111_1110010100010100_1010001110111000"; -- -0.1051538157365873
	pesos_i(8573) := b"0000000000000000_0000000000000000_0000000100111011_0010110100001011"; -- 0.004809203330623926
	pesos_i(8574) := b"1111111111111111_1111111111111111_1110101000110101_0100001010010100"; -- -0.08512481584028725
	pesos_i(8575) := b"0000000000000000_0000000000000000_0001111100001010_1000111101001000"; -- 0.12125487804366512
	pesos_i(8576) := b"1111111111111111_1111111111111111_1111010001011110_1110111001000100"; -- -0.04542647216908655
	pesos_i(8577) := b"1111111111111111_1111111111111111_1110110011010010_0011000001011000"; -- -0.0749177728641839
	pesos_i(8578) := b"1111111111111111_1111111111111111_1110110000000000_1100010110001111"; -- -0.07811322450856893
	pesos_i(8579) := b"0000000000000000_0000000000000000_0001100111001010_1111000010000110"; -- 0.10075286165268033
	pesos_i(8580) := b"1111111111111111_1111111111111111_1110100101110100_1110010101110001"; -- -0.08806005463028971
	pesos_i(8581) := b"0000000000000000_0000000000000000_0001100000000101_0111001101110110"; -- 0.09383317603926679
	pesos_i(8582) := b"1111111111111111_1111111111111111_1111100011101011_0110101100100000"; -- -0.02765779946027277
	pesos_i(8583) := b"0000000000000000_0000000000000000_0001100110101000_1011110101100100"; -- 0.10023101521623842
	pesos_i(8584) := b"0000000000000000_0000000000000000_0000111001010100_0001000001000100"; -- 0.05597020789778197
	pesos_i(8585) := b"0000000000000000_0000000000000000_0000111010110110_0011101111010001"; -- 0.05746816494080215
	pesos_i(8586) := b"1111111111111111_1111111111111111_1110100010111100_1111010010111110"; -- -0.09086675990486522
	pesos_i(8587) := b"1111111111111111_1111111111111111_1111000010000010_1111100111011010"; -- -0.06050146521719961
	pesos_i(8588) := b"0000000000000000_0000000000000000_0000111000010111_0111110111111001"; -- 0.055045960604206225
	pesos_i(8589) := b"0000000000000000_0000000000000000_0000010110000100_1101011100001010"; -- 0.02155822746318975
	pesos_i(8590) := b"0000000000000000_0000000000000000_0000001011001000_1111101111111001"; -- 0.0108792764669416
	pesos_i(8591) := b"1111111111111111_1111111111111111_1110101111011110_1111101100011001"; -- -0.07862883222559737
	pesos_i(8592) := b"0000000000000000_0000000000000000_0010011001011101_0101011100101100"; -- 0.1498617631235775
	pesos_i(8593) := b"1111111111111111_1111111111111111_1110000001101111_0001110010011011"; -- -0.12330456945300591
	pesos_i(8594) := b"0000000000000000_0000000000000000_0010000110001010_0011000011010001"; -- 0.13101487264152956
	pesos_i(8595) := b"1111111111111111_1111111111111111_1110000110011100_0110100101110111"; -- -0.118707092756761
	pesos_i(8596) := b"0000000000000000_0000000000000000_0001011010101001_1011101010011011"; -- 0.08852735795716582
	pesos_i(8597) := b"0000000000000000_0000000000000000_0001111011110101_1111100011101001"; -- 0.12094073948845797
	pesos_i(8598) := b"1111111111111111_1111111111111111_1110000011011011_1101100000111001"; -- -0.12164543738184606
	pesos_i(8599) := b"0000000000000000_0000000000000000_0010000010000101_0001001111001110"; -- 0.1270305994438396
	pesos_i(8600) := b"1111111111111111_1111111111111111_1101011110111100_0100110110001010"; -- -0.15728297605365352
	pesos_i(8601) := b"1111111111111111_1111111111111111_1110001011100001_0100011100100010"; -- -0.11375003266997803
	pesos_i(8602) := b"0000000000000000_0000000000000000_0001011111011001_0000011000010000"; -- 0.09315526857554554
	pesos_i(8603) := b"1111111111111111_1111111111111111_1111101110100000_1101010110111010"; -- -0.017077104666497252
	pesos_i(8604) := b"1111111111111111_1111111111111111_1110000110010000_1001010011111001"; -- -0.11888760486825868
	pesos_i(8605) := b"0000000000000000_0000000000000000_0000100111000000_0110000110111101"; -- 0.03809176310142139
	pesos_i(8606) := b"1111111111111111_1111111111111111_1111110000010001_0011011110111100"; -- -0.015362278634204614
	pesos_i(8607) := b"1111111111111111_1111111111111111_1110111110011001_1001111010111101"; -- -0.06406219379671423
	pesos_i(8608) := b"0000000000000000_0000000000000000_0000000011110111_1101110100110010"; -- 0.0037821051271546683
	pesos_i(8609) := b"0000000000000000_0000000000000000_0001111100011110_1100100101110010"; -- 0.12156352076102703
	pesos_i(8610) := b"0000000000000000_0000000000000000_0010010000001101_0001110001011100"; -- 0.14082505457228314
	pesos_i(8611) := b"1111111111111111_1111111111111111_1110110000010100_0011100110011110"; -- -0.077816389969856
	pesos_i(8612) := b"1111111111111111_1111111111111111_1101110111111111_0001111000100010"; -- -0.13282596282760542
	pesos_i(8613) := b"1111111111111111_1111111111111111_1110010101000101_0111001010101011"; -- -0.10440905872205662
	pesos_i(8614) := b"1111111111111111_1111111111111111_1111111110101011_1100110111000000"; -- -0.0012847333159550583
	pesos_i(8615) := b"0000000000000000_0000000000000000_0010011100001111_0100100110101101"; -- 0.15257702327743078
	pesos_i(8616) := b"1111111111111111_1111111111111111_1110000110011001_1101011111010011"; -- -0.11874629112928406
	pesos_i(8617) := b"1111111111111111_1111111111111111_1110100111011110_1101110010110101"; -- -0.0864431435502297
	pesos_i(8618) := b"0000000000000000_0000000000000000_0000100011100001_1010011111000100"; -- 0.034693227104878634
	pesos_i(8619) := b"1111111111111111_1111111111111111_1111000111001000_1100010101000001"; -- -0.055530234859762384
	pesos_i(8620) := b"1111111111111111_1111111111111111_1110101111101001_0010111010111000"; -- -0.07847316752049151
	pesos_i(8621) := b"0000000000000000_0000000000000000_0000011000101001_0000101010100011"; -- 0.02406374442147033
	pesos_i(8622) := b"0000000000000000_0000000000000000_0000010100000001_1100111110110110"; -- 0.01955888927895768
	pesos_i(8623) := b"0000000000000000_0000000000000000_0001010011000011_1101111101101101"; -- 0.08111378117867932
	pesos_i(8624) := b"0000000000000000_0000000000000000_0001000010110110_0100000101110101"; -- 0.06528100114874516
	pesos_i(8625) := b"1111111111111111_1111111111111111_1111110010010110_0101101100000101"; -- -0.013330756554318103
	pesos_i(8626) := b"1111111111111111_1111111111111111_1110001100110101_1111101001101111"; -- -0.11245760718513167
	pesos_i(8627) := b"1111111111111111_1111111111111111_1111010110011101_1011010101101111"; -- -0.0405623058201102
	pesos_i(8628) := b"0000000000000000_0000000000000000_0000100000111101_1100001010010100"; -- 0.032192383941202066
	pesos_i(8629) := b"1111111111111111_1111111111111111_1101110000101011_1110001000000100"; -- -0.13995540044605717
	pesos_i(8630) := b"1111111111111111_1111111111111111_1110110001100000_1100111001110100"; -- -0.07664785058175388
	pesos_i(8631) := b"1111111111111111_1111111111111111_1111001110110101_0101011110000101"; -- -0.04801419249913595
	pesos_i(8632) := b"1111111111111111_1111111111111111_1111111011001001_0110100010010110"; -- -0.004739249535725328
	pesos_i(8633) := b"0000000000000000_0000000000000000_0010011111000001_1010000010100100"; -- 0.1552982713289612
	pesos_i(8634) := b"0000000000000000_0000000000000000_0010001001101010_0111000101111111"; -- 0.13443669663757746
	pesos_i(8635) := b"1111111111111111_1111111111111111_1111100101100101_0101000001010100"; -- -0.02579782441479006
	pesos_i(8636) := b"0000000000000000_0000000000000000_0000110000100011_0100110101101011"; -- 0.04741367213134888
	pesos_i(8637) := b"1111111111111111_1111111111111111_1110011110000000_0011011000011111"; -- -0.09569989920959214
	pesos_i(8638) := b"0000000000000000_0000000000000000_0001000100010101_0000101011101011"; -- 0.06672733541873369
	pesos_i(8639) := b"1111111111111111_1111111111111111_1111000111010010_1101010110100101"; -- -0.05537667007092055
	pesos_i(8640) := b"1111111111111111_1111111111111111_1110010001111011_1100110111100010"; -- -0.1074858973726406
	pesos_i(8641) := b"0000000000000000_0000000000000000_0001001110000000_0001011110010111"; -- 0.07617328105067524
	pesos_i(8642) := b"1111111111111111_1111111111111111_1111101000111111_1011101111111001"; -- -0.022464992333845513
	pesos_i(8643) := b"0000000000000000_0000000000000000_0000000000101001_1011010100110111"; -- 0.000636411483809025
	pesos_i(8644) := b"0000000000000000_0000000000000000_0001110100011011_0110101111111010"; -- 0.11369967324055537
	pesos_i(8645) := b"1111111111111111_1111111111111111_1101110110001010_0010111111111001"; -- -0.13461017766430403
	pesos_i(8646) := b"1111111111111111_1111111111111111_1111100001001110_0010111110001001"; -- -0.030056981234988563
	pesos_i(8647) := b"1111111111111111_1111111111111111_1111110110111101_0010010010111010"; -- -0.008832649812772536
	pesos_i(8648) := b"1111111111111111_1111111111111111_1110010011110101_1111111111111110"; -- -0.10562133824615073
	pesos_i(8649) := b"1111111111111111_1111111111111111_1111110000111000_0001101111110011"; -- -0.014768842018508579
	pesos_i(8650) := b"0000000000000000_0000000000000000_0001110000101110_1011111110000100"; -- 0.11008831953806755
	pesos_i(8651) := b"0000000000000000_0000000000000000_0001110001110010_0000010001010011"; -- 0.11111475980643366
	pesos_i(8652) := b"0000000000000000_0000000000000000_0010001001000100_1001011100100001"; -- 0.1338591056256542
	pesos_i(8653) := b"1111111111111111_1111111111111111_1110100001110000_0010010011010100"; -- -0.09203882050101364
	pesos_i(8654) := b"1111111111111111_1111111111111111_1110000010101111_0011100001011110"; -- -0.12232635206746907
	pesos_i(8655) := b"1111111111111111_1111111111111111_1111111001000001_0110000100110011"; -- -0.0068148852647256595
	pesos_i(8656) := b"1111111111111111_1111111111111111_1110101001110010_1101011110011110"; -- -0.08418514632591177
	pesos_i(8657) := b"0000000000000000_0000000000000000_0010010001011001_1111101011001011"; -- 0.14199798060846702
	pesos_i(8658) := b"0000000000000000_0000000000000000_0000010111001100_1001011100111011"; -- 0.022653057038958733
	pesos_i(8659) := b"1111111111111111_1111111111111111_1110011111101100_0010110100011011"; -- -0.09405248738729227
	pesos_i(8660) := b"1111111111111111_1111111111111111_1110111001111110_1010100011100100"; -- -0.06837982598345328
	pesos_i(8661) := b"0000000000000000_0000000000000000_0000011100000011_0111110011011100"; -- 0.027396968630961586
	pesos_i(8662) := b"0000000000000000_0000000000000000_0000101001101101_0011000000101111"; -- 0.040728579878227845
	pesos_i(8663) := b"0000000000000000_0000000000000000_0001010011101110_0010101000110111"; -- 0.08175910792856926
	pesos_i(8664) := b"0000000000000000_0000000000000000_0010001001110110_0010001111001010"; -- 0.13461517018827776
	pesos_i(8665) := b"0000000000000000_0000000000000000_0001111100001110_0010001010000000"; -- 0.12130942943688477
	pesos_i(8666) := b"0000000000000000_0000000000000000_0001111000111111_0010011000000111"; -- 0.11815107024046792
	pesos_i(8667) := b"0000000000000000_0000000000000000_0000001110111011_0001000100001111"; -- 0.014573160274712001
	pesos_i(8668) := b"0000000000000000_0000000000000000_0010000100100000_0011011011011011"; -- 0.12939780079122937
	pesos_i(8669) := b"1111111111111111_1111111111111111_1101111110001000_0010100101110001"; -- -0.1268285845799452
	pesos_i(8670) := b"0000000000000000_0000000000000000_0001011101100011_1100011110011011"; -- 0.09136626744310301
	pesos_i(8671) := b"1111111111111111_1111111111111111_1111100001001111_1100101110010111"; -- -0.030032420751109595
	pesos_i(8672) := b"1111111111111111_1111111111111111_1111000010111001_1000001111100110"; -- -0.059669262339699394
	pesos_i(8673) := b"1111111111111111_1111111111111111_1110111010010111_0110011011011100"; -- -0.06800229205123433
	pesos_i(8674) := b"0000000000000000_0000000000000000_0010010001001011_1100110110100100"; -- 0.14178166633038042
	pesos_i(8675) := b"0000000000000000_0000000000000000_0001011011100001_0101111111011001"; -- 0.08937644056472298
	pesos_i(8676) := b"1111111111111111_1111111111111111_1101101001000111_1011111001111100"; -- -0.14734277223376585
	pesos_i(8677) := b"1111111111111111_1111111111111111_1101101000101110_1100000110100100"; -- -0.14772405391301835
	pesos_i(8678) := b"0000000000000000_0000000000000000_0001100111010110_0101001000000011"; -- 0.1009265190674352
	pesos_i(8679) := b"1111111111111111_1111111111111111_1110100001001110_1101001011110010"; -- -0.09254724101988666
	pesos_i(8680) := b"0000000000000000_0000000000000000_0001100010101000_0111111101001101"; -- 0.09632106438379967
	pesos_i(8681) := b"1111111111111111_1111111111111111_1111100011101001_1110100001111011"; -- -0.02768084531977543
	pesos_i(8682) := b"1111111111111111_1111111111111111_1110111001101100_0010010010011100"; -- -0.06866236879605479
	pesos_i(8683) := b"1111111111111111_1111111111111111_1111001010001011_0001000101111111"; -- -0.05256548547769115
	pesos_i(8684) := b"0000000000000000_0000000000000000_0000010100000000_1111110100001100"; -- 0.019546332747435988
	pesos_i(8685) := b"1111111111111111_1111111111111111_1111010011100001_0110001101001011"; -- -0.043435854228234226
	pesos_i(8686) := b"1111111111111111_1111111111111111_1111001000111000_0101011001111101"; -- -0.0538278526866824
	pesos_i(8687) := b"1111111111111111_1111111111111111_1111111101111001_1010110101010001"; -- -0.002049605978585319
	pesos_i(8688) := b"0000000000000000_0000000000000000_0000010010011101_0000101000011010"; -- 0.018021231868725743
	pesos_i(8689) := b"0000000000000000_0000000000000000_0010011011010100_0100111100000101"; -- 0.15167707317547197
	pesos_i(8690) := b"0000000000000000_0000000000000000_0000100001110111_1001011011110101"; -- 0.03307479369158931
	pesos_i(8691) := b"0000000000000000_0000000000000000_0000100110100001_0101100110100000"; -- 0.03761825714384302
	pesos_i(8692) := b"0000000000000000_0000000000000000_0000011000111010_0101110000011111"; -- 0.024328000597641262
	pesos_i(8693) := b"0000000000000000_0000000000000000_0001001100010010_1000110011110001"; -- 0.07450180907369719
	pesos_i(8694) := b"0000000000000000_0000000000000000_0000110011101101_1101111100100111"; -- 0.050504633903670534
	pesos_i(8695) := b"1111111111111111_1111111111111111_1111110000010101_0101001110100101"; -- -0.015299579791941575
	pesos_i(8696) := b"1111111111111111_1111111111111111_1110000011111001_1111000111010111"; -- -0.12118614664026703
	pesos_i(8697) := b"1111111111111111_1111111111111111_1110101000011010_1010110110110101"; -- -0.08553041772024676
	pesos_i(8698) := b"0000000000000000_0000000000000000_0001001011100000_1001010111010000"; -- 0.07373939830954118
	pesos_i(8699) := b"1111111111111111_1111111111111111_1101111101100111_1111010010001110"; -- -0.12732001810475066
	pesos_i(8700) := b"0000000000000000_0000000000000000_0001110101000110_1010010010111001"; -- 0.11435918340241036
	pesos_i(8701) := b"1111111111111111_1111111111111111_1111110011000010_0011100011110011"; -- -0.012661400582912095
	pesos_i(8702) := b"0000000000000000_0000000000000000_0001000001101111_0110111000010100"; -- 0.06420028683198492
	pesos_i(8703) := b"0000000000000000_0000000000000000_0010011011010001_1111010011011001"; -- 0.15164118102842078
	pesos_i(8704) := b"0000000000000000_0000000000000000_0000010101110000_0111100011111110"; -- 0.021247446183102175
	pesos_i(8705) := b"0000000000000000_0000000000000000_0010001101010010_1111001101000100"; -- 0.13798447035390748
	pesos_i(8706) := b"0000000000000000_0000000000000000_0010010010110011_0011101010010100"; -- 0.14335981471404527
	pesos_i(8707) := b"1111111111111111_1111111111111111_1111110010000011_1111011101101001"; -- -0.013611351839651436
	pesos_i(8708) := b"0000000000000000_0000000000000000_0001000111000110_1000000010000110"; -- 0.0694351508307817
	pesos_i(8709) := b"1111111111111111_1111111111111111_1111000000101000_1110101001000100"; -- -0.06187568511713677
	pesos_i(8710) := b"0000000000000000_0000000000000000_0000000000010110_1000100011001011"; -- 0.00034384681458116194
	pesos_i(8711) := b"0000000000000000_0000000000000000_0010000011101100_0010001010101101"; -- 0.1286031410257542
	pesos_i(8712) := b"1111111111111111_1111111111111111_1110010010110111_1101110000101110"; -- -0.10656951798086789
	pesos_i(8713) := b"0000000000000000_0000000000000000_0000101101001111_0000010011011111"; -- 0.0441744846473045
	pesos_i(8714) := b"0000000000000000_0000000000000000_0000011111011101_1110011000100101"; -- 0.030729660156420476
	pesos_i(8715) := b"1111111111111111_1111111111111111_1111110100010110_0110011010010101"; -- -0.011376942289666403
	pesos_i(8716) := b"1111111111111111_1111111111111111_1110101100101111_0010111010100110"; -- -0.08131130642191595
	pesos_i(8717) := b"0000000000000000_0000000000000000_0000101101011110_0101100010001111"; -- 0.044408354718003924
	pesos_i(8718) := b"0000000000000000_0000000000000000_0010001011100110_0011001000111000"; -- 0.13632501483963394
	pesos_i(8719) := b"0000000000000000_0000000000000000_0000000011011010_1010001101100000"; -- 0.0033361538300446664
	pesos_i(8720) := b"1111111111111111_1111111111111111_1110011111111101_0001101100001010"; -- -0.09379416471984185
	pesos_i(8721) := b"1111111111111111_1111111111111111_1111101100010101_0100000110110111"; -- -0.01920689847947472
	pesos_i(8722) := b"1111111111111111_1111111111111111_1110001000000111_0001010001011011"; -- -0.11707947526084918
	pesos_i(8723) := b"1111111111111111_1111111111111111_1111110010001111_1011101000111101"; -- -0.013431892604854521
	pesos_i(8724) := b"0000000000000000_0000000000000000_0000000111100100_0101111101011010"; -- 0.007390937202912048
	pesos_i(8725) := b"0000000000000000_0000000000000000_0001110100111011_0011010000111011"; -- 0.11418463178422476
	pesos_i(8726) := b"0000000000000000_0000000000000000_0001010001110011_0101011100110100"; -- 0.07988495839445044
	pesos_i(8727) := b"1111111111111111_1111111111111111_1111010110100100_0100000100010011"; -- -0.04046242993472859
	pesos_i(8728) := b"1111111111111111_1111111111111111_1110010101101101_0011101001000011"; -- -0.10380206924508983
	pesos_i(8729) := b"0000000000000000_0000000000000000_0000000110110010_0001001011110010"; -- 0.006623443583891392
	pesos_i(8730) := b"0000000000000000_0000000000000000_0001001111111111_1111011000001101"; -- 0.07812440689081078
	pesos_i(8731) := b"1111111111111111_1111111111111111_1111000010010100_0000000011101001"; -- -0.060241644870162224
	pesos_i(8732) := b"1111111111111111_1111111111111111_1101100101001101_0111001110110000"; -- -0.15116192777032403
	pesos_i(8733) := b"1111111111111111_1111111111111111_1110001110100110_0011110111011101"; -- -0.11074460359122752
	pesos_i(8734) := b"0000000000000000_0000000000000000_0001001101101010_1000111111100111"; -- 0.07584475889087533
	pesos_i(8735) := b"1111111111111111_1111111111111111_1110001100011101_1010100001110000"; -- -0.11282870544169564
	pesos_i(8736) := b"0000000000000000_0000000000000000_0000100000111100_1110011001001000"; -- 0.03217925325647903
	pesos_i(8737) := b"1111111111111111_1111111111111111_1111001000110111_0011111111111011"; -- -0.053844452992034456
	pesos_i(8738) := b"0000000000000000_0000000000000000_0000011011000011_0011110010111011"; -- 0.02641658380049115
	pesos_i(8739) := b"0000000000000000_0000000000000000_0000000101101011_1000001110110110"; -- 0.005546790904833037
	pesos_i(8740) := b"1111111111111111_1111111111111111_1111111001100011_1100000000011111"; -- -0.006290428515240666
	pesos_i(8741) := b"1111111111111111_1111111111111111_1101100010010110_0011010001101110"; -- -0.15395805665553955
	pesos_i(8742) := b"1111111111111111_1111111111111111_1111011001000001_1110000110001001"; -- -0.0380572357556282
	pesos_i(8743) := b"0000000000000000_0000000000000000_0000000101010100_0001000111101011"; -- 0.005189056310197529
	pesos_i(8744) := b"1111111111111111_1111111111111111_1110111111001111_0100010111010111"; -- -0.06324351798928371
	pesos_i(8745) := b"0000000000000000_0000000000000000_0000110101100111_0110001010100101"; -- 0.05235878497803681
	pesos_i(8746) := b"1111111111111111_1111111111111111_1101101001000101_0101001001011110"; -- -0.1473797340517625
	pesos_i(8747) := b"0000000000000000_0000000000000000_0001001010110000_1101101110111010"; -- 0.0730111436140665
	pesos_i(8748) := b"0000000000000000_0000000000000000_0001010000001110_0011101011110111"; -- 0.07834213764822354
	pesos_i(8749) := b"0000000000000000_0000000000000000_0000000011000111_0100001100100101"; -- 0.003040501222570373
	pesos_i(8750) := b"0000000000000000_0000000000000000_0001100000101010_0111101110000101"; -- 0.09439823159130377
	pesos_i(8751) := b"1111111111111111_1111111111111111_1111011111010011_1001010001110110"; -- -0.03192779657427238
	pesos_i(8752) := b"1111111111111111_1111111111111111_1110000100111111_1110001101101101"; -- -0.12011889071409954
	pesos_i(8753) := b"0000000000000000_0000000000000000_0000001011100000_1110000001011000"; -- 0.01124384073084029
	pesos_i(8754) := b"1111111111111111_1111111111111111_1111011101000001_1011010010110010"; -- -0.03415365835346992
	pesos_i(8755) := b"0000000000000000_0000000000000000_0001000001000011_0011110101001100"; -- 0.06352599245306711
	pesos_i(8756) := b"1111111111111111_1111111111111111_1111111111100001_0001011100110010"; -- -0.0004716398742532906
	pesos_i(8757) := b"1111111111111111_1111111111111111_1101110111101110_0101001010100000"; -- -0.13308223344169254
	pesos_i(8758) := b"1111111111111111_1111111111111111_1110111110000100_1010110110110110"; -- -0.06438173588029694
	pesos_i(8759) := b"1111111111111111_1111111111111111_1111100011110000_1111001010101000"; -- -0.02757342724749303
	pesos_i(8760) := b"1111111111111111_1111111111111111_1101101100110011_0000110101111011"; -- -0.14375224822018043
	pesos_i(8761) := b"1111111111111111_1111111111111111_1111110100011110_1001111010000010"; -- -0.011251538413954433
	pesos_i(8762) := b"0000000000000000_0000000000000000_0000000111010000_1010111001001101"; -- 0.007090467263423981
	pesos_i(8763) := b"0000000000000000_0000000000000000_0001100010010011_1101000011111110"; -- 0.09600549881069018
	pesos_i(8764) := b"1111111111111111_1111111111111111_1111101100011110_0011001101011110"; -- -0.019070424686328052
	pesos_i(8765) := b"0000000000000000_0000000000000000_0000011011111101_1000001000001100"; -- 0.027305725048157228
	pesos_i(8766) := b"1111111111111111_1111111111111111_1111100000000010_0101011011101010"; -- -0.031214301911024932
	pesos_i(8767) := b"1111111111111111_1111111111111111_1110000001101000_0101101011110000"; -- -0.12340766557833424
	pesos_i(8768) := b"0000000000000000_0000000000000000_0001010100001101_1100110010111011"; -- 0.08224181706762543
	pesos_i(8769) := b"1111111111111111_1111111111111111_1101110100110001_1111000110000011"; -- -0.13595667416188154
	pesos_i(8770) := b"1111111111111111_1111111111111111_1101111001110001_1111000101010111"; -- -0.13107387189535188
	pesos_i(8771) := b"1111111111111111_1111111111111111_1110001000111101_0101001100101110"; -- -0.11625175587621893
	pesos_i(8772) := b"1111111111111111_1111111111111111_1111011001100100_1001101101100100"; -- -0.03752735915303356
	pesos_i(8773) := b"1111111111111111_1111111111111111_1111010001110010_1100100111001101"; -- -0.04512346983352031
	pesos_i(8774) := b"1111111111111111_1111111111111111_1111011110011100_1001100111110101"; -- -0.032766702333924196
	pesos_i(8775) := b"1111111111111111_1111111111111111_1110011110111001_1010001100100010"; -- -0.09482365049385824
	pesos_i(8776) := b"0000000000000000_0000000000000000_0010000000100000_0100101100010111"; -- 0.12549275699980836
	pesos_i(8777) := b"0000000000000000_0000000000000000_0000011101111110_0001110011101000"; -- 0.029268080311657167
	pesos_i(8778) := b"1111111111111111_1111111111111111_1111111110101110_0110110000001110"; -- -0.0012447801632184136
	pesos_i(8779) := b"1111111111111111_1111111111111111_1111001010010010_0001010010010100"; -- -0.05245849027937238
	pesos_i(8780) := b"1111111111111111_1111111111111111_1111010101111100_0111001011110110"; -- -0.0410698078532639
	pesos_i(8781) := b"1111111111111111_1111111111111111_1111101000100011_1101001100101111"; -- -0.022890854857710075
	pesos_i(8782) := b"1111111111111111_1111111111111111_1111111110111010_1100011111111101"; -- -0.0010561950226997106
	pesos_i(8783) := b"1111111111111111_1111111111111111_1110110010101011_1000100111011000"; -- -0.07550753090750638
	pesos_i(8784) := b"1111111111111111_1111111111111111_1111000000111110_0101001110010110"; -- -0.0615489728759976
	pesos_i(8785) := b"1111111111111111_1111111111111111_1110101110111100_1011100010001110"; -- -0.07915159742158254
	pesos_i(8786) := b"0000000000000000_0000000000000000_0000001101001101_0100100011111110"; -- 0.01289802750034911
	pesos_i(8787) := b"0000000000000000_0000000000000000_0000110010000111_0100101000100010"; -- 0.04893935513323072
	pesos_i(8788) := b"0000000000000000_0000000000000000_0001100110001000_0000011010110010"; -- 0.09973184434855259
	pesos_i(8789) := b"1111111111111111_1111111111111111_1111011010000000_1000001100001000"; -- -0.037101564970330396
	pesos_i(8790) := b"1111111111111111_1111111111111111_1111010011010001_0010001000100100"; -- -0.043683878199780944
	pesos_i(8791) := b"0000000000000000_0000000000000000_0001111000001100_1110110010110101"; -- 0.11738471440499311
	pesos_i(8792) := b"0000000000000000_0000000000000000_0000111100111111_0010100100110001"; -- 0.05955750879639414
	pesos_i(8793) := b"1111111111111111_1111111111111111_1111110101010011_0001011110100100"; -- -0.010450861497107998
	pesos_i(8794) := b"1111111111111111_1111111111111111_1111010111011010_1011111000011100"; -- -0.0396310025214733
	pesos_i(8795) := b"0000000000000000_0000000000000000_0001010100001101_0001001101111111"; -- 0.08223077632128545
	pesos_i(8796) := b"0000000000000000_0000000000000000_0001111110111111_1011100111010100"; -- 0.12401925502660321
	pesos_i(8797) := b"1111111111111111_1111111111111111_1110000011101100_1000000111001110"; -- -0.12139118888479015
	pesos_i(8798) := b"1111111111111111_1111111111111111_1110000111011011_1010101010111110"; -- -0.11774189812299941
	pesos_i(8799) := b"0000000000000000_0000000000000000_0001100111001111_1000111111100000"; -- 0.10082339499887877
	pesos_i(8800) := b"1111111111111111_1111111111111111_1111101110100011_0000010000110010"; -- -0.01704381736959022
	pesos_i(8801) := b"0000000000000000_0000000000000000_0001101111101111_0000011101000010"; -- 0.10911603323605538
	pesos_i(8802) := b"1111111111111111_1111111111111111_1111110001111011_0000111101010001"; -- -0.013747256036506703
	pesos_i(8803) := b"0000000000000000_0000000000000000_0000111001100100_0110000111001100"; -- 0.056219208072581496
	pesos_i(8804) := b"1111111111111111_1111111111111111_1101101010010111_1111010100100001"; -- -0.14611881203401547
	pesos_i(8805) := b"1111111111111111_1111111111111111_1111000110001111_1100011000010011"; -- -0.05639993711322809
	pesos_i(8806) := b"0000000000000000_0000000000000000_0000011110000100_0111001111111111"; -- 0.029364824105575626
	pesos_i(8807) := b"1111111111111111_1111111111111111_1111100100111100_0011000001111100"; -- -0.026425332708704622
	pesos_i(8808) := b"1111111111111111_1111111111111111_1111111110101110_0010001111010110"; -- -0.0012490846736289557
	pesos_i(8809) := b"1111111111111111_1111111111111111_1110000001011110_0001100001010100"; -- -0.12356422374944784
	pesos_i(8810) := b"1111111111111111_1111111111111111_1110100100001010_0010001110111011"; -- -0.08968903243741311
	pesos_i(8811) := b"0000000000000000_0000000000000000_0000011010100100_0001001101001101"; -- 0.025941091774390027
	pesos_i(8812) := b"1111111111111111_1111111111111111_1111111011101101_0100100111111011"; -- -0.004191757397885075
	pesos_i(8813) := b"0000000000000000_0000000000000000_0001001111111111_0111100011110111"; -- 0.07811695134687156
	pesos_i(8814) := b"1111111111111111_1111111111111111_1111101011011101_0110011001111011"; -- -0.020059199281486185
	pesos_i(8815) := b"0000000000000000_0000000000000000_0000110000111101_1001010000000101"; -- 0.047814608883434306
	pesos_i(8816) := b"0000000000000000_0000000000000000_0000110010000101_1000001000011110"; -- 0.04891217455526898
	pesos_i(8817) := b"1111111111111111_1111111111111111_1111000101101011_0101110010111000"; -- -0.0569555330307969
	pesos_i(8818) := b"0000000000000000_0000000000000000_0001100110011101_0110110110001000"; -- 0.10005840833832826
	pesos_i(8819) := b"0000000000000000_0000000000000000_0000000111010110_1110101011110010"; -- 0.00718563474165499
	pesos_i(8820) := b"1111111111111111_1111111111111111_1111111010111101_0011001110101100"; -- -0.0049255089764430535
	pesos_i(8821) := b"1111111111111111_1111111111111111_1110100101000001_1100010101100110"; -- -0.08884016276331604
	pesos_i(8822) := b"0000000000000000_0000000000000000_0000010001101000_1111110001111000"; -- 0.017226962359352824
	pesos_i(8823) := b"1111111111111111_1111111111111111_1111001000101011_0111111100000001"; -- -0.054023801981622724
	pesos_i(8824) := b"0000000000000000_0000000000000000_0000100101000000_1010010100111000"; -- 0.036142660255244964
	pesos_i(8825) := b"1111111111111111_1111111111111111_1111110001010000_1101110010010010"; -- -0.014391149891507915
	pesos_i(8826) := b"0000000000000000_0000000000000000_0001011010110111_1000011110010010"; -- 0.08873793901581914
	pesos_i(8827) := b"1111111111111111_1111111111111111_1111011011000111_0010001001100101"; -- -0.03602395097650525
	pesos_i(8828) := b"0000000000000000_0000000000000000_0000111000100010_0100000111000100"; -- 0.055210218810617134
	pesos_i(8829) := b"1111111111111111_1111111111111111_1111111110111011_1010110001010100"; -- -0.0010425848554265558
	pesos_i(8830) := b"0000000000000000_0000000000000000_0001111000100010_0011111010011011"; -- 0.1177100303139077
	pesos_i(8831) := b"1111111111111111_1111111111111111_1111100110011001_1001001101010001"; -- -0.025000374540296723
	pesos_i(8832) := b"0000000000000000_0000000000000000_0010010100010110_1011000010010010"; -- 0.14487746773195845
	pesos_i(8833) := b"1111111111111111_1111111111111111_1111000011111011_0000000110101100"; -- -0.058669944316196584
	pesos_i(8834) := b"1111111111111111_1111111111111111_1111001101101100_1010111110010011"; -- -0.049122835638383926
	pesos_i(8835) := b"0000000000000000_0000000000000000_0001100001001000_1011011111010001"; -- 0.09485958920043719
	pesos_i(8836) := b"1111111111111111_1111111111111111_1111110001100100_1101100000001111"; -- -0.014086242929007663
	pesos_i(8837) := b"0000000000000000_0000000000000000_0001111101010100_0110111100101011"; -- 0.12238211449080667
	pesos_i(8838) := b"0000000000000000_0000000000000000_0001001101011101_1000101101010011"; -- 0.0756461217268995
	pesos_i(8839) := b"1111111111111111_1111111111111111_1111011000000000_0000000100110111"; -- -0.03906242759313222
	pesos_i(8840) := b"1111111111111111_1111111111111111_1111110011111100_0100010100101110"; -- -0.01177566169745441
	pesos_i(8841) := b"0000000000000000_0000000000000000_0001010110010011_0010110100001010"; -- 0.08427697643898857
	pesos_i(8842) := b"1111111111111111_1111111111111111_1110011110111100_0101101001100101"; -- -0.0947822096930838
	pesos_i(8843) := b"1111111111111111_1111111111111111_1110101000111010_1001101001100000"; -- -0.0850432887460505
	pesos_i(8844) := b"1111111111111111_1111111111111111_1110001111010111_0001001100011100"; -- -0.10999947126927781
	pesos_i(8845) := b"0000000000000000_0000000000000000_0000000100001110_1001010101010000"; -- 0.004128772811777084
	pesos_i(8846) := b"1111111111111111_1111111111111111_1111011011110101_1000011010010111"; -- -0.03531607457547517
	pesos_i(8847) := b"0000000000000000_0000000000000000_0001101001010011_1110011000101010"; -- 0.10284269828955725
	pesos_i(8848) := b"0000000000000000_0000000000000000_0001001011101101_0111100011001110"; -- 0.07393603356654999
	pesos_i(8849) := b"1111111111111111_1111111111111111_1111011001011100_1111011000000100"; -- -0.0376440276320219
	pesos_i(8850) := b"1111111111111111_1111111111111111_1110101011011101_1011101110000000"; -- -0.08255413166309382
	pesos_i(8851) := b"1111111111111111_1111111111111111_1110110100010011_0100111100101110"; -- -0.07392411361883344
	pesos_i(8852) := b"1111111111111111_1111111111111111_1101111110100111_1010100110101101"; -- -0.12634791879411827
	pesos_i(8853) := b"1111111111111111_1111111111111111_1110011101110001_1100011101011001"; -- -0.09592012467469456
	pesos_i(8854) := b"0000000000000000_0000000000000000_0000011101000110_1110100000110101"; -- 0.028425705913149135
	pesos_i(8855) := b"0000000000000000_0000000000000000_0001101101110110_0111001111001110"; -- 0.10727618956369186
	pesos_i(8856) := b"1111111111111111_1111111111111111_1110100000001110_0011000101101001"; -- -0.09353343181631266
	pesos_i(8857) := b"1111111111111111_1111111111111111_1101110111011010_0110011111011101"; -- -0.13338614324506645
	pesos_i(8858) := b"0000000000000000_0000000000000000_0000011001101001_1011100110000111"; -- 0.02505073110354792
	pesos_i(8859) := b"0000000000000000_0000000000000000_0001011110011000_0000011100111101"; -- 0.0921635172709925
	pesos_i(8860) := b"0000000000000000_0000000000000000_0000111000101001_0011110111000011"; -- 0.05531679156016444
	pesos_i(8861) := b"1111111111111111_1111111111111111_1111000011100110_0111001011001001"; -- -0.0589836367181716
	pesos_i(8862) := b"1111111111111111_1111111111111111_1111100101000010_1101110010010010"; -- -0.02632352293518954
	pesos_i(8863) := b"1111111111111111_1111111111111111_1101100111110011_1110110011010101"; -- -0.1486217480224453
	pesos_i(8864) := b"1111111111111111_1111111111111111_1110101100111101_0000110111000001"; -- -0.08109964413211307
	pesos_i(8865) := b"1111111111111111_1111111111111111_1110000011011001_0010101010110100"; -- -0.12168629740502811
	pesos_i(8866) := b"0000000000000000_0000000000000000_0010000000111011_1000010111110011"; -- 0.1259082526564797
	pesos_i(8867) := b"0000000000000000_0000000000000000_0001100111010010_1110010011000011"; -- 0.10087423094715639
	pesos_i(8868) := b"0000000000000000_0000000000000000_0010001110111100_0010000011010100"; -- 0.1395893591048113
	pesos_i(8869) := b"1111111111111111_1111111111111111_1111001000001110_1010101100100101"; -- -0.054463675875931636
	pesos_i(8870) := b"1111111111111111_1111111111111111_1111011101110000_0100111110110101"; -- -0.03344251468420695
	pesos_i(8871) := b"0000000000000000_0000000000000000_0000001000000001_0001001001000001"; -- 0.007828846819916056
	pesos_i(8872) := b"1111111111111111_1111111111111111_1101111001010011_1001100100101000"; -- -0.13153689169467334
	pesos_i(8873) := b"0000000000000000_0000000000000000_0010001110010110_0001101010011100"; -- 0.13900915428868393
	pesos_i(8874) := b"0000000000000000_0000000000000000_0000001101101011_0110100001101111"; -- 0.013357665058863504
	pesos_i(8875) := b"0000000000000000_0000000000000000_0010100001001101_0000001100110101"; -- 0.15742511780713206
	pesos_i(8876) := b"1111111111111111_1111111111111111_1101111100010001_1100010010100100"; -- -0.1286351299834845
	pesos_i(8877) := b"1111111111111111_1111111111111111_1111001001010000_0100001001011011"; -- -0.05346284171755712
	pesos_i(8878) := b"1111111111111111_1111111111111111_1110000000001010_1001100100101011"; -- -0.1248382825888438
	pesos_i(8879) := b"0000000000000000_0000000000000000_0000011100000100_0010000000110010"; -- 0.02740670424839801
	pesos_i(8880) := b"0000000000000000_0000000000000000_0000111100101011_0000001000100010"; -- 0.059250005075148805
	pesos_i(8881) := b"1111111111111111_1111111111111111_1101111100110100_1100000111011011"; -- -0.12810123824044137
	pesos_i(8882) := b"1111111111111111_1111111111111111_1111101010100101_1110100110111101"; -- -0.02090586789551332
	pesos_i(8883) := b"1111111111111111_1111111111111111_1111100011111001_1111100000100110"; -- -0.027435770827418236
	pesos_i(8884) := b"1111111111111111_1111111111111111_1111111000110111_0001101000000100"; -- -0.006971715896201082
	pesos_i(8885) := b"1111111111111111_1111111111111111_1111010011001101_1100100101110000"; -- -0.043734941520567235
	pesos_i(8886) := b"1111111111111111_1111111111111111_1111000101101001_0110100111110011"; -- -0.05698526198661924
	pesos_i(8887) := b"0000000000000000_0000000000000000_0001111111101001_0101100001101011"; -- 0.12465431795684405
	pesos_i(8888) := b"1111111111111111_1111111111111111_1111100010011111_1100100100111011"; -- -0.02881185825978955
	pesos_i(8889) := b"0000000000000000_0000000000000000_0001111011001011_1001100101000101"; -- 0.12029416973798096
	pesos_i(8890) := b"1111111111111111_1111111111111111_1101111000100111_0010111110001000"; -- -0.1322145740482656
	pesos_i(8891) := b"0000000000000000_0000000000000000_0001011101000001_0111110000000101"; -- 0.09084296352759309
	pesos_i(8892) := b"1111111111111111_1111111111111111_1111100011101010_1110011100001100"; -- -0.027665671934646755
	pesos_i(8893) := b"1111111111111111_1111111111111111_1111001011001100_1001001011110011"; -- -0.051565948092155346
	pesos_i(8894) := b"1111111111111111_1111111111111111_1110101101100101_0101110000110010"; -- -0.08048461705103828
	pesos_i(8895) := b"0000000000000000_0000000000000000_0000111000001011_1111110110101000"; -- 0.05487046576127964
	pesos_i(8896) := b"1111111111111111_1111111111111111_1111010000101100_1100001101011011"; -- -0.046191969226732785
	pesos_i(8897) := b"0000000000000000_0000000000000000_0001111111111110_1111101111011000"; -- 0.12498449350680635
	pesos_i(8898) := b"0000000000000000_0000000000000000_0001100000001010_0111001101100010"; -- 0.09390946528809137
	pesos_i(8899) := b"0000000000000000_0000000000000000_0001010111000011_1010110110011000"; -- 0.0850170607759648
	pesos_i(8900) := b"1111111111111111_1111111111111111_1101111010100110_0010101000100100"; -- -0.13027702918145626
	pesos_i(8901) := b"0000000000000000_0000000000000000_0010010100100000_1100010011101010"; -- 0.1450312682864548
	pesos_i(8902) := b"1111111111111111_1111111111111111_1111111011000111_1011000111100010"; -- -0.004765398223914177
	pesos_i(8903) := b"1111111111111111_1111111111111111_1111110101000110_1001011111000111"; -- -0.010641588059608508
	pesos_i(8904) := b"0000000000000000_0000000000000000_0010001100011011_1011010110101001"; -- 0.1371415650818473
	pesos_i(8905) := b"0000000000000000_0000000000000000_0000000110100110_1000000001001111"; -- 0.0064468568605321784
	pesos_i(8906) := b"0000000000000000_0000000000000000_0000010011111001_0100100011011000"; -- 0.019428780230250492
	pesos_i(8907) := b"0000000000000000_0000000000000000_0001100110110001_0000001001011101"; -- 0.10035719648679552
	pesos_i(8908) := b"0000000000000000_0000000000000000_0001101110011010_0000101010110000"; -- 0.10781924044292027
	pesos_i(8909) := b"1111111111111111_1111111111111111_1110110100100001_0010010111110101"; -- -0.07371294745550215
	pesos_i(8910) := b"1111111111111111_1111111111111111_1110000001101111_1100000000101001"; -- -0.12329482078854292
	pesos_i(8911) := b"0000000000000000_0000000000000000_0000101000110011_1111001111111011"; -- 0.03985524060155527
	pesos_i(8912) := b"0000000000000000_0000000000000000_0001111000100000_1001111100010000"; -- 0.1176852621236036
	pesos_i(8913) := b"1111111111111111_1111111111111111_1111101111101001_1111110101011011"; -- -0.015960850907358725
	pesos_i(8914) := b"0000000000000000_0000000000000000_0000100010101110_1101000011111100"; -- 0.03391748581990466
	pesos_i(8915) := b"0000000000000000_0000000000000000_0000100011110100_0011011110100001"; -- 0.03497646037290743
	pesos_i(8916) := b"1111111111111111_1111111111111111_1110010001001001_1100100111101010"; -- -0.1082490733258111
	pesos_i(8917) := b"0000000000000000_0000000000000000_0001111100111001_1110000111010011"; -- 0.121976961233479
	pesos_i(8918) := b"1111111111111111_1111111111111111_1110111011101111_1001110110001011"; -- -0.0666562590696291
	pesos_i(8919) := b"0000000000000000_0000000000000000_0010011011001000_0100011100011100"; -- 0.1514934962668477
	pesos_i(8920) := b"0000000000000000_0000000000000000_0000011100011010_1010010010001000"; -- 0.02775028540684628
	pesos_i(8921) := b"0000000000000000_0000000000000000_0000010001010100_1111111011010111"; -- 0.01692192801955464
	pesos_i(8922) := b"1111111111111111_1111111111111111_1111011010101011_1101100010111000"; -- -0.036440329658734616
	pesos_i(8923) := b"0000000000000000_0000000000000000_0001100010000010_0010011000111001"; -- 0.09573592091649995
	pesos_i(8924) := b"0000000000000000_0000000000000000_0010010110011111_1110001101001000"; -- 0.14697094442671013
	pesos_i(8925) := b"1111111111111111_1111111111111111_1111001000001011_0011001100110100"; -- -0.05451660134481592
	pesos_i(8926) := b"0000000000000000_0000000000000000_0010000001011100_1001010101010011"; -- 0.12641270906496094
	pesos_i(8927) := b"0000000000000000_0000000000000000_0000011011001010_1100000101110111"; -- 0.026531306728273144
	pesos_i(8928) := b"0000000000000000_0000000000000000_0000111111110010_1110010110001100"; -- 0.06230005891056956
	pesos_i(8929) := b"1111111111111111_1111111111111111_1111001101101000_0111011101101011"; -- -0.04918721812844095
	pesos_i(8930) := b"0000000000000000_0000000000000000_0000101111010000_0101110000101011"; -- 0.04614807172598676
	pesos_i(8931) := b"1111111111111111_1111111111111111_1111101000001010_0111100000010111"; -- -0.023277754183574122
	pesos_i(8932) := b"0000000000000000_0000000000000000_0000001000101111_0110010000000011"; -- 0.008535624351703281
	pesos_i(8933) := b"0000000000000000_0000000000000000_0000001011011110_1000010111100001"; -- 0.011207930948153706
	pesos_i(8934) := b"1111111111111111_1111111111111111_1101101000001110_1000101001100111"; -- -0.14821562759253595
	pesos_i(8935) := b"1111111111111111_1111111111111111_1101111110010111_1111110101110101"; -- -0.12658706565708994
	pesos_i(8936) := b"1111111111111111_1111111111111111_1101100011100000_1000100100111111"; -- -0.1528238508090677
	pesos_i(8937) := b"0000000000000000_0000000000000000_0000001111101000_1111010100110000"; -- 0.015273403349580562
	pesos_i(8938) := b"0000000000000000_0000000000000000_0001110001110100_1101011111101111"; -- 0.11115789010242556
	pesos_i(8939) := b"1111111111111111_1111111111111111_1110100100000101_0111000011000011"; -- -0.08976073490483394
	pesos_i(8940) := b"1111111111111111_1111111111111111_1110011101000111_1000000011100111"; -- -0.09656519285900614
	pesos_i(8941) := b"0000000000000000_0000000000000000_0001110011110000_1100110110001001"; -- 0.11304936014719846
	pesos_i(8942) := b"1111111111111111_1111111111111111_1110100100101100_0101111110010110"; -- -0.08916666589760767
	pesos_i(8943) := b"0000000000000000_0000000000000000_0001000101011001_0111101101011000"; -- 0.06777163419797058
	pesos_i(8944) := b"1111111111111111_1111111111111111_1111001011101101_0011111111001000"; -- -0.05106736538813782
	pesos_i(8945) := b"0000000000000000_0000000000000000_0001011001101010_0000001000010010"; -- 0.08755505511638671
	pesos_i(8946) := b"0000000000000000_0000000000000000_0001000010111101_0100000000110101"; -- 0.06538773818502615
	pesos_i(8947) := b"1111111111111111_1111111111111111_1111111000001000_1101011110011111"; -- -0.007677577643186927
	pesos_i(8948) := b"0000000000000000_0000000000000000_0010000101101111_1111111101000000"; -- 0.1306151896392078
	pesos_i(8949) := b"1111111111111111_1111111111111111_1110011100101000_1100011011101010"; -- -0.09703404222743425
	pesos_i(8950) := b"0000000000000000_0000000000000000_0010010110011000_1011001100000100"; -- 0.1468612560256799
	pesos_i(8951) := b"1111111111111111_1111111111111111_1111001111010001_0011000001011111"; -- -0.047589280017665374
	pesos_i(8952) := b"1111111111111111_1111111111111111_1111011111001000_0001101110011010"; -- -0.03210284701755238
	pesos_i(8953) := b"0000000000000000_0000000000000000_0001010000100110_1110100001000110"; -- 0.07871867845676134
	pesos_i(8954) := b"0000000000000000_0000000000000000_0001011011011010_0100100110101110"; -- 0.08926830768395246
	pesos_i(8955) := b"0000000000000000_0000000000000000_0000001111101000_1100111011001111"; -- 0.015271115800082192
	pesos_i(8956) := b"0000000000000000_0000000000000000_0000101000010010_0110101110101111"; -- 0.03934357657107616
	pesos_i(8957) := b"1111111111111111_1111111111111111_1111110111110101_1011011111011010"; -- -0.007969388303854486
	pesos_i(8958) := b"1111111111111111_1111111111111111_1111010100100110_0000100000101111"; -- -0.04238842813414738
	pesos_i(8959) := b"0000000000000000_0000000000000000_0010000011001101_0110100100011011"; -- 0.1281343165591406
	pesos_i(8960) := b"0000000000000000_0000000000000000_0010000111111001_0101100111011010"; -- 0.13271104403738349
	pesos_i(8961) := b"1111111111111111_1111111111111111_1111001111000110_1110001100111000"; -- -0.047746466392254244
	pesos_i(8962) := b"0000000000000000_0000000000000000_0001111110011011_1111100100010001"; -- 0.1234737079071877
	pesos_i(8963) := b"1111111111111111_1111111111111111_1111000111001100_0100010001001011"; -- -0.05547688643578816
	pesos_i(8964) := b"1111111111111111_1111111111111111_1111001100001011_0000111110001010"; -- -0.05061247710522235
	pesos_i(8965) := b"0000000000000000_0000000000000000_0000010000111110_1011010001101111"; -- 0.01658179966007154
	pesos_i(8966) := b"0000000000000000_0000000000000000_0001011111100101_1100100101111101"; -- 0.09335002224854325
	pesos_i(8967) := b"1111111111111111_1111111111111111_1110101000001101_1101000111010110"; -- -0.08572662858289531
	pesos_i(8968) := b"1111111111111111_1111111111111111_1111101010110110_1010110000000001"; -- -0.020650148062501514
	pesos_i(8969) := b"1111111111111111_1111111111111111_1111101010101111_0110011000110011"; -- -0.020761120406240858
	pesos_i(8970) := b"1111111111111111_1111111111111111_1110010111010111_1001011100001010"; -- -0.10217910776444239
	pesos_i(8971) := b"0000000000000000_0000000000000000_0001001100110001_1101001010011100"; -- 0.07497898396485443
	pesos_i(8972) := b"1111111111111111_1111111111111111_1111011000101010_1001101000111011"; -- -0.03841243792612278
	pesos_i(8973) := b"1111111111111111_1111111111111111_1111010100000101_1111100010000010"; -- -0.04287764393201009
	pesos_i(8974) := b"0000000000000000_0000000000000000_0000000011111001_1111010011100110"; -- 0.0038140355165745808
	pesos_i(8975) := b"0000000000000000_0000000000000000_0000000110001000_1111111010101100"; -- 0.005996624851458347
	pesos_i(8976) := b"0000000000000000_0000000000000000_0000101100101110_0000101110001101"; -- 0.04367134284415252
	pesos_i(8977) := b"1111111111111111_1111111111111111_1111101000001101_0000001111000111"; -- -0.023238910620436336
	pesos_i(8978) := b"1111111111111111_1111111111111111_1111000110101011_1100010000111001"; -- -0.055972801329356905
	pesos_i(8979) := b"0000000000000000_0000000000000000_0001000011000100_1100000001000000"; -- 0.0655021815339476
	pesos_i(8980) := b"1111111111111111_1111111111111111_1111000010000011_0011100000101101"; -- -0.06049775021889131
	pesos_i(8981) := b"1111111111111111_1111111111111111_1110001011011010_0111100010000001"; -- -0.11385390145150184
	pesos_i(8982) := b"1111111111111111_1111111111111111_1110100001100001_0111011001001010"; -- -0.09226284677282892
	pesos_i(8983) := b"1111111111111111_1111111111111111_1111001111010110_0100011001110101"; -- -0.04751166967418243
	pesos_i(8984) := b"1111111111111111_1111111111111111_1101110001101101_1010000001001101"; -- -0.13895223729651476
	pesos_i(8985) := b"0000000000000000_0000000000000000_0000010100100001_1100000101100011"; -- 0.020046316682773686
	pesos_i(8986) := b"0000000000000000_0000000000000000_0000100010110001_1001000000111110"; -- 0.033959403136967305
	pesos_i(8987) := b"0000000000000000_0000000000000000_0010000100011111_1110111010000110"; -- 0.12939348953735585
	pesos_i(8988) := b"0000000000000000_0000000000000000_0000100011101111_1101101011110111"; -- 0.034909901909770315
	pesos_i(8989) := b"1111111111111111_1111111111111111_1111111011111110_0000110000001000"; -- -0.003936050454608878
	pesos_i(8990) := b"0000000000000000_0000000000000000_0010001101011001_0110101111100101"; -- 0.13808321335042953
	pesos_i(8991) := b"1111111111111111_1111111111111111_1111011111000101_0111010001011001"; -- -0.032143333779727216
	pesos_i(8992) := b"0000000000000000_0000000000000000_0010000101111110_1100101011000010"; -- 0.13084094281626676
	pesos_i(8993) := b"0000000000000000_0000000000000000_0001000101110110_0110101010101111"; -- 0.06821314584192002
	pesos_i(8994) := b"0000000000000000_0000000000000000_0001001100000100_1111000001001011"; -- 0.07429410764372711
	pesos_i(8995) := b"1111111111111111_1111111111111111_1101100001001001_1100110111110000"; -- -0.15512383360122928
	pesos_i(8996) := b"1111111111111111_1111111111111111_1110001100110100_1110000010110001"; -- -0.11247440030462968
	pesos_i(8997) := b"0000000000000000_0000000000000000_0000000100111010_0000000111010111"; -- 0.004791369420425611
	pesos_i(8998) := b"1111111111111111_1111111111111111_1110000100111110_0000010101101000"; -- -0.12014738294529824
	pesos_i(8999) := b"1111111111111111_1111111111111111_1111000000000011_1011111000110101"; -- -0.06244288643831714
	pesos_i(9000) := b"1111111111111111_1111111111111111_1111001001010001_0000011111111000"; -- -0.053451063157441164
	pesos_i(9001) := b"1111111111111111_1111111111111111_1111110101001100_1001010010010010"; -- -0.01055022658806927
	pesos_i(9002) := b"1111111111111111_1111111111111111_1111010111001100_0110111100000100"; -- -0.03984933998765103
	pesos_i(9003) := b"1111111111111111_1111111111111111_1101011010010001_0010100111011011"; -- -0.16184748079490552
	pesos_i(9004) := b"0000000000000000_0000000000000000_0010001001110101_1000100011001101"; -- 0.13460593234386997
	pesos_i(9005) := b"0000000000000000_0000000000000000_0001100111101010_0101010001111111"; -- 0.10123184298029497
	pesos_i(9006) := b"0000000000000000_0000000000000000_0000011111101101_1000011011111001"; -- 0.030968128104449204
	pesos_i(9007) := b"0000000000000000_0000000000000000_0000111111101011_0111000010000101"; -- 0.062186272178051234
	pesos_i(9008) := b"0000000000000000_0000000000000000_0001011110100000_0000110011011010"; -- 0.09228592225590401
	pesos_i(9009) := b"1111111111111111_1111111111111111_1111000011100001_0110010001001110"; -- -0.05906079388181577
	pesos_i(9010) := b"1111111111111111_1111111111111111_1110011100100000_1011000011111001"; -- -0.09715742043820635
	pesos_i(9011) := b"0000000000000000_0000000000000000_0001000100100101_1001110010110000"; -- 0.06698016458358713
	pesos_i(9012) := b"1111111111111111_1111111111111111_1101100011100111_1110100110001011"; -- -0.15271129954377108
	pesos_i(9013) := b"0000000000000000_0000000000000000_0010001011010100_1100000011010101"; -- 0.1360588569409033
	pesos_i(9014) := b"0000000000000000_0000000000000000_0000001101100001_1101110110001110"; -- 0.013212058222293393
	pesos_i(9015) := b"0000000000000000_0000000000000000_0001101101100110_0011000001100110"; -- 0.10702803122145739
	pesos_i(9016) := b"1111111111111111_1111111111111111_1111100110001000_1011000011100101"; -- -0.025258011058514163
	pesos_i(9017) := b"0000000000000000_0000000000000000_0001111100000101_1001110100011011"; -- 0.12117940817093806
	pesos_i(9018) := b"0000000000000000_0000000000000000_0001101101111101_1101000011000111"; -- 0.10738854279627291
	pesos_i(9019) := b"1111111111111111_1111111111111111_1110011100010011_1011110110011011"; -- -0.09735503174109024
	pesos_i(9020) := b"0000000000000000_0000000000000000_0001000000011100_1000010110101100"; -- 0.06293521346006885
	pesos_i(9021) := b"1111111111111111_1111111111111111_1110011101011110_0111000110101100"; -- -0.0962151484254013
	pesos_i(9022) := b"1111111111111111_1111111111111111_1110110000110000_1001100001000101"; -- -0.07738350219299042
	pesos_i(9023) := b"1111111111111111_1111111111111111_1110000000001101_1110100101001101"; -- -0.1247877300106489
	pesos_i(9024) := b"0000000000000000_0000000000000000_0001111000001010_1010110111100000"; -- 0.1173504517468308
	pesos_i(9025) := b"0000000000000000_0000000000000000_0001000111100100_0010010001000101"; -- 0.06988741563156743
	pesos_i(9026) := b"1111111111111111_1111111111111111_1101101010000000_1100110110100100"; -- -0.14647211778749758
	pesos_i(9027) := b"1111111111111111_1111111111111111_1111001111011000_0101100101110001"; -- -0.047480020404512026
	pesos_i(9028) := b"0000000000000000_0000000000000000_0001001010011111_0000010110111100"; -- 0.07273898924857762
	pesos_i(9029) := b"1111111111111111_1111111111111111_1110001110111110_1111101111010000"; -- -0.11036707086924995
	pesos_i(9030) := b"0000000000000000_0000000000000000_0001000000011101_0110010110101100"; -- 0.06294856505494846
	pesos_i(9031) := b"0000000000000000_0000000000000000_0001111100111010_1111001111100110"; -- 0.12199329724275453
	pesos_i(9032) := b"1111111111111111_1111111111111111_1111001010001001_0010110100011110"; -- -0.052594356674414616
	pesos_i(9033) := b"1111111111111111_1111111111111111_1110111100111000_0101011110100011"; -- -0.06554653435599418
	pesos_i(9034) := b"1111111111111111_1111111111111111_1101101000011110_1010010101011000"; -- -0.1479698811687068
	pesos_i(9035) := b"1111111111111111_1111111111111111_1110001000100000_0110011010010110"; -- -0.11669310405040433
	pesos_i(9036) := b"1111111111111111_1111111111111111_1111100011110100_1110001000001100"; -- -0.027513382000412426
	pesos_i(9037) := b"1111111111111111_1111111111111111_1111011100101000_0110010011101100"; -- -0.03453988297850662
	pesos_i(9038) := b"0000000000000000_0000000000000000_0000111100011100_0011110101000010"; -- 0.05902464735441529
	pesos_i(9039) := b"1111111111111111_1111111111111111_1110111111100110_1011101111010000"; -- -0.0628855339962253
	pesos_i(9040) := b"1111111111111111_1111111111111111_1101111000111101_0010001001100010"; -- -0.131879664560601
	pesos_i(9041) := b"1111111111111111_1111111111111111_1101100000100100_1010001100111101"; -- -0.15569095384393003
	pesos_i(9042) := b"0000000000000000_0000000000000000_0001001010100101_1101111010101110"; -- 0.07284347288279847
	pesos_i(9043) := b"0000000000000000_0000000000000000_0000110111000000_0011000000100101"; -- 0.05371380709261524
	pesos_i(9044) := b"1111111111111111_1111111111111111_1111100001101010_0001010011110111"; -- -0.029631318677821476
	pesos_i(9045) := b"1111111111111111_1111111111111111_1110000010101011_0101111111001111"; -- -0.12238503632877556
	pesos_i(9046) := b"0000000000000000_0000000000000000_0001111001101110_0101001010000110"; -- 0.11887088555522948
	pesos_i(9047) := b"1111111111111111_1111111111111111_1111100010111111_0011000000111101"; -- -0.028332695962003933
	pesos_i(9048) := b"0000000000000000_0000000000000000_0000010000010100_0001111011001110"; -- 0.015932011994541796
	pesos_i(9049) := b"0000000000000000_0000000000000000_0001000110100100_1110010111000011"; -- 0.068922386363577
	pesos_i(9050) := b"1111111111111111_1111111111111111_1101011110001011_1110011000100100"; -- -0.15802156080230492
	pesos_i(9051) := b"1111111111111111_1111111111111111_1111001110000000_1100000110111101"; -- -0.0488165773356393
	pesos_i(9052) := b"0000000000000000_0000000000000000_0001101010000001_0110011010000100"; -- 0.10353699417447783
	pesos_i(9053) := b"0000000000000000_0000000000000000_0010011101001101_1111110001011001"; -- 0.15353371791646156
	pesos_i(9054) := b"1111111111111111_1111111111111111_1110101001011000_1101011010101011"; -- -0.08458193128494622
	pesos_i(9055) := b"0000000000000000_0000000000000000_0000010110111101_0101010111110000"; -- 0.02242028347776029
	pesos_i(9056) := b"1111111111111111_1111111111111111_1110010101000101_0010101110111111"; -- -0.10441328600665943
	pesos_i(9057) := b"0000000000000000_0000000000000000_0000101100000101_0011010010001000"; -- 0.043048175152546025
	pesos_i(9058) := b"0000000000000000_0000000000000000_0000101010111110_0000010010011010"; -- 0.04196194417948119
	pesos_i(9059) := b"1111111111111111_1111111111111111_1111000000110100_1100011111100110"; -- -0.0616946280884611
	pesos_i(9060) := b"0000000000000000_0000000000000000_0001000100111101_0011010011111000"; -- 0.06734019324569078
	pesos_i(9061) := b"1111111111111111_1111111111111111_1111101001001000_0111101001111010"; -- -0.02233156695451302
	pesos_i(9062) := b"1111111111111111_1111111111111111_1110100111011111_0001111001101001"; -- -0.08643922738654448
	pesos_i(9063) := b"1111111111111111_1111111111111111_1111100101111100_1010101001111101"; -- -0.025441498260246883
	pesos_i(9064) := b"0000000000000000_0000000000000000_0000001111100101_0000011001001110"; -- 0.015213388452616123
	pesos_i(9065) := b"0000000000000000_0000000000000000_0001000001101001_0010001101011000"; -- 0.06410427943471912
	pesos_i(9066) := b"1111111111111111_1111111111111111_1110100110111001_0110101011001101"; -- -0.08701450831395138
	pesos_i(9067) := b"1111111111111111_1111111111111111_1110111000011101_0001110110001010"; -- -0.06986823448510861
	pesos_i(9068) := b"0000000000000000_0000000000000000_0010011011111001_0010001010010101"; -- 0.15223899975719443
	pesos_i(9069) := b"1111111111111111_1111111111111111_1111100000000101_0110000110101110"; -- -0.03116788379977976
	pesos_i(9070) := b"1111111111111111_1111111111111111_1101101100000110_0101110111011111"; -- -0.14443410201401388
	pesos_i(9071) := b"0000000000000000_0000000000000000_0001011111100110_1101000101011111"; -- 0.09336575089799658
	pesos_i(9072) := b"1111111111111111_1111111111111111_1110100010101010_0111000001001000"; -- -0.09114931348636099
	pesos_i(9073) := b"1111111111111111_1111111111111111_1110100101010110_0000010010010101"; -- -0.0885312209702629
	pesos_i(9074) := b"1111111111111111_1111111111111111_1111111011001001_1101000010101111"; -- -0.004733044998417323
	pesos_i(9075) := b"1111111111111111_1111111111111111_1111000111110000_0111010001011111"; -- -0.054924704357736484
	pesos_i(9076) := b"1111111111111111_1111111111111111_1110000111000110_1101000011001110"; -- -0.11806006395923735
	pesos_i(9077) := b"0000000000000000_0000000000000000_0000111011001101_1110010101101011"; -- 0.057829226063068985
	pesos_i(9078) := b"0000000000000000_0000000000000000_0010010111101101_1011011011011010"; -- 0.14815848178087326
	pesos_i(9079) := b"1111111111111111_1111111111111111_1111101110101111_0110011100010011"; -- -0.016854818138341825
	pesos_i(9080) := b"0000000000000000_0000000000000000_0000000011010011_1111100000010011"; -- 0.0032343908127757982
	pesos_i(9081) := b"0000000000000000_0000000000000000_0001111011111101_0101000111011100"; -- 0.12105285290248052
	pesos_i(9082) := b"0000000000000000_0000000000000000_0001001000001011_0001011100000001"; -- 0.07048171782790996
	pesos_i(9083) := b"0000000000000000_0000000000000000_0001101110000001_1001111101010010"; -- 0.10744663006141027
	pesos_i(9084) := b"1111111111111111_1111111111111111_1110111001101111_0000110010100100"; -- -0.06861802092482502
	pesos_i(9085) := b"0000000000000000_0000000000000000_0010000100000000_1011101001100110"; -- 0.12891736019743485
	pesos_i(9086) := b"1111111111111111_1111111111111111_1110010011100111_1011101011111011"; -- -0.10583907478400315
	pesos_i(9087) := b"0000000000000000_0000000000000000_0010000101100001_0111100011010011"; -- 0.13039355424203317
	pesos_i(9088) := b"0000000000000000_0000000000000000_0000101001011110_0110010100101010"; -- 0.04050285608892726
	pesos_i(9089) := b"1111111111111111_1111111111111111_1101111000010101_1100100100010101"; -- -0.13248008007192985
	pesos_i(9090) := b"0000000000000000_0000000000000000_0000001000000110_1111110101010011"; -- 0.007919151938731958
	pesos_i(9091) := b"1111111111111111_1111111111111111_1111101100100100_1000000100101001"; -- -0.01897423514017897
	pesos_i(9092) := b"1111111111111111_1111111111111111_1110000111101100_0000001111100111"; -- -0.11749244314136933
	pesos_i(9093) := b"1111111111111111_1111111111111111_1111100110001111_0010100100001000"; -- -0.02515929743145027
	pesos_i(9094) := b"0000000000000000_0000000000000000_0000010110011010_1111001101100101"; -- 0.02189561107278357
	pesos_i(9095) := b"1111111111111111_1111111111111111_1110010011100001_1110100011110111"; -- -0.10592788662968913
	pesos_i(9096) := b"1111111111111111_1111111111111111_1110010000100010_1001101010101010"; -- -0.1088469823831195
	pesos_i(9097) := b"0000000000000000_0000000000000000_0001001100011001_1001010010001110"; -- 0.0746090741867601
	pesos_i(9098) := b"0000000000000000_0000000000000000_0000001110110010_1001110010111110"; -- 0.014444157045255398
	pesos_i(9099) := b"1111111111111111_1111111111111111_1101110011110011_1100100001101010"; -- -0.13690516867350147
	pesos_i(9100) := b"0000000000000000_0000000000000000_0000001111010010_0110011100111111"; -- 0.014929249548328532
	pesos_i(9101) := b"1111111111111111_1111111111111111_1111110010101010_0001000100111101"; -- -0.013029978396451434
	pesos_i(9102) := b"0000000000000000_0000000000000000_0010011010100100_1000001010001011"; -- 0.15094772226453865
	pesos_i(9103) := b"0000000000000000_0000000000000000_0000100100111001_1000111000111111"; -- 0.03603447944122969
	pesos_i(9104) := b"0000000000000000_0000000000000000_0001000111010010_0010001111111010"; -- 0.06961274007024616
	pesos_i(9105) := b"1111111111111111_1111111111111111_1110110010101101_1000110001111110"; -- -0.07547685548315355
	pesos_i(9106) := b"0000000000000000_0000000000000000_0001010110001001_0000111011110000"; -- 0.08412259453616647
	pesos_i(9107) := b"1111111111111111_1111111111111111_1110111001011001_1101001110111010"; -- -0.06894184781695037
	pesos_i(9108) := b"1111111111111111_1111111111111111_1110101001101010_1000101011010100"; -- -0.08431179362529238
	pesos_i(9109) := b"0000000000000000_0000000000000000_0001011100001101_1001011000100010"; -- 0.09005106293606613
	pesos_i(9110) := b"0000000000000000_0000000000000000_0010001000100011_0100100010100101"; -- 0.1333508875123492
	pesos_i(9111) := b"0000000000000000_0000000000000000_0001101110111001_1010000101110100"; -- 0.1083012494357361
	pesos_i(9112) := b"1111111111111111_1111111111111111_1111001011011001_0111001111001110"; -- -0.05136944024003151
	pesos_i(9113) := b"1111111111111111_1111111111111111_1111000000001000_1001011111011000"; -- -0.062368878979632114
	pesos_i(9114) := b"0000000000000000_0000000000000000_0000011011010100_1101101100000000"; -- 0.026685416785784125
	pesos_i(9115) := b"1111111111111111_1111111111111111_1111110111011110_0001001001111000"; -- -0.008330198092725722
	pesos_i(9116) := b"1111111111111111_1111111111111111_1110101101110101_1011101011100101"; -- -0.08023483181664111
	pesos_i(9117) := b"1111111111111111_1111111111111111_1111100001000111_1001001100000110"; -- -0.030157862580782718
	pesos_i(9118) := b"0000000000000000_0000000000000000_0010000010001111_1011001000100011"; -- 0.12719262463357114
	pesos_i(9119) := b"1111111111111111_1111111111111111_1101110100011110_1001110100100100"; -- -0.13625161997491037
	pesos_i(9120) := b"1111111111111111_1111111111111111_1101111100100001_0111001111010001"; -- -0.1283958068167597
	pesos_i(9121) := b"0000000000000000_0000000000000000_0001000000100010_0101001000100101"; -- 0.06302369505028742
	pesos_i(9122) := b"1111111111111111_1111111111111111_1111010110010010_0011111111000010"; -- -0.040737166528864485
	pesos_i(9123) := b"0000000000000000_0000000000000000_0001101011000110_1001001110100100"; -- 0.10459254034861866
	pesos_i(9124) := b"0000000000000000_0000000000000000_0001101100111010_1011011111101101"; -- 0.10636472265041937
	pesos_i(9125) := b"0000000000000000_0000000000000000_0010011101010001_1111010010000110"; -- 0.1535942867541417
	pesos_i(9126) := b"1111111111111111_1111111111111111_1111101001101011_0011011110010000"; -- -0.02180149786285122
	pesos_i(9127) := b"1111111111111111_1111111111111111_1101111100110010_1011010011101000"; -- -0.12813252763086316
	pesos_i(9128) := b"1111111111111111_1111111111111111_1110101000110111_1000010000011111"; -- -0.08509039146669028
	pesos_i(9129) := b"1111111111111111_1111111111111111_1111001111101010_1101010011101011"; -- -0.047198002514194363
	pesos_i(9130) := b"1111111111111111_1111111111111111_1111000001111011_0101111111111111"; -- -0.060617447085472106
	pesos_i(9131) := b"0000000000000000_0000000000000000_0000111010111001_0001110101010011"; -- 0.05751212375240787
	pesos_i(9132) := b"0000000000000000_0000000000000000_0001010011011000_0010111101010111"; -- 0.0814237200251625
	pesos_i(9133) := b"1111111111111111_1111111111111111_1101110000101011_1100011001101011"; -- -0.13995704547051213
	pesos_i(9134) := b"0000000000000000_0000000000000000_0000000111101110_1100010100011001"; -- 0.007549589802558922
	pesos_i(9135) := b"0000000000000000_0000000000000000_0010010111011110_0001001011001111"; -- 0.1479198222188893
	pesos_i(9136) := b"0000000000000000_0000000000000000_0001101111000110_1101111111100100"; -- 0.10850333516728468
	pesos_i(9137) := b"0000000000000000_0000000000000000_0001111010100001_0010000100101111"; -- 0.11964614293315129
	pesos_i(9138) := b"1111111111111111_1111111111111111_1110100101011011_0110100110111010"; -- -0.0884488983115689
	pesos_i(9139) := b"1111111111111111_1111111111111111_1111101001101101_1001011100010101"; -- -0.021765286695091722
	pesos_i(9140) := b"1111111111111111_1111111111111111_1101101010101001_1110101010001101"; -- -0.1458447844434048
	pesos_i(9141) := b"1111111111111111_1111111111111111_1111011010001111_1100100111110111"; -- -0.036868455172381506
	pesos_i(9142) := b"1111111111111111_1111111111111111_1111010010100101_0101110001011011"; -- -0.04435179504427609
	pesos_i(9143) := b"0000000000000000_0000000000000000_0001011101111101_0101110110111011"; -- 0.09175668538618449
	pesos_i(9144) := b"0000000000000000_0000000000000000_0000100111000100_1111100101110100"; -- 0.0381618412204786
	pesos_i(9145) := b"1111111111111111_1111111111111111_1111111110111010_0001111011100111"; -- -0.0010662733132726088
	pesos_i(9146) := b"1111111111111111_1111111111111111_1111101011000010_1111110111111100"; -- -0.020462156305315032
	pesos_i(9147) := b"0000000000000000_0000000000000000_0010001111110100_1000110110011101"; -- 0.14045033540764423
	pesos_i(9148) := b"1111111111111111_1111111111111111_1110110110100100_0110101101011011"; -- -0.07170990979392383
	pesos_i(9149) := b"1111111111111111_1111111111111111_1110001110111000_0000011010100100"; -- -0.11047323705765909
	pesos_i(9150) := b"1111111111111111_1111111111111111_1110110100111111_0111110110000101"; -- -0.07324996464723055
	pesos_i(9151) := b"0000000000000000_0000000000000000_0001000000011110_1110000110000011"; -- 0.06297120518766658
	pesos_i(9152) := b"0000000000000000_0000000000000000_0001011000000011_0001110010000111"; -- 0.08598497669612665
	pesos_i(9153) := b"0000000000000000_0000000000000000_0001101001001010_0001001100001001"; -- 0.10269278486861225
	pesos_i(9154) := b"1111111111111111_1111111111111111_1111000000100100_1110001000011010"; -- -0.06193720679182522
	pesos_i(9155) := b"1111111111111111_1111111111111111_1110010011011011_0011000110100111"; -- -0.10603036567811608
	pesos_i(9156) := b"0000000000000000_0000000000000000_0001000111110010_1100101001001000"; -- 0.07011093393282203
	pesos_i(9157) := b"1111111111111111_1111111111111111_1101100010001111_1100100000011011"; -- -0.15405606595757884
	pesos_i(9158) := b"0000000000000000_0000000000000000_0000000110001100_1001101001111010"; -- 0.006051688014686797
	pesos_i(9159) := b"0000000000000000_0000000000000000_0010001000011111_0111010110110001"; -- 0.13329253741060906
	pesos_i(9160) := b"1111111111111111_1111111111111111_1110000110001100_1000111001001110"; -- -0.11894903748579892
	pesos_i(9161) := b"0000000000000000_0000000000000000_0000101011101110_1111000011000000"; -- 0.04270844169966778
	pesos_i(9162) := b"0000000000000000_0000000000000000_0001110000011111_0100111000000100"; -- 0.10985267256404527
	pesos_i(9163) := b"1111111111111111_1111111111111111_1111011010111100_1001011011101000"; -- -0.03618485284392611
	pesos_i(9164) := b"0000000000000000_0000000000000000_0001011110111111_1010001011011111"; -- 0.09276788656473503
	pesos_i(9165) := b"1111111111111111_1111111111111111_1111011001001100_0111011110000101"; -- -0.03789570800178147
	pesos_i(9166) := b"0000000000000000_0000000000000000_0010011001011101_0010011111111111"; -- 0.14985895127972457
	pesos_i(9167) := b"1111111111111111_1111111111111111_1111110100111100_1000100001101010"; -- -0.010795091743302105
	pesos_i(9168) := b"0000000000000000_0000000000000000_0010010100111110_0101011100010101"; -- 0.14548248550418771
	pesos_i(9169) := b"1111111111111111_1111111111111111_1101100011011110_0100000000000111"; -- -0.15285873245558707
	pesos_i(9170) := b"0000000000000000_0000000000000000_0010001011000011_0001111110101000"; -- 0.13578985078312564
	pesos_i(9171) := b"1111111111111111_1111111111111111_1111010101000001_0111101010010101"; -- -0.041969622180589736
	pesos_i(9172) := b"0000000000000000_0000000000000000_0001110110001000_1011100111101100"; -- 0.1153675270122541
	pesos_i(9173) := b"0000000000000000_0000000000000000_0000000010001100_0010001100100101"; -- 0.0021383251795624924
	pesos_i(9174) := b"0000000000000000_0000000000000000_0001111011101011_0000101010110001"; -- 0.12077395276637841
	pesos_i(9175) := b"0000000000000000_0000000000000000_0001011000100001_1110111001101001"; -- 0.08645525031356989
	pesos_i(9176) := b"1111111111111111_1111111111111111_1110001010000110_0101100011111000"; -- -0.115137519331842
	pesos_i(9177) := b"1111111111111111_1111111111111111_1111101101000001_0111000101111001"; -- -0.018532665236374337
	pesos_i(9178) := b"1111111111111111_1111111111111111_1110111000101001_1100101011110000"; -- -0.0696747935858929
	pesos_i(9179) := b"1111111111111111_1111111111111111_1110001110011000_0010010010000111"; -- -0.1109597368760721
	pesos_i(9180) := b"1111111111111111_1111111111111111_1111110111101010_1100101001100110"; -- -0.008136129416915864
	pesos_i(9181) := b"1111111111111111_1111111111111111_1101111001001110_0110010000111110"; -- -0.13161633963179095
	pesos_i(9182) := b"0000000000000000_0000000000000000_0000111111110001_1110111011000000"; -- 0.062285348746012145
	pesos_i(9183) := b"0000000000000000_0000000000000000_0000111010010010_0111101101100101"; -- 0.05692263811505931
	pesos_i(9184) := b"1111111111111111_1111111111111111_1111110111101101_1101000000000110"; -- -0.008090017798559113
	pesos_i(9185) := b"1111111111111111_1111111111111111_1110101010001011_0101010100111000"; -- -0.08381144888521065
	pesos_i(9186) := b"1111111111111111_1111111111111111_1110111110001110_0001011010110001"; -- -0.06423814949804557
	pesos_i(9187) := b"1111111111111111_1111111111111111_1101110010111001_1111010101101101"; -- -0.13778749560704323
	pesos_i(9188) := b"0000000000000000_0000000000000000_0000001101000001_1000011110101110"; -- 0.012718658369586999
	pesos_i(9189) := b"1111111111111111_1111111111111111_1101011010110010_0010100100111001"; -- -0.16134397841015075
	pesos_i(9190) := b"0000000000000000_0000000000000000_0000110010000000_0011001011110100"; -- 0.04883116200258622
	pesos_i(9191) := b"0000000000000000_0000000000000000_0001101110000101_0000010011110001"; -- 0.10749846340812678
	pesos_i(9192) := b"1111111111111111_1111111111111111_1111111000011001_1100000110001001"; -- -0.007419494641603978
	pesos_i(9193) := b"0000000000000000_0000000000000000_0001110100001111_0101110110000000"; -- 0.11351570483175122
	pesos_i(9194) := b"0000000000000000_0000000000000000_0000100001011000_0101101000010000"; -- 0.032598141504720596
	pesos_i(9195) := b"1111111111111111_1111111111111111_1101011111000110_0010010111101111"; -- -0.15713274880767625
	pesos_i(9196) := b"1111111111111111_1111111111111111_1111111011100100_1111101110111010"; -- -0.004318491972403198
	pesos_i(9197) := b"0000000000000000_0000000000000000_0001101110011111_1010101100101010"; -- 0.10790509955513398
	pesos_i(9198) := b"1111111111111111_1111111111111111_1111000100001111_1000110100101010"; -- -0.05835645412638074
	pesos_i(9199) := b"0000000000000000_0000000000000000_0001101001001110_0111100010110010"; -- 0.10275987949213683
	pesos_i(9200) := b"0000000000000000_0000000000000000_0001100100001100_1011111111111001"; -- 0.09785079782363042
	pesos_i(9201) := b"1111111111111111_1111111111111111_1110100111101011_1100110010100100"; -- -0.08624573708043587
	pesos_i(9202) := b"0000000000000000_0000000000000000_0000100100101011_1100101100010001"; -- 0.035824481577579316
	pesos_i(9203) := b"1111111111111111_1111111111111111_1111100000001111_0010011010110111"; -- -0.03101881058302915
	pesos_i(9204) := b"1111111111111111_1111111111111111_1111100110111000_0010101010110111"; -- -0.024533586744155938
	pesos_i(9205) := b"1111111111111111_1111111111111111_1110010110111000_0011110111110011"; -- -0.10265744030161786
	pesos_i(9206) := b"1111111111111111_1111111111111111_1110110010011000_0011101110100000"; -- -0.07580211015185997
	pesos_i(9207) := b"0000000000000000_0000000000000000_0001010100000010_1101000101000001"; -- 0.08207424011992867
	pesos_i(9208) := b"1111111111111111_1111111111111111_1101111100010100_0011010001101001"; -- -0.12859795043344227
	pesos_i(9209) := b"1111111111111111_1111111111111111_1111010101110000_1110011111110000"; -- -0.04124594109392493
	pesos_i(9210) := b"0000000000000000_0000000000000000_0001010101001010_1000010011100100"; -- 0.08316832135615666
	pesos_i(9211) := b"1111111111111111_1111111111111111_1111010000000001_0011111010000001"; -- -0.04685601577355045
	pesos_i(9212) := b"1111111111111111_1111111111111111_1110111110011001_1000100011000111"; -- -0.0640635026929056
	pesos_i(9213) := b"1111111111111111_1111111111111111_1110000011010101_0101000001001110"; -- -0.12174509150490175
	pesos_i(9214) := b"0000000000000000_0000000000000000_0001111011101001_1010100010010011"; -- 0.12075284559795181
	pesos_i(9215) := b"0000000000000000_0000000000000000_0010010101101010_0100111011000010"; -- 0.14615337605159473
	pesos_i(9216) := b"0000000000000000_0000000000000000_0001111111011110_1011010111100100"; -- 0.12449204263228332
	pesos_i(9217) := b"0000000000000000_0000000000000000_0001101110000000_1101101101111111"; -- 0.1074349579156318
	pesos_i(9218) := b"0000000000000000_0000000000000000_0010000110001011_1001000111010010"; -- 0.1310359132509085
	pesos_i(9219) := b"1111111111111111_1111111111111111_1110000110011000_0101000010110111"; -- -0.11876960300112215
	pesos_i(9220) := b"1111111111111111_1111111111111111_1111100101101001_1000011101101011"; -- -0.02573350551465371
	pesos_i(9221) := b"1111111111111111_1111111111111111_1101110100011010_0010111001001100"; -- -0.13631926196399455
	pesos_i(9222) := b"1111111111111111_1111111111111111_1110000110000111_1110100001011110"; -- -0.11901996332828252
	pesos_i(9223) := b"0000000000000000_0000000000000000_0001100001000000_1101011000110101"; -- 0.0947393303310574
	pesos_i(9224) := b"0000000000000000_0000000000000000_0000111101000001_1000100100001110"; -- 0.05959374044931171
	pesos_i(9225) := b"1111111111111111_1111111111111111_1110110010101010_1110100111010101"; -- -0.07551706829284542
	pesos_i(9226) := b"0000000000000000_0000000000000000_0001101101111100_0010000111100100"; -- 0.10736285998797705
	pesos_i(9227) := b"1111111111111111_1111111111111111_1111000011101110_1000111000001101"; -- -0.05885994139640083
	pesos_i(9228) := b"0000000000000000_0000000000000000_0000000110000010_1101100001010011"; -- 0.005902786578470107
	pesos_i(9229) := b"1111111111111111_1111111111111111_1110111111000101_0110010110100110"; -- -0.06339420976910286
	pesos_i(9230) := b"0000000000000000_0000000000000000_0000010101100111_0100101000111001"; -- 0.021107329203667806
	pesos_i(9231) := b"1111111111111111_1111111111111111_1110100110101000_0101110111101110"; -- -0.08727467490105452
	pesos_i(9232) := b"0000000000000000_0000000000000000_0001101101110101_1011010110101000"; -- 0.10726485591586317
	pesos_i(9233) := b"1111111111111111_1111111111111111_1111001111111000_0101001110000011"; -- -0.04699209273142875
	pesos_i(9234) := b"1111111111111111_1111111111111111_1111100111111011_0010001110100000"; -- -0.02351167042528797
	pesos_i(9235) := b"0000000000000000_0000000000000000_0000111100000001_1111111000111010"; -- 0.05862416189606176
	pesos_i(9236) := b"1111111111111111_1111111111111111_1110111011101001_1100000100100011"; -- -0.0667456903704451
	pesos_i(9237) := b"0000000000000000_0000000000000000_0001111100100100_1000011001001011"; -- 0.12165107094719324
	pesos_i(9238) := b"0000000000000000_0000000000000000_0010001110011000_1101010110001000"; -- 0.13905081334174502
	pesos_i(9239) := b"1111111111111111_1111111111111111_1111111100111001_1011100000111011"; -- -0.0030255181475157588
	pesos_i(9240) := b"0000000000000000_0000000000000000_0010010100011001_1111001010011010"; -- 0.14492717982882952
	pesos_i(9241) := b"1111111111111111_1111111111111111_1111111010111100_0000010100111101"; -- -0.004943535436668091
	pesos_i(9242) := b"1111111111111111_1111111111111111_1110101111101101_1100010000010100"; -- -0.07840322992205664
	pesos_i(9243) := b"0000000000000000_0000000000000000_0000010100010001_0000101111111111"; -- 0.019791364492403807
	pesos_i(9244) := b"1111111111111111_1111111111111111_1111110001100001_1101111110001100"; -- -0.01413157301581256
	pesos_i(9245) := b"0000000000000000_0000000000000000_0001000000100010_1000110010101100"; -- 0.06302718346553328
	pesos_i(9246) := b"1111111111111111_1111111111111111_1110010000011010_0100101000110010"; -- -0.10897384915059286
	pesos_i(9247) := b"0000000000000000_0000000000000000_0000011000010001_1010100100111000"; -- 0.02370698559355649
	pesos_i(9248) := b"0000000000000000_0000000000000000_0001000111001110_1011001011100111"; -- 0.06956022400170099
	pesos_i(9249) := b"1111111111111111_1111111111111111_1101011100011010_1011110101100010"; -- -0.15974823347642772
	pesos_i(9250) := b"0000000000000000_0000000000000000_0000101011101010_0101011000011110"; -- 0.04263818973013295
	pesos_i(9251) := b"0000000000000000_0000000000000000_0000111110001010_0010000011111101"; -- 0.060701429242412994
	pesos_i(9252) := b"1111111111111111_1111111111111111_1110100110011001_1100001000001001"; -- -0.08749758988288996
	pesos_i(9253) := b"1111111111111111_1111111111111111_1111110101110110_1101110100001000"; -- -0.00990503848519173
	pesos_i(9254) := b"1111111111111111_1111111111111111_1110110010111000_1010011000101101"; -- -0.07530747786665637
	pesos_i(9255) := b"1111111111111111_1111111111111111_1111000010111001_1001111101011001"; -- -0.05966762622442124
	pesos_i(9256) := b"0000000000000000_0000000000000000_0001111100110100_1100111110011001"; -- 0.12189958081698041
	pesos_i(9257) := b"1111111111111111_1111111111111111_1110010110100110_1111110000000101"; -- -0.1029207694486722
	pesos_i(9258) := b"1111111111111111_1111111111111111_1110011111000001_1000010100101000"; -- -0.0947033670548089
	pesos_i(9259) := b"0000000000000000_0000000000000000_0001000011010001_1001000110011111"; -- 0.06569776655637087
	pesos_i(9260) := b"1111111111111111_1111111111111111_1110100100101111_0110110101011110"; -- -0.08912006814588068
	pesos_i(9261) := b"0000000000000000_0000000000000000_0010000001010100_0111110110100101"; -- 0.12628922717471044
	pesos_i(9262) := b"0000000000000000_0000000000000000_0010000110100010_0000111000110011"; -- 0.13137902015779002
	pesos_i(9263) := b"0000000000000000_0000000000000000_0010001000101001_1101101100001011"; -- 0.13345116622419348
	pesos_i(9264) := b"0000000000000000_0000000000000000_0001100001101010_1110000010000011"; -- 0.0953808135200665
	pesos_i(9265) := b"0000000000000000_0000000000000000_0000001110000000_1100110000111011"; -- 0.013684048083758534
	pesos_i(9266) := b"1111111111111111_1111111111111111_1111010101100101_0111001001011100"; -- -0.04142079592703653
	pesos_i(9267) := b"0000000000000000_0000000000000000_0001111011101110_0101010101100101"; -- 0.1208241816036788
	pesos_i(9268) := b"0000000000000000_0000000000000000_0000110000001101_1111000010011100"; -- 0.0470877055904295
	pesos_i(9269) := b"1111111111111111_1111111111111111_1111111100110101_1100010101111101"; -- -0.0030857630627470294
	pesos_i(9270) := b"0000000000000000_0000000000000000_0001110100001101_1110011111110110"; -- 0.1134934401136184
	pesos_i(9271) := b"0000000000000000_0000000000000000_0010111011111110_0111010000100100"; -- 0.18357015499874968
	pesos_i(9272) := b"0000000000000000_0000000000000000_0000000111100000_1001000010001000"; -- 0.007332833428684448
	pesos_i(9273) := b"0000000000000000_0000000000000000_0010100000011011_0000011101100000"; -- 0.15666242690949292
	pesos_i(9274) := b"0000000000000000_0000000000000000_0000110111100011_1001000110011001"; -- 0.05425367347455705
	pesos_i(9275) := b"1111111111111111_1111111111111111_1111101110010101_1101101101111110"; -- -0.01724460760005859
	pesos_i(9276) := b"1111111111111111_1111111111111111_1110100101000111_1101000101100100"; -- -0.08874789540607003
	pesos_i(9277) := b"0000000000000000_0000000000000000_0010100101110000_1101110100111000"; -- 0.16187842011817288
	pesos_i(9278) := b"1111111111111111_1111111111111111_1111010000100100_0001111100001000"; -- -0.04632383398393916
	pesos_i(9279) := b"0000000000000000_0000000000000000_0001101010111110_0010100100011111"; -- 0.10446412081669768
	pesos_i(9280) := b"0000000000000000_0000000000000000_0000101011001110_0001011010100011"; -- 0.0422071598744867
	pesos_i(9281) := b"1111111111111111_1111111111111111_1110001010010000_0101100110101001"; -- -0.11498489031890888
	pesos_i(9282) := b"0000000000000000_0000000000000000_0010000111110100_0101111011010010"; -- 0.1326350462135761
	pesos_i(9283) := b"1111111111111111_1111111111111111_1111110100010011_0111000111101001"; -- -0.011422043457473741
	pesos_i(9284) := b"1111111111111111_1111111111111111_1110001011001010_0010101000101100"; -- -0.11410271106109796
	pesos_i(9285) := b"0000000000000000_0000000000000000_0000101101001101_0011100100000010"; -- 0.044147074800049646
	pesos_i(9286) := b"1111111111111111_1111111111111111_1111001001111110_1111101011001011"; -- -0.05274994409529649
	pesos_i(9287) := b"0000000000000000_0000000000000000_0000100100110000_1011101000001010"; -- 0.035899760679408636
	pesos_i(9288) := b"0000000000000000_0000000000000000_0000010100111000_0111000101011101"; -- 0.02039249911369142
	pesos_i(9289) := b"1111111111111111_1111111111111111_1111011110010010_1110010100101100"; -- -0.032914807057986994
	pesos_i(9290) := b"0000000000000000_0000000000000000_0000111011011010_1010010111000001"; -- 0.05802379573011035
	pesos_i(9291) := b"1111111111111111_1111111111111111_1101100100011110_1111010110000011"; -- -0.1518713526263162
	pesos_i(9292) := b"1111111111111111_1111111111111111_1110100111110111_1010100000011011"; -- -0.08606480932316193
	pesos_i(9293) := b"0000000000000000_0000000000000000_0001010100000101_1010101001011001"; -- 0.08211769747752372
	pesos_i(9294) := b"1111111111111111_1111111111111111_1101100110101001_1101010111001000"; -- -0.14975227233661362
	pesos_i(9295) := b"1111111111111111_1111111111111111_1111011110000010_1000011111001101"; -- -0.03316451307895046
	pesos_i(9296) := b"0000000000000000_0000000000000000_0000000100001011_1000110100101101"; -- 0.004082511475010717
	pesos_i(9297) := b"0000000000000000_0000000000000000_0000010010000010_0110101101001110"; -- 0.01761503847465797
	pesos_i(9298) := b"0000000000000000_0000000000000000_0000010001111001_1011000000110000"; -- 0.017481815181410055
	pesos_i(9299) := b"1111111111111111_1111111111111111_1110001010011011_0010110001010001"; -- -0.11481974621750905
	pesos_i(9300) := b"1111111111111111_1111111111111111_1111011101111010_0110001001001001"; -- -0.033288819556638344
	pesos_i(9301) := b"1111111111111111_1111111111111111_1110010100111110_1111100000010111"; -- -0.10450791782098451
	pesos_i(9302) := b"1111111111111111_1111111111111111_1111101000111100_1100101000100111"; -- -0.022509923355950017
	pesos_i(9303) := b"0000000000000000_0000000000000000_0001110110110000_0010001100000000"; -- 0.11596888312624111
	pesos_i(9304) := b"0000000000000000_0000000000000000_0001110011000101_0111100101111011"; -- 0.11238822235641051
	pesos_i(9305) := b"0000000000000000_0000000000000000_0001110010110101_1100000111111111"; -- 0.11214840380242316
	pesos_i(9306) := b"1111111111111111_1111111111111111_1111101110001111_0100000010100001"; -- -0.017345390867428243
	pesos_i(9307) := b"1111111111111111_1111111111111111_1111001001111100_1010110100001111"; -- -0.052785094989711755
	pesos_i(9308) := b"0000000000000000_0000000000000000_0001111000101100_0011001000010000"; -- 0.11786187075399608
	pesos_i(9309) := b"0000000000000000_0000000000000000_0000110100000000_1111000101001010"; -- 0.050795631862671574
	pesos_i(9310) := b"0000000000000000_0000000000000000_0010001011001001_1110010101001110"; -- 0.13589318434208972
	pesos_i(9311) := b"0000000000000000_0000000000000000_0010001011101000_0000111110001110"; -- 0.1363534661923535
	pesos_i(9312) := b"1111111111111111_1111111111111111_1110011011111001_0000010011100100"; -- -0.09776277012725525
	pesos_i(9313) := b"1111111111111111_1111111111111111_1111111000000001_0100010111011110"; -- -0.00779307691361072
	pesos_i(9314) := b"0000000000000000_0000000000000000_0001000000100011_0101011101011000"; -- 0.06303926376431378
	pesos_i(9315) := b"0000000000000000_0000000000000000_0010001100011110_1110101111100100"; -- 0.13719057392856795
	pesos_i(9316) := b"1111111111111111_1111111111111111_1101111111111011_1000110010100110"; -- -0.125067910603659
	pesos_i(9317) := b"1111111111111111_1111111111111111_1101111000011010_1000011001000110"; -- -0.13240776817620853
	pesos_i(9318) := b"1111111111111111_1111111111111111_1110110101010101_0000101000101110"; -- -0.0729211460686359
	pesos_i(9319) := b"1111111111111111_1111111111111111_1111101111001010_0110101000111001"; -- -0.016442643323463804
	pesos_i(9320) := b"0000000000000000_0000000000000000_0000011001100011_0001001001010100"; -- 0.024949212629681774
	pesos_i(9321) := b"1111111111111111_1111111111111111_1111100011010100_1010011110101000"; -- -0.02800514368985497
	pesos_i(9322) := b"1111111111111111_1111111111111111_1111000111111110_1110010100010110"; -- -0.05470436305446477
	pesos_i(9323) := b"0000000000000000_0000000000000000_0000100000010111_1000001110010010"; -- 0.031608794432414024
	pesos_i(9324) := b"1111111111111111_1111111111111111_1111100100011110_0010011100110000"; -- -0.026883650633110046
	pesos_i(9325) := b"1111111111111111_1111111111111111_1101111110001000_0011011011001010"; -- -0.12682778893612606
	pesos_i(9326) := b"1111111111111111_1111111111111111_1101111001100000_0101101101000000"; -- -0.13134221728368342
	pesos_i(9327) := b"0000000000000000_0000000000000000_0001100010110010_0001100010110101"; -- 0.09646753717830751
	pesos_i(9328) := b"0000000000000000_0000000000000000_0000010111100010_0101110001110111"; -- 0.022985247578452266
	pesos_i(9329) := b"1111111111111111_1111111111111111_1111001000011000_1011001100100011"; -- -0.054310611610976126
	pesos_i(9330) := b"1111111111111111_1111111111111111_1110000110000101_0001001010011000"; -- -0.11906322282335234
	pesos_i(9331) := b"1111111111111111_1111111111111111_1111110011011011_0111000011001000"; -- -0.012276602858089543
	pesos_i(9332) := b"0000000000000000_0000000000000000_0001100101110110_0001100000100000"; -- 0.09945822503290469
	pesos_i(9333) := b"0000000000000000_0000000000000000_0001001111100100_0010101010010110"; -- 0.07770029214367141
	pesos_i(9334) := b"0000000000000000_0000000000000000_0000111000111100_0101010100100011"; -- 0.05560810180939578
	pesos_i(9335) := b"1111111111111111_1111111111111111_1111010100111010_1000010101000001"; -- -0.0420757977180426
	pesos_i(9336) := b"0000000000000000_0000000000000000_0010011000101110_1000110101100011"; -- 0.1491478316341981
	pesos_i(9337) := b"0000000000000000_0000000000000000_0010000001111110_0111101010110010"; -- 0.12692992063206238
	pesos_i(9338) := b"0000000000000000_0000000000000000_0001111010101011_0110101110000100"; -- 0.11980316137824866
	pesos_i(9339) := b"0000000000000000_0000000000000000_0000100110111011_0100011101100001"; -- 0.038013898074341815
	pesos_i(9340) := b"1111111111111111_1111111111111111_1111010000011010_1100100100110011"; -- -0.04646627916682203
	pesos_i(9341) := b"0000000000000000_0000000000000000_0010100001101000_0001111000100110"; -- 0.15783871113178782
	pesos_i(9342) := b"0000000000000000_0000000000000000_0000001111110001_1011011011111100"; -- 0.01540702485287672
	pesos_i(9343) := b"1111111111111111_1111111111111111_1101100110001011_0001111101101101"; -- -0.15022090511782413
	pesos_i(9344) := b"0000000000000000_0000000000000000_0000010100100000_1110010010110011"; -- 0.02003316289830804
	pesos_i(9345) := b"0000000000000000_0000000000000000_0001011011101101_1111000111001100"; -- 0.08956824513331045
	pesos_i(9346) := b"1111111111111111_1111111111111111_1110100001100100_1111000011010001"; -- -0.09220976729613975
	pesos_i(9347) := b"1111111111111111_1111111111111111_1110000011010101_0110011001011101"; -- -0.12174377665851988
	pesos_i(9348) := b"0000000000000000_0000000000000000_0001100110010001_0011110110110110"; -- 0.09987245274374999
	pesos_i(9349) := b"1111111111111111_1111111111111111_1110000111100010_0001010100111101"; -- -0.11764399777082477
	pesos_i(9350) := b"1111111111111111_1111111111111111_1111001011101011_1101001010010001"; -- -0.05108913381648367
	pesos_i(9351) := b"0000000000000000_0000000000000000_0001000000001000_0101000000001011"; -- 0.06262684122781778
	pesos_i(9352) := b"1111111111111111_1111111111111111_1111110010010010_1111001110111101"; -- -0.013382688794443844
	pesos_i(9353) := b"0000000000000000_0000000000000000_0000010101101110_1011100011111110"; -- 0.02122074319894827
	pesos_i(9354) := b"0000000000000000_0000000000000000_0000111010011000_0010110011011111"; -- 0.057009510446362655
	pesos_i(9355) := b"0000000000000000_0000000000000000_0001010111100111_0101010101010111"; -- 0.08556111687243909
	pesos_i(9356) := b"0000000000000000_0000000000000000_0010001101101010_1100100101100100"; -- 0.1383481855696569
	pesos_i(9357) := b"0000000000000000_0000000000000000_0001011101001100_0010100010111100"; -- 0.09100584598233316
	pesos_i(9358) := b"0000000000000000_0000000000000000_0000010101001101_1001101000111100"; -- 0.020715369729474888
	pesos_i(9359) := b"0000000000000000_0000000000000000_0001011111001010_1011011110001010"; -- 0.09293696513661485
	pesos_i(9360) := b"1111111111111111_1111111111111111_1110110001000101_1011010011011000"; -- -0.07706136440811491
	pesos_i(9361) := b"1111111111111111_1111111111111111_1111001001001000_0101000111001100"; -- -0.05358399171578329
	pesos_i(9362) := b"1111111111111111_1111111111111111_1111101110010000_0011001100001000"; -- -0.01733094259415905
	pesos_i(9363) := b"1111111111111111_1111111111111111_1110110011011010_1011010011100101"; -- -0.07478780171562592
	pesos_i(9364) := b"0000000000000000_0000000000000000_0000010100110011_0100101110010110"; -- 0.020313953562117737
	pesos_i(9365) := b"0000000000000000_0000000000000000_0001100100111101_0011010101011010"; -- 0.09859021611053446
	pesos_i(9366) := b"1111111111111111_1111111111111111_1110010011011110_1101001110000101"; -- -0.10597494121695945
	pesos_i(9367) := b"0000000000000000_0000000000000000_0000010011110010_0001001101111010"; -- 0.019318787777523886
	pesos_i(9368) := b"0000000000000000_0000000000000000_0001110000000001_1011100001100110"; -- 0.10940124987659802
	pesos_i(9369) := b"0000000000000000_0000000000000000_0010010011110010_0011111101001111"; -- 0.14432140050096234
	pesos_i(9370) := b"0000000000000000_0000000000000000_0001010111011111_0001011100001111"; -- 0.08543533432912712
	pesos_i(9371) := b"1111111111111111_1111111111111111_1110101001110000_0001001001101100"; -- -0.08422741757367991
	pesos_i(9372) := b"0000000000000000_0000000000000000_0000111010101100_0100010101111111"; -- 0.05731615401887141
	pesos_i(9373) := b"0000000000000000_0000000000000000_0001101010111100_1001110010010101"; -- 0.10444048540961598
	pesos_i(9374) := b"0000000000000000_0000000000000000_0001001101011000_0111001011001110"; -- 0.07556836635129151
	pesos_i(9375) := b"0000000000000000_0000000000000000_0001010010000001_0000000110101000"; -- 0.08009348253086543
	pesos_i(9376) := b"1111111111111111_1111111111111111_1101100111000110_1010101111001111"; -- -0.14931226914586487
	pesos_i(9377) := b"0000000000000000_0000000000000000_0010001000100010_1110100111010011"; -- 0.13334523592506772
	pesos_i(9378) := b"1111111111111111_1111111111111111_1110001110010011_0101010101000111"; -- -0.11103312509158454
	pesos_i(9379) := b"0000000000000000_0000000000000000_0001110100011010_1110110010000000"; -- 0.11369207508592558
	pesos_i(9380) := b"0000000000000000_0000000000000000_0001110011001000_1111100011011110"; -- 0.11244159137363105
	pesos_i(9381) := b"1111111111111111_1111111111111111_1111010110111100_1010000010001011"; -- -0.040090528452462124
	pesos_i(9382) := b"1111111111111111_1111111111111111_1111010101101100_1001110101010010"; -- -0.04131142386756984
	pesos_i(9383) := b"0000000000000000_0000000000000000_0010000011110100_0001000011111110"; -- 0.12872415728852493
	pesos_i(9384) := b"0000000000000000_0000000000000000_0001001011101010_0011100101011110"; -- 0.07388647590089416
	pesos_i(9385) := b"0000000000000000_0000000000000000_0001001011100001_0110010100000101"; -- 0.07375174877204337
	pesos_i(9386) := b"0000000000000000_0000000000000000_0000010111100011_0000011111110011"; -- 0.022995469002945162
	pesos_i(9387) := b"1111111111111111_1111111111111111_1101101111001001_1001100110110001"; -- -0.14145507274161515
	pesos_i(9388) := b"1111111111111111_1111111111111111_1110011101001111_1011111010010011"; -- -0.09643944656014725
	pesos_i(9389) := b"1111111111111111_1111111111111111_1111000110010010_0100000000110100"; -- -0.05636213994767945
	pesos_i(9390) := b"1111111111111111_1111111111111111_1110011101111101_1010101110000010"; -- -0.09573867876190066
	pesos_i(9391) := b"1111111111111111_1111111111111111_1110000000001000_0111101100100010"; -- -0.12487059043843828
	pesos_i(9392) := b"0000000000000000_0000000000000000_0001101100101100_0001010110000001"; -- 0.10614141844428777
	pesos_i(9393) := b"1111111111111111_1111111111111111_1110000011001010_0100101000001001"; -- -0.12191331169265258
	pesos_i(9394) := b"0000000000000000_0000000000000000_0000001000111100_1101100011000001"; -- 0.008740946935023168
	pesos_i(9395) := b"1111111111111111_1111111111111111_1110111011000100_0111010101111010"; -- -0.06731477517819458
	pesos_i(9396) := b"1111111111111111_1111111111111111_1111001011101110_1101110110101101"; -- -0.05104269519596204
	pesos_i(9397) := b"1111111111111111_1111111111111111_1111001000001111_0110110010101000"; -- -0.05445214166554775
	pesos_i(9398) := b"0000000000000000_0000000000000000_0001001011110101_0001111010100000"; -- 0.07405272875660635
	pesos_i(9399) := b"1111111111111111_1111111111111111_1101111001011100_0100010111011100"; -- -0.1314045274850938
	pesos_i(9400) := b"1111111111111111_1111111111111111_1111011010010010_0001111000000000"; -- -0.0368329285596192
	pesos_i(9401) := b"1111111111111111_1111111111111111_1110011011100111_0110011100001010"; -- -0.09803157810690023
	pesos_i(9402) := b"0000000000000000_0000000000000000_0000001000011001_1101001110011111"; -- 0.008206583427770487
	pesos_i(9403) := b"0000000000000000_0000000000000000_0000100001010101_1101000110010111"; -- 0.03255948966890024
	pesos_i(9404) := b"0000000000000000_0000000000000000_0000011111001100_0101100101110000"; -- 0.030461873807215958
	pesos_i(9405) := b"0000000000000000_0000000000000000_0000110010110011_0101011111001100"; -- 0.04961155635317203
	pesos_i(9406) := b"0000000000000000_0000000000000000_0001000000111000_1110100110110100"; -- 0.06336842198207941
	pesos_i(9407) := b"0000000000000000_0000000000000000_0000001011000111_0011111110010110"; -- 0.010852789099973463
	pesos_i(9408) := b"0000000000000000_0000000000000000_0010010011001101_0001101100001111"; -- 0.14375466461590636
	pesos_i(9409) := b"1111111111111111_1111111111111111_1110001001000111_0111011100000110"; -- -0.11609703168949749
	pesos_i(9410) := b"0000000000000000_0000000000000000_0001011001011010_0101100001101100"; -- 0.08731606145131439
	pesos_i(9411) := b"1111111111111111_1111111111111111_1101100110100010_1001010100001110"; -- -0.14986294172714193
	pesos_i(9412) := b"0000000000000000_0000000000000000_0001111100001000_0011101000101010"; -- 0.121219287148956
	pesos_i(9413) := b"1111111111111111_1111111111111111_1111110000110001_0010111111001010"; -- -0.01487447090804459
	pesos_i(9414) := b"0000000000000000_0000000000000000_0001011010101000_0000101101111110"; -- 0.08850166163375052
	pesos_i(9415) := b"0000000000000000_0000000000000000_0001010010110111_0100110011011011"; -- 0.08092193923484221
	pesos_i(9416) := b"0000000000000000_0000000000000000_0000110101011110_1000011001110001"; -- 0.052223589470130956
	pesos_i(9417) := b"1111111111111111_1111111111111111_1101100001000101_0100110100011011"; -- -0.15519254769921562
	pesos_i(9418) := b"0000000000000000_0000000000000000_0010011011010100_0001010100001100"; -- 0.15167361782980324
	pesos_i(9419) := b"0000000000000000_0000000000000000_0010010000100011_0111001010101100"; -- 0.14116589251225048
	pesos_i(9420) := b"1111111111111111_1111111111111111_1111110011011100_1010110100011001"; -- -0.012257749003646764
	pesos_i(9421) := b"0000000000000000_0000000000000000_0000100110010100_0101101001100001"; -- 0.037419937890770597
	pesos_i(9422) := b"1111111111111111_1111111111111111_1111000011000111_0010001100010100"; -- -0.05946141014817458
	pesos_i(9423) := b"0000000000000000_0000000000000000_0001101110101000_1001101101111110"; -- 0.10804149454073382
	pesos_i(9424) := b"1111111111111111_1111111111111111_1101101100000100_1010100111101100"; -- -0.1444600867798049
	pesos_i(9425) := b"0000000000000000_0000000000000000_0000000111011110_0110000011111110"; -- 0.007299482310393646
	pesos_i(9426) := b"0000000000000000_0000000000000000_0001101111001101_1010010110101110"; -- 0.10860667703732393
	pesos_i(9427) := b"1111111111111111_1111111111111111_1111110101101010_1110011100011001"; -- -0.010087543761545435
	pesos_i(9428) := b"0000000000000000_0000000000000000_0001011110001011_0110100011000101"; -- 0.0919709665123758
	pesos_i(9429) := b"1111111111111111_1111111111111111_1110010010000001_1000010101101101"; -- -0.10739866348987404
	pesos_i(9430) := b"1111111111111111_1111111111111111_1101101100111001_0100010010010000"; -- -0.14365741237611004
	pesos_i(9431) := b"0000000000000000_0000000000000000_0001101001110100_1110111111100011"; -- 0.1033468179066035
	pesos_i(9432) := b"1111111111111111_1111111111111111_1111011111100100_1000000011110110"; -- -0.03166955938873753
	pesos_i(9433) := b"1111111111111111_1111111111111111_1110001101111111_0011111100100101"; -- -0.11133962017602271
	pesos_i(9434) := b"1111111111111111_1111111111111111_1111100111100111_1110001010010111"; -- -0.023805463815529598
	pesos_i(9435) := b"0000000000000000_0000000000000000_0001000010010000_0111000011101011"; -- 0.06470399607995779
	pesos_i(9436) := b"0000000000000000_0000000000000000_0010001110010000_1001111011010101"; -- 0.1389254827142972
	pesos_i(9437) := b"0000000000000000_0000000000000000_0000011011010111_0110101111100100"; -- 0.026724570394460787
	pesos_i(9438) := b"0000000000000000_0000000000000000_0000001111111001_0100010110110001"; -- 0.01552234244114675
	pesos_i(9439) := b"1111111111111111_1111111111111111_1101111100001000_0100001101010100"; -- -0.12878016668576986
	pesos_i(9440) := b"1111111111111111_1111111111111111_1101100001011011_1101000100010110"; -- -0.1548489876056893
	pesos_i(9441) := b"1111111111111111_1111111111111111_1110100101100000_0001001101101011"; -- -0.08837774889708279
	pesos_i(9442) := b"1111111111111111_1111111111111111_1111011111110011_0000000000110111"; -- -0.03144835147413223
	pesos_i(9443) := b"0000000000000000_0000000000000000_0000111110111001_0111111000000110"; -- 0.06142413752282814
	pesos_i(9444) := b"1111111111111111_1111111111111111_1110111101100101_0010001001100111"; -- -0.0648630617729179
	pesos_i(9445) := b"0000000000000000_0000000000000000_0000001111011110_1100100100000010"; -- 0.015118182194452745
	pesos_i(9446) := b"1111111111111111_1111111111111111_1110110010100010_0110000111110000"; -- -0.0756472387565443
	pesos_i(9447) := b"0000000000000000_0000000000000000_0001011110011000_0011111011111100"; -- 0.09216684010993728
	pesos_i(9448) := b"0000000000000000_0000000000000000_0000000100110010_0100100111101011"; -- 0.0046735953645603975
	pesos_i(9449) := b"0000000000000000_0000000000000000_0000001111000000_1111101000000101"; -- 0.014663339817690876
	pesos_i(9450) := b"0000000000000000_0000000000000000_0000110110011110_1101100010100110"; -- 0.05320505198153192
	pesos_i(9451) := b"0000000000000000_0000000000000000_0000001000000010_0010011100111100"; -- 0.007845356087534257
	pesos_i(9452) := b"0000000000000000_0000000000000000_0000111000010110_1001011010011010"; -- 0.05503216999376179
	pesos_i(9453) := b"1111111111111111_1111111111111111_1110110011011001_0011001111110001"; -- -0.07481074678611767
	pesos_i(9454) := b"0000000000000000_0000000000000000_0001011110100100_1110011001000010"; -- 0.09235991576374981
	pesos_i(9455) := b"1111111111111111_1111111111111111_1101110110001110_0101100001110100"; -- -0.13454672964585032
	pesos_i(9456) := b"0000000000000000_0000000000000000_0000011000110001_1011011001010101"; -- 0.02419604838462731
	pesos_i(9457) := b"0000000000000000_0000000000000000_0010000101110001_0010011000000111"; -- 0.13063275983942182
	pesos_i(9458) := b"1111111111111111_1111111111111111_1111001011010101_1101100001101010"; -- -0.051424478559712515
	pesos_i(9459) := b"0000000000000000_0000000000000000_0010011100101100_0111010110011001"; -- 0.15302214607679074
	pesos_i(9460) := b"0000000000000000_0000000000000000_0000000001011010_1110100011111000"; -- 0.0013871769418726636
	pesos_i(9461) := b"0000000000000000_0000000000000000_0000110001011011_0110101001110001"; -- 0.048269894119997915
	pesos_i(9462) := b"1111111111111111_1111111111111111_1111000011010111_0110100011101011"; -- -0.05921310667131582
	pesos_i(9463) := b"1111111111111111_1111111111111111_1111010010010011_0000010111011001"; -- -0.04463160934930337
	pesos_i(9464) := b"0000000000000000_0000000000000000_0010000010111101_0000101010111100"; -- 0.12788455089598907
	pesos_i(9465) := b"1111111111111111_1111111111111111_1111010100101010_1100101110001101"; -- -0.042315748211048027
	pesos_i(9466) := b"0000000000000000_0000000000000000_0000101110011000_1100101110010010"; -- 0.045300219616926124
	pesos_i(9467) := b"0000000000000000_0000000000000000_0010000000111001_1101001110001001"; -- 0.12588235951370513
	pesos_i(9468) := b"0000000000000000_0000000000000000_0010001001100010_0001111101101100"; -- 0.13430973422226908
	pesos_i(9469) := b"1111111111111111_1111111111111111_1111001100101100_0110011101111101"; -- -0.050103694825784056
	pesos_i(9470) := b"0000000000000000_0000000000000000_0000111011001010_0100111101110111"; -- 0.057774511975338214
	pesos_i(9471) := b"1111111111111111_1111111111111111_1111101011111011_1111100011011000"; -- -0.01959271177474737
	pesos_i(9472) := b"1111111111111111_1111111111111111_1101100011100010_1001001000101001"; -- -0.15279280188920058
	pesos_i(9473) := b"0000000000000000_0000000000000000_0001010001101100_0100011011101111"; -- 0.07977717730453415
	pesos_i(9474) := b"0000000000000000_0000000000000000_0001101011111110_1000111000111111"; -- 0.10544671092981595
	pesos_i(9475) := b"0000000000000000_0000000000000000_0001001101010000_1001100011001010"; -- 0.07544856009402764
	pesos_i(9476) := b"0000000000000000_0000000000000000_0010011001001101_1110000001101100"; -- 0.14962580344562854
	pesos_i(9477) := b"1111111111111111_1111111111111111_1111000111110010_0010011010000000"; -- -0.05489882838308068
	pesos_i(9478) := b"1111111111111111_1111111111111111_1111000001100000_0000101001101010"; -- -0.06103453547218017
	pesos_i(9479) := b"1111111111111111_1111111111111111_1101100100111011_1101100001101110"; -- -0.15143058127911307
	pesos_i(9480) := b"1111111111111111_1111111111111111_1110000000101110_1100111110011101"; -- -0.12428572095752473
	pesos_i(9481) := b"1111111111111111_1111111111111111_1111111000010011_0101100101000101"; -- -0.007517262129186391
	pesos_i(9482) := b"0000000000000000_0000000000000000_0010001011000000_0011001001010011"; -- 0.13574518695740903
	pesos_i(9483) := b"0000000000000000_0000000000000000_0010010101000110_0011011010001000"; -- 0.14560261550872358
	pesos_i(9484) := b"1111111111111111_1111111111111111_1110011001001100_1001100010101110"; -- -0.10039373160294297
	pesos_i(9485) := b"1111111111111111_1111111111111111_1101111100101001_1100010111011010"; -- -0.12826884677841635
	pesos_i(9486) := b"0000000000000000_0000000000000000_0000100010011010_0010100110011011"; -- 0.033602333471143324
	pesos_i(9487) := b"1111111111111111_1111111111111111_1111010111001011_1100101010110001"; -- -0.039859134381058724
	pesos_i(9488) := b"1111111111111111_1111111111111111_1110110101001100_1111100100010011"; -- -0.07304423610740182
	pesos_i(9489) := b"1111111111111111_1111111111111111_1111100000000010_1001011100011001"; -- -0.03121047619355062
	pesos_i(9490) := b"1111111111111111_1111111111111111_1111011000110110_0010100010000000"; -- -0.038236111518611574
	pesos_i(9491) := b"1111111111111111_1111111111111111_1111111011000000_0000111111111110"; -- -0.004881859217634917
	pesos_i(9492) := b"1111111111111111_1111111111111111_1110001110101101_0111111001110011"; -- -0.11063394264531448
	pesos_i(9493) := b"0000000000000000_0000000000000000_0001101111111001_1100001101110000"; -- 0.10927983735766558
	pesos_i(9494) := b"0000000000000000_0000000000000000_0000011010110011_0111111100011100"; -- 0.026176399459042154
	pesos_i(9495) := b"0000000000000000_0000000000000000_0001000100110101_1000100011010111"; -- 0.06722312207199035
	pesos_i(9496) := b"0000000000000000_0000000000000000_0000001010100101_0011001110001101"; -- 0.010333272886531492
	pesos_i(9497) := b"1111111111111111_1111111111111111_1101110010000011_0101000110101000"; -- -0.13862123142602462
	pesos_i(9498) := b"1111111111111111_1111111111111111_1101100111111101_1001100111101000"; -- -0.14847410295166347
	pesos_i(9499) := b"1111111111111111_1111111111111111_1101110101000110_0000101011110100"; -- -0.1356499819623321
	pesos_i(9500) := b"1111111111111111_1111111111111111_1101111111110011_0010001101001001"; -- -0.12519626120773164
	pesos_i(9501) := b"0000000000000000_0000000000000000_0000111000001010_0001001001000010"; -- 0.05484117603688321
	pesos_i(9502) := b"1111111111111111_1111111111111111_1101100101100111_0001001111110000"; -- -0.15077090627718068
	pesos_i(9503) := b"1111111111111111_1111111111111111_1111111010111100_0000010101001010"; -- -0.0049435324469334
	pesos_i(9504) := b"1111111111111111_1111111111111111_1111001110101110_0000000101100100"; -- -0.048126137763013464
	pesos_i(9505) := b"1111111111111111_1111111111111111_1101110000010101_0101000110110001"; -- -0.14029969619961494
	pesos_i(9506) := b"1111111111111111_1111111111111111_1111001011011011_0001110000011000"; -- -0.05134415077860957
	pesos_i(9507) := b"1111111111111111_1111111111111111_1110001011110100_0110110111001001"; -- -0.11345781174415584
	pesos_i(9508) := b"1111111111111111_1111111111111111_1111011000100111_1001111000001101"; -- -0.03845798670247453
	pesos_i(9509) := b"1111111111111111_1111111111111111_1111100010001011_0111110100011110"; -- -0.029121570775384947
	pesos_i(9510) := b"1111111111111111_1111111111111111_1110111110001100_0001011101100011"; -- -0.06426862560860583
	pesos_i(9511) := b"1111111111111111_1111111111111111_1110111001110100_1101000001100011"; -- -0.06853005966191951
	pesos_i(9512) := b"1111111111111111_1111111111111111_1110111100100110_1010010000110110"; -- -0.06581662820675704
	pesos_i(9513) := b"1111111111111111_1111111111111111_1110101111111111_0011011011000010"; -- -0.07813699490261239
	pesos_i(9514) := b"0000000000000000_0000000000000000_0001011111100011_0011111100011110"; -- 0.09331125716489204
	pesos_i(9515) := b"0000000000000000_0000000000000000_0001111101100111_0100100100101010"; -- 0.12266976611246053
	pesos_i(9516) := b"0000000000000000_0000000000000000_0001110011000001_1001101001111111"; -- 0.11232915488331079
	pesos_i(9517) := b"0000000000000000_0000000000000000_0000100011010100_0011001100011111"; -- 0.03448791034058911
	pesos_i(9518) := b"1111111111111111_1111111111111111_1110101000100011_0011111110111010"; -- -0.08539964393067412
	pesos_i(9519) := b"1111111111111111_1111111111111111_1111000110001001_1010010110101001"; -- -0.056493421782893044
	pesos_i(9520) := b"1111111111111111_1111111111111111_1111010101111101_1111010000111001"; -- -0.04104684463268067
	pesos_i(9521) := b"0000000000000000_0000000000000000_0000111100101001_1101100000111000"; -- 0.059232248084210785
	pesos_i(9522) := b"1111111111111111_1111111111111111_1110011011001110_0000101011001010"; -- -0.09841854627769984
	pesos_i(9523) := b"1111111111111111_1111111111111111_1110101001101110_1100100101010111"; -- -0.08424703232866433
	pesos_i(9524) := b"0000000000000000_0000000000000000_0001000011000000_0010100010010011"; -- 0.06543210581754752
	pesos_i(9525) := b"0000000000000000_0000000000000000_0000010110111101_0101001011011110"; -- 0.022420100511876453
	pesos_i(9526) := b"0000000000000000_0000000000000000_0000011001001100_0011001011100001"; -- 0.02460020047347951
	pesos_i(9527) := b"0000000000000000_0000000000000000_0001100100010100_1010011010000101"; -- 0.09797135111053075
	pesos_i(9528) := b"1111111111111111_1111111111111111_1101110111000010_0111010001100000"; -- -0.13375160833395947
	pesos_i(9529) := b"0000000000000000_0000000000000000_0010000001101001_1000101111101111"; -- 0.12661051349780297
	pesos_i(9530) := b"0000000000000000_0000000000000000_0000010001001011_1111101110000101"; -- 0.016784400861463475
	pesos_i(9531) := b"1111111111111111_1111111111111111_1110100100011100_0001011101001010"; -- -0.08941511586108654
	pesos_i(9532) := b"0000000000000000_0000000000000000_0000100101110100_1011111101100011"; -- 0.03693767715523151
	pesos_i(9533) := b"1111111111111111_1111111111111111_1110011110111011_0100000101100010"; -- -0.09479895933504826
	pesos_i(9534) := b"1111111111111111_1111111111111111_1101110010000010_0000110000100000"; -- -0.13864063479858743
	pesos_i(9535) := b"0000000000000000_0000000000000000_0001100010011111_0111110000001110"; -- 0.09618354177741824
	pesos_i(9536) := b"0000000000000000_0000000000000000_0000110001000001_0110011011000100"; -- 0.04787294650708712
	pesos_i(9537) := b"1111111111111111_1111111111111111_1111010001010100_0000011111011100"; -- -0.045592793187558815
	pesos_i(9538) := b"0000000000000000_0000000000000000_0001111101100010_1000000000111001"; -- 0.12259675406801576
	pesos_i(9539) := b"1111111111111111_1111111111111111_1111010010100101_0100010101000000"; -- -0.04435317227220056
	pesos_i(9540) := b"0000000000000000_0000000000000000_0000010001000011_0000110000110111"; -- 0.01664806699129967
	pesos_i(9541) := b"0000000000000000_0000000000000000_0001101010000011_0001110001000100"; -- 0.10356308608130785
	pesos_i(9542) := b"1111111111111111_1111111111111111_1111000100111001_1011111101010010"; -- -0.05771259540868793
	pesos_i(9543) := b"0000000000000000_0000000000000000_0000010110010010_0001100010001000"; -- 0.021760495493715653
	pesos_i(9544) := b"0000000000000000_0000000000000000_0000011000000100_0101000000001101"; -- 0.023503306475377548
	pesos_i(9545) := b"1111111111111111_1111111111111111_1111110100100011_1011110010010110"; -- -0.011173451739665918
	pesos_i(9546) := b"1111111111111111_1111111111111111_1110110101111000_0010100001011011"; -- -0.07238528999093292
	pesos_i(9547) := b"1111111111111111_1111111111111111_1110000011111100_1110011101101010"; -- -0.12114099174130989
	pesos_i(9548) := b"1111111111111111_1111111111111111_1110101000000110_0110000110100101"; -- -0.08584012727125431
	pesos_i(9549) := b"0000000000000000_0000000000000000_0010001000100110_0010100011110000"; -- 0.1333947741555945
	pesos_i(9550) := b"0000000000000000_0000000000000000_0001001000111010_1100011111110000"; -- 0.07120942685767742
	pesos_i(9551) := b"1111111111111111_1111111111111111_1110100101101101_0010001110111011"; -- -0.08817841236137894
	pesos_i(9552) := b"0000000000000000_0000000000000000_0000001000111011_0000111100100011"; -- 0.00871367087702605
	pesos_i(9553) := b"0000000000000000_0000000000000000_0010010010011011_1100000101011000"; -- 0.14300163638425709
	pesos_i(9554) := b"0000000000000000_0000000000000000_0010010010110000_0110010000111000"; -- 0.14331652036201023
	pesos_i(9555) := b"1111111111111111_1111111111111111_1101100100000010_0010000101010101"; -- -0.15231124559679685
	pesos_i(9556) := b"0000000000000000_0000000000000000_0001110100010001_1010011011001100"; -- 0.11355059132525551
	pesos_i(9557) := b"1111111111111111_1111111111111111_1110100000111011_1111101000111001"; -- -0.09283481699008718
	pesos_i(9558) := b"0000000000000000_0000000000000000_0000101111001100_1111010011011011"; -- 0.046096137531112524
	pesos_i(9559) := b"0000000000000000_0000000000000000_0000100110110101_1001010101100001"; -- 0.03792699453712551
	pesos_i(9560) := b"0000000000000000_0000000000000000_0010100010001110_0000100000011010"; -- 0.15841723088048892
	pesos_i(9561) := b"1111111111111111_1111111111111111_1111101011100010_0010011011111011"; -- -0.01998669031643817
	pesos_i(9562) := b"1111111111111111_1111111111111111_1101110100100110_1000100011111011"; -- -0.13613075123522042
	pesos_i(9563) := b"0000000000000000_0000000000000000_0000010010000110_1010011001111101"; -- 0.01767960115084338
	pesos_i(9564) := b"0000000000000000_0000000000000000_0001111111110001_0010000110110001"; -- 0.12477312629031646
	pesos_i(9565) := b"1111111111111111_1111111111111111_1110000111101001_0110100111001100"; -- -0.11753214606816563
	pesos_i(9566) := b"1111111111111111_1111111111111111_1110011000010000_0010011100101000"; -- -0.10131602556401023
	pesos_i(9567) := b"1111111111111111_1111111111111111_1111010000001000_1010111110000010"; -- -0.04674246849904162
	pesos_i(9568) := b"1111111111111111_1111111111111111_1111000111100101_0000101001000010"; -- -0.05509887586561322
	pesos_i(9569) := b"0000000000000000_0000000000000000_0000111110101100_0011110000100100"; -- 0.06122184638527197
	pesos_i(9570) := b"0000000000000000_0000000000000000_0000011101010101_1111100111110100"; -- 0.028655645373501237
	pesos_i(9571) := b"1111111111111111_1111111111111111_1110101000111010_1011010101011011"; -- -0.08504168052823424
	pesos_i(9572) := b"1111111111111111_1111111111111111_1110101100001110_0011010100111101"; -- -0.08181445370783201
	pesos_i(9573) := b"1111111111111111_1111111111111111_1110111101100010_1100010111001111"; -- -0.06489909826795905
	pesos_i(9574) := b"0000000000000000_0000000000000000_0000110011000011_1011101000111001"; -- 0.04986156361082219
	pesos_i(9575) := b"1111111111111111_1111111111111111_1111000001110000_0101100001011101"; -- -0.060785748861273685
	pesos_i(9576) := b"1111111111111111_1111111111111111_1101111100001000_0101110101111011"; -- -0.1287786077075477
	pesos_i(9577) := b"1111111111111111_1111111111111111_1111110101100110_0010001010101000"; -- -0.010160287900093408
	pesos_i(9578) := b"0000000000000000_0000000000000000_0010011000000011_1001001100100101"; -- 0.14849204695289442
	pesos_i(9579) := b"1111111111111111_1111111111111111_1111001100001100_1001110110001110"; -- -0.05058875344204849
	pesos_i(9580) := b"0000000000000000_0000000000000000_0001001000111000_0100011000010011"; -- 0.07117116904803394
	pesos_i(9581) := b"0000000000000000_0000000000000000_0001101001100111_0000000010001000"; -- 0.10313418697626336
	pesos_i(9582) := b"1111111111111111_1111111111111111_1111101010110101_0001100110110110"; -- -0.02067412657833122
	pesos_i(9583) := b"1111111111111111_1111111111111111_1111001011100111_1110111011000011"; -- -0.05114848845009457
	pesos_i(9584) := b"0000000000000000_0000000000000000_0000000001011110_1111011001100101"; -- 0.0014490125092394641
	pesos_i(9585) := b"0000000000000000_0000000000000000_0001100010101011_0010001100100110"; -- 0.09636134798380515
	pesos_i(9586) := b"1111111111111111_1111111111111111_1111000101010111_0111000100010011"; -- -0.05725949548775073
	pesos_i(9587) := b"0000000000000000_0000000000000000_0010000101110010_0100000010001001"; -- 0.13064959861551728
	pesos_i(9588) := b"1111111111111111_1111111111111111_1111101111010110_1110011000011011"; -- -0.016252153702572148
	pesos_i(9589) := b"0000000000000000_0000000000000000_0010000011111010_1010101100100011"; -- 0.12882489791178658
	pesos_i(9590) := b"1111111111111111_1111111111111111_1111000010100100_0110100110111000"; -- -0.05999125733955273
	pesos_i(9591) := b"0000000000000000_0000000000000000_0000101110111110_0000110010101010"; -- 0.045868674668622315
	pesos_i(9592) := b"1111111111111111_1111111111111111_1111101010001001_0010101000001110"; -- -0.02134453927792225
	pesos_i(9593) := b"0000000000000000_0000000000000000_0000110100110100_1010101110100000"; -- 0.05158493660983307
	pesos_i(9594) := b"0000000000000000_0000000000000000_0001100001111001_0000010101011000"; -- 0.09559663199535041
	pesos_i(9595) := b"1111111111111111_1111111111111111_1111000000000000_0111010111010110"; -- -0.06249297643144796
	pesos_i(9596) := b"0000000000000000_0000000000000000_0001101100100111_0010101100011100"; -- 0.1060664122838777
	pesos_i(9597) := b"1111111111111111_1111111111111111_1110110001000000_0111111110000111"; -- -0.07714083632657372
	pesos_i(9598) := b"1111111111111111_1111111111111111_1110111111000001_0101111000010001"; -- -0.06345569692540544
	pesos_i(9599) := b"0000000000000000_0000000000000000_0000011101101101_0000000110000110"; -- 0.029007048872423245
	pesos_i(9600) := b"1111111111111111_1111111111111111_1110111100001101_1111011100111010"; -- -0.06619314993509086
	pesos_i(9601) := b"0000000000000000_0000000000000000_0001110001010100_0000110111100110"; -- 0.1106575665884918
	pesos_i(9602) := b"1111111111111111_1111111111111111_1110101001000001_0100001011010101"; -- -0.08494169525014819
	pesos_i(9603) := b"1111111111111111_1111111111111111_1101110001111011_0011011001100110"; -- -0.138744926466591
	pesos_i(9604) := b"1111111111111111_1111111111111111_1101110010110001_0011011101010000"; -- -0.1379208974257565
	pesos_i(9605) := b"0000000000000000_0000000000000000_0001110010111001_0111011011100010"; -- 0.11220496183551674
	pesos_i(9606) := b"0000000000000000_0000000000000000_0000011000100001_1111110001101010"; -- 0.023956085085595644
	pesos_i(9607) := b"1111111111111111_1111111111111111_1110000100110000_1111000011001010"; -- -0.12034697593218124
	pesos_i(9608) := b"1111111111111111_1111111111111111_1110000101111000_0111101001001111"; -- -0.11925540522491518
	pesos_i(9609) := b"0000000000000000_0000000000000000_0000010110111110_1110111011011100"; -- 0.022444657081122452
	pesos_i(9610) := b"0000000000000000_0000000000000000_0010011011110100_1110101100100010"; -- 0.1521746594459174
	pesos_i(9611) := b"0000000000000000_0000000000000000_0000011010001101_1100101001001001"; -- 0.025601046441151805
	pesos_i(9612) := b"1111111111111111_1111111111111111_1110010011101010_1100000001110101"; -- -0.10579297194033328
	pesos_i(9613) := b"0000000000000000_0000000000000000_0000110011100101_0000011100000111"; -- 0.050369681607091946
	pesos_i(9614) := b"1111111111111111_1111111111111111_1111010101111011_1010011000110111"; -- -0.04108201166390185
	pesos_i(9615) := b"1111111111111111_1111111111111111_1110011111001001_1010010111011101"; -- -0.09457934726166925
	pesos_i(9616) := b"0000000000000000_0000000000000000_0001101011100101_1101111001000110"; -- 0.10507001126573298
	pesos_i(9617) := b"1111111111111111_1111111111111111_1110000110001100_1011110011101111"; -- -0.1189462582419126
	pesos_i(9618) := b"0000000000000000_0000000000000000_0000100011010001_1011101011110110"; -- 0.034450230625628644
	pesos_i(9619) := b"0000000000000000_0000000000000000_0001011110010111_1111111100000010"; -- 0.09216302684902923
	pesos_i(9620) := b"0000000000000000_0000000000000000_0001010111011000_1000101111001010"; -- 0.08533548051813168
	pesos_i(9621) := b"1111111111111111_1111111111111111_1101101101110110_1010110000101011"; -- -0.14272045080563459
	pesos_i(9622) := b"1111111111111111_1111111111111111_1110100010011110_0100011011100101"; -- -0.09133488565772117
	pesos_i(9623) := b"1111111111111111_1111111111111111_1111100011001001_0010000000000010"; -- -0.02818107568732108
	pesos_i(9624) := b"0000000000000000_0000000000000000_0001110001110100_0001001101000101"; -- 0.11114616807999098
	pesos_i(9625) := b"0000000000000000_0000000000000000_0001001111101101_1100101110100011"; -- 0.07784722080490493
	pesos_i(9626) := b"1111111111111111_1111111111111111_1110000101100100_0110111001001101"; -- -0.11956129677092434
	pesos_i(9627) := b"1111111111111111_1111111111111111_1101100000001101_0010011010111010"; -- -0.15604932739210764
	pesos_i(9628) := b"1111111111111111_1111111111111111_1110101111000000_1100100000101000"; -- -0.07908963233381053
	pesos_i(9629) := b"0000000000000000_0000000000000000_0001110011011110_0000011001001100"; -- 0.11276282645734317
	pesos_i(9630) := b"1111111111111111_1111111111111111_1110000110000100_1000101100001111"; -- -0.11907130122521023
	pesos_i(9631) := b"0000000000000000_0000000000000000_0000100011101001_1100110110101001"; -- 0.034817556091820946
	pesos_i(9632) := b"1111111111111111_1111111111111111_1110111011100001_0010100101100001"; -- -0.066876806190498
	pesos_i(9633) := b"1111111111111111_1111111111111111_1101101110111000_0110000100110011"; -- -0.14171783926915918
	pesos_i(9634) := b"1111111111111111_1111111111111111_1110001010101011_0010000111100110"; -- -0.11457622664346795
	pesos_i(9635) := b"0000000000000000_0000000000000000_0000000001010111_1000110111111001"; -- 0.0013359768612435608
	pesos_i(9636) := b"1111111111111111_1111111111111111_1110001011100111_1111110110101111"; -- -0.1136475989426621
	pesos_i(9637) := b"1111111111111111_1111111111111111_1111011100010100_0000010101010011"; -- -0.03485075693116697
	pesos_i(9638) := b"1111111111111111_1111111111111111_1110101011100111_0000010011100110"; -- -0.08241242776957165
	pesos_i(9639) := b"1111111111111111_1111111111111111_1110010011101100_1100011000100011"; -- -0.10576211598081518
	pesos_i(9640) := b"0000000000000000_0000000000000000_0010101100110000_1000100101001111"; -- 0.1687093561859988
	pesos_i(9641) := b"0000000000000000_0000000000000000_0000010011000100_1100001000001010"; -- 0.01862728835291756
	pesos_i(9642) := b"1111111111111111_1111111111111111_1111110001100010_0011011000000101"; -- -0.014126418880553474
	pesos_i(9643) := b"0000000000000000_0000000000000000_0001100100010011_1110110101101101"; -- 0.09796031874221334
	pesos_i(9644) := b"1111111111111111_1111111111111111_1111010011001010_0101011000010101"; -- -0.043787593634891916
	pesos_i(9645) := b"0000000000000000_0000000000000000_0001110101100111_1001001110010100"; -- 0.11486170159085232
	pesos_i(9646) := b"0000000000000000_0000000000000000_0001100100100101_1111001101000111"; -- 0.09823532564565628
	pesos_i(9647) := b"0000000000000000_0000000000000000_0000001011101011_1010010111111101"; -- 0.011408209117654054
	pesos_i(9648) := b"0000000000000000_0000000000000000_0001000000111111_0011001101000100"; -- 0.06346435941430219
	pesos_i(9649) := b"0000000000000000_0000000000000000_0000001100000110_0111100111011010"; -- 0.011817565588680913
	pesos_i(9650) := b"1111111111111111_1111111111111111_1110011111100110_0101110111000010"; -- -0.0941411400161936
	pesos_i(9651) := b"0000000000000000_0000000000000000_0010100000110100_1101000011000101"; -- 0.1570559005988452
	pesos_i(9652) := b"1111111111111111_1111111111111111_1110010010010011_0101101101011000"; -- -0.10712651358800254
	pesos_i(9653) := b"0000000000000000_0000000000000000_0001101010001111_0010000001001101"; -- 0.1037464321048854
	pesos_i(9654) := b"0000000000000000_0000000000000000_0000100001011010_1000101000001000"; -- 0.03263151842408759
	pesos_i(9655) := b"0000000000000000_0000000000000000_0000110110001111_0100101001000011"; -- 0.05296768319020461
	pesos_i(9656) := b"1111111111111111_1111111111111111_1110101010011111_0011111100001110"; -- -0.08350759423498162
	pesos_i(9657) := b"1111111111111111_1111111111111111_1111111101111100_0100110100111010"; -- -0.0020095571279662755
	pesos_i(9658) := b"0000000000000000_0000000000000000_0001111000111001_1010010100001000"; -- 0.11806708753212722
	pesos_i(9659) := b"0000000000000000_0000000000000000_0001101110001100_1001010001011010"; -- 0.1076138229005371
	pesos_i(9660) := b"1111111111111111_1111111111111111_1111101101100010_0100000101110100"; -- -0.018031987463433242
	pesos_i(9661) := b"0000000000000000_0000000000000000_0000110101100110_0011001011100111"; -- 0.05234068040198608
	pesos_i(9662) := b"0000000000000000_0000000000000000_0001010010100001_0110111001011010"; -- 0.08058824240313592
	pesos_i(9663) := b"0000000000000000_0000000000000000_0000001000010011_0101110000111111"; -- 0.008107915172115943
	pesos_i(9664) := b"1111111111111111_1111111111111111_1111010101000001_1011001001010011"; -- -0.04196629983788774
	pesos_i(9665) := b"0000000000000000_0000000000000000_0000100101110011_1110100100100100"; -- 0.036924907022783324
	pesos_i(9666) := b"1111111111111111_1111111111111111_1111001101100001_1010001000011110"; -- -0.04929148442048887
	pesos_i(9667) := b"0000000000000000_0000000000000000_0001111011101000_1100010001111110"; -- 0.12073925091077685
	pesos_i(9668) := b"0000000000000000_0000000000000000_0000111100000011_0111000000100100"; -- 0.05864621045812514
	pesos_i(9669) := b"1111111111111111_1111111111111111_1110101111000011_0011110010110011"; -- -0.07905216823373035
	pesos_i(9670) := b"0000000000000000_0000000000000000_0010011010010011_1010000111001010"; -- 0.15069018542474694
	pesos_i(9671) := b"1111111111111111_1111111111111111_1101110111000010_1101010000101000"; -- -0.13374589939854886
	pesos_i(9672) := b"0000000000000000_0000000000000000_0001011100111001_0000010010101100"; -- 0.09071377955399554
	pesos_i(9673) := b"0000000000000000_0000000000000000_0000110100010000_1001010011001000"; -- 0.051034258686475896
	pesos_i(9674) := b"1111111111111111_1111111111111111_1110101010111110_0000000001110100"; -- -0.08303830302161515
	pesos_i(9675) := b"0000000000000000_0000000000000000_0000000101001001_0011101110001111"; -- 0.0050236916248315696
	pesos_i(9676) := b"1111111111111111_1111111111111111_1110111111010111_0010101001101001"; -- -0.06312308253714874
	pesos_i(9677) := b"0000000000000000_0000000000000000_0001111111011110_1011111010010100"; -- 0.12449256047612962
	pesos_i(9678) := b"1111111111111111_1111111111111111_1110000111000110_0110101001010010"; -- -0.11806617246697317
	pesos_i(9679) := b"1111111111111111_1111111111111111_1101110100101001_1011111010001011"; -- -0.13608178235798093
	pesos_i(9680) := b"0000000000000000_0000000000000000_0010000001011011_1101111000111100"; -- 0.12640179607398616
	pesos_i(9681) := b"1111111111111111_1111111111111111_1111100010010011_1100001011011110"; -- -0.02899534303305289
	pesos_i(9682) := b"0000000000000000_0000000000000000_0001010110001111_1011111010010000"; -- 0.08422461517336408
	pesos_i(9683) := b"0000000000000000_0000000000000000_0000100111101111_0000011100001101"; -- 0.03880352092339135
	pesos_i(9684) := b"0000000000000000_0000000000000000_0001101111000110_0000000000011001"; -- 0.10848999600665046
	pesos_i(9685) := b"1111111111111111_1111111111111111_1111000010010000_1010000001111110"; -- -0.06029316818075655
	pesos_i(9686) := b"0000000000000000_0000000000000000_0001011101000110_1001101101010011"; -- 0.09092112336992644
	pesos_i(9687) := b"1111111111111111_1111111111111111_1110011101111101_1010010011000110"; -- -0.09573908013314968
	pesos_i(9688) := b"0000000000000000_0000000000000000_0010100100010110_0011000100011100"; -- 0.16049487050992875
	pesos_i(9689) := b"1111111111111111_1111111111111111_1101110001000111_0010101011111001"; -- -0.13953906462953625
	pesos_i(9690) := b"1111111111111111_1111111111111111_1110001001101101_1011010101101011"; -- -0.11551347858024939
	pesos_i(9691) := b"0000000000000000_0000000000000000_0010000101011010_0000011111100110"; -- 0.13028001186826046
	pesos_i(9692) := b"0000000000000000_0000000000000000_0001001000011011_1100011110101011"; -- 0.07073638834211425
	pesos_i(9693) := b"1111111111111111_1111111111111111_1111010000010111_0011110011011101"; -- -0.04652042001858991
	pesos_i(9694) := b"1111111111111111_1111111111111111_1110101011101111_1001011010101111"; -- -0.08228166793229248
	pesos_i(9695) := b"1111111111111111_1111111111111111_1110000011110100_0011101010101100"; -- -0.12127335843500175
	pesos_i(9696) := b"0000000000000000_0000000000000000_0001011011111010_1100000011011001"; -- 0.08976369183830886
	pesos_i(9697) := b"0000000000000000_0000000000000000_0010001111000011_1100100001011000"; -- 0.1397061552739271
	pesos_i(9698) := b"0000000000000000_0000000000000000_0010000001010110_1010101001110011"; -- 0.1263224154153251
	pesos_i(9699) := b"1111111111111111_1111111111111111_1111000111100100_0001010110011111"; -- -0.05511345729596159
	pesos_i(9700) := b"1111111111111111_1111111111111111_1111110100100000_0101011100101111"; -- -0.011225272160923113
	pesos_i(9701) := b"0000000000000000_0000000000000000_0001001101110010_1100101101100110"; -- 0.0759703755217938
	pesos_i(9702) := b"0000000000000000_0000000000000000_0001100010000110_1010010100111100"; -- 0.09580452635714287
	pesos_i(9703) := b"1111111111111111_1111111111111111_1110110011101000_0010001000000101"; -- -0.0745829332195261
	pesos_i(9704) := b"1111111111111111_1111111111111111_1101110001001100_1111110000100101"; -- -0.13945030310883716
	pesos_i(9705) := b"0000000000000000_0000000000000000_0001001110101100_1011001000100111"; -- 0.07685388042820132
	pesos_i(9706) := b"0000000000000000_0000000000000000_0001101000000101_0011110000001100"; -- 0.10164237305995166
	pesos_i(9707) := b"0000000000000000_0000000000000000_0000011101001010_1011110100001101"; -- 0.02848416866263977
	pesos_i(9708) := b"1111111111111111_1111111111111111_1110110001101100_1101100001101011"; -- -0.07646415126559637
	pesos_i(9709) := b"1111111111111111_1111111111111111_1111110000100000_1111101111110011"; -- -0.015121701372598072
	pesos_i(9710) := b"0000000000000000_0000000000000000_0001111001110101_0110110100111001"; -- 0.11897928849866117
	pesos_i(9711) := b"0000000000000000_0000000000000000_0010001011110111_1001011100100010"; -- 0.13659042905516056
	pesos_i(9712) := b"1111111111111111_1111111111111111_1110011110000110_0001100000111011"; -- -0.09561012800367544
	pesos_i(9713) := b"1111111111111111_1111111111111111_1111100111010100_1000101110111101"; -- -0.02410055767393271
	pesos_i(9714) := b"1111111111111111_1111111111111111_1101111001100111_0100111011001111"; -- -0.13123614733418262
	pesos_i(9715) := b"1111111111111111_1111111111111111_1111111100111110_1000110110000001"; -- -0.002951770805952842
	pesos_i(9716) := b"1111111111111111_1111111111111111_1110111001010100_0100111110111100"; -- -0.06902600927791604
	pesos_i(9717) := b"1111111111111111_1111111111111111_1101111001111110_0011110011001010"; -- -0.13088626931454728
	pesos_i(9718) := b"1111111111111111_1111111111111111_1110100010101001_1101001010010101"; -- -0.0911587129395983
	pesos_i(9719) := b"0000000000000000_0000000000000000_0000101101110000_0100010011011000"; -- 0.04468183788106741
	pesos_i(9720) := b"1111111111111111_1111111111111111_1110101000101100_0001010011101110"; -- -0.085264865827523
	pesos_i(9721) := b"0000000000000000_0000000000000000_0001111000011101_0101110000101101"; -- 0.1176354990464451
	pesos_i(9722) := b"0000000000000000_0000000000000000_0010010100111001_0100100111101110"; -- 0.1454054075495321
	pesos_i(9723) := b"0000000000000000_0000000000000000_0000101111111001_1100110111001100"; -- 0.04678045493344439
	pesos_i(9724) := b"1111111111111111_1111111111111111_1111001110010101_1111010111110111"; -- -0.048493029818069584
	pesos_i(9725) := b"1111111111111111_1111111111111111_1110011010001100_1101011100101001"; -- -0.09941344498481026
	pesos_i(9726) := b"1111111111111111_1111111111111111_1110011110100010_1110101001000001"; -- -0.09517036343932181
	pesos_i(9727) := b"0000000000000000_0000000000000000_0000001010110010_0101001101111000"; -- 0.010533539511056367
	pesos_i(9728) := b"0000000000000000_0000000000000000_0001110111000001_0000101101010011"; -- 0.11622687115499503
	pesos_i(9729) := b"0000000000000000_0000000000000000_0000001100001010_1101000110011110"; -- 0.011883831969934621
	pesos_i(9730) := b"0000000000000000_0000000000000000_0001001100111011_1010101011000101"; -- 0.07512919709663701
	pesos_i(9731) := b"0000000000000000_0000000000000000_0010001011111001_0001100110001110"; -- 0.13661346158868046
	pesos_i(9732) := b"1111111111111111_1111111111111111_1101111110000100_1111010010100111"; -- -0.1268775073337974
	pesos_i(9733) := b"1111111111111111_1111111111111111_1110010100101111_1011101110111010"; -- -0.10474039751593525
	pesos_i(9734) := b"0000000000000000_0000000000000000_0001010100001100_0101011110110001"; -- 0.08221958239497605
	pesos_i(9735) := b"0000000000000000_0000000000000000_0000011011111110_0100110100111001"; -- 0.027317835337571306
	pesos_i(9736) := b"1111111111111111_1111111111111111_1101100100000110_1011001000110001"; -- -0.15224157633971397
	pesos_i(9737) := b"0000000000000000_0000000000000000_0000000011100011_0100101100011010"; -- 0.0034682214455683986
	pesos_i(9738) := b"1111111111111111_1111111111111111_1101010111010111_0001010011010101"; -- -0.1646868686094821
	pesos_i(9739) := b"0000000000000000_0000000000000000_0000000011100101_0010100000111011"; -- 0.0034966607206760357
	pesos_i(9740) := b"0000000000000000_0000000000000000_0001000000010010_1011011100000110"; -- 0.06278556728365438
	pesos_i(9741) := b"0000000000000000_0000000000000000_0001100101000000_1101110111111010"; -- 0.0986460432283175
	pesos_i(9742) := b"0000000000000000_0000000000000000_0010000010011001_1111010000110011"; -- 0.12734915017970327
	pesos_i(9743) := b"1111111111111111_1111111111111111_1110010000111001_1110101000100000"; -- -0.10849129403961412
	pesos_i(9744) := b"1111111111111111_1111111111111111_1111000001111111_0001001110100011"; -- -0.060560963285694276
	pesos_i(9745) := b"1111111111111111_1111111111111111_1111011110010101_1101011110000111"; -- -0.0328698440040894
	pesos_i(9746) := b"1111111111111111_1111111111111111_1111111110000111_0001100001010001"; -- -0.0018448640973103443
	pesos_i(9747) := b"1111111111111111_1111111111111111_1110111011111111_1100100011111000"; -- -0.06640953000629674
	pesos_i(9748) := b"1111111111111111_1111111111111111_1110101110110110_1011110100000000"; -- -0.07924288518700509
	pesos_i(9749) := b"1111111111111111_1111111111111111_1101111100111000_0000011011011010"; -- -0.12805134942603624
	pesos_i(9750) := b"1111111111111111_1111111111111111_1111100001000111_1000011101000001"; -- -0.03015856428690535
	pesos_i(9751) := b"0000000000000000_0000000000000000_0001111100110010_1010101001010010"; -- 0.12186684138070877
	pesos_i(9752) := b"1111111111111111_1111111111111111_1110010011111011_0100110000000111"; -- -0.10554051238866798
	pesos_i(9753) := b"1111111111111111_1111111111111111_1110100010011110_1001101100010100"; -- -0.0913298680510925
	pesos_i(9754) := b"0000000000000000_0000000000000000_0001011000011100_1000100010111000"; -- 0.08637289520195503
	pesos_i(9755) := b"1111111111111111_1111111111111111_1101111101100011_1000000101000110"; -- -0.12738792461051948
	pesos_i(9756) := b"1111111111111111_1111111111111111_1101101111010111_0010000101010100"; -- -0.14124862384881479
	pesos_i(9757) := b"1111111111111111_1111111111111111_1111101110100010_1100001101000010"; -- -0.01704768792358797
	pesos_i(9758) := b"0000000000000000_0000000000000000_0000111100000011_0110111100011011"; -- 0.05864614870303587
	pesos_i(9759) := b"0000000000000000_0000000000000000_0010001101101010_0001100011111110"; -- 0.1383376712977284
	pesos_i(9760) := b"1111111111111111_1111111111111111_1110000100100011_0000111001000110"; -- -0.12055884157106864
	pesos_i(9761) := b"0000000000000000_0000000000000000_0001000111000010_1010010011111101"; -- 0.06937628921033526
	pesos_i(9762) := b"0000000000000000_0000000000000000_0000010000010100_1000110100110011"; -- 0.0159385918643962
	pesos_i(9763) := b"0000000000000000_0000000000000000_0001101111110001_1001010000101010"; -- 0.10915494947742123
	pesos_i(9764) := b"1111111111111111_1111111111111111_1110010001001010_1111001110111111"; -- -0.10823132125875859
	pesos_i(9765) := b"1111111111111111_1111111111111111_1111111001011001_0010111011001110"; -- -0.006451678053399725
	pesos_i(9766) := b"0000000000000000_0000000000000000_0001001011001001_1011111010011100"; -- 0.07339087772578215
	pesos_i(9767) := b"0000000000000000_0000000000000000_0001010111000001_1111101000100100"; -- 0.08499110577916681
	pesos_i(9768) := b"1111111111111111_1111111111111111_1110100111001100_1010010000001011"; -- -0.08672117928525616
	pesos_i(9769) := b"0000000000000000_0000000000000000_0001100001010010_1100110000111011"; -- 0.09501339376331601
	pesos_i(9770) := b"0000000000000000_0000000000000000_0000101101001111_1110011101101001"; -- 0.044187987525531096
	pesos_i(9771) := b"1111111111111111_1111111111111111_1111001110010100_1101010100010001"; -- -0.04851024956521593
	pesos_i(9772) := b"1111111111111111_1111111111111111_1111011011000011_0100001101101111"; -- -0.03608301680298437
	pesos_i(9773) := b"1111111111111111_1111111111111111_1111101101011100_0010111100000100"; -- -0.018124639058305508
	pesos_i(9774) := b"1111111111111111_1111111111111111_1111100011111111_1101110001001101"; -- -0.02734587788722805
	pesos_i(9775) := b"1111111111111111_1111111111111111_1101111011110001_1100111010100100"; -- -0.12912281518893132
	pesos_i(9776) := b"1111111111111111_1111111111111111_1110011111000010_1001001100101010"; -- -0.094687273224736
	pesos_i(9777) := b"1111111111111111_1111111111111111_1110010010000010_0100010001101111"; -- -0.10738727855280074
	pesos_i(9778) := b"0000000000000000_0000000000000000_0000100010001100_0010111101001111"; -- 0.033389050216516676
	pesos_i(9779) := b"1111111111111111_1111111111111111_1110111101111010_1000011111010011"; -- -0.06453658195899159
	pesos_i(9780) := b"1111111111111111_1111111111111111_1111111101011101_1000001111110000"; -- -0.0024793185563947995
	pesos_i(9781) := b"0000000000000000_0000000000000000_0010011011000110_1110010101111100"; -- 0.15147241862754263
	pesos_i(9782) := b"0000000000000000_0000000000000000_0000101000100110_0111001010011001"; -- 0.039649164542497575
	pesos_i(9783) := b"0000000000000000_0000000000000000_0001111110010010_0110011101111101"; -- 0.12332770168931884
	pesos_i(9784) := b"1111111111111111_1111111111111111_1101111010010111_0101001110000100"; -- -0.13050344485663357
	pesos_i(9785) := b"1111111111111111_1111111111111111_1111000000000100_0111101110001001"; -- -0.0624316015108132
	pesos_i(9786) := b"1111111111111111_1111111111111111_1110001000000110_1010011100110010"; -- -0.11708598171195579
	pesos_i(9787) := b"1111111111111111_1111111111111111_1101011001100101_0001101110000100"; -- -0.16251972235413706
	pesos_i(9788) := b"0000000000000000_0000000000000000_0001101101100010_1000000110010001"; -- 0.10697183417805084
	pesos_i(9789) := b"0000000000000000_0000000000000000_0001110100001010_1011010111101010"; -- 0.1134446808711787
	pesos_i(9790) := b"1111111111111111_1111111111111111_1110011101110001_1101001100010010"; -- -0.09591942600844278
	pesos_i(9791) := b"1111111111111111_1111111111111111_1111101000001110_1000011101101100"; -- -0.0232158052489098
	pesos_i(9792) := b"1111111111111111_1111111111111111_1111010001110110_0000011110011111"; -- -0.045074008590342475
	pesos_i(9793) := b"0000000000000000_0000000000000000_0000010111001000_1101110101100010"; -- 0.022596203316352634
	pesos_i(9794) := b"1111111111111111_1111111111111111_1110010011011001_1100010010111100"; -- -0.10605211638459763
	pesos_i(9795) := b"0000000000000000_0000000000000000_0000000100001010_1010100000110011"; -- 0.004068863458998035
	pesos_i(9796) := b"0000000000000000_0000000000000000_0000110110010011_1101000100000101"; -- 0.053036750521463075
	pesos_i(9797) := b"1111111111111111_1111111111111111_1111010100011000_1001110001001011"; -- -0.04259322334009011
	pesos_i(9798) := b"1111111111111111_1111111111111111_1101101000001110_0000011001010000"; -- -0.14822350076931884
	pesos_i(9799) := b"1111111111111111_1111111111111111_1111111101001111_0100100000111000"; -- -0.0026965011679725213
	pesos_i(9800) := b"0000000000000000_0000000000000000_0001001000100100_1011001101001101"; -- 0.07087250367884419
	pesos_i(9801) := b"0000000000000000_0000000000000000_0001000011011000_1100010010100001"; -- 0.06580761835075273
	pesos_i(9802) := b"0000000000000000_0000000000000000_0001010000001111_1011110111100011"; -- 0.07836520006385185
	pesos_i(9803) := b"0000000000000000_0000000000000000_0000110100100010_1111110111111111"; -- 0.051315188205315415
	pesos_i(9804) := b"1111111111111111_1111111111111111_1111100001101100_1101111101110110"; -- -0.02958873150588399
	pesos_i(9805) := b"0000000000000000_0000000000000000_0001010100000010_0101111100111011"; -- 0.08206744372119
	pesos_i(9806) := b"1111111111111111_1111111111111111_1101111110010110_1111111111010011"; -- -0.12660218327973666
	pesos_i(9807) := b"0000000000000000_0000000000000000_0001100111011011_0101001111000010"; -- 0.1010029172695414
	pesos_i(9808) := b"0000000000000000_0000000000000000_0010001101110010_0111011101011111"; -- 0.13846536691007064
	pesos_i(9809) := b"0000000000000000_0000000000000000_0000000111111011_0011000011011001"; -- 0.007739117620298756
	pesos_i(9810) := b"0000000000000000_0000000000000000_0000001111001000_1010111111011010"; -- 0.014780989357690141
	pesos_i(9811) := b"0000000000000000_0000000000000000_0000000001110001_0101011000100000"; -- 0.001729376619021707
	pesos_i(9812) := b"0000000000000000_0000000000000000_0000101101101011_1100011011010001"; -- 0.04461329086243674
	pesos_i(9813) := b"0000000000000000_0000000000000000_0000011101011011_1011111111001100"; -- 0.02874373172223501
	pesos_i(9814) := b"1111111111111111_1111111111111111_1111011010011010_1110100101010001"; -- -0.036698739712447755
	pesos_i(9815) := b"0000000000000000_0000000000000000_0001111111110110_0001110100101110"; -- 0.1248491512449573
	pesos_i(9816) := b"1111111111111111_1111111111111111_1101011100011000_0101110101011110"; -- -0.1597844738756898
	pesos_i(9817) := b"1111111111111111_1111111111111111_1111000010100010_1000001010001110"; -- -0.06002029460150941
	pesos_i(9818) := b"1111111111111111_1111111111111111_1110100110110101_0111001111101000"; -- -0.08707500064783368
	pesos_i(9819) := b"0000000000000000_0000000000000000_0000000000011011_1101010110100110"; -- 0.0004247216425017143
	pesos_i(9820) := b"0000000000000000_0000000000000000_0000111001101001_0110110001011011"; -- 0.05629613135977985
	pesos_i(9821) := b"0000000000000000_0000000000000000_0001101011011011_1101111001011101"; -- 0.10491742857744205
	pesos_i(9822) := b"1111111111111111_1111111111111111_1110001001001101_0011011110111101"; -- -0.11600925096095348
	pesos_i(9823) := b"1111111111111111_1111111111111111_1101111101110001_0001000010100000"; -- -0.12718101587856478
	pesos_i(9824) := b"1111111111111111_1111111111111111_1101110011000010_1010010011000010"; -- -0.13765497456389847
	pesos_i(9825) := b"0000000000000000_0000000000000000_0001111101111000_1011000011001000"; -- 0.12293534164567844
	pesos_i(9826) := b"1111111111111111_1111111111111111_1111010010010101_1100011000010010"; -- -0.04458963455296387
	pesos_i(9827) := b"0000000000000000_0000000000000000_0001010100101111_0010101101100001"; -- 0.08275099865406349
	pesos_i(9828) := b"0000000000000000_0000000000000000_0000001100110010_0111111000000111"; -- 0.012489201212020542
	pesos_i(9829) := b"1111111111111111_1111111111111111_1111101001000100_0101010011010010"; -- -0.02239484662151052
	pesos_i(9830) := b"1111111111111111_1111111111111111_1101011110101100_0000111110111001"; -- -0.15753080113290294
	pesos_i(9831) := b"1111111111111111_1111111111111111_1111101101011001_1110110110001011"; -- -0.01815905907624878
	pesos_i(9832) := b"1111111111111111_1111111111111111_1111101010101101_0100100010011000"; -- -0.020793402622297886
	pesos_i(9833) := b"1111111111111111_1111111111111111_1110011111111000_0100101010011011"; -- -0.09386762345605976
	pesos_i(9834) := b"0000000000000000_0000000000000000_0001101111111010_0111100001100100"; -- 0.10929062301703099
	pesos_i(9835) := b"0000000000000000_0000000000000000_0001011100001010_1010111011000010"; -- 0.09000675415725201
	pesos_i(9836) := b"1111111111111111_1111111111111111_1111110101100110_0001001101011111"; -- -0.010161198872224487
	pesos_i(9837) := b"0000000000000000_0000000000000000_0000000011001110_0000011000010011"; -- 0.0031436725711171667
	pesos_i(9838) := b"0000000000000000_0000000000000000_0000100000010111_0110100001110010"; -- 0.03160717751551246
	pesos_i(9839) := b"0000000000000000_0000000000000000_0001100100101000_1111101000010100"; -- 0.09828150730632672
	pesos_i(9840) := b"1111111111111111_1111111111111111_1101111100000011_1100001110010001"; -- -0.12884881697696007
	pesos_i(9841) := b"0000000000000000_0000000000000000_0001101000010001_1100010110110001"; -- 0.1018336827208017
	pesos_i(9842) := b"0000000000000000_0000000000000000_0000001100110001_1010011010011000"; -- 0.012476360525727568
	pesos_i(9843) := b"0000000000000000_0000000000000000_0000101000100111_1110110101010011"; -- 0.039671738310776763
	pesos_i(9844) := b"0000000000000000_0000000000000000_0010000001100000_1111010010111100"; -- 0.12647943114399002
	pesos_i(9845) := b"0000000000000000_0000000000000000_0001111100101001_0000001010100101"; -- 0.12171951801320575
	pesos_i(9846) := b"0000000000000000_0000000000000000_0001010000101010_1001001010100110"; -- 0.07877460996440984
	pesos_i(9847) := b"1111111111111111_1111111111111111_1111110010001111_0010101010111110"; -- -0.013440445640658324
	pesos_i(9848) := b"1111111111111111_1111111111111111_1111101101100101_1111001100101111"; -- -0.017975617512858963
	pesos_i(9849) := b"0000000000000000_0000000000000000_0010000101101011_0110001001010001"; -- 0.13054480055147363
	pesos_i(9850) := b"0000000000000000_0000000000000000_0000101000010110_1100111110000100"; -- 0.03941056221628896
	pesos_i(9851) := b"0000000000000000_0000000000000000_0000101001000110_0001110000111010"; -- 0.04013229760751563
	pesos_i(9852) := b"0000000000000000_0000000000000000_0001101110110101_0011100100001011"; -- 0.10823399082092786
	pesos_i(9853) := b"1111111111111111_1111111111111111_1101110000110111_0111100101100000"; -- -0.1397785320940886
	pesos_i(9854) := b"1111111111111111_1111111111111111_1110100011100011_1001000110101110"; -- -0.09027757168681089
	pesos_i(9855) := b"1111111111111111_1111111111111111_1111101101000010_1100000110111011"; -- -0.01851262257847304
	pesos_i(9856) := b"0000000000000000_0000000000000000_0000110011110111_0001110101001001"; -- 0.050645666407551554
	pesos_i(9857) := b"0000000000000000_0000000000000000_0000010110110111_0110111100010010"; -- 0.022330228595024683
	pesos_i(9858) := b"1111111111111111_1111111111111111_1110010100011001_0010011000000100"; -- -0.10508501425897131
	pesos_i(9859) := b"0000000000000000_0000000000000000_0000111101001100_0110100100111000"; -- 0.05975968953236724
	pesos_i(9860) := b"0000000000000000_0000000000000000_0001111010000110_1101000101010101"; -- 0.11924465499728937
	pesos_i(9861) := b"0000000000000000_0000000000000000_0000000000001111_1101100110111110"; -- 0.00024186036387502982
	pesos_i(9862) := b"0000000000000000_0000000000000000_0000100010101000_1001000101010111"; -- 0.03382213944378023
	pesos_i(9863) := b"1111111111111111_1111111111111111_1110011110100100_0100110100011001"; -- -0.09514921328979827
	pesos_i(9864) := b"1111111111111111_1111111111111111_1110100101010110_1101101101110011"; -- -0.08851841396832925
	pesos_i(9865) := b"1111111111111111_1111111111111111_1101110111111011_0101110000110101"; -- -0.13288329794444176
	pesos_i(9866) := b"0000000000000000_0000000000000000_0010100010110010_1110100100011010"; -- 0.15897995848644886
	pesos_i(9867) := b"0000000000000000_0000000000000000_0000101100111110_1110011111010101"; -- 0.043928613089895964
	pesos_i(9868) := b"1111111111111111_1111111111111111_1110100100110010_0100011000111011"; -- -0.08907662455300117
	pesos_i(9869) := b"1111111111111111_1111111111111111_1110000001000001_1111001100111010"; -- -0.12399368130817082
	pesos_i(9870) := b"0000000000000000_0000000000000000_0010010011011010_1000111110101101"; -- 0.14395997977159913
	pesos_i(9871) := b"1111111111111111_1111111111111111_1111001100000110_0111110011001001"; -- -0.050682259571465285
	pesos_i(9872) := b"1111111111111111_1111111111111111_1110100010011101_1101111101111111"; -- -0.09134104869519412
	pesos_i(9873) := b"1111111111111111_1111111111111111_1110110011101101_1010100000011110"; -- -0.07449864650860152
	pesos_i(9874) := b"0000000000000000_0000000000000000_0010010000011001_1011000110100111"; -- 0.14101705865750447
	pesos_i(9875) := b"0000000000000000_0000000000000000_0001101001001001_0111010100000110"; -- 0.10268336665833382
	pesos_i(9876) := b"0000000000000000_0000000000000000_0000100010001101_0101000000110001"; -- 0.03340626897344309
	pesos_i(9877) := b"0000000000000000_0000000000000000_0000110111000101_1111101101000011"; -- 0.05380220771820645
	pesos_i(9878) := b"1111111111111111_1111111111111111_1111011111110011_1110101111010100"; -- -0.0314343079083433
	pesos_i(9879) := b"0000000000000000_0000000000000000_0000010100011101_0111010001110001"; -- 0.019980695418519608
	pesos_i(9880) := b"1111111111111111_1111111111111111_1111101001011100_1000010100010100"; -- -0.02202575939999782
	pesos_i(9881) := b"0000000000000000_0000000000000000_0000000001111001_0111110111101011"; -- 0.001853818823895282
	pesos_i(9882) := b"0000000000000000_0000000000000000_0000101110011100_0000011101010001"; -- 0.04534955712236701
	pesos_i(9883) := b"0000000000000000_0000000000000000_0001100111110010_0000010110111110"; -- 0.1013492192830722
	pesos_i(9884) := b"0000000000000000_0000000000000000_0000110100001001_1100111110110000"; -- 0.05093095826687742
	pesos_i(9885) := b"0000000000000000_0000000000000000_0001111011110011_0101001001111000"; -- 0.12090030136846465
	pesos_i(9886) := b"1111111111111111_1111111111111111_1111011100110100_1100011111101111"; -- -0.0343508761082001
	pesos_i(9887) := b"1111111111111111_1111111111111111_1101110100000011_0111110011100011"; -- -0.1366655298568259
	pesos_i(9888) := b"0000000000000000_0000000000000000_0000000111000000_0010111110111011"; -- 0.006838782491880641
	pesos_i(9889) := b"0000000000000000_0000000000000000_0000010010011110_1001100110101001"; -- 0.01804504760692073
	pesos_i(9890) := b"1111111111111111_1111111111111111_1111110011001110_1000100011111011"; -- -0.012473524850591895
	pesos_i(9891) := b"1111111111111111_1111111111111111_1111111001001000_1111110001011110"; -- -0.006698824844336332
	pesos_i(9892) := b"0000000000000000_0000000000000000_0000111110101111_1111011100100001"; -- 0.06127876811134514
	pesos_i(9893) := b"1111111111111111_1111111111111111_1101100010000100_0001101110101011"; -- -0.1542341906578629
	pesos_i(9894) := b"0000000000000000_0000000000000000_0001001001101110_1101001100000110"; -- 0.07200354488235812
	pesos_i(9895) := b"0000000000000000_0000000000000000_0001111111101100_0111110001100101"; -- 0.1247022386248283
	pesos_i(9896) := b"1111111111111111_1111111111111111_1110110100001001_1001101101001000"; -- -0.07407216545023881
	pesos_i(9897) := b"0000000000000000_0000000000000000_0010011101011010_0001110001110011"; -- 0.15371873678915568
	pesos_i(9898) := b"0000000000000000_0000000000000000_0000011111011110_1100010010001000"; -- 0.030742915402200033
	pesos_i(9899) := b"1111111111111111_1111111111111111_1110101001000110_1010011100010110"; -- -0.08485942560916451
	pesos_i(9900) := b"0000000000000000_0000000000000000_0001011010010110_0101100011011000"; -- 0.08823161376564106
	pesos_i(9901) := b"1111111111111111_1111111111111111_1110101111101011_0100010011001001"; -- -0.07844133463005441
	pesos_i(9902) := b"0000000000000000_0000000000000000_0000011011001010_0100100110110111"; -- 0.0265241691226707
	pesos_i(9903) := b"0000000000000000_0000000000000000_0000100101111011_0111001111010000"; -- 0.03703998398497417
	pesos_i(9904) := b"0000000000000000_0000000000000000_0001010101110000_1111011101100100"; -- 0.0837549801007641
	pesos_i(9905) := b"0000000000000000_0000000000000000_0000001011001011_0110010101010011"; -- 0.010916073558278878
	pesos_i(9906) := b"1111111111111111_1111111111111111_1111111000110110_1100001010100101"; -- -0.006976923779071312
	pesos_i(9907) := b"1111111111111111_1111111111111111_1111111111011000_0110101001101011"; -- -0.0006040085367010673
	pesos_i(9908) := b"1111111111111111_1111111111111111_1111010110011011_0110011011001100"; -- -0.04059751055021008
	pesos_i(9909) := b"1111111111111111_1111111111111111_1110000101011011_1100000111101101"; -- -0.11969364138762564
	pesos_i(9910) := b"0000000000000000_0000000000000000_0001110110101000_1011001100101111"; -- 0.11585540663365167
	pesos_i(9911) := b"0000000000000000_0000000000000000_0000100100010100_1110100010100111"; -- 0.035475292882538034
	pesos_i(9912) := b"0000000000000000_0000000000000000_0001110000001111_1000000111111111"; -- 0.10961163025996783
	pesos_i(9913) := b"1111111111111111_1111111111111111_1110100000101111_0000110011000010"; -- -0.09303207647748021
	pesos_i(9914) := b"1111111111111111_1111111111111111_1111010001001000_1101111010110110"; -- -0.045763092637840765
	pesos_i(9915) := b"1111111111111111_1111111111111111_1110000101100011_1111100100011001"; -- -0.11956828247856222
	pesos_i(9916) := b"1111111111111111_1111111111111111_1111000100101001_1101011010110000"; -- -0.05795534318686605
	pesos_i(9917) := b"0000000000000000_0000000000000000_0000101011011101_0101110100100101"; -- 0.042440244153426745
	pesos_i(9918) := b"1111111111111111_1111111111111111_1101111100111100_0011000110001101"; -- -0.1279877692647574
	pesos_i(9919) := b"0000000000000000_0000000000000000_0000100011000011_1111101110001111"; -- 0.03424045781675311
	pesos_i(9920) := b"0000000000000000_0000000000000000_0000001010111000_1111011100001111"; -- 0.010634843079122686
	pesos_i(9921) := b"1111111111111111_1111111111111111_1111010001110101_0101001100111010"; -- -0.04508476094967302
	pesos_i(9922) := b"1111111111111111_1111111111111111_1110100010000111_0100000001010110"; -- -0.09168622869528885
	pesos_i(9923) := b"1111111111111111_1111111111111111_1111101110001110_1100110110110100"; -- -0.017352241097175605
	pesos_i(9924) := b"1111111111111111_1111111111111111_1111100100101001_1010000010000111"; -- -0.026708571414823475
	pesos_i(9925) := b"1111111111111111_1111111111111111_1111010100100010_1011101011101101"; -- -0.042438809509747516
	pesos_i(9926) := b"0000000000000000_0000000000000000_0000111010111000_1011010111111101"; -- 0.05750596453532835
	pesos_i(9927) := b"0000000000000000_0000000000000000_0000100001011111_0111111111101101"; -- 0.03270720994263131
	pesos_i(9928) := b"1111111111111111_1111111111111111_1111011001100111_1001011001100111"; -- -0.0374818799818874
	pesos_i(9929) := b"1111111111111111_1111111111111111_1101101001001100_1001101110001110"; -- -0.14726856019288637
	pesos_i(9930) := b"1111111111111111_1111111111111111_1111000011100011_1011110110010010"; -- -0.05902495557605939
	pesos_i(9931) := b"0000000000000000_0000000000000000_0010000001011010_0110100100001011"; -- 0.12637955210732568
	pesos_i(9932) := b"1111111111111111_1111111111111111_1101110110111111_0000000011010000"; -- -0.13380427291341027
	pesos_i(9933) := b"0000000000000000_0000000000000000_0010010101000000_0111100101011111"; -- 0.1455150468944749
	pesos_i(9934) := b"1111111111111111_1111111111111111_1101110000110100_1000001100000011"; -- -0.13982373401725107
	pesos_i(9935) := b"1111111111111111_1111111111111111_1111100101000001_0011000010101000"; -- -0.026349028548111608
	pesos_i(9936) := b"1111111111111111_1111111111111111_1101101111001100_1010000001001110"; -- -0.14140890203991038
	pesos_i(9937) := b"0000000000000000_0000000000000000_0001110011000011_1010111011010101"; -- 0.11236088470752156
	pesos_i(9938) := b"1111111111111111_1111111111111111_1110111101100011_0101011010111110"; -- -0.06489045960180473
	pesos_i(9939) := b"1111111111111111_1111111111111111_1111011111000110_0011010111110001"; -- -0.03213179457850801
	pesos_i(9940) := b"1111111111111111_1111111111111111_1110110101001100_0001000111000000"; -- -0.07305802400104476
	pesos_i(9941) := b"1111111111111111_1111111111111111_1110100100001001_1111101001101001"; -- -0.0896914953762944
	pesos_i(9942) := b"0000000000000000_0000000000000000_0001000010101111_1011010110111000"; -- 0.06518111941372715
	pesos_i(9943) := b"1111111111111111_1111111111111111_1101101111001010_0111000000111101"; -- -0.1414422847213707
	pesos_i(9944) := b"1111111111111111_1111111111111111_1111111110010100_0110011000101010"; -- -0.0016418598343608311
	pesos_i(9945) := b"1111111111111111_1111111111111111_1111111011110011_1000110110101000"; -- -0.00409617079836621
	pesos_i(9946) := b"1111111111111111_1111111111111111_1110101111010001_1000011101000010"; -- -0.07883410119231846
	pesos_i(9947) := b"0000000000000000_0000000000000000_0001010011101101_1000111011010001"; -- 0.0817498454879448
	pesos_i(9948) := b"1111111111111111_1111111111111111_1111101010010011_1101100111101100"; -- -0.021181468742331237
	pesos_i(9949) := b"0000000000000000_0000000000000000_0000010110111000_0101000000001110"; -- 0.022343638932456476
	pesos_i(9950) := b"1111111111111111_1111111111111111_1110011111110011_1110111100110000"; -- -0.09393410760641788
	pesos_i(9951) := b"0000000000000000_0000000000000000_0001001101001111_0010000000000101"; -- 0.07542610280716722
	pesos_i(9952) := b"1111111111111111_1111111111111111_1111010101010000_0110110000001011"; -- -0.04174160700358859
	pesos_i(9953) := b"0000000000000000_0000000000000000_0000000111111001_0010000101111010"; -- 0.007707683909589587
	pesos_i(9954) := b"0000000000000000_0000000000000000_0000011100001101_1010110001011101"; -- 0.02755238797369
	pesos_i(9955) := b"0000000000000000_0000000000000000_0010001110011101_0110010100011100"; -- 0.139120406361466
	pesos_i(9956) := b"1111111111111111_1111111111111111_1111101001000111_0011000101011110"; -- -0.0223511833816229
	pesos_i(9957) := b"0000000000000000_0000000000000000_0001101000111000_0011101111001010"; -- 0.10242055599581819
	pesos_i(9958) := b"0000000000000000_0000000000000000_0000111100011100_0100110001001011"; -- 0.05902554353446613
	pesos_i(9959) := b"1111111111111111_1111111111111111_1111001011100000_1001011111001001"; -- -0.05126048410442245
	pesos_i(9960) := b"1111111111111111_1111111111111111_1101101110010010_1000100101001110"; -- -0.1422952828182054
	pesos_i(9961) := b"1111111111111111_1111111111111111_1110110100110100_1111101011110101"; -- -0.07341033488007427
	pesos_i(9962) := b"0000000000000000_0000000000000000_0000110000010111_0101000110010010"; -- 0.04723081404040462
	pesos_i(9963) := b"0000000000000000_0000000000000000_0001000100001011_1110001001110011"; -- 0.06658759405307046
	pesos_i(9964) := b"0000000000000000_0000000000000000_0000111110011111_1010001110000001"; -- 0.061029643057334965
	pesos_i(9965) := b"0000000000000000_0000000000000000_0001110101110000_0010100100011001"; -- 0.11499268391985958
	pesos_i(9966) := b"1111111111111111_1111111111111111_1110011101111000_0110010011111010"; -- -0.0958191767001175
	pesos_i(9967) := b"1111111111111111_1111111111111111_1111110111100001_1010100110001001"; -- -0.008275417311798153
	pesos_i(9968) := b"1111111111111111_1111111111111111_1101101111011011_0100000011010011"; -- -0.14118571138637262
	pesos_i(9969) := b"1111111111111111_1111111111111111_1110100111011011_1011111111101000"; -- -0.08649063662358934
	pesos_i(9970) := b"1111111111111111_1111111111111111_1111011000011101_1100000001011011"; -- -0.03860852989083868
	pesos_i(9971) := b"0000000000000000_0000000000000000_0001010011110000_1011100001110011"; -- 0.08179810329023846
	pesos_i(9972) := b"1111111111111111_1111111111111111_1110010010000100_1011010111010100"; -- -0.10735000209451559
	pesos_i(9973) := b"0000000000000000_0000000000000000_0000010110000100_0011111001110011"; -- 0.02154913245957819
	pesos_i(9974) := b"1111111111111111_1111111111111111_1111111111000000_0010110100100100"; -- -0.0009738718328705386
	pesos_i(9975) := b"0000000000000000_0000000000000000_0010011101001000_0010011111101100"; -- 0.15344476240869057
	pesos_i(9976) := b"0000000000000000_0000000000000000_0001001111111010_0000010111101000"; -- 0.07803379922503711
	pesos_i(9977) := b"0000000000000000_0000000000000000_0010000101001110_0001100100111000"; -- 0.13009793866477606
	pesos_i(9978) := b"0000000000000000_0000000000000000_0001010001111001_1110100011010101"; -- 0.0799851913223928
	pesos_i(9979) := b"0000000000000000_0000000000000000_0001100000010101_1101110110000010"; -- 0.09408363756400896
	pesos_i(9980) := b"1111111111111111_1111111111111111_1110000001001110_1001110000110000"; -- -0.12380050505873305
	pesos_i(9981) := b"1111111111111111_1111111111111111_1101110101000101_1110011010011010"; -- -0.1356521487172947
	pesos_i(9982) := b"1111111111111111_1111111111111111_1111111100100111_0101100001010111"; -- -0.003305891677592325
	pesos_i(9983) := b"1111111111111111_1111111111111111_1110110011101100_1000000110110011"; -- -0.0745161950601602
	pesos_i(9984) := b"0000000000000000_0000000000000000_0001110000110011_0110000101100111"; -- 0.11015900386064899
	pesos_i(9985) := b"0000000000000000_0000000000000000_0001000111001001_0010110011111101"; -- 0.06947594818906842
	pesos_i(9986) := b"1111111111111111_1111111111111111_1111100110001100_0010001100110010"; -- -0.02520542181472068
	pesos_i(9987) := b"1111111111111111_1111111111111111_1111010101011010_0000100010100000"; -- -0.041594944924975126
	pesos_i(9988) := b"1111111111111111_1111111111111111_1110100001101110_1100101001000100"; -- -0.09205947728273497
	pesos_i(9989) := b"1111111111111111_1111111111111111_1110101000000100_1111001011101100"; -- -0.08586198565942725
	pesos_i(9990) := b"1111111111111111_1111111111111111_1111000100000111_1110101100110001"; -- -0.05847292005522056
	pesos_i(9991) := b"1111111111111111_1111111111111111_1110100000101000_0011001001010100"; -- -0.09313664866768241
	pesos_i(9992) := b"0000000000000000_0000000000000000_0010100001100111_1110100001110001"; -- 0.15783550975898553
	pesos_i(9993) := b"0000000000000000_0000000000000000_0000001110011000_0101001110001110"; -- 0.01404306615770836
	pesos_i(9994) := b"0000000000000000_0000000000000000_0000100000110000_0111110100001011"; -- 0.03198987490751102
	pesos_i(9995) := b"0000000000000000_0000000000000000_0001000010001000_0011110001101100"; -- 0.06457879675768484
	pesos_i(9996) := b"1111111111111111_1111111111111111_1111001100001010_0101010100110000"; -- -0.050623584467978724
	pesos_i(9997) := b"1111111111111111_1111111111111111_1110000001000101_0011011101010010"; -- -0.12394384610598842
	pesos_i(9998) := b"0000000000000000_0000000000000000_0000110011101111_0100000011011111"; -- 0.05052571724321654
	pesos_i(9999) := b"0000000000000000_0000000000000000_0001011011001110_0001000100100110"; -- 0.08908183268265274
	pesos_i(10000) := b"1111111111111111_1111111111111111_1111000111101101_0010101101001001"; -- -0.0549748369272287
	pesos_i(10001) := b"0000000000000000_0000000000000000_0010010101010100_0110010001000010"; -- 0.145818964083847
	pesos_i(10002) := b"1111111111111111_1111111111111111_1111010000110010_1110001001110011"; -- -0.046098563224368484
	pesos_i(10003) := b"0000000000000000_0000000000000000_0000100101001011_1011010101100110"; -- 0.03631147140949492
	pesos_i(10004) := b"1111111111111111_1111111111111111_1111101110110001_1111000010010111"; -- -0.016816104067723398
	pesos_i(10005) := b"0000000000000000_0000000000000000_0000100011010011_1010110010011010"; -- 0.03447989237033481
	pesos_i(10006) := b"1111111111111111_1111111111111111_1110001011011100_1001010100100000"; -- -0.1138216778613623
	pesos_i(10007) := b"1111111111111111_1111111111111111_1101110101001110_0110110101001000"; -- -0.13552205082374952
	pesos_i(10008) := b"0000000000000000_0000000000000000_0000101100110000_0111010001101000"; -- 0.04370811019143923
	pesos_i(10009) := b"0000000000000000_0000000000000000_0001000111101111_0011000111011011"; -- 0.07005607229556488
	pesos_i(10010) := b"0000000000000000_0000000000000000_0000111100111111_0001111101100011"; -- 0.059556924599243326
	pesos_i(10011) := b"1111111111111111_1111111111111111_1111001000100010_1001110100010110"; -- -0.05415933813125528
	pesos_i(10012) := b"0000000000000000_0000000000000000_0001110001101100_1100110111011110"; -- 0.11103521976502005
	pesos_i(10013) := b"1111111111111111_1111111111111111_1111010100000100_1001001000100000"; -- -0.04289900519354884
	pesos_i(10014) := b"1111111111111111_1111111111111111_1111111001100010_0000110011011100"; -- -0.0063163721648862815
	pesos_i(10015) := b"1111111111111111_1111111111111111_1110100110011100_0111111100100100"; -- -0.08745580067642224
	pesos_i(10016) := b"1111111111111111_1111111111111111_1110100001001100_0110001110010001"; -- -0.09258439747269016
	pesos_i(10017) := b"1111111111111111_1111111111111111_1111110010001010_1100111001001101"; -- -0.013506990519107144
	pesos_i(10018) := b"1111111111111111_1111111111111111_1111101111001100_1011101011011101"; -- -0.01640731903580618
	pesos_i(10019) := b"1111111111111111_1111111111111111_1111111110101011_1110111000010010"; -- -0.001282807043629832
	pesos_i(10020) := b"0000000000000000_0000000000000000_0001010100100110_0001110010111000"; -- 0.08261279564698314
	pesos_i(10021) := b"1111111111111111_1111111111111111_1101111100100100_1110001110000010"; -- -0.12834337300831292
	pesos_i(10022) := b"0000000000000000_0000000000000000_0010010100101010_0010111010100011"; -- 0.1451748988372787
	pesos_i(10023) := b"0000000000000000_0000000000000000_0000011100000110_1101110101011111"; -- 0.02744849737309199
	pesos_i(10024) := b"1111111111111111_1111111111111111_1110011011000010_1000101111001111"; -- -0.09859396176530316
	pesos_i(10025) := b"0000000000000000_0000000000000000_0001011110110001_1000101001111110"; -- 0.09255281036529926
	pesos_i(10026) := b"1111111111111111_1111111111111111_1110110101111010_0011000010000110"; -- -0.07235428561308499
	pesos_i(10027) := b"1111111111111111_1111111111111111_1111101010000011_1101000010011001"; -- -0.021426165268830902
	pesos_i(10028) := b"0000000000000000_0000000000000000_0000111001010011_0100101111110000"; -- 0.055958505785228936
	pesos_i(10029) := b"1111111111111111_1111111111111111_1110010010111010_0010011001010000"; -- -0.10653458158945708
	pesos_i(10030) := b"0000000000000000_0000000000000000_0010010011011010_0110101000001110"; -- 0.14395773731762465
	pesos_i(10031) := b"1111111111111111_1111111111111111_1101111001000101_1110010000011110"; -- -0.13174604672747972
	pesos_i(10032) := b"1111111111111111_1111111111111111_1101111011101000_0010100001000100"; -- -0.12927006091643115
	pesos_i(10033) := b"0000000000000000_0000000000000000_0001111101010101_1000011111100110"; -- 0.12239884732728412
	pesos_i(10034) := b"1111111111111111_1111111111111111_1111100100110000_0100010011011010"; -- -0.02660722429578091
	pesos_i(10035) := b"0000000000000000_0000000000000000_0000011101001001_0010101001111010"; -- 0.028460173292936757
	pesos_i(10036) := b"0000000000000000_0000000000000000_0010000111010101_0110101100011100"; -- 0.1321627562171223
	pesos_i(10037) := b"0000000000000000_0000000000000000_0001010010110111_1011101101000100"; -- 0.08092852018623245
	pesos_i(10038) := b"0000000000000000_0000000000000000_0001011100001011_0110000010111001"; -- 0.09001736189294374
	pesos_i(10039) := b"0000000000000000_0000000000000000_0000011101000000_0000101000010000"; -- 0.02832091224909437
	pesos_i(10040) := b"1111111111111111_1111111111111111_1111101100000010_1001001011111110"; -- -0.019491971088992654
	pesos_i(10041) := b"0000000000000000_0000000000000000_0000111110111010_1000000010000001"; -- 0.061439544233188356
	pesos_i(10042) := b"0000000000000000_0000000000000000_0001110101000010_1001101100110111"; -- 0.11429758172006414
	pesos_i(10043) := b"0000000000000000_0000000000000000_0000000000011101_0111101110010100"; -- 0.0004498707662420685
	pesos_i(10044) := b"0000000000000000_0000000000000000_0000110000010101_0011001100111101"; -- 0.04719848851957601
	pesos_i(10045) := b"1111111111111111_1111111111111111_1110101110100011_1111011011011001"; -- -0.07952935411093719
	pesos_i(10046) := b"0000000000000000_0000000000000000_0000101110010000_0101101011011110"; -- 0.04517143183620911
	pesos_i(10047) := b"0000000000000000_0000000000000000_0010010100000001_0100101000111100"; -- 0.1445509334797608
	pesos_i(10048) := b"0000000000000000_0000000000000000_0001111011111110_1111010011000101"; -- 0.12107782180772353
	pesos_i(10049) := b"0000000000000000_0000000000000000_0000001111100010_0111000000111101"; -- 0.015173926282029605
	pesos_i(10050) := b"1111111111111111_1111111111111111_1111001001011010_1101110010010101"; -- -0.053301061309476955
	pesos_i(10051) := b"0000000000000000_0000000000000000_0001010011000110_0000010011111000"; -- 0.08114653647155548
	pesos_i(10052) := b"1111111111111111_1111111111111111_1110110110110111_1010010000000100"; -- -0.07141661549476347
	pesos_i(10053) := b"0000000000000000_0000000000000000_0000010011000111_0001011011011111"; -- 0.018662862251414378
	pesos_i(10054) := b"1111111111111111_1111111111111111_1111100000000101_1000101110100110"; -- -0.031165382367980877
	pesos_i(10055) := b"1111111111111111_1111111111111111_1101111101101010_1100001111101010"; -- -0.12727714104140242
	pesos_i(10056) := b"1111111111111111_1111111111111111_1110110101010000_0111110110111010"; -- -0.07299055295756143
	pesos_i(10057) := b"0000000000000000_0000000000000000_0001110000100101_1001101011110111"; -- 0.1099488117644794
	pesos_i(10058) := b"0000000000000000_0000000000000000_0001110111000100_1000111001010111"; -- 0.1162804567208489
	pesos_i(10059) := b"1111111111111111_1111111111111111_1101100101101101_0101101001111111"; -- -0.15067514792563755
	pesos_i(10060) := b"1111111111111111_1111111111111111_1110000100111001_1101000111001001"; -- -0.12021149482807023
	pesos_i(10061) := b"0000000000000000_0000000000000000_0000111000100101_1001010101011011"; -- 0.05526097742486643
	pesos_i(10062) := b"0000000000000000_0000000000000000_0001010110001000_1010011011111100"; -- 0.08411639831328489
	pesos_i(10063) := b"1111111111111111_1111111111111111_1111101111110010_1111000110111010"; -- -0.015824214972341183
	pesos_i(10064) := b"0000000000000000_0000000000000000_0010011100100000_1100000010001001"; -- 0.15284350712812722
	pesos_i(10065) := b"0000000000000000_0000000000000000_0001111000011010_1100011011001101"; -- 0.11759607808118534
	pesos_i(10066) := b"1111111111111111_1111111111111111_1110001001011010_0101000110001010"; -- -0.11580934889675787
	pesos_i(10067) := b"1111111111111111_1111111111111111_1110100110000001_0011101110111011"; -- -0.08787180599921765
	pesos_i(10068) := b"1111111111111111_1111111111111111_1110100011001000_0000100001000011"; -- -0.09069774982652677
	pesos_i(10069) := b"1111111111111111_1111111111111111_1111100100110000_1010110110101010"; -- -0.02660097690086889
	pesos_i(10070) := b"0000000000000000_0000000000000000_0001111010110001_1000100001110000"; -- 0.11989643807793518
	pesos_i(10071) := b"0000000000000000_0000000000000000_0000110000010111_1110000001000011"; -- 0.0472393190819715
	pesos_i(10072) := b"1111111111111111_1111111111111111_1110011100111001_0011111100010000"; -- -0.09678274015199072
	pesos_i(10073) := b"0000000000000000_0000000000000000_0001000001011010_0010100011010011"; -- 0.06387572436036923
	pesos_i(10074) := b"0000000000000000_0000000000000000_0000000010010010_0111101001111100"; -- 0.002235083805954857
	pesos_i(10075) := b"0000000000000000_0000000000000000_0010100001000100_0100100010001110"; -- 0.1572919221678741
	pesos_i(10076) := b"0000000000000000_0000000000000000_0001001111000111_0110001011101100"; -- 0.07726114525580262
	pesos_i(10077) := b"1111111111111111_1111111111111111_1111101100011100_0100110110101111"; -- -0.01909937369845553
	pesos_i(10078) := b"0000000000000000_0000000000000000_0001011011100011_0101010001011000"; -- 0.08940627235265383
	pesos_i(10079) := b"0000000000000000_0000000000000000_0010010010011110_1101110101101101"; -- 0.14304908679240416
	pesos_i(10080) := b"1111111111111111_1111111111111111_1110000000100010_1110011110011110"; -- -0.12446739582321478
	pesos_i(10081) := b"1111111111111111_1111111111111111_1111110111011000_1101111100101100"; -- -0.008409549380458658
	pesos_i(10082) := b"1111111111111111_1111111111111111_1110100101100100_1110100101111010"; -- -0.08830395470669572
	pesos_i(10083) := b"0000000000000000_0000000000000000_0001000010010110_0100111010111111"; -- 0.06479351189511806
	pesos_i(10084) := b"0000000000000000_0000000000000000_0000111100110100_1100110110110001"; -- 0.05939946714422631
	pesos_i(10085) := b"1111111111111111_1111111111111111_1111011110001001_0111011110101011"; -- -0.033058663239946356
	pesos_i(10086) := b"1111111111111111_1111111111111111_1111000011000101_1111010101011010"; -- -0.05947939438171871
	pesos_i(10087) := b"1111111111111111_1111111111111111_1101100110001011_1110110110100100"; -- -0.15020861391344942
	pesos_i(10088) := b"1111111111111111_1111111111111111_1101110001001100_1111011111011101"; -- -0.13945055831300485
	pesos_i(10089) := b"1111111111111111_1111111111111111_1110100110000001_0101010101101101"; -- -0.08787027453227028
	pesos_i(10090) := b"1111111111111111_1111111111111111_1101101111001001_1001101100001101"; -- -0.1414549915472287
	pesos_i(10091) := b"0000000000000000_0000000000000000_0000111001100001_1011000100000110"; -- 0.056178154056609794
	pesos_i(10092) := b"0000000000000000_0000000000000000_0000011101110000_0011001010001100"; -- 0.029055747291659974
	pesos_i(10093) := b"0000000000000000_0000000000000000_0001111100001011_0001110101001001"; -- 0.12126334229427396
	pesos_i(10094) := b"1111111111111111_1111111111111111_1110101101100101_0000100101001001"; -- -0.08048955878105613
	pesos_i(10095) := b"1111111111111111_1111111111111111_1111000010110101_1010011011000101"; -- -0.059728219028952166
	pesos_i(10096) := b"1111111111111111_1111111111111111_1110011010111100_0111000110110111"; -- -0.09868706975749432
	pesos_i(10097) := b"1111111111111111_1111111111111111_1110110111000011_0111110011100011"; -- -0.07123584221835152
	pesos_i(10098) := b"1111111111111111_1111111111111111_1110011011001001_0101010011001101"; -- -0.09849042890273056
	pesos_i(10099) := b"0000000000000000_0000000000000000_0001011100111000_1100011000110111"; -- 0.0907100565971051
	pesos_i(10100) := b"1111111111111111_1111111111111111_1110000101110010_0001010101111000"; -- -0.11935296835157702
	pesos_i(10101) := b"0000000000000000_0000000000000000_0000100011110011_0011100000100101"; -- 0.03496123212819366
	pesos_i(10102) := b"0000000000000000_0000000000000000_0000110001000110_0001001111011001"; -- 0.047944298262772855
	pesos_i(10103) := b"1111111111111111_1111111111111111_1110100001011001_1111010111101010"; -- -0.09237731014773325
	pesos_i(10104) := b"0000000000000000_0000000000000000_0001110100101100_1000001010010010"; -- 0.1139604193765999
	pesos_i(10105) := b"1111111111111111_1111111111111111_1111111011011011_1001010100111011"; -- -0.004461930434310048
	pesos_i(10106) := b"1111111111111111_1111111111111111_1111101011110100_0111100010011001"; -- -0.01970716729468194
	pesos_i(10107) := b"0000000000000000_0000000000000000_0000000010100110_1110101010101111"; -- 0.00254694726474455
	pesos_i(10108) := b"0000000000000000_0000000000000000_0010000010011001_1100010001110001"; -- 0.127346303464283
	pesos_i(10109) := b"1111111111111111_1111111111111111_1110010101010110_0110001000100110"; -- -0.10415064404170751
	pesos_i(10110) := b"1111111111111111_1111111111111111_1110010101100110_1101011101101001"; -- -0.1038995141252231
	pesos_i(10111) := b"1111111111111111_1111111111111111_1111111011001101_0011110001001110"; -- -0.004680853827994086
	pesos_i(10112) := b"1111111111111111_1111111111111111_1101111111111000_1011101011110101"; -- -0.12511092688465508
	pesos_i(10113) := b"1111111111111111_1111111111111111_1101100111100111_1101101100001010"; -- -0.14880591403843058
	pesos_i(10114) := b"1111111111111111_1111111111111111_1110111101100101_1100001110110001"; -- -0.06485344820650144
	pesos_i(10115) := b"1111111111111111_1111111111111111_1111100111010011_1111010101101010"; -- -0.024109517633929173
	pesos_i(10116) := b"1111111111111111_1111111111111111_1111110101000001_0111111010100010"; -- -0.010719380695912344
	pesos_i(10117) := b"1111111111111111_1111111111111111_1101101101100110_0011010001101000"; -- -0.14297172991929702
	pesos_i(10118) := b"0000000000000000_0000000000000000_0010010111001110_1100011000000101"; -- 0.14768636347117706
	pesos_i(10119) := b"0000000000000000_0000000000000000_0001111000110111_1100111010101000"; -- 0.11803905107055376
	pesos_i(10120) := b"0000000000000000_0000000000000000_0001001010101100_1111100000011010"; -- 0.07295179975147065
	pesos_i(10121) := b"1111111111111111_1111111111111111_1111010011011010_1100101001011010"; -- -0.043536522802493906
	pesos_i(10122) := b"1111111111111111_1111111111111111_1110010101010101_1010100000111100"; -- -0.10416172549215483
	pesos_i(10123) := b"0000000000000000_0000000000000000_0000111101001100_1101010000101011"; -- 0.05976606417794995
	pesos_i(10124) := b"0000000000000000_0000000000000000_0001100110111100_0011000111111111"; -- 0.1005278823323227
	pesos_i(10125) := b"0000000000000000_0000000000000000_0010001100001101_0101000100010111"; -- 0.13692194756687343
	pesos_i(10126) := b"0000000000000000_0000000000000000_0010001000101001_1100011101111100"; -- 0.13345000056905268
	pesos_i(10127) := b"0000000000000000_0000000000000000_0001100101100111_0100110010110100"; -- 0.09923247702777546
	pesos_i(10128) := b"1111111111111111_1111111111111111_1110110110011111_0100010101001001"; -- -0.07178847275662081
	pesos_i(10129) := b"1111111111111111_1111111111111111_1111000010001100_1001110100010111"; -- -0.06035440613452454
	pesos_i(10130) := b"1111111111111111_1111111111111111_1101101101011001_0111110001101000"; -- -0.14316580264062703
	pesos_i(10131) := b"0000000000000000_0000000000000000_0001101111011110_0111001101001101"; -- 0.10886307354578742
	pesos_i(10132) := b"0000000000000000_0000000000000000_0001001100001101_0100000100010100"; -- 0.07442099311373959
	pesos_i(10133) := b"1111111111111111_1111111111111111_1110111110100010_0001111001111100"; -- -0.06393250916929172
	pesos_i(10134) := b"0000000000000000_0000000000000000_0001000011110100_0100000101011011"; -- 0.06622703992268626
	pesos_i(10135) := b"0000000000000000_0000000000000000_0000111110100110_1010011111100111"; -- 0.061136716843530975
	pesos_i(10136) := b"1111111111111111_1111111111111111_1110001110001000_0011101110001101"; -- -0.11120250524648492
	pesos_i(10137) := b"1111111111111111_1111111111111111_1110011011000001_0100000000110001"; -- -0.09861372764262265
	pesos_i(10138) := b"1111111111111111_1111111111111111_1110100101001111_1001100011101001"; -- -0.08862919160849889
	pesos_i(10139) := b"0000000000000000_0000000000000000_0001111010100001_0111001101010100"; -- 0.11965103909763715
	pesos_i(10140) := b"1111111111111111_1111111111111111_1111001101101110_1100110101000100"; -- -0.049090548352303996
	pesos_i(10141) := b"1111111111111111_1111111111111111_1101111101110110_0010111111111010"; -- -0.12710285323102258
	pesos_i(10142) := b"0000000000000000_0000000000000000_0000110010010101_0001010111101100"; -- 0.04914986622146448
	pesos_i(10143) := b"0000000000000000_0000000000000000_0001100101110100_1000001000100011"; -- 0.09943402622922817
	pesos_i(10144) := b"1111111111111111_1111111111111111_1110001011111010_0000000100010001"; -- -0.11337273914596839
	pesos_i(10145) := b"1111111111111111_1111111111111111_1110011100001100_0000101101111100"; -- -0.09747245997507645
	pesos_i(10146) := b"0000000000000000_0000000000000000_0010000101001101_0110000110011011"; -- 0.13008699459436673
	pesos_i(10147) := b"1111111111111111_1111111111111111_1110110011110110_0111100110101000"; -- -0.07436408665068363
	pesos_i(10148) := b"1111111111111111_1111111111111111_1110100111111110_0000011111001110"; -- -0.0859675524072905
	pesos_i(10149) := b"1111111111111111_1111111111111111_1111010101011110_0100001101011101"; -- -0.04153040861862421
	pesos_i(10150) := b"1111111111111111_1111111111111111_1111100111010101_1011010111010000"; -- -0.0240827910481812
	pesos_i(10151) := b"0000000000000000_0000000000000000_0000010011011011_1010111011101010"; -- 0.01897710055774859
	pesos_i(10152) := b"0000000000000000_0000000000000000_0001100110100000_1110010011101100"; -- 0.1001113011437948
	pesos_i(10153) := b"1111111111111111_1111111111111111_1111001000011010_1010101110100110"; -- -0.05428054053137617
	pesos_i(10154) := b"0000000000000000_0000000000000000_0000111010101000_0110100000111000"; -- 0.0572571883777684
	pesos_i(10155) := b"1111111111111111_1111111111111111_1110101100111101_0101101000111010"; -- -0.08109508589611589
	pesos_i(10156) := b"0000000000000000_0000000000000000_0001000111000011_1111100010010111"; -- 0.0693965308903651
	pesos_i(10157) := b"1111111111111111_1111111111111111_1110011100110101_0000101111100101"; -- -0.09684682530934097
	pesos_i(10158) := b"0000000000000000_0000000000000000_0001000111100011_1010010111011010"; -- 0.06987988063098724
	pesos_i(10159) := b"1111111111111111_1111111111111111_1110111000110110_1000011001101000"; -- -0.06948051412151494
	pesos_i(10160) := b"0000000000000000_0000000000000000_0001100111101111_1111111101000011"; -- 0.10131831542005174
	pesos_i(10161) := b"0000000000000000_0000000000000000_0001001010001010_1100000101010010"; -- 0.07242973558521208
	pesos_i(10162) := b"0000000000000000_0000000000000000_0001101101000011_0000010101100010"; -- 0.10649140967601747
	pesos_i(10163) := b"0000000000000000_0000000000000000_0010010011011001_1110111111010010"; -- 0.14395045174579243
	pesos_i(10164) := b"0000000000000000_0000000000000000_0001000111110101_0010101111110011"; -- 0.07014727283316163
	pesos_i(10165) := b"0000000000000000_0000000000000000_0000101110101001_1000100111110100"; -- 0.045555708006543974
	pesos_i(10166) := b"0000000000000000_0000000000000000_0001111111110010_0010110111011011"; -- 0.12478911023806054
	pesos_i(10167) := b"1111111111111111_1111111111111111_1110011100101111_0101010000001100"; -- -0.09693407721600944
	pesos_i(10168) := b"1111111111111111_1111111111111111_1110110011010000_0000000010001111"; -- -0.0749511385073849
	pesos_i(10169) := b"0000000000000000_0000000000000000_0001010001000000_1100111110110000"; -- 0.07911394173441673
	pesos_i(10170) := b"1111111111111111_1111111111111111_1110000110001010_1101010111100110"; -- -0.11897528779805723
	pesos_i(10171) := b"1111111111111111_1111111111111111_1110010001011111_0001101001000000"; -- -0.10792385039294283
	pesos_i(10172) := b"1111111111111111_1111111111111111_1110010010000111_0011000011000011"; -- -0.10731215712517572
	pesos_i(10173) := b"0000000000000000_0000000000000000_0001011000011010_0000101010111111"; -- 0.08633486904333262
	pesos_i(10174) := b"1111111111111111_1111111111111111_1101111100000110_1100011010110110"; -- -0.12880285320332757
	pesos_i(10175) := b"1111111111111111_1111111111111111_1111001010010111_0011010001101101"; -- -0.05238029794896772
	pesos_i(10176) := b"1111111111111111_1111111111111111_1110011010101011_1101110001110100"; -- -0.09894010707475624
	pesos_i(10177) := b"0000000000000000_0000000000000000_0000111000110101_1110000110100110"; -- 0.05550966557374441
	pesos_i(10178) := b"1111111111111111_1111111111111111_1111101111010111_0110000010001011"; -- -0.01624485592604711
	pesos_i(10179) := b"0000000000000000_0000000000000000_0000100110001000_1000001110001100"; -- 0.03723928617360737
	pesos_i(10180) := b"1111111111111111_1111111111111111_1111000000001110_0001111111111101"; -- -0.06228447039627313
	pesos_i(10181) := b"0000000000000000_0000000000000000_0001100010100001_0111010110011101"; -- 0.09621367542068723
	pesos_i(10182) := b"0000000000000000_0000000000000000_0010000010100011_1001010110110001"; -- 0.12749610499284733
	pesos_i(10183) := b"1111111111111111_1111111111111111_1110110010011001_1101011000010101"; -- -0.0757776450053377
	pesos_i(10184) := b"0000000000000000_0000000000000000_0000101010000111_0001000110000001"; -- 0.041123479796598854
	pesos_i(10185) := b"1111111111111111_1111111111111111_1111010000000101_1100000101011011"; -- -0.046787181226752114
	pesos_i(10186) := b"1111111111111111_1111111111111111_1110011100100111_1100001101000101"; -- -0.09704951817316745
	pesos_i(10187) := b"1111111111111111_1111111111111111_1111100010100000_0011010010110010"; -- -0.028805452782410715
	pesos_i(10188) := b"1111111111111111_1111111111111111_1110011010100010_1011111101000101"; -- -0.0990791756490848
	pesos_i(10189) := b"1111111111111111_1111111111111111_1111010001010110_1101111011011110"; -- -0.04554946030906078
	pesos_i(10190) := b"1111111111111111_1111111111111111_1110111001001010_1111011010110110"; -- -0.06916864438606746
	pesos_i(10191) := b"0000000000000000_0000000000000000_0001010110101111_1110111110010000"; -- 0.0847158171602847
	pesos_i(10192) := b"0000000000000000_0000000000000000_0000010001010101_1011110001111101"; -- 0.016933231810999566
	pesos_i(10193) := b"1111111111111111_1111111111111111_1111011011011111_0111110100100100"; -- -0.0356523309700351
	pesos_i(10194) := b"0000000000000000_0000000000000000_0010000001100011_0100101110111111"; -- 0.1265151348518522
	pesos_i(10195) := b"0000000000000000_0000000000000000_0001101001111100_1110111100110111"; -- 0.10346884807808587
	pesos_i(10196) := b"1111111111111111_1111111111111111_1111010101011001_1101101011010010"; -- -0.041597675081818754
	pesos_i(10197) := b"0000000000000000_0000000000000000_0010010110011110_1001001100110110"; -- 0.1469509130810773
	pesos_i(10198) := b"1111111111111111_1111111111111111_1101101101100110_0000100110011010"; -- -0.14297428124540076
	pesos_i(10199) := b"1111111111111111_1111111111111111_1101100111011001_1001000101000010"; -- -0.1490239346854049
	pesos_i(10200) := b"1111111111111111_1111111111111111_1110001110110100_1001001111001100"; -- -0.1105258586724708
	pesos_i(10201) := b"0000000000000000_0000000000000000_0001000100010000_0001000010001010"; -- 0.06665137640528263
	pesos_i(10202) := b"0000000000000000_0000000000000000_0010001100011110_1111010001100011"; -- 0.13719108025240195
	pesos_i(10203) := b"0000000000000000_0000000000000000_0001010011110100_1111100000001110"; -- 0.0818629298420219
	pesos_i(10204) := b"0000000000000000_0000000000000000_0001011110110101_0011100111111011"; -- 0.09260904671523466
	pesos_i(10205) := b"0000000000000000_0000000000000000_0000100000010100_0111111100011010"; -- 0.031562751715390525
	pesos_i(10206) := b"0000000000000000_0000000000000000_0001001011101100_1100000000100000"; -- 0.07392502580048223
	pesos_i(10207) := b"1111111111111111_1111111111111111_1101011000011010_0110001110011100"; -- -0.1636598341876841
	pesos_i(10208) := b"0000000000000000_0000000000000000_0000110010111001_0000010100010101"; -- 0.0496981787796488
	pesos_i(10209) := b"1111111111111111_1111111111111111_1110011000101100_0101001011101010"; -- -0.10088617110669408
	pesos_i(10210) := b"0000000000000000_0000000000000000_0000101101111110_1100001010101010"; -- 0.04490296024000366
	pesos_i(10211) := b"1111111111111111_1111111111111111_1111000101000011_0100000110011110"; -- -0.05756750008791148
	pesos_i(10212) := b"1111111111111111_1111111111111111_1111010010110001_1000110000000010"; -- -0.04416584920830643
	pesos_i(10213) := b"1111111111111111_1111111111111111_1111101000010101_1101000000111100"; -- -0.02310465369070332
	pesos_i(10214) := b"0000000000000000_0000000000000000_0001011010011010_0001101100010110"; -- 0.08828896788940657
	pesos_i(10215) := b"0000000000000000_0000000000000000_0001101001110100_1111100101010011"; -- 0.10334738045007309
	pesos_i(10216) := b"1111111111111111_1111111111111111_1111110100101101_1100101001110011"; -- -0.011020037549107953
	pesos_i(10217) := b"1111111111111111_1111111111111111_1111010000111000_1110110110001001"; -- -0.046006349650005794
	pesos_i(10218) := b"1111111111111111_1111111111111111_1110011000001000_1111010010111110"; -- -0.10142584201982235
	pesos_i(10219) := b"0000000000000000_0000000000000000_0001001000101001_0000100110110000"; -- 0.07093868782840075
	pesos_i(10220) := b"1111111111111111_1111111111111111_1110000000011010_1011111010000010"; -- -0.12459191632008736
	pesos_i(10221) := b"1111111111111111_1111111111111111_1110001100100001_1101111001011000"; -- -0.11276445729269502
	pesos_i(10222) := b"1111111111111111_1111111111111111_1110011110000001_1001100110101110"; -- -0.09567870614850223
	pesos_i(10223) := b"1111111111111111_1111111111111111_1111010001000011_1000000100001010"; -- -0.045844969847405555
	pesos_i(10224) := b"1111111111111111_1111111111111111_1110101110000011_0111011110011010"; -- -0.08002521985827785
	pesos_i(10225) := b"0000000000000000_0000000000000000_0000111101010101_1000110110101010"; -- 0.05989919087624815
	pesos_i(10226) := b"0000000000000000_0000000000000000_0001011001100001_1010000011010011"; -- 0.08742718845848631
	pesos_i(10227) := b"0000000000000000_0000000000000000_0010000100011010_1100110101110100"; -- 0.12931522440987028
	pesos_i(10228) := b"1111111111111111_1111111111111111_1110011001111001_0100011100100101"; -- -0.09971194594147997
	pesos_i(10229) := b"1111111111111111_1111111111111111_1111100111001011_0100110000000011"; -- -0.024241685144430616
	pesos_i(10230) := b"0000000000000000_0000000000000000_0000100101100010_1000010010101110"; -- 0.036659519642863084
	pesos_i(10231) := b"1111111111111111_1111111111111111_1111111010000000_0011111011111010"; -- -0.005855621372386867
	pesos_i(10232) := b"1111111111111111_1111111111111111_1101110110010011_1100110111110101"; -- -0.13446343205858788
	pesos_i(10233) := b"0000000000000000_0000000000000000_0000000001010100_0001010010001010"; -- 0.0012829626083829726
	pesos_i(10234) := b"1111111111111111_1111111111111111_1111100000000000_1111100110010011"; -- -0.031235124294040725
	pesos_i(10235) := b"0000000000000000_0000000000000000_0000011010110000_1110110001101011"; -- 0.026137138383346362
	pesos_i(10236) := b"0000000000000000_0000000000000000_0001000101011101_1000110011011010"; -- 0.0678337128313867
	pesos_i(10237) := b"0000000000000000_0000000000000000_0001110001001100_1000101011101011"; -- 0.11054294814104243
	pesos_i(10238) := b"0000000000000000_0000000000000000_0000000011000101_1001111101111100"; -- 0.0030154874565083605
	pesos_i(10239) := b"0000000000000000_0000000000000000_0000101101110100_1101000101010100"; -- 0.044751246552067594
	pesos_i(10240) := b"1111111111111111_1111111111111111_1110010101101000_0101000010011110"; -- -0.10387703077222966
	pesos_i(10241) := b"0000000000000000_0000000000000000_0000101110000000_0010010100011110"; -- 0.0449240873832917
	pesos_i(10242) := b"0000000000000000_0000000000000000_0000001101010100_1101101000001100"; -- 0.013013484980709675
	pesos_i(10243) := b"1111111111111111_1111111111111111_1111110100000001_1000101011010011"; -- -0.011695216552844048
	pesos_i(10244) := b"1111111111111111_1111111111111111_1111010110101010_1010110000000010"; -- -0.04036450342032287
	pesos_i(10245) := b"0000000000000000_0000000000000000_0000101101011100_0110000010010001"; -- 0.04437831432887734
	pesos_i(10246) := b"1111111111111111_1111111111111111_1111100100010110_0011101010111111"; -- -0.02700455506499271
	pesos_i(10247) := b"0000000000000000_0000000000000000_0001110001110011_1101110000000000"; -- 0.1111428737948189
	pesos_i(10248) := b"0000000000000000_0000000000000000_0000000111001110_1001001011011100"; -- 0.00705831407923267
	pesos_i(10249) := b"0000000000000000_0000000000000000_0001110111110101_0111110100000011"; -- 0.11702710455408656
	pesos_i(10250) := b"1111111111111111_1111111111111111_1111001000000111_0010000011010011"; -- -0.05457873207131055
	pesos_i(10251) := b"0000000000000000_0000000000000000_0001010101011001_1111110100011101"; -- 0.08340436904300219
	pesos_i(10252) := b"0000000000000000_0000000000000000_0000010000000101_1110110011000111"; -- 0.015715407047525616
	pesos_i(10253) := b"1111111111111111_1111111111111111_1110111000110101_1000101010010000"; -- -0.06949552511066885
	pesos_i(10254) := b"0000000000000000_0000000000000000_0000110010101100_1011010011000010"; -- 0.049510285701291505
	pesos_i(10255) := b"0000000000000000_0000000000000000_0001011000010000_0010110100100111"; -- 0.08618433193993044
	pesos_i(10256) := b"0000000000000000_0000000000000000_0000011101011001_0001011011110100"; -- 0.02870315041803512
	pesos_i(10257) := b"0000000000000000_0000000000000000_0010000110101100_0110011111111000"; -- 0.13153695866630563
	pesos_i(10258) := b"0000000000000000_0000000000000000_0001101110001011_1100001100101110"; -- 0.10760135533194307
	pesos_i(10259) := b"1111111111111111_1111111111111111_1101101011010110_1010001000100110"; -- -0.14516245430507715
	pesos_i(10260) := b"0000000000000000_0000000000000000_0001000000010000_0000001001000101"; -- 0.06274427580866757
	pesos_i(10261) := b"1111111111111111_1111111111111111_1110110001001100_1110000111001010"; -- -0.07695187397006091
	pesos_i(10262) := b"0000000000000000_0000000000000000_0001101111100001_1001101010110110"; -- 0.10891119901690098
	pesos_i(10263) := b"1111111111111111_1111111111111111_1110001111101010_1110110010010100"; -- -0.10969659216769566
	pesos_i(10264) := b"1111111111111111_1111111111111111_1111000100101000_1001011100110101"; -- -0.057974385901535974
	pesos_i(10265) := b"1111111111111111_1111111111111111_1110000110010001_0110100010010000"; -- -0.1188749930670979
	pesos_i(10266) := b"1111111111111111_1111111111111111_1111111011010010_0110000000111100"; -- -0.004602418302217479
	pesos_i(10267) := b"0000000000000000_0000000000000000_0000100010011000_0010000001001010"; -- 0.03357126058979076
	pesos_i(10268) := b"0000000000000000_0000000000000000_0010010001011111_1010110001010001"; -- 0.14208485580409114
	pesos_i(10269) := b"0000000000000000_0000000000000000_0000010000110000_1000000010011101"; -- 0.01636508773765101
	pesos_i(10270) := b"0000000000000000_0000000000000000_0001100111101011_1100011111111001"; -- 0.10125398482684161
	pesos_i(10271) := b"0000000000000000_0000000000000000_0010010100010100_0101000011100001"; -- 0.14484124648815494
	pesos_i(10272) := b"1111111111111111_1111111111111111_1110101011010001_1011100101001111"; -- -0.08273736793891077
	pesos_i(10273) := b"1111111111111111_1111111111111111_1111111100000011_0100011111010000"; -- -0.003856193228741549
	pesos_i(10274) := b"0000000000000000_0000000000000000_0001001110000001_0111001100011101"; -- 0.07619399513093364
	pesos_i(10275) := b"0000000000000000_0000000000000000_0001001011000111_1000101100011001"; -- 0.07335728990224143
	pesos_i(10276) := b"0000000000000000_0000000000000000_0001110011111001_1111110111100010"; -- 0.11318957118282796
	pesos_i(10277) := b"1111111111111111_1111111111111111_1110010000011111_1011110111101011"; -- -0.10889065744278636
	pesos_i(10278) := b"0000000000000000_0000000000000000_0000101000011100_0110010001101000"; -- 0.03949573082315158
	pesos_i(10279) := b"0000000000000000_0000000000000000_0010011101001000_1110111101110110"; -- 0.15345665583899948
	pesos_i(10280) := b"1111111111111111_1111111111111111_1101111010001101_1111110110100000"; -- -0.13064589342711985
	pesos_i(10281) := b"1111111111111111_1111111111111111_1111010100110011_1110101010100101"; -- -0.04217656576470526
	pesos_i(10282) := b"1111111111111111_1111111111111111_1101101011101101_0001100000111000"; -- -0.14481972353630132
	pesos_i(10283) := b"0000000000000000_0000000000000000_0010001001010100_1111000110110101"; -- 0.13410864508243558
	pesos_i(10284) := b"0000000000000000_0000000000000000_0010001011110011_1100111001101100"; -- 0.13653268938724636
	pesos_i(10285) := b"1111111111111111_1111111111111111_1111010100111011_1111001000001101"; -- -0.04205405401403361
	pesos_i(10286) := b"0000000000000000_0000000000000000_0001111111100110_1000110101001010"; -- 0.12461169299760132
	pesos_i(10287) := b"0000000000000000_0000000000000000_0001011110010101_1001110001100011"; -- 0.09212663086099138
	pesos_i(10288) := b"0000000000000000_0000000000000000_0000111110100010_1111100010110000"; -- 0.06108049684824354
	pesos_i(10289) := b"0000000000000000_0000000000000000_0010000000001010_0000101110000110"; -- 0.1251532746342177
	pesos_i(10290) := b"1111111111111111_1111111111111111_1101101001011010_1110101101001010"; -- -0.14705018463726924
	pesos_i(10291) := b"0000000000000000_0000000000000000_0000101100100011_0010101000100111"; -- 0.04350532013321792
	pesos_i(10292) := b"1111111111111111_1111111111111111_1110111101101011_1000010111011101"; -- -0.06476558065813193
	pesos_i(10293) := b"1111111111111111_1111111111111111_1110101010010110_0111000110100101"; -- -0.08364190793642796
	pesos_i(10294) := b"0000000000000000_0000000000000000_0001011011101001_1111100000010100"; -- 0.08950758446343078
	pesos_i(10295) := b"0000000000000000_0000000000000000_0000011001100111_0100101110111101"; -- 0.02501366966178531
	pesos_i(10296) := b"1111111111111111_1111111111111111_1110111000001100_0010110001111100"; -- -0.07012674314252489
	pesos_i(10297) := b"0000000000000000_0000000000000000_0000100101000101_0000011111111101"; -- 0.03620958261070683
	pesos_i(10298) := b"1111111111111111_1111111111111111_1110101011000110_1011100000101011"; -- -0.08290528254958127
	pesos_i(10299) := b"1111111111111111_1111111111111111_1101111110101011_0011000111000001"; -- -0.12629403159194674
	pesos_i(10300) := b"0000000000000000_0000000000000000_0000011111100001_0001000000001110"; -- 0.030777934454477834
	pesos_i(10301) := b"0000000000000000_0000000000000000_0010010100011000_1011001010011010"; -- 0.1449081065114115
	pesos_i(10302) := b"0000000000000000_0000000000000000_0001110111100001_1110100000001110"; -- 0.11672830909786494
	pesos_i(10303) := b"1111111111111111_1111111111111111_1111011010001011_0110011011101000"; -- -0.036935394691751486
	pesos_i(10304) := b"0000000000000000_0000000000000000_0000111110000101_1000111101100010"; -- 0.06063171522173994
	pesos_i(10305) := b"0000000000000000_0000000000000000_0000100111001011_0100001101110111"; -- 0.038257805338204776
	pesos_i(10306) := b"0000000000000000_0000000000000000_0000111010001111_0001101001010100"; -- 0.05687107619819867
	pesos_i(10307) := b"0000000000000000_0000000000000000_0000100000000011_1111111111101111"; -- 0.031311031151394664
	pesos_i(10308) := b"0000000000000000_0000000000000000_0010001100011110_1000010111100001"; -- 0.13718449357293538
	pesos_i(10309) := b"0000000000000000_0000000000000000_0010001101111000_0100011101101101"; -- 0.13855406195379832
	pesos_i(10310) := b"1111111111111111_1111111111111111_1110111111111111_1100010110111111"; -- -0.0625034722382522
	pesos_i(10311) := b"1111111111111111_1111111111111111_1110010000110011_0000000011011000"; -- -0.10859675140578715
	pesos_i(10312) := b"1111111111111111_1111111111111111_1111010001010001_1010000001010110"; -- -0.0456294813098323
	pesos_i(10313) := b"1111111111111111_1111111111111111_1111111001010100_0111011110000000"; -- -0.006523638903534889
	pesos_i(10314) := b"1111111111111111_1111111111111111_1110010101011101_0010111011010100"; -- -0.10404689143230987
	pesos_i(10315) := b"1111111111111111_1111111111111111_1111111100111110_1011011101110011"; -- -0.0029492707633389766
	pesos_i(10316) := b"0000000000000000_0000000000000000_0000000011100010_1001010110110101"; -- 0.0034574094686883683
	pesos_i(10317) := b"0000000000000000_0000000000000000_0000111011011110_0011101100101100"; -- 0.05807847816344693
	pesos_i(10318) := b"0000000000000000_0000000000000000_0000010110100100_0101000000110000"; -- 0.022038470895832638
	pesos_i(10319) := b"0000000000000000_0000000000000000_0001000000000111_1100110110101001"; -- 0.06261906991394398
	pesos_i(10320) := b"1111111111111111_1111111111111111_1110001001000110_0111101000010101"; -- -0.1161121080402562
	pesos_i(10321) := b"1111111111111111_1111111111111111_1111101001101000_1010100111111001"; -- -0.02184045489014034
	pesos_i(10322) := b"0000000000000000_0000000000000000_0010010110111000_0000110101111011"; -- 0.14733967069173878
	pesos_i(10323) := b"0000000000000000_0000000000000000_0000100100100101_1100001101111110"; -- 0.035732477506468616
	pesos_i(10324) := b"0000000000000000_0000000000000000_0001011111011100_0000010001001001"; -- 0.09320093904943313
	pesos_i(10325) := b"0000000000000000_0000000000000000_0001010111001101_1110101101011000"; -- 0.08517332940868472
	pesos_i(10326) := b"1111111111111111_1111111111111111_1110001000011110_1000000101001101"; -- -0.11672202942790433
	pesos_i(10327) := b"1111111111111111_1111111111111111_1110100101010100_0111111000110001"; -- -0.08855449004965861
	pesos_i(10328) := b"1111111111111111_1111111111111111_1110010101100101_1111101100111000"; -- -0.10391263847115544
	pesos_i(10329) := b"1111111111111111_1111111111111111_1110101101111001_0100101111000000"; -- -0.08018042141876416
	pesos_i(10330) := b"0000000000000000_0000000000000000_0010000010010000_1000101010000001"; -- 0.12720552111302078
	pesos_i(10331) := b"1111111111111111_1111111111111111_1110011011101101_0100101111100100"; -- -0.09794164352732733
	pesos_i(10332) := b"1111111111111111_1111111111111111_1110001001110111_0101010001110011"; -- -0.11536667051856173
	pesos_i(10333) := b"0000000000000000_0000000000000000_0001001001110000_1000110111000111"; -- 0.07202993484758308
	pesos_i(10334) := b"1111111111111111_1111111111111111_1101111000011101_0000010111011101"; -- -0.13236964564623113
	pesos_i(10335) := b"1111111111111111_1111111111111111_1110100010000010_1000001000010000"; -- -0.09175860502872195
	pesos_i(10336) := b"0000000000000000_0000000000000000_0001000011101101_1001110010100110"; -- 0.06612566994586995
	pesos_i(10337) := b"0000000000000000_0000000000000000_0000111111010001_1100111110111010"; -- 0.06179521839140521
	pesos_i(10338) := b"0000000000000000_0000000000000000_0001000001010011_0011111111100110"; -- 0.06377028816323747
	pesos_i(10339) := b"1111111111111111_1111111111111111_1110011101101100_1110111111111101"; -- -0.09599399639925739
	pesos_i(10340) := b"1111111111111111_1111111111111111_1101101100011001_0010111001101100"; -- -0.1441470132382385
	pesos_i(10341) := b"1111111111111111_1111111111111111_1110000001100110_1100111100101111"; -- -0.12343125435937012
	pesos_i(10342) := b"1111111111111111_1111111111111111_1110110000101010_0010010110000110"; -- -0.07748189425723226
	pesos_i(10343) := b"1111111111111111_1111111111111111_1101100100011111_0010000100111000"; -- -0.1518687475286723
	pesos_i(10344) := b"1111111111111111_1111111111111111_1110011010010101_0010001101100111"; -- -0.09928683027413733
	pesos_i(10345) := b"1111111111111111_1111111111111111_1111110111011011_0000110000111100"; -- -0.00837634600647673
	pesos_i(10346) := b"1111111111111111_1111111111111111_1111110010111000_0100000010011101"; -- -0.012813531461390686
	pesos_i(10347) := b"1111111111111111_1111111111111111_1110100101000100_1110110001101000"; -- -0.08879206144603262
	pesos_i(10348) := b"1111111111111111_1111111111111111_1111100011010111_0111010001001011"; -- -0.02796242886410701
	pesos_i(10349) := b"1111111111111111_1111111111111111_1110010000110101_0000011001101011"; -- -0.10856590163889472
	pesos_i(10350) := b"0000000000000000_0000000000000000_0001001111010100_1111011011010111"; -- 0.0774683260069435
	pesos_i(10351) := b"0000000000000000_0000000000000000_0010011110001010_0011010111001001"; -- 0.15445266863972362
	pesos_i(10352) := b"1111111111111111_1111111111111111_1110011011000111_0111011001011011"; -- -0.0985189464364967
	pesos_i(10353) := b"0000000000000000_0000000000000000_0001000010000110_0010011010101101"; -- 0.06454698305381384
	pesos_i(10354) := b"1111111111111111_1111111111111111_1110110010010111_1000000010101001"; -- -0.07581325412303666
	pesos_i(10355) := b"0000000000000000_0000000000000000_0010001111011001_1101001100101011"; -- 0.14004249371874344
	pesos_i(10356) := b"0000000000000000_0000000000000000_0000001100100111_0000000010011101"; -- 0.012313879313059146
	pesos_i(10357) := b"1111111111111111_1111111111111111_1111101100000110_1011000000011010"; -- -0.019429200685029683
	pesos_i(10358) := b"1111111111111111_1111111111111111_1110101011001001_0001110001110110"; -- -0.08286878710856681
	pesos_i(10359) := b"1111111111111111_1111111111111111_1110000101000110_1110101101100010"; -- -0.12001160483886521
	pesos_i(10360) := b"0000000000000000_0000000000000000_0001000100111000_1001010011000101"; -- 0.06726960948294901
	pesos_i(10361) := b"0000000000000000_0000000000000000_0001100011001110_0100011100110100"; -- 0.0968975546470633
	pesos_i(10362) := b"1111111111111111_1111111111111111_1110001111001101_0111111011001011"; -- -0.11014564082988963
	pesos_i(10363) := b"1111111111111111_1111111111111111_1110001001000101_0011000001000110"; -- -0.11613176616726305
	pesos_i(10364) := b"0000000000000000_0000000000000000_0000010010000000_1110101011101110"; -- 0.017592127803920467
	pesos_i(10365) := b"0000000000000000_0000000000000000_0010000000101001_1111001110101000"; -- 0.12564013329539014
	pesos_i(10366) := b"0000000000000000_0000000000000000_0000100011011010_0000100000100101"; -- 0.03457690147796371
	pesos_i(10367) := b"1111111111111111_1111111111111111_1110100011101111_1100000111011110"; -- -0.0900915939499771
	pesos_i(10368) := b"0000000000000000_0000000000000000_0000010010000000_1101010100010000"; -- 0.01759082442187956
	pesos_i(10369) := b"1111111111111111_1111111111111111_1110001111001100_0110010010101010"; -- -0.11016245705814788
	pesos_i(10370) := b"0000000000000000_0000000000000000_0000111000100100_0001000110001000"; -- 0.055237861236899936
	pesos_i(10371) := b"0000000000000000_0000000000000000_0000000100100110_0100000000011110"; -- 0.004489905647245871
	pesos_i(10372) := b"1111111111111111_1111111111111111_1110111100101001_0101110110001000"; -- -0.06577506473188749
	pesos_i(10373) := b"0000000000000000_0000000000000000_0001010010010110_1101110100000010"; -- 0.08042699151287747
	pesos_i(10374) := b"0000000000000000_0000000000000000_0001111110111101_0110101101100011"; -- 0.12398406191232604
	pesos_i(10375) := b"1111111111111111_1111111111111111_1111110000010111_0000010011010011"; -- -0.015273760323165499
	pesos_i(10376) := b"1111111111111111_1111111111111111_1111111000100000_0111101110101101"; -- -0.007316846985812423
	pesos_i(10377) := b"0000000000000000_0000000000000000_0001001011001111_1101110011110100"; -- 0.0734842391320819
	pesos_i(10378) := b"1111111111111111_1111111111111111_1101101100101000_0101010010010101"; -- -0.14391585704759585
	pesos_i(10379) := b"0000000000000000_0000000000000000_0001010111010010_0000110101101011"; -- 0.0852363954742464
	pesos_i(10380) := b"0000000000000000_0000000000000000_0000100101010110_1010101010100100"; -- 0.03647867674446602
	pesos_i(10381) := b"1111111111111111_1111111111111111_1110110111011000_1111110111100100"; -- -0.0709077184129898
	pesos_i(10382) := b"1111111111111111_1111111111111111_1111001000000001_1100111101111101"; -- -0.054659873997210756
	pesos_i(10383) := b"1111111111111111_1111111111111111_1110111001001001_0010100111010111"; -- -0.06919611453285225
	pesos_i(10384) := b"0000000000000000_0000000000000000_0010011110011111_0101100111000001"; -- 0.1547752472409401
	pesos_i(10385) := b"1111111111111111_1111111111111111_1111000000110100_1000101001010000"; -- -0.06169829887856745
	pesos_i(10386) := b"0000000000000000_0000000000000000_0000001101010001_1100011101110101"; -- 0.012966600476245514
	pesos_i(10387) := b"1111111111111111_1111111111111111_1110111110110100_0100011111000001"; -- -0.06365539105058612
	pesos_i(10388) := b"1111111111111111_1111111111111111_1111101111011101_0011101100010010"; -- -0.01615553683270258
	pesos_i(10389) := b"1111111111111111_1111111111111111_1110101100011010_0000010000111110"; -- -0.08163426861424855
	pesos_i(10390) := b"1111111111111111_1111111111111111_1110001010011000_0001100000010010"; -- -0.11486672945246666
	pesos_i(10391) := b"0000000000000000_0000000000000000_0001000100001011_1010010101010111"; -- 0.06658395167531694
	pesos_i(10392) := b"1111111111111111_1111111111111111_1101101100011010_0011001111011011"; -- -0.14413143071046247
	pesos_i(10393) := b"1111111111111111_1111111111111111_1111101111101110_1111001111111111"; -- -0.015885114989065273
	pesos_i(10394) := b"1111111111111111_1111111111111111_1111010001010100_1011111001011101"; -- -0.045581915265268926
	pesos_i(10395) := b"1111111111111111_1111111111111111_1101111111010010_0000101000101001"; -- -0.12570129876152658
	pesos_i(10396) := b"1111111111111111_1111111111111111_1110110011100011_0010000100000110"; -- -0.07465928655662106
	pesos_i(10397) := b"0000000000000000_0000000000000000_0000101111101011_0001001010110111"; -- 0.04655568085910501
	pesos_i(10398) := b"0000000000000000_0000000000000000_0001100000000100_0100101111001110"; -- 0.09381555358337348
	pesos_i(10399) := b"1111111111111111_1111111111111111_1110000001010110_0010010011010011"; -- -0.12368554923547766
	pesos_i(10400) := b"1111111111111111_1111111111111111_1110100000100101_1100001111000101"; -- -0.09317375613627658
	pesos_i(10401) := b"1111111111111111_1111111111111111_1111101101101111_0110100011000101"; -- -0.017831279678963214
	pesos_i(10402) := b"1111111111111111_1111111111111111_1101111001011110_0100110010111100"; -- -0.13137360014715355
	pesos_i(10403) := b"1111111111111111_1111111111111111_1110011011000011_0000111101001010"; -- -0.09858612479888523
	pesos_i(10404) := b"0000000000000000_0000000000000000_0000110000110011_0110010110101001"; -- 0.04765925768716943
	pesos_i(10405) := b"1111111111111111_1111111111111111_1111101001010111_0101110101111001"; -- -0.022104413874673795
	pesos_i(10406) := b"0000000000000000_0000000000000000_0001001111101111_1110111111101000"; -- 0.07787990020252546
	pesos_i(10407) := b"0000000000000000_0000000000000000_0000001100011101_0110011010011101"; -- 0.012167371133158298
	pesos_i(10408) := b"0000000000000000_0000000000000000_0001001001110001_0101100010101110"; -- 0.072042028779742
	pesos_i(10409) := b"0000000000000000_0000000000000000_0001111001010100_1111111110111111"; -- 0.11848448191827601
	pesos_i(10410) := b"0000000000000000_0000000000000000_0000000000111111_1100111011010000"; -- 0.0009736305953256117
	pesos_i(10411) := b"0000000000000000_0000000000000000_0001010011001101_1001000000011001"; -- 0.08126164057607893
	pesos_i(10412) := b"0000000000000000_0000000000000000_0000011011001101_0010011011010010"; -- 0.02656786557940345
	pesos_i(10413) := b"1111111111111111_1111111111111111_1111011101000100_1100101011110110"; -- -0.03410655499483623
	pesos_i(10414) := b"1111111111111111_1111111111111111_1110011101010100_0100010100101010"; -- -0.09637038915400249
	pesos_i(10415) := b"1111111111111111_1111111111111111_1110000001111001_0110100111011101"; -- -0.12314737662499661
	pesos_i(10416) := b"1111111111111111_1111111111111111_1101110001010010_0011000100001011"; -- -0.139370856003621
	pesos_i(10417) := b"0000000000000000_0000000000000000_0000110010010010_1001010100010010"; -- 0.049111668483470414
	pesos_i(10418) := b"1111111111111111_1111111111111111_1111100100101110_0111100011101000"; -- -0.026634639062487482
	pesos_i(10419) := b"0000000000000000_0000000000000000_0001000100010001_0001001111011110"; -- 0.06666683353528034
	pesos_i(10420) := b"1111111111111111_1111111111111111_1101101001001110_1011111101001111"; -- -0.14723591158154908
	pesos_i(10421) := b"1111111111111111_1111111111111111_1111010001000010_0000100111000100"; -- -0.045867337786483976
	pesos_i(10422) := b"1111111111111111_1111111111111111_1101111100111111_0000111111010110"; -- -0.12794400245662668
	pesos_i(10423) := b"0000000000000000_0000000000000000_0000001011010110_1111001111111111"; -- 0.011092424203553702
	pesos_i(10424) := b"0000000000000000_0000000000000000_0010000010111000_0111011000011111"; -- 0.1278146577183991
	pesos_i(10425) := b"0000000000000000_0000000000000000_0001000101111110_1000011011010011"; -- 0.06833689363768244
	pesos_i(10426) := b"0000000000000000_0000000000000000_0010000010011010_1100010110100100"; -- 0.12736163392948763
	pesos_i(10427) := b"1111111111111111_1111111111111111_1110000000110100_1010011100001111"; -- -0.12419658545778298
	pesos_i(10428) := b"0000000000000000_0000000000000000_0000111110010100_0011000111010001"; -- 0.06085502009831786
	pesos_i(10429) := b"0000000000000000_0000000000000000_0010011000011100_1000110100101001"; -- 0.14887315992501868
	pesos_i(10430) := b"0000000000000000_0000000000000000_0001110110100111_1101010110000010"; -- 0.11584219374874079
	pesos_i(10431) := b"0000000000000000_0000000000000000_0001001011011001_1100110101001110"; -- 0.07363589438694605
	pesos_i(10432) := b"0000000000000000_0000000000000000_0000101100000110_0100100011111111"; -- 0.043064653670583944
	pesos_i(10433) := b"0000000000000000_0000000000000000_0001001101010000_1000011010110010"; -- 0.07544748168823068
	pesos_i(10434) := b"1111111111111111_1111111111111111_1110111100000011_0010001000000110"; -- -0.06635844575547785
	pesos_i(10435) := b"0000000000000000_0000000000000000_0000010001010001_0110100111110110"; -- 0.01686727763863937
	pesos_i(10436) := b"1111111111111111_1111111111111111_1101100010001100_1010110111111001"; -- -0.15410340002807613
	pesos_i(10437) := b"0000000000000000_0000000000000000_0000100100011101_0101001111000000"; -- 0.03560374672940628
	pesos_i(10438) := b"0000000000000000_0000000000000000_0001100111110110_0011100111110111"; -- 0.10141336715662991
	pesos_i(10439) := b"1111111111111111_1111111111111111_1111101111000001_0000111101100000"; -- -0.016585387228294925
	pesos_i(10440) := b"1111111111111111_1111111111111111_1110010100111100_0101010101000010"; -- -0.10454814081679574
	pesos_i(10441) := b"1111111111111111_1111111111111111_1111101110000001_1101101010010111"; -- -0.017549837140126034
	pesos_i(10442) := b"1111111111111111_1111111111111111_1111110010000011_1101111101000011"; -- -0.013612791238470583
	pesos_i(10443) := b"1111111111111111_1111111111111111_1110101101000001_1111000000000110"; -- -0.08102512226853785
	pesos_i(10444) := b"0000000000000000_0000000000000000_0010000110000000_1111010111111100"; -- 0.13087403685289295
	pesos_i(10445) := b"0000000000000000_0000000000000000_0000111011000101_1111001001011101"; -- 0.05770792737162629
	pesos_i(10446) := b"1111111111111111_1111111111111111_1111110111110100_0000110101001110"; -- -0.00799481240555472
	pesos_i(10447) := b"1111111111111111_1111111111111111_1111100000100101_0110110100000111"; -- -0.03067892628687203
	pesos_i(10448) := b"1111111111111111_1111111111111111_1110010110101111_0111011010000011"; -- -0.10279139805965533
	pesos_i(10449) := b"1111111111111111_1111111111111111_1101111100110001_0100011111100011"; -- -0.12815428464272532
	pesos_i(10450) := b"0000000000000000_0000000000000000_0001100110000010_1101000110101110"; -- 0.09965239056009831
	pesos_i(10451) := b"0000000000000000_0000000000000000_0000010111001011_0010110100001001"; -- 0.022631468442776925
	pesos_i(10452) := b"1111111111111111_1111111111111111_1111010010000100_0100110110101001"; -- -0.044856210858546075
	pesos_i(10453) := b"1111111111111111_1111111111111111_1111101110011010_1001011110100011"; -- -0.017172358284810077
	pesos_i(10454) := b"1111111111111111_1111111111111111_1111111100100000_1100101110111000"; -- -0.0034058262295919538
	pesos_i(10455) := b"0000000000000000_0000000000000000_0000011000011000_0000111101001111"; -- 0.02380462340574106
	pesos_i(10456) := b"1111111111111111_1111111111111111_1110110011101011_1000110100111000"; -- -0.07453076730704662
	pesos_i(10457) := b"1111111111111111_1111111111111111_1110100001110010_0000011011000001"; -- -0.09201009537442795
	pesos_i(10458) := b"1111111111111111_1111111111111111_1111011100110000_1110010000000001"; -- -0.034410238012905076
	pesos_i(10459) := b"0000000000000000_0000000000000000_0000011110011111_1101111000111111"; -- 0.02978314434358867
	pesos_i(10460) := b"0000000000000000_0000000000000000_0001000101000000_1110111100100101"; -- 0.06739706663869502
	pesos_i(10461) := b"0000000000000000_0000000000000000_0010010111011001_1001101111101101"; -- 0.14785170115400734
	pesos_i(10462) := b"0000000000000000_0000000000000000_0001000000111001_1011100111011000"; -- 0.06338082801464295
	pesos_i(10463) := b"0000000000000000_0000000000000000_0010000011110101_0000001101010111"; -- 0.12873860250497532
	pesos_i(10464) := b"1111111111111111_1111111111111111_1111101111101010_1111000100000111"; -- -0.015946327115903682
	pesos_i(10465) := b"1111111111111111_1111111111111111_1111110010011100_1010011010001011"; -- -0.01323470225010023
	pesos_i(10466) := b"1111111111111111_1111111111111111_1101110000001110_0101001111111101"; -- -0.14040637080095883
	pesos_i(10467) := b"1111111111111111_1111111111111111_1111101011110111_0000111010110110"; -- -0.019667702372929634
	pesos_i(10468) := b"0000000000000000_0000000000000000_0001101001000000_0110011100001111"; -- 0.10254520523301242
	pesos_i(10469) := b"0000000000000000_0000000000000000_0000010101000010_0111100111011110"; -- 0.020545593906540843
	pesos_i(10470) := b"0000000000000000_0000000000000000_0010101001011001_0010011101010101"; -- 0.16542287670545477
	pesos_i(10471) := b"0000000000000000_0000000000000000_0000100001001011_1010111111011100"; -- 0.032404891276198174
	pesos_i(10472) := b"1111111111111111_1111111111111111_1110100011011101_0010000000011010"; -- -0.0903758942788145
	pesos_i(10473) := b"1111111111111111_1111111111111111_1111111011000100_1011000000100101"; -- -0.004811278264809985
	pesos_i(10474) := b"0000000000000000_0000000000000000_0010001111001110_0111101110110011"; -- 0.13986943356748716
	pesos_i(10475) := b"0000000000000000_0000000000000000_0010010011100000_0001101010101010"; -- 0.14404455808895406
	pesos_i(10476) := b"1111111111111111_1111111111111111_1101100111000010_1101000111011111"; -- -0.1493710356691604
	pesos_i(10477) := b"0000000000000000_0000000000000000_0000001010100000_1100101001001110"; -- 0.010265964654396775
	pesos_i(10478) := b"0000000000000000_0000000000000000_0001000010110101_1100001010111001"; -- 0.06527344720499409
	pesos_i(10479) := b"0000000000000000_0000000000000000_0000001000111011_0101011101011111"; -- 0.008717976351103749
	pesos_i(10480) := b"0000000000000000_0000000000000000_0001011001000000_1111010000110010"; -- 0.0869286176312939
	pesos_i(10481) := b"0000000000000000_0000000000000000_0000011000101011_0001100111011001"; -- 0.024095168481899354
	pesos_i(10482) := b"0000000000000000_0000000000000000_0010000000111000_1101010000000011"; -- 0.1258671290415209
	pesos_i(10483) := b"1111111111111111_1111111111111111_1101110100111111_1111110110100011"; -- -0.13574232834771036
	pesos_i(10484) := b"1111111111111111_1111111111111111_1111011110101110_0011001000111110"; -- -0.03249822601973864
	pesos_i(10485) := b"1111111111111111_1111111111111111_1111011110001101_1111110101011001"; -- -0.03298965996192108
	pesos_i(10486) := b"0000000000000000_0000000000000000_0000000000000001_1101000111000100"; -- 2.7761826548372383e-05
	pesos_i(10487) := b"0000000000000000_0000000000000000_0001010010010110_0110100001100101"; -- 0.0804200407371532
	pesos_i(10488) := b"0000000000000000_0000000000000000_0010001101100001_0101100010001110"; -- 0.13820413087135835
	pesos_i(10489) := b"0000000000000000_0000000000000000_0000111101001101_0111111111111000"; -- 0.05977630423798344
	pesos_i(10490) := b"0000000000000000_0000000000000000_0000111100010001_1111111110101011"; -- 0.058868388314390736
	pesos_i(10491) := b"1111111111111111_1111111111111111_1110010100110111_1011000100100001"; -- -0.10461895893007345
	pesos_i(10492) := b"0000000000000000_0000000000000000_0001001111100011_0001000111001111"; -- 0.07768355652355784
	pesos_i(10493) := b"1111111111111111_1111111111111111_1111000001010000_0100111111111101"; -- -0.06127452921720891
	pesos_i(10494) := b"1111111111111111_1111111111111111_1110101011111011_0110001000001110"; -- -0.08210169953491712
	pesos_i(10495) := b"1111111111111111_1111111111111111_1101111110010100_1111000010110100"; -- -0.12663360220185493
	pesos_i(10496) := b"1111111111111111_1111111111111111_1111001100111010_1001011010011110"; -- -0.04988726273583273
	pesos_i(10497) := b"0000000000000000_0000000000000000_0000101110010100_0000110010011110"; -- 0.04522780285738968
	pesos_i(10498) := b"0000000000000000_0000000000000000_0000011000110001_0000101101100110"; -- 0.024185860059797355
	pesos_i(10499) := b"1111111111111111_1111111111111111_1110101010111111_0001111110101100"; -- -0.08302118351290004
	pesos_i(10500) := b"1111111111111111_1111111111111111_1110111000000011_0011011100001101"; -- -0.07026344230601685
	pesos_i(10501) := b"0000000000000000_0000000000000000_0000101101111001_1001111100001000"; -- 0.04482454245181992
	pesos_i(10502) := b"1111111111111111_1111111111111111_1111110000001010_0101110101001011"; -- -0.01546685136545092
	pesos_i(10503) := b"1111111111111111_1111111111111111_1110001110011110_0110010110111001"; -- -0.11086429823844615
	pesos_i(10504) := b"1111111111111111_1111111111111111_1110011000111000_1001110101111111"; -- -0.10069862033630289
	pesos_i(10505) := b"1111111111111111_1111111111111111_1110001000101110_1011011001110110"; -- -0.11647472012448003
	pesos_i(10506) := b"0000000000000000_0000000000000000_0001000011110110_1111110111011110"; -- 0.06626879366878498
	pesos_i(10507) := b"0000000000000000_0000000000000000_0000011001000111_1000011110011000"; -- 0.024528956080104157
	pesos_i(10508) := b"0000000000000000_0000000000000000_0001111101100100_0010111110101111"; -- 0.12262247102981211
	pesos_i(10509) := b"0000000000000000_0000000000000000_0010000100001001_1101111000010010"; -- 0.12905681558463
	pesos_i(10510) := b"1111111111111111_1111111111111111_1111011110010110_1000011111111000"; -- -0.032859327382813115
	pesos_i(10511) := b"0000000000000000_0000000000000000_0001000101110100_0000100001001001"; -- 0.06817676334218627
	pesos_i(10512) := b"1111111111111111_1111111111111111_1111010111000110_0101010110100011"; -- -0.0399424054704132
	pesos_i(10513) := b"1111111111111111_1111111111111111_1110010000011101_1110000111011001"; -- -0.10891903362458255
	pesos_i(10514) := b"0000000000000000_0000000000000000_0001110100011010_1001110010010001"; -- 0.11368731066893072
	pesos_i(10515) := b"1111111111111111_1111111111111111_1111110010001100_0101011010100111"; -- -0.013483604732540271
	pesos_i(10516) := b"0000000000000000_0000000000000000_0001000111001000_0101111100011100"; -- 0.06946367669005482
	pesos_i(10517) := b"1111111111111111_1111111111111111_1101111100101111_0110111110011110"; -- -0.1281824341212859
	pesos_i(10518) := b"0000000000000000_0000000000000000_0010111011011010_1111000000000011"; -- 0.1830282218457044
	pesos_i(10519) := b"1111111111111111_1111111111111111_1110110101100110_0101001001111010"; -- -0.07265743762736128
	pesos_i(10520) := b"1111111111111111_1111111111111111_1111001000110010_0100100000101000"; -- -0.05392025971036331
	pesos_i(10521) := b"1111111111111111_1111111111111111_1111001001001011_1000010101001011"; -- -0.0535351460088776
	pesos_i(10522) := b"1111111111111111_1111111111111111_1101100001011111_1001100111000011"; -- -0.15479125020915513
	pesos_i(10523) := b"1111111111111111_1111111111111111_1101111000001100_0110000100010011"; -- -0.13262360843163767
	pesos_i(10524) := b"1111111111111111_1111111111111111_1111010100011100_0001111000010100"; -- -0.04253971100818047
	pesos_i(10525) := b"1111111111111111_1111111111111111_1111000010111000_1010001101001111"; -- -0.05968264893864603
	pesos_i(10526) := b"0000000000000000_0000000000000000_0001010011101011_0110100101100000"; -- 0.08171709619770276
	pesos_i(10527) := b"0000000000000000_0000000000000000_0001010011111110_0010111011100111"; -- 0.082003527993938
	pesos_i(10528) := b"1111111111111111_1111111111111111_1110000001110111_0000000101101101"; -- -0.12318411909648551
	pesos_i(10529) := b"0000000000000000_0000000000000000_0001010000010011_1001101001011001"; -- 0.07842411682495029
	pesos_i(10530) := b"1111111111111111_1111111111111111_1111001110011011_1101110101011100"; -- -0.04840294370447897
	pesos_i(10531) := b"1111111111111111_1111111111111111_1101011010010010_1001100110001101"; -- -0.16182556448271698
	pesos_i(10532) := b"0000000000000000_0000000000000000_0001001111000101_1111000001100110"; -- 0.07723906022776228
	pesos_i(10533) := b"1111111111111111_1111111111111111_1110100100010100_0011101001101111"; -- -0.08953509129949053
	pesos_i(10534) := b"1111111111111111_1111111111111111_1111010001100000_0001000101101000"; -- -0.04540911867771258
	pesos_i(10535) := b"1111111111111111_1111111111111111_1110011111100111_0001111110001010"; -- -0.09412958977487214
	pesos_i(10536) := b"0000000000000000_0000000000000000_0001110011100001_1110011000110010"; -- 0.11282194829414356
	pesos_i(10537) := b"0000000000000000_0000000000000000_0010001111011011_0100001110111111"; -- 0.14006446273087914
	pesos_i(10538) := b"0000000000000000_0000000000000000_0001010101001001_1000101110011111"; -- 0.08315346359455345
	pesos_i(10539) := b"0000000000000000_0000000000000000_0000010001101001_1001100010101010"; -- 0.01723627238687436
	pesos_i(10540) := b"1111111111111111_1111111111111111_1111011010111101_0101111110100110"; -- -0.036172887721455625
	pesos_i(10541) := b"1111111111111111_1111111111111111_1110010101001100_1110111010010000"; -- -0.1042948626485982
	pesos_i(10542) := b"1111111111111111_1111111111111111_1101110101010101_1100111100100100"; -- -0.13540940629867118
	pesos_i(10543) := b"1111111111111111_1111111111111111_1101111011000111_0001010010010000"; -- -0.1297747754562747
	pesos_i(10544) := b"1111111111111111_1111111111111111_1110101000101100_0100011111001011"; -- -0.08526183409982338
	pesos_i(10545) := b"0000000000000000_0000000000000000_0000111001100000_1010111110100010"; -- 0.05616281220449291
	pesos_i(10546) := b"1111111111111111_1111111111111111_1110100110010000_0011010111100001"; -- -0.08764327298732046
	pesos_i(10547) := b"1111111111111111_1111111111111111_1111111101010010_0101000110100000"; -- -0.002650164137856987
	pesos_i(10548) := b"0000000000000000_0000000000000000_0010101000010111_1010110000100110"; -- 0.1644237129432065
	pesos_i(10549) := b"1111111111111111_1111111111111111_1110111011111100_1011111100100111"; -- -0.06645589161172057
	pesos_i(10550) := b"0000000000000000_0000000000000000_0001101100101110_0000110011100111"; -- 0.1061714234464844
	pesos_i(10551) := b"0000000000000000_0000000000000000_0001011111011100_0000100101101010"; -- 0.09320124475587335
	pesos_i(10552) := b"1111111111111111_1111111111111111_1111000000100101_0010010001100101"; -- -0.06193325543740656
	pesos_i(10553) := b"0000000000000000_0000000000000000_0001101000101011_1001000001011000"; -- 0.10222723141632324
	pesos_i(10554) := b"1111111111111111_1111111111111111_1111101101110010_0010111111101111"; -- -0.01778889098236779
	pesos_i(10555) := b"1111111111111111_1111111111111111_1101111010111110_0011110010000111"; -- -0.1299097223900456
	pesos_i(10556) := b"1111111111111111_1111111111111111_1110001001100001_0101100110100001"; -- -0.11570205517486586
	pesos_i(10557) := b"0000000000000000_0000000000000000_0000011111011011_0110100001101001"; -- 0.030691648161664312
	pesos_i(10558) := b"0000000000000000_0000000000000000_0000111001000101_0111001011011010"; -- 0.05574720208790888
	pesos_i(10559) := b"0000000000000000_0000000000000000_0000001111000011_1111110001110101"; -- 0.01470926138418163
	pesos_i(10560) := b"1111111111111111_1111111111111111_1101111110001101_1100111011100110"; -- -0.12674242868761806
	pesos_i(10561) := b"0000000000000000_0000000000000000_0000100001111011_0010111101001010"; -- 0.03312964981394603
	pesos_i(10562) := b"1111111111111111_1111111111111111_1101011111100111_1000111101110010"; -- -0.15662291982052565
	pesos_i(10563) := b"1111111111111111_1111111111111111_1110001010010010_1110100100000100"; -- -0.11494582790891918
	pesos_i(10564) := b"0000000000000000_0000000000000000_0000000011011010_1001011100101110"; -- 0.003335427016017909
	pesos_i(10565) := b"1111111111111111_1111111111111111_1110101001011011_0110001001100110"; -- -0.0845430852406321
	pesos_i(10566) := b"0000000000000000_0000000000000000_0010011010110010_0110011000000011"; -- 0.15115964491607753
	pesos_i(10567) := b"1111111111111111_1111111111111111_1101101001101110_0010111111110100"; -- -0.14675617499499102
	pesos_i(10568) := b"1111111111111111_1111111111111111_1110100001011011_1111001111011011"; -- -0.09234691525023003
	pesos_i(10569) := b"1111111111111111_1111111111111111_1110101010010111_0111100000100001"; -- -0.0836262626918405
	pesos_i(10570) := b"0000000000000000_0000000000000000_0001111111001011_1111110000010101"; -- 0.12420630942932118
	pesos_i(10571) := b"0000000000000000_0000000000000000_0001010110101100_0101010101101111"; -- 0.08466085405591536
	pesos_i(10572) := b"0000000000000000_0000000000000000_0010000010101111_0100000111100100"; -- 0.12767421555731148
	pesos_i(10573) := b"0000000000000000_0000000000000000_0000000110001110_1101110110110001"; -- 0.006086211850365119
	pesos_i(10574) := b"0000000000000000_0000000000000000_0000110011101111_0101100111000000"; -- 0.05052720008875197
	pesos_i(10575) := b"0000000000000000_0000000000000000_0001100001001111_1111001101110100"; -- 0.09496995537812204
	pesos_i(10576) := b"1111111111111111_1111111111111111_1111100011100111_0111011111110100"; -- -0.027718069861807814
	pesos_i(10577) := b"1111111111111111_1111111111111111_1111001000001111_1101101101001110"; -- -0.0544455466832285
	pesos_i(10578) := b"1111111111111111_1111111111111111_1111001011101100_1000011010011100"; -- -0.05107840254331019
	pesos_i(10579) := b"1111111111111111_1111111111111111_1110001011100010_1011001110100111"; -- -0.11372830550266633
	pesos_i(10580) := b"1111111111111111_1111111111111111_1101111101101100_1000111010111101"; -- -0.12724979283449822
	pesos_i(10581) := b"1111111111111111_1111111111111111_1101111110000110_1110101011001110"; -- -0.12684757676041372
	pesos_i(10582) := b"1111111111111111_1111111111111111_1110101000101101_0000001001101110"; -- -0.08525070977928578
	pesos_i(10583) := b"0000000000000000_0000000000000000_0000001001100111_1101001110111111"; -- 0.009396776215877166
	pesos_i(10584) := b"1111111111111111_1111111111111111_1101101000110100_0011101101101111"; -- -0.14764050048790947
	pesos_i(10585) := b"0000000000000000_0000000000000000_0001011000100000_0111010011001000"; -- 0.08643274188843877
	pesos_i(10586) := b"1111111111111111_1111111111111111_1111111010010101_1010001010001100"; -- -0.00552925189457237
	pesos_i(10587) := b"1111111111111111_1111111111111111_1110101000111100_1001100101101010"; -- -0.0850128283505181
	pesos_i(10588) := b"1111111111111111_1111111111111111_1111101000111001_0101101101110110"; -- -0.0225622974559755
	pesos_i(10589) := b"0000000000000000_0000000000000000_0001010111010110_1000001101100100"; -- 0.08530446228739944
	pesos_i(10590) := b"1111111111111111_1111111111111111_1101111100000010_0100011001000000"; -- -0.12887154508674922
	pesos_i(10591) := b"1111111111111111_1111111111111111_1110100110110101_1110111000001100"; -- -0.08706772041055547
	pesos_i(10592) := b"0000000000000000_0000000000000000_0001011001010111_1010011010000101"; -- 0.08727493993174776
	pesos_i(10593) := b"1111111111111111_1111111111111111_1110101000010001_1000101111111100"; -- -0.08566975694284894
	pesos_i(10594) := b"1111111111111111_1111111111111111_1110000111101000_0110100101001101"; -- -0.11754743463020687
	pesos_i(10595) := b"1111111111111111_1111111111111111_1110010100011101_1101111010010110"; -- -0.10501297791365287
	pesos_i(10596) := b"0000000000000000_0000000000000000_0010001010001000_1011010010010100"; -- 0.1348984586598935
	pesos_i(10597) := b"0000000000000000_0000000000000000_0000000011010111_0011101111100110"; -- 0.0032842097634871526
	pesos_i(10598) := b"1111111111111111_1111111111111111_1101110010111001_0011110011010011"; -- -0.13779849854091825
	pesos_i(10599) := b"1111111111111111_1111111111111111_1110010001001111_0110100100000000"; -- -0.1081632971178452
	pesos_i(10600) := b"0000000000000000_0000000000000000_0001001111110101_0111110010000101"; -- 0.07796457515829532
	pesos_i(10601) := b"1111111111111111_1111111111111111_1101111110101010_1111100010110111"; -- -0.12629743138063168
	pesos_i(10602) := b"0000000000000000_0000000000000000_0000000110011100_1010001111100001"; -- 0.0062963890407915935
	pesos_i(10603) := b"0000000000000000_0000000000000000_0001011111101111_0110111011010100"; -- 0.09349720656924833
	pesos_i(10604) := b"0000000000000000_0000000000000000_0000101001011001_0100100100110011"; -- 0.04042489535076344
	pesos_i(10605) := b"1111111111111111_1111111111111111_1101110111001101_1000001010000001"; -- -0.13358291971462083
	pesos_i(10606) := b"0000000000000000_0000000000000000_0000011010111001_0000010101001110"; -- 0.026260692270202626
	pesos_i(10607) := b"1111111111111111_1111111111111111_1110010111100100_1100100011100111"; -- -0.10197777147958895
	pesos_i(10608) := b"0000000000000000_0000000000000000_0010001111111011_1100000100110011"; -- 0.14056022156725087
	pesos_i(10609) := b"1111111111111111_1111111111111111_1101111100110011_0111110110001110"; -- -0.12812056811482578
	pesos_i(10610) := b"0000000000000000_0000000000000000_0000101001001111_0111111011011111"; -- 0.04027550654036009
	pesos_i(10611) := b"0000000000000000_0000000000000000_0001010011011100_1111001100110010"; -- 0.08149642915822936
	pesos_i(10612) := b"0000000000000000_0000000000000000_0000010101001000_0011011011101001"; -- 0.02063315570546525
	pesos_i(10613) := b"0000000000000000_0000000000000000_0010011110110111_1110011100001010"; -- 0.15514987945468758
	pesos_i(10614) := b"1111111111111111_1111111111111111_1110000111011101_0100101100100010"; -- -0.11771707938780629
	pesos_i(10615) := b"1111111111111111_1111111111111111_1110010001011101_0111000000000100"; -- -0.10794925587071753
	pesos_i(10616) := b"1111111111111111_1111111111111111_1110011010110111_0011111011000010"; -- -0.09876640095298729
	pesos_i(10617) := b"0000000000000000_0000000000000000_0001111011010001_0001011100010100"; -- 0.1203779624586384
	pesos_i(10618) := b"1111111111111111_1111111111111111_1110010101100110_0100100101010001"; -- -0.1039079835826187
	pesos_i(10619) := b"1111111111111111_1111111111111111_1110000111111000_0000111100100010"; -- -0.11730866833516766
	pesos_i(10620) := b"0000000000000000_0000000000000000_0001001111000001_1011101001011011"; -- 0.0771748038601782
	pesos_i(10621) := b"1111111111111111_1111111111111111_1111111111101011_1001011111101110"; -- -0.0003113788281615048
	pesos_i(10622) := b"1111111111111111_1111111111111111_1101110010111101_1000000011110011"; -- -0.137733402872921
	pesos_i(10623) := b"1111111111111111_1111111111111111_1111001010110100_0100001100110101"; -- -0.05193691220465826
	pesos_i(10624) := b"1111111111111111_1111111111111111_1101100011010111_0100110011001001"; -- -0.15296478369429742
	pesos_i(10625) := b"0000000000000000_0000000000000000_0010001110100001_1010001010111111"; -- 0.13918511553715152
	pesos_i(10626) := b"1111111111111111_1111111111111111_1110010110110010_1111000111010101"; -- -0.10273827133111156
	pesos_i(10627) := b"1111111111111111_1111111111111111_1110110000011110_0000011110110100"; -- -0.07766677715480735
	pesos_i(10628) := b"0000000000000000_0000000000000000_0001011001000010_0000100100111010"; -- 0.08694513000193259
	pesos_i(10629) := b"1111111111111111_1111111111111111_1101110111011011_1001110100001110"; -- -0.13336771399019917
	pesos_i(10630) := b"1111111111111111_1111111111111111_1110001000010111_1000000111111001"; -- -0.1168288009823252
	pesos_i(10631) := b"1111111111111111_1111111111111111_1111000100010100_0100111010011000"; -- -0.058283889569014855
	pesos_i(10632) := b"0000000000000000_0000000000000000_0001110011011010_1100111011100011"; -- 0.1127137473799656
	pesos_i(10633) := b"1111111111111111_1111111111111111_1111001110110011_1101110100100001"; -- -0.04803674641896685
	pesos_i(10634) := b"1111111111111111_1111111111111111_1111001010011011_1010110001001010"; -- -0.05231211854419166
	pesos_i(10635) := b"1111111111111111_1111111111111111_1111001110101000_0100011001011110"; -- -0.04821357912507127
	pesos_i(10636) := b"1111111111111111_1111111111111111_1110001110001100_0010001110000110"; -- -0.11114290213541134
	pesos_i(10637) := b"1111111111111111_1111111111111111_1111011011000110_0101010010001011"; -- -0.036036220580847475
	pesos_i(10638) := b"0000000000000000_0000000000000000_0000111011011111_1000001101111001"; -- 0.05809804628085468
	pesos_i(10639) := b"1111111111111111_1111111111111111_1110110001101000_0100010110101111"; -- -0.07653393249511532
	pesos_i(10640) := b"0000000000000000_0000000000000000_0001011111111011_1111011110001011"; -- 0.09368846084427696
	pesos_i(10641) := b"1111111111111111_1111111111111111_1110001011000010_0111000110110100"; -- -0.11422051769496205
	pesos_i(10642) := b"1111111111111111_1111111111111111_1111100111000001_0110100001011101"; -- -0.02439258321048986
	pesos_i(10643) := b"0000000000000000_0000000000000000_0000010100001100_1111110010111110"; -- 0.019729420185063826
	pesos_i(10644) := b"1111111111111111_1111111111111111_1101111000011110_0001000111110000"; -- -0.1323536672656405
	pesos_i(10645) := b"0000000000000000_0000000000000000_0000101010010101_0100000100011101"; -- 0.04133994055010862
	pesos_i(10646) := b"1111111111111111_1111111111111111_1110001011000100_1110101000110010"; -- -0.11418281819869346
	pesos_i(10647) := b"1111111111111111_1111111111111111_1101111000001110_1000000111111100"; -- -0.13259112926251468
	pesos_i(10648) := b"0000000000000000_0000000000000000_0000000100100111_0100001110010100"; -- 0.004505370744877941
	pesos_i(10649) := b"0000000000000000_0000000000000000_0000001101000010_1110001101111111"; -- 0.01273938986885703
	pesos_i(10650) := b"0000000000000000_0000000000000000_0001101011000001_0100100111101110"; -- 0.10451185275160645
	pesos_i(10651) := b"1111111111111111_1111111111111111_1101101111000010_0110110100110010"; -- -0.14156453642194602
	pesos_i(10652) := b"1111111111111111_1111111111111111_1101101110111010_1001001001100001"; -- -0.14168439044208578
	pesos_i(10653) := b"0000000000000000_0000000000000000_0000000011100000_0101111110010110"; -- 0.0034236660944359787
	pesos_i(10654) := b"1111111111111111_1111111111111111_1110110101101110_0101010001001011"; -- -0.07253525905768894
	pesos_i(10655) := b"0000000000000000_0000000000000000_0001110100110111_1011101001001110"; -- 0.1141315879708027
	pesos_i(10656) := b"1111111111111111_1111111111111111_1110111001011000_0000100011101101"; -- -0.06896919452645764
	pesos_i(10657) := b"1111111111111111_1111111111111111_1110100000100001_1101111011110100"; -- -0.09323317102998797
	pesos_i(10658) := b"1111111111111111_1111111111111111_1111101101110011_1010000100000110"; -- -0.017766891598028096
	pesos_i(10659) := b"0000000000000000_0000000000000000_0001010111000111_1000000000010111"; -- 0.08507538367940212
	pesos_i(10660) := b"1111111111111111_1111111111111111_1110100001110101_1001000011000001"; -- -0.09195609360913791
	pesos_i(10661) := b"0000000000000000_0000000000000000_0000111101010001_1100101110101000"; -- 0.05984185078992468
	pesos_i(10662) := b"0000000000000000_0000000000000000_0001011100010000_0111110101110001"; -- 0.09009536753601705
	pesos_i(10663) := b"1111111111111111_1111111111111111_1101111100010110_0001010110101110"; -- -0.12856926451122136
	pesos_i(10664) := b"1111111111111111_1111111111111111_1110011010011010_1100001110100110"; -- -0.09920098483357616
	pesos_i(10665) := b"0000000000000000_0000000000000000_0001111101001100_0000000011011010"; -- 0.12225346882346085
	pesos_i(10666) := b"0000000000000000_0000000000000000_0000011001100111_0110111100101100"; -- 0.0250157816647109
	pesos_i(10667) := b"1111111111111111_1111111111111111_1110011101001000_0000111011011001"; -- -0.09655673226756356
	pesos_i(10668) := b"1111111111111111_1111111111111111_1111001011001110_0000100010000100"; -- -0.05154368199699497
	pesos_i(10669) := b"1111111111111111_1111111111111111_1110100010010001_0101000010111100"; -- -0.09153266349722389
	pesos_i(10670) := b"0000000000000000_0000000000000000_0001000001000111_1100011100000010"; -- 0.06359523578345755
	pesos_i(10671) := b"1111111111111111_1111111111111111_1111100110101110_0111100101110011"; -- -0.024681481657209115
	pesos_i(10672) := b"1111111111111111_1111111111111111_1101110100010100_1001110000110000"; -- -0.13640426469210906
	pesos_i(10673) := b"0000000000000000_0000000000000000_0001000100001100_1100100010010010"; -- 0.06660131034575384
	pesos_i(10674) := b"0000000000000000_0000000000000000_0001110001110010_1011010101011101"; -- 0.11112531215766679
	pesos_i(10675) := b"0000000000000000_0000000000000000_0000110010101111_0101011011000010"; -- 0.04955045922231694
	pesos_i(10676) := b"1111111111111111_1111111111111111_1110110111111100_1101011100000110"; -- -0.0703607187414945
	pesos_i(10677) := b"0000000000000000_0000000000000000_0000101100101110_0010001110011000"; -- 0.043672775903927645
	pesos_i(10678) := b"0000000000000000_0000000000000000_0010001100111110_0011011110011000"; -- 0.13766810845537095
	pesos_i(10679) := b"0000000000000000_0000000000000000_0000000010111101_0101100101000010"; -- 0.0028892313650729787
	pesos_i(10680) := b"1111111111111111_1111111111111111_1111000110010110_0110110111010110"; -- -0.056298384973218554
	pesos_i(10681) := b"0000000000000000_0000000000000000_0000110111111110_0111011011010001"; -- 0.05466406442940842
	pesos_i(10682) := b"0000000000000000_0000000000000000_0000011100100100_0110111100000100"; -- 0.027899683448670633
	pesos_i(10683) := b"0000000000000000_0000000000000000_0000110010111010_1111000101101111"; -- 0.04972752524097766
	pesos_i(10684) := b"0000000000000000_0000000000000000_0001111101010010_1110101101110101"; -- 0.12235900507446308
	pesos_i(10685) := b"1111111111111111_1111111111111111_1111101001000111_0110101001010101"; -- -0.022347788174902416
	pesos_i(10686) := b"0000000000000000_0000000000000000_0001111000000001_0010110001111110"; -- 0.11720541081919245
	pesos_i(10687) := b"0000000000000000_0000000000000000_0000011000011111_0000111111101111"; -- 0.023911472168141674
	pesos_i(10688) := b"0000000000000000_0000000000000000_0000100001000011_0111011101110110"; -- 0.03227945937941576
	pesos_i(10689) := b"1111111111111111_1111111111111111_1101101011111010_1011100001011001"; -- -0.14461181479865334
	pesos_i(10690) := b"0000000000000000_0000000000000000_0001011011001000_1001111101100011"; -- 0.08899875794443944
	pesos_i(10691) := b"1111111111111111_1111111111111111_1111000111000100_1000000000101111"; -- -0.05559538696336933
	pesos_i(10692) := b"1111111111111111_1111111111111111_1111001001001000_0001010001100000"; -- -0.053587652642618694
	pesos_i(10693) := b"0000000000000000_0000000000000000_0001101000111010_0101100000111000"; -- 0.10245276804876327
	pesos_i(10694) := b"0000000000000000_0000000000000000_0000011001111000_1010101110101111"; -- 0.025278787795148402
	pesos_i(10695) := b"0000000000000000_0000000000000000_0000100111000110_1111100101111000"; -- 0.03819235971866329
	pesos_i(10696) := b"1111111111111111_1111111111111111_1111101111101100_1101010011100000"; -- -0.015917487552761553
	pesos_i(10697) := b"0000000000000000_0000000000000000_0001011111000111_0110100000110111"; -- 0.09288646072341816
	pesos_i(10698) := b"0000000000000000_0000000000000000_0001110011000010_0000101010001100"; -- 0.11233583378758907
	pesos_i(10699) := b"0000000000000000_0000000000000000_0000000001111110_1001010100011000"; -- 0.001931494175741357
	pesos_i(10700) := b"0000000000000000_0000000000000000_0000010001101100_1111001001110011"; -- 0.017287400227626037
	pesos_i(10701) := b"1111111111111111_1111111111111111_1101100111111010_1001010100010111"; -- -0.14852016629851003
	pesos_i(10702) := b"0000000000000000_0000000000000000_0010010000001001_0011101011000010"; -- 0.14076583137007684
	pesos_i(10703) := b"0000000000000000_0000000000000000_0001101111010101_1110001101110000"; -- 0.1087324285131567
	pesos_i(10704) := b"0000000000000000_0000000000000000_0001111111110010_0110000101010111"; -- 0.12479217883859589
	pesos_i(10705) := b"1111111111111111_1111111111111111_1110000011111100_1111001110010011"; -- -0.12114026705631832
	pesos_i(10706) := b"0000000000000000_0000000000000000_0001011101110011_1111000101010001"; -- 0.09161289432798492
	pesos_i(10707) := b"0000000000000000_0000000000000000_0000100011110111_1001101010101000"; -- 0.03502813909603654
	pesos_i(10708) := b"1111111111111111_1111111111111111_1110001101100100_0000101010110100"; -- -0.111754733105913
	pesos_i(10709) := b"0000000000000000_0000000000000000_0000010010101010_0111001000000100"; -- 0.0182257899987464
	pesos_i(10710) := b"1111111111111111_1111111111111111_1101111111110110_1001000110011100"; -- -0.12514390892324853
	pesos_i(10711) := b"0000000000000000_0000000000000000_0000000111011001_1101111001001110"; -- 0.007230657709492147
	pesos_i(10712) := b"0000000000000000_0000000000000000_0001110101011101_0111111010101100"; -- 0.11470786764915147
	pesos_i(10713) := b"1111111111111111_1111111111111111_1110000111101100_0000111110001110"; -- -0.11749174865868947
	pesos_i(10714) := b"0000000000000000_0000000000000000_0001110000001011_1101000101001101"; -- 0.10955532199121641
	pesos_i(10715) := b"1111111111111111_1111111111111111_1111011000010100_0010111011110011"; -- -0.03875452585358255
	pesos_i(10716) := b"1111111111111111_1111111111111111_1111001010000110_0100010010001010"; -- -0.05263873700079218
	pesos_i(10717) := b"1111111111111111_1111111111111111_1110001010000100_0011011110101000"; -- -0.11517002244472183
	pesos_i(10718) := b"1111111111111111_1111111111111111_1110001110010111_0110010010001101"; -- -0.11097117956963069
	pesos_i(10719) := b"0000000000000000_0000000000000000_0010000101101100_1100100000100001"; -- 0.1305661279009875
	pesos_i(10720) := b"0000000000000000_0000000000000000_0001100010100100_0011110011001111"; -- 0.09625606589443243
	pesos_i(10721) := b"1111111111111111_1111111111111111_1110011100010011_0001100010001100"; -- -0.09736486996855177
	pesos_i(10722) := b"1111111111111111_1111111111111111_1110101101001111_0111000001111101"; -- -0.08081910077586636
	pesos_i(10723) := b"0000000000000000_0000000000000000_0001010001011001_0100010111101001"; -- 0.07948719923466713
	pesos_i(10724) := b"0000000000000000_0000000000000000_0010001101101001_0000111100001011"; -- 0.13832181936719695
	pesos_i(10725) := b"1111111111111111_1111111111111111_1101011011111110_0010001111001000"; -- -0.16018463486904722
	pesos_i(10726) := b"0000000000000000_0000000000000000_0001011100111001_1101101100111100"; -- 0.09072656832560416
	pesos_i(10727) := b"0000000000000000_0000000000000000_0001101000010011_0011001000010011"; -- 0.10185540159255516
	pesos_i(10728) := b"1111111111111111_1111111111111111_1110001101111000_1111111110100001"; -- -0.11143495869553328
	pesos_i(10729) := b"1111111111111111_1111111111111111_1111011110000101_1000110011011010"; -- -0.03311843566177174
	pesos_i(10730) := b"0000000000000000_0000000000000000_0000101110011110_1110110011110100"; -- 0.04539376220109065
	pesos_i(10731) := b"1111111111111111_1111111111111111_1111110101000011_0010001001011110"; -- -0.010694362704219708
	pesos_i(10732) := b"1111111111111111_1111111111111111_1110000011001010_1111100010100101"; -- -0.12190290426917641
	pesos_i(10733) := b"0000000000000000_0000000000000000_0010000011010000_1110111011101010"; -- 0.1281880686192765
	pesos_i(10734) := b"1111111111111111_1111111111111111_1110111000011011_1100001110001101"; -- -0.06988885700598346
	pesos_i(10735) := b"1111111111111111_1111111111111111_1110110100011110_1100110010011011"; -- -0.0737487909705582
	pesos_i(10736) := b"0000000000000000_0000000000000000_0001011000000010_1000111010000111"; -- 0.08597651280094463
	pesos_i(10737) := b"1111111111111111_1111111111111111_1101100100111010_1000000110111001"; -- -0.15145100824527533
	pesos_i(10738) := b"0000000000000000_0000000000000000_0010010100010010_1110010001101010"; -- 0.14481952284145824
	pesos_i(10739) := b"1111111111111111_1111111111111111_1111001011110001_0001010010000000"; -- -0.0510089100552754
	pesos_i(10740) := b"1111111111111111_1111111111111111_1111110101110111_1011110110000000"; -- -0.009891659115910409
	pesos_i(10741) := b"0000000000000000_0000000000000000_0010010000101111_1010100011000010"; -- 0.14135222177934342
	pesos_i(10742) := b"0000000000000000_0000000000000000_0001100000101101_1101110110000010"; -- 0.09444984828635136
	pesos_i(10743) := b"0000000000000000_0000000000000000_0001100100110111_1100010100001111"; -- 0.09850722897964143
	pesos_i(10744) := b"0000000000000000_0000000000000000_0000110101001101_1011000010101010"; -- 0.051966706742929004
	pesos_i(10745) := b"1111111111111111_1111111111111111_1111011110111101_1011100110100000"; -- -0.032261274821821666
	pesos_i(10746) := b"0000000000000000_0000000000000000_0001110001100011_0010100000100100"; -- 0.11088801258634337
	pesos_i(10747) := b"0000000000000000_0000000000000000_0010000011000001_1000101001110101"; -- 0.1279531989742064
	pesos_i(10748) := b"1111111111111111_1111111111111111_1111010101001000_0011001000110010"; -- -0.041867125414522796
	pesos_i(10749) := b"0000000000000000_0000000000000000_0000001101110010_1110010000011111"; -- 0.013471849130038908
	pesos_i(10750) := b"0000000000000000_0000000000000000_0001101011101011_0011111010111111"; -- 0.10515205550444882
	pesos_i(10751) := b"1111111111111111_1111111111111111_1110000100100000_0011111010010001"; -- -0.12060173942502642
	pesos_i(10752) := b"0000000000000000_0000000000000000_0010001100000011_1010001010010111"; -- 0.1367742175863897
	pesos_i(10753) := b"0000000000000000_0000000000000000_0001011001111101_1001000010001011"; -- 0.0878534640767473
	pesos_i(10754) := b"1111111111111111_1111111111111111_1110000000100110_1000101000111000"; -- -0.12441192750640674
	pesos_i(10755) := b"0000000000000000_0000000000000000_0010011000011110_0111110101011000"; -- 0.14890273479703758
	pesos_i(10756) := b"0000000000000000_0000000000000000_0000111110001100_1000100101111000"; -- 0.060738174148981236
	pesos_i(10757) := b"0000000000000000_0000000000000000_0001001111011100_0011111011011100"; -- 0.0775794302447638
	pesos_i(10758) := b"0000000000000000_0000000000000000_0001010110101000_1101000101011110"; -- 0.08460720582717901
	pesos_i(10759) := b"0000000000000000_0000000000000000_0001011010001101_0010010110001101"; -- 0.08809122751360249
	pesos_i(10760) := b"1111111111111111_1111111111111111_1101111111011101_1101011011001001"; -- -0.12552125533001307
	pesos_i(10761) := b"1111111111111111_1111111111111111_1111011100010100_0101000010011011"; -- -0.03484626985748887
	pesos_i(10762) := b"1111111111111111_1111111111111111_1110001101100011_0001100100011110"; -- -0.11176913285678153
	pesos_i(10763) := b"1111111111111111_1111111111111111_1110001101101001_0011110111000001"; -- -0.11167539622938992
	pesos_i(10764) := b"0000000000000000_0000000000000000_0001010110111101_1010010111111011"; -- 0.08492505429213146
	pesos_i(10765) := b"1111111111111111_1111111111111111_1101100010100010_1101010110101011"; -- -0.15376534066040712
	pesos_i(10766) := b"0000000000000000_0000000000000000_0001100110010010_0100110111011101"; -- 0.09988867431265921
	pesos_i(10767) := b"1111111111111111_1111111111111111_1110110110000001_0010100101100011"; -- -0.07224789940414722
	pesos_i(10768) := b"0000000000000000_0000000000000000_0001000010001101_0100110000111001"; -- 0.06465603257324391
	pesos_i(10769) := b"1111111111111111_1111111111111111_1110111110000010_0011110111110110"; -- -0.06441891421223564
	pesos_i(10770) := b"1111111111111111_1111111111111111_1110110110100010_0011110010011110"; -- -0.07174321317455942
	pesos_i(10771) := b"1111111111111111_1111111111111111_1110011100011110_0001111001101101"; -- -0.09719667285005974
	pesos_i(10772) := b"1111111111111111_1111111111111111_1101110110010110_1100100101001110"; -- -0.13441793303771998
	pesos_i(10773) := b"1111111111111111_1111111111111111_1111111000100001_1010000100010011"; -- -0.007299359148707704
	pesos_i(10774) := b"1111111111111111_1111111111111111_1110110110111011_1000111111010011"; -- -0.07135678390011545
	pesos_i(10775) := b"0000000000000000_0000000000000000_0001110001010001_1111111000111001"; -- 0.1106261147761014
	pesos_i(10776) := b"1111111111111111_1111111111111111_1101101001100000_0101011111111001"; -- -0.14696741256360427
	pesos_i(10777) := b"0000000000000000_0000000000000000_0001100001100100_0110001111000101"; -- 0.09528182562882584
	pesos_i(10778) := b"0000000000000000_0000000000000000_0000011111101000_0000110010101010"; -- 0.030884543839096616
	pesos_i(10779) := b"1111111111111111_1111111111111111_1111001001010011_0000001001000001"; -- -0.05342088611793654
	pesos_i(10780) := b"1111111111111111_1111111111111111_1101100010111011_1100100010001011"; -- -0.1533846532100492
	pesos_i(10781) := b"0000000000000000_0000000000000000_0000101100111010_1100101111111011"; -- 0.04386591789310484
	pesos_i(10782) := b"1111111111111111_1111111111111111_1111111000010000_0010010001111001"; -- -0.007566185443657876
	pesos_i(10783) := b"0000000000000000_0000000000000000_0000111100100101_0100010110001100"; -- 0.05916247058626804
	pesos_i(10784) := b"0000000000000000_0000000000000000_0000000100111000_0100011000111000"; -- 0.004764927445599797
	pesos_i(10785) := b"0000000000000000_0000000000000000_0001110001011100_1011000010100110"; -- 0.11078933776358618
	pesos_i(10786) := b"0000000000000000_0000000000000000_0001111001011100_0111000101101000"; -- 0.11859806822624012
	pesos_i(10787) := b"1111111111111111_1111111111111111_1110000101111101_0011100110111000"; -- -0.11918296114990831
	pesos_i(10788) := b"0000000000000000_0000000000000000_0001101010011110_1100101001100100"; -- 0.10398545199249253
	pesos_i(10789) := b"1111111111111111_1111111111111111_1101101111001101_1000010001001011"; -- -0.1413953129869888
	pesos_i(10790) := b"0000000000000000_0000000000000000_0001010101000110_0110101111110100"; -- 0.08310579966257653
	pesos_i(10791) := b"1111111111111111_1111111111111111_1110111110111000_1010011101011111"; -- -0.0635886567751491
	pesos_i(10792) := b"1111111111111111_1111111111111111_1111010010011111_1010001101101100"; -- -0.04443911186978609
	pesos_i(10793) := b"0000000000000000_0000000000000000_0000100011100110_0000110100101110"; -- 0.03476030701825078
	pesos_i(10794) := b"0000000000000000_0000000000000000_0000111101111000_0000100011000011"; -- 0.06042532697051708
	pesos_i(10795) := b"0000000000000000_0000000000000000_0000001010011110_0001110100010000"; -- 0.010225120877661694
	pesos_i(10796) := b"1111111111111111_1111111111111111_1110110101001000_1111001100001100"; -- -0.07310563052520982
	pesos_i(10797) := b"0000000000000000_0000000000000000_0001010010010011_0000100001010111"; -- 0.08036853903996663
	pesos_i(10798) := b"1111111111111111_1111111111111111_1110001001001101_1001011010000100"; -- -0.11600360172334605
	pesos_i(10799) := b"0000000000000000_0000000000000000_0001101011000110_1111110100010110"; -- 0.10459882541169574
	pesos_i(10800) := b"1111111111111111_1111111111111111_1111001001101101_1001011110010101"; -- -0.053015257071088874
	pesos_i(10801) := b"0000000000000000_0000000000000000_0001100010011010_1010110011000001"; -- 0.09611015040666558
	pesos_i(10802) := b"1111111111111111_1111111111111111_1101111100010010_0000101010010100"; -- -0.12863096126999646
	pesos_i(10803) := b"0000000000000000_0000000000000000_0001000100111011_1001001101000111"; -- 0.06731529700163551
	pesos_i(10804) := b"0000000000000000_0000000000000000_0000000100111111_1011010001100011"; -- 0.004878305713285479
	pesos_i(10805) := b"0000000000000000_0000000000000000_0000110011101110_0111000000101110"; -- 0.05051327813914467
	pesos_i(10806) := b"1111111111111111_1111111111111111_1111100010110011_0000101001100010"; -- -0.028518057855658575
	pesos_i(10807) := b"1111111111111111_1111111111111111_1101110111101100_0011111001001101"; -- -0.1331139623147788
	pesos_i(10808) := b"1111111111111111_1111111111111111_1110001011101000_1011011011100011"; -- -0.11363656013097168
	pesos_i(10809) := b"0000000000000000_0000000000000000_0010010011101000_1011101001111001"; -- 0.14417615377000167
	pesos_i(10810) := b"0000000000000000_0000000000000000_0000100000100111_1000101110110111"; -- 0.03185342034308026
	pesos_i(10811) := b"0000000000000000_0000000000000000_0001101101001001_0000101011110010"; -- 0.10658329388632805
	pesos_i(10812) := b"1111111111111111_1111111111111111_1111000001001101_1110100001000001"; -- -0.06131122988223809
	pesos_i(10813) := b"0000000000000000_0000000000000000_0000101110100000_0000001011010010"; -- 0.04541032442547569
	pesos_i(10814) := b"1111111111111111_1111111111111111_1110001100000001_0010110010001010"; -- -0.11326333644071579
	pesos_i(10815) := b"1111111111111111_1111111111111111_1110010100011101_0100110101011000"; -- -0.10502163510794987
	pesos_i(10816) := b"0000000000000000_0000000000000000_0001000010100111_0110001100110000"; -- 0.06505412977963951
	pesos_i(10817) := b"1111111111111111_1111111111111111_1111110000000010_0001001011110000"; -- -0.015593353560867046
	pesos_i(10818) := b"1111111111111111_1111111111111111_1110011111101100_1000000110010000"; -- -0.09404745331356355
	pesos_i(10819) := b"1111111111111111_1111111111111111_1111110100000001_1011001001100010"; -- -0.01169285886336849
	pesos_i(10820) := b"0000000000000000_0000000000000000_0001111001011000_1010100001111010"; -- 0.11854031535813664
	pesos_i(10821) := b"1111111111111111_1111111111111111_1110110011110111_1001101110101010"; -- -0.07434680088919972
	pesos_i(10822) := b"1111111111111111_1111111111111111_1110100011111001_0011000001100011"; -- -0.08994767738193188
	pesos_i(10823) := b"0000000000000000_0000000000000000_0001110001110100_0011011000100010"; -- 0.11114824610764922
	pesos_i(10824) := b"1111111111111111_1111111111111111_1111001010111010_1010011100010101"; -- -0.05183940646475957
	pesos_i(10825) := b"1111111111111111_1111111111111111_1110111101101011_0011001101011000"; -- -0.06477049921305106
	pesos_i(10826) := b"0000000000000000_0000000000000000_0010001001001001_0011100100111000"; -- 0.1339298020539441
	pesos_i(10827) := b"1111111111111111_1111111111111111_1101101101100010_1111111010100011"; -- -0.14302071109647396
	pesos_i(10828) := b"0000000000000000_0000000000000000_0000001010111111_1010111110001011"; -- 0.010737391940317614
	pesos_i(10829) := b"1111111111111111_1111111111111111_1101111100001100_0000011010011000"; -- -0.1287227514304742
	pesos_i(10830) := b"0000000000000000_0000000000000000_0000101001000110_1010010111010001"; -- 0.04014049872616343
	pesos_i(10831) := b"0000000000000000_0000000000000000_0000010111010100_0111111111111101"; -- 0.022773742047396833
	pesos_i(10832) := b"0000000000000000_0000000000000000_0000000010101101_0100001011100110"; -- 0.002643758072593677
	pesos_i(10833) := b"1111111111111111_1111111111111111_1110001111110101_1000111111000011"; -- -0.10953427775025283
	pesos_i(10834) := b"1111111111111111_1111111111111111_1111001001110110_0011001110111001"; -- -0.052883879991360745
	pesos_i(10835) := b"1111111111111111_1111111111111111_1110000011110101_1100011101000001"; -- -0.12124972012324071
	pesos_i(10836) := b"0000000000000000_0000000000000000_0000000110111111_0100001111010011"; -- 0.006824721401650284
	pesos_i(10837) := b"0000000000000000_0000000000000000_0000101100111100_0010111111001011"; -- 0.043887126042161106
	pesos_i(10838) := b"1111111111111111_1111111111111111_1101110101100000_1100110011010010"; -- -0.13524169805014022
	pesos_i(10839) := b"0000000000000000_0000000000000000_0000100011010000_0110111101110110"; -- 0.034430471691298425
	pesos_i(10840) := b"0000000000000000_0000000000000000_0001010001110000_0111010111111010"; -- 0.07984101629119111
	pesos_i(10841) := b"1111111111111111_1111111111111111_1111111101011111_1001001110001100"; -- -0.002447870516793653
	pesos_i(10842) := b"0000000000000000_0000000000000000_0010000101100011_1001010001001000"; -- 0.13042570829794956
	pesos_i(10843) := b"1111111111111111_1111111111111111_1111110101010110_0010001010111111"; -- -0.010404423185704297
	pesos_i(10844) := b"0000000000000000_0000000000000000_0001010101111000_1110101010001101"; -- 0.08387628492596232
	pesos_i(10845) := b"0000000000000000_0000000000000000_0001101010110110_0000010000001110"; -- 0.10433984119808559
	pesos_i(10846) := b"1111111111111111_1111111111111111_1110110011001001_1110111011100011"; -- -0.07504374463255219
	pesos_i(10847) := b"1111111111111111_1111111111111111_1110110110001111_1001100111010110"; -- -0.0720275737961885
	pesos_i(10848) := b"1111111111111111_1111111111111111_1110010010110100_0100001010100110"; -- -0.10662444536692929
	pesos_i(10849) := b"0000000000000000_0000000000000000_0001101111001100_1111111111110100"; -- 0.10859679906268122
	pesos_i(10850) := b"0000000000000000_0000000000000000_0000001101010001_1001010000100010"; -- 0.012963541319594171
	pesos_i(10851) := b"1111111111111111_1111111111111111_1111011111101001_0001111111111010"; -- -0.03159904610007309
	pesos_i(10852) := b"0000000000000000_0000000000000000_0000110011110100_0110101010011101"; -- 0.05060449908719733
	pesos_i(10853) := b"1111111111111111_1111111111111111_1110000000010100_1101010110110000"; -- -0.12468208749286272
	pesos_i(10854) := b"1111111111111111_1111111111111111_1111000010011110_0010100100100110"; -- -0.060086658620712816
	pesos_i(10855) := b"0000000000000000_0000000000000000_0000000011110001_0001100000100010"; -- 0.0036788065092058135
	pesos_i(10856) := b"1111111111111111_1111111111111111_1111011100010001_1010100110111111"; -- -0.034886732951860455
	pesos_i(10857) := b"0000000000000000_0000000000000000_0001010100000110_1100011110010110"; -- 0.08213469905562902
	pesos_i(10858) := b"1111111111111111_1111111111111111_1110000100000000_1000100100011100"; -- -0.12108557772330533
	pesos_i(10859) := b"1111111111111111_1111111111111111_1111101011100000_0011010010010011"; -- -0.020016397692695562
	pesos_i(10860) := b"0000000000000000_0000000000000000_0001011001011000_1000101100100000"; -- 0.08728856599842758
	pesos_i(10861) := b"0000000000000000_0000000000000000_0001111110010000_1110101010100001"; -- 0.12330500058126304
	pesos_i(10862) := b"0000000000000000_0000000000000000_0000110001011100_1010110011101011"; -- 0.04828911529194229
	pesos_i(10863) := b"0000000000000000_0000000000000000_0001000110000100_1010010010101101"; -- 0.0684302256106724
	pesos_i(10864) := b"1111111111111111_1111111111111111_1101101100011111_0100100000000111"; -- -0.14405393436526429
	pesos_i(10865) := b"1111111111111111_1111111111111111_1110001000100111_0000110101000101"; -- -0.11659161632750077
	pesos_i(10866) := b"0000000000000000_0000000000000000_0010001010111011_0000111100001101"; -- 0.13566679069031426
	pesos_i(10867) := b"0000000000000000_0000000000000000_0001110010100100_1101111101110011"; -- 0.1118907600493629
	pesos_i(10868) := b"0000000000000000_0000000000000000_0000010110001111_1011101011110010"; -- 0.021724399548435733
	pesos_i(10869) := b"1111111111111111_1111111111111111_1110111100111001_1110001010000000"; -- -0.06552299852046423
	pesos_i(10870) := b"1111111111111111_1111111111111111_1111001100010100_0100011110000110"; -- -0.05047181110330254
	pesos_i(10871) := b"1111111111111111_1111111111111111_1111010101000010_0000001011000011"; -- -0.04196150529512275
	pesos_i(10872) := b"0000000000000000_0000000000000000_0010010100000101_0100101001011110"; -- 0.14461197646190568
	pesos_i(10873) := b"1111111111111111_1111111111111111_1101101001001000_1100001001001010"; -- -0.14732728658676883
	pesos_i(10874) := b"1111111111111111_1111111111111111_1101111011111011_0111001010111111"; -- -0.12897570445809245
	pesos_i(10875) := b"1111111111111111_1111111111111111_1111110111110100_1100100101001011"; -- -0.007983607546154457
	pesos_i(10876) := b"1111111111111111_1111111111111111_1110111001101100_0101011110111000"; -- -0.0686593223836003
	pesos_i(10877) := b"0000000000000000_0000000000000000_0001110110101010_1001001110011111"; -- 0.11588404307247417
	pesos_i(10878) := b"1111111111111111_1111111111111111_1110111011111000_1111000000010010"; -- -0.06651401103731956
	pesos_i(10879) := b"1111111111111111_1111111111111111_1111101111011001_1000011110010110"; -- -0.016212011280977434
	pesos_i(10880) := b"1111111111111111_1111111111111111_1110011100011110_1001101101011000"; -- -0.09718922717428677
	pesos_i(10881) := b"0000000000000000_0000000000000000_0010001011001000_0000101111110110"; -- 0.13586497063847858
	pesos_i(10882) := b"0000000000000000_0000000000000000_0000101011000010_1100111100101111"; -- 0.04203505417190535
	pesos_i(10883) := b"1111111111111111_1111111111111111_1111111011011011_1001001000001000"; -- -0.004462121087662454
	pesos_i(10884) := b"1111111111111111_1111111111111111_1111000100001110_0011001101000100"; -- -0.05837707134861494
	pesos_i(10885) := b"1111111111111111_1111111111111111_1101110110111010_1111011001001110"; -- -0.13386593427182125
	pesos_i(10886) := b"1111111111111111_1111111111111111_1110110101101101_1011101000010111"; -- -0.07254445025934349
	pesos_i(10887) := b"0000000000000000_0000000000000000_0000101001000110_0100000000100110"; -- 0.04013443879128389
	pesos_i(10888) := b"0000000000000000_0000000000000000_0010001110010111_0101100101010101"; -- 0.13902815184025571
	pesos_i(10889) := b"1111111111111111_1111111111111111_1111000111111101_1011010111101000"; -- -0.05472243394520389
	pesos_i(10890) := b"0000000000000000_0000000000000000_0001100010111111_1001111011010011"; -- 0.09667389532627754
	pesos_i(10891) := b"0000000000000000_0000000000000000_0010011100001101_0110101010100010"; -- 0.15254847002851435
	pesos_i(10892) := b"1111111111111111_1111111111111111_1111111001011110_1001110111010101"; -- -0.006368766203748149
	pesos_i(10893) := b"1111111111111111_1111111111111111_1111010111111011_0111100000000011"; -- -0.039131640579319386
	pesos_i(10894) := b"1111111111111111_1111111111111111_1111110110000110_0101101001011101"; -- -0.009668686161211491
	pesos_i(10895) := b"0000000000000000_0000000000000000_0001010001001100_1011101101100001"; -- 0.07929583668707313
	pesos_i(10896) := b"0000000000000000_0000000000000000_0000000011111111_1101100010001001"; -- 0.003903897781753449
	pesos_i(10897) := b"0000000000000000_0000000000000000_0000100011100011_1100001001110011"; -- 0.03472533509555245
	pesos_i(10898) := b"1111111111111111_1111111111111111_1111101101000010_1111011001111101"; -- -0.018509478151596495
	pesos_i(10899) := b"0000000000000000_0000000000000000_0001001111110001_1100111001111011"; -- 0.07790842535198851
	pesos_i(10900) := b"1111111111111111_1111111111111111_1110000011001010_0011101011010000"; -- -0.12191421917861345
	pesos_i(10901) := b"1111111111111111_1111111111111111_1101110110110101_1111000110110010"; -- -0.1339425030167086
	pesos_i(10902) := b"0000000000000000_0000000000000000_0000101000100101_0111010111001001"; -- 0.039634095624244095
	pesos_i(10903) := b"0000000000000000_0000000000000000_0010010001110010_1100000011100011"; -- 0.1423759989846298
	pesos_i(10904) := b"1111111111111111_1111111111111111_1111011010110000_1101000110001101"; -- -0.03636446292071748
	pesos_i(10905) := b"0000000000000000_0000000000000000_0001111011111001_0001011001000110"; -- 0.12098826610683598
	pesos_i(10906) := b"0000000000000000_0000000000000000_0000010011011010_0100010101010001"; -- 0.018955547598494465
	pesos_i(10907) := b"1111111111111111_1111111111111111_1111010010011000_1101110000000000"; -- -0.04454255094073801
	pesos_i(10908) := b"0000000000000000_0000000000000000_0010100010101110_1010100000100011"; -- 0.158915051042318
	pesos_i(10909) := b"0000000000000000_0000000000000000_0010000111101111_1111011001011101"; -- 0.13256778495726987
	pesos_i(10910) := b"1111111111111111_1111111111111111_1111001101101010_1111100101101001"; -- -0.04914895241558863
	pesos_i(10911) := b"0000000000000000_0000000000000000_0000110001111111_1110000100101001"; -- 0.04882628681896677
	pesos_i(10912) := b"1111111111111111_1111111111111111_1111011000010010_1111011000011110"; -- -0.03877317212256787
	pesos_i(10913) := b"1111111111111111_1111111111111111_1101011111011111_1111111010110100"; -- -0.15673835852403564
	pesos_i(10914) := b"1111111111111111_1111111111111111_1110000110011000_0110101101110110"; -- -0.11876800897731213
	pesos_i(10915) := b"0000000000000000_0000000000000000_0000100111011101_1101000001000011"; -- 0.03854085574400519
	pesos_i(10916) := b"1111111111111111_1111111111111111_1110011100111101_1101011000010110"; -- -0.09671270333937718
	pesos_i(10917) := b"0000000000000000_0000000000000000_0000111001100111_1110110100010111"; -- 0.05627328698597428
	pesos_i(10918) := b"1111111111111111_1111111111111111_1101110001100001_0111110001000111"; -- -0.13913749004070053
	pesos_i(10919) := b"1111111111111111_1111111111111111_1110000001010101_0100101001110010"; -- -0.12369856569813947
	pesos_i(10920) := b"1111111111111111_1111111111111111_1110000111010001_0110011110100010"; -- -0.11789848601645751
	pesos_i(10921) := b"1111111111111111_1111111111111111_1101100010100110_1111000110100000"; -- -0.15370263897408873
	pesos_i(10922) := b"0000000000000000_0000000000000000_0001110000111110_0010001111010100"; -- 0.11032318039426793
	pesos_i(10923) := b"1111111111111111_1111111111111111_1111111111101101_1101100010001011"; -- -0.00027700995281387233
	pesos_i(10924) := b"0000000000000000_0000000000000000_0001100000000111_0101011110001000"; -- 0.09386202887450314
	pesos_i(10925) := b"1111111111111111_1111111111111111_1111100000101000_1011101110101011"; -- -0.0306284625320225
	pesos_i(10926) := b"0000000000000000_0000000000000000_0001011000010011_1001101111010100"; -- 0.08623670502670304
	pesos_i(10927) := b"1111111111111111_1111111111111111_1101101010101011_0111111010001011"; -- -0.14582070446608755
	pesos_i(10928) := b"0000000000000000_0000000000000000_0010000001100010_0000100110010010"; -- 0.12649593172993487
	pesos_i(10929) := b"0000000000000000_0000000000000000_0001111110111100_1010101100011001"; -- 0.12397260059799256
	pesos_i(10930) := b"1111111111111111_1111111111111111_1110000000111011_1111100000100010"; -- -0.12408494162381806
	pesos_i(10931) := b"0000000000000000_0000000000000000_0001000000010111_1000111111101110"; -- 0.06285953102265482
	pesos_i(10932) := b"1111111111111111_1111111111111111_1111010101001100_1101011000010111"; -- -0.04179632134104665
	pesos_i(10933) := b"1111111111111111_1111111111111111_1111101100111001_1010010011000110"; -- -0.018651677816079692
	pesos_i(10934) := b"0000000000000000_0000000000000000_0000001101010100_1001011010111110"; -- 0.013009473317028244
	pesos_i(10935) := b"1111111111111111_1111111111111111_1111011111111100_0011000010110100"; -- -0.031308132258535765
	pesos_i(10936) := b"1111111111111111_1111111111111111_1101111011101000_1000000100101011"; -- -0.12926476200441958
	pesos_i(10937) := b"1111111111111111_1111111111111111_1110011110000011_1110000101010110"; -- -0.09564391752678857
	pesos_i(10938) := b"0000000000000000_0000000000000000_0000010111010110_0011001110111010"; -- 0.022799714074737784
	pesos_i(10939) := b"0000000000000000_0000000000000000_0001011100100100_0000101011101011"; -- 0.09039371714212575
	pesos_i(10940) := b"1111111111111111_1111111111111111_1110010111110110_1011111101110001"; -- -0.10170367714436361
	pesos_i(10941) := b"0000000000000000_0000000000000000_0001010000000000_0100011011000010"; -- 0.07812921751772546
	pesos_i(10942) := b"0000000000000000_0000000000000000_0001001110010000_0001010010011111"; -- 0.07641724462565234
	pesos_i(10943) := b"1111111111111111_1111111111111111_1110111111111100_0000000001000001"; -- -0.0625610200185638
	pesos_i(10944) := b"0000000000000000_0000000000000000_0000010010000100_0010110110111010"; -- 0.017641885715075623
	pesos_i(10945) := b"1111111111111111_1111111111111111_1110001100011010_1100101000100101"; -- -0.11287247264946236
	pesos_i(10946) := b"1111111111111111_1111111111111111_1111011111100101_1101010001000101"; -- -0.031649334976965794
	pesos_i(10947) := b"1111111111111111_1111111111111111_1111001100010111_1000100100101011"; -- -0.05042212200827446
	pesos_i(10948) := b"0000000000000000_0000000000000000_0000001101100100_0001111001110110"; -- 0.013246444580710117
	pesos_i(10949) := b"1111111111111111_1111111111111111_1110001011101010_1010111111011001"; -- -0.1136064619942349
	pesos_i(10950) := b"0000000000000000_0000000000000000_0000001000111000_0000111001001010"; -- 0.008667843949442465
	pesos_i(10951) := b"1111111111111111_1111111111111111_1110001111011011_0010100100001000"; -- -0.10993712952502223
	pesos_i(10952) := b"0000000000000000_0000000000000000_0010000010011110_0111110010100001"; -- 0.12741831714698731
	pesos_i(10953) := b"0000000000000000_0000000000000000_0010011000111011_1000001111001001"; -- 0.14934562350234135
	pesos_i(10954) := b"0000000000000000_0000000000000000_0000101100110010_1001010110110111"; -- 0.043740613038504385
	pesos_i(10955) := b"0000000000000000_0000000000000000_0000010101101100_1100100010010010"; -- 0.021191154135036763
	pesos_i(10956) := b"1111111111111111_1111111111111111_1111101000101001_0011100010010011"; -- -0.022808517673742767
	pesos_i(10957) := b"0000000000000000_0000000000000000_0001100110011010_0101111001101110"; -- 0.1000117319699434
	pesos_i(10958) := b"1111111111111111_1111111111111111_1111111101101000_0010001001111101"; -- -0.002317280174604779
	pesos_i(10959) := b"0000000000000000_0000000000000000_0001100110000010_1111110111111111"; -- 0.09965503203709075
	pesos_i(10960) := b"0000000000000000_0000000000000000_0010011100111110_0001110110101010"; -- 0.1532915630242516
	pesos_i(10961) := b"1111111111111111_1111111111111111_1110011011001010_1010110110111110"; -- -0.09846986877633519
	pesos_i(10962) := b"1111111111111111_1111111111111111_1101100110000111_0111100110100100"; -- -0.15027656312873328
	pesos_i(10963) := b"0000000000000000_0000000000000000_0001110001111110_0001111010011011"; -- 0.11129943171017158
	pesos_i(10964) := b"0000000000000000_0000000000000000_0010011000111010_1110101000100010"; -- 0.149336465065024
	pesos_i(10965) := b"1111111111111111_1111111111111111_1101010111011011_0101100111000110"; -- -0.1646217241779113
	pesos_i(10966) := b"0000000000000000_0000000000000000_0001110011001100_0110101101001011"; -- 0.11249418811283787
	pesos_i(10967) := b"0000000000000000_0000000000000000_0010001110010011_0010101100100100"; -- 0.13896436342729637
	pesos_i(10968) := b"1111111111111111_1111111111111111_1111100010110000_0000100001111010"; -- -0.02856394792594201
	pesos_i(10969) := b"0000000000000000_0000000000000000_0010001100100011_0010101111001010"; -- 0.13725541764471813
	pesos_i(10970) := b"1111111111111111_1111111111111111_1110010001010000_1111000011110000"; -- -0.10813993598024711
	pesos_i(10971) := b"1111111111111111_1111111111111111_1111000111100011_0000110111110000"; -- -0.055129174185209656
	pesos_i(10972) := b"0000000000000000_0000000000000000_0000000010100001_0001100111010111"; -- 0.0024582052140104393
	pesos_i(10973) := b"1111111111111111_1111111111111111_1110100010011110_0010000111111100"; -- -0.09133708573016368
	pesos_i(10974) := b"0000000000000000_0000000000000000_0010010101010101_0101101010010110"; -- 0.14583364650653585
	pesos_i(10975) := b"0000000000000000_0000000000000000_0001110001110000_1100110010001100"; -- 0.11109617627290332
	pesos_i(10976) := b"0000000000000000_0000000000000000_0010000110101000_0001000110110111"; -- 0.13147078248601415
	pesos_i(10977) := b"1111111111111111_1111111111111111_1111110010101111_0100111001101010"; -- -0.012950038061817916
	pesos_i(10978) := b"0000000000000000_0000000000000000_0001110110100000_1001101100000010"; -- 0.11573189552962412
	pesos_i(10979) := b"1111111111111111_1111111111111111_1111110101001110_0011101100000101"; -- -0.010525046709214265
	pesos_i(10980) := b"0000000000000000_0000000000000000_0001101000001000_1011010110111110"; -- 0.10169540299634361
	pesos_i(10981) := b"0000000000000000_0000000000000000_0010100001101011_0011111011110100"; -- 0.1578864428020336
	pesos_i(10982) := b"0000000000000000_0000000000000000_0010001000010011_0001001011101111"; -- 0.13310354550588877
	pesos_i(10983) := b"0000000000000000_0000000000000000_0010010001011110_0110101010010000"; -- 0.14206567776647683
	pesos_i(10984) := b"0000000000000000_0000000000000000_0000011100010010_0010110001010000"; -- 0.02762104932164369
	pesos_i(10985) := b"1111111111111111_1111111111111111_1110001111101100_0011011000001111"; -- -0.10967695357150252
	pesos_i(10986) := b"0000000000000000_0000000000000000_0000000010001001_0101100100110010"; -- 0.002095770533805718
	pesos_i(10987) := b"0000000000000000_0000000000000000_0010000010001111_0111001011110100"; -- 0.12718885847883565
	pesos_i(10988) := b"1111111111111111_1111111111111111_1111111100001011_0000101010011001"; -- -0.0037377716231603766
	pesos_i(10989) := b"1111111111111111_1111111111111111_1110100001001110_1101110010010111"; -- -0.09254666631041517
	pesos_i(10990) := b"1111111111111111_1111111111111111_1111000110000000_0000111111100001"; -- -0.05663967847778009
	pesos_i(10991) := b"1111111111111111_1111111111111111_1111000001111101_0010100011001110"; -- -0.06059021916987924
	pesos_i(10992) := b"0000000000000000_0000000000000000_0000000111100000_0101110010101001"; -- 0.007329741681672517
	pesos_i(10993) := b"1111111111111111_1111111111111111_1101111010010101_0000011110111110"; -- -0.130538479002292
	pesos_i(10994) := b"1111111111111111_1111111111111111_1110101100110010_0111100011011001"; -- -0.08126110756804612
	pesos_i(10995) := b"1111111111111111_1111111111111111_1110001011001110_0100111111100111"; -- -0.11403942696194876
	pesos_i(10996) := b"0000000000000000_0000000000000000_0001111110011111_1001110011111011"; -- 0.1235292541515514
	pesos_i(10997) := b"0000000000000000_0000000000000000_0000101011011001_0000110110000101"; -- 0.042374462964191034
	pesos_i(10998) := b"1111111111111111_1111111111111111_1110111001101100_1010111111001101"; -- -0.06865407229032636
	pesos_i(10999) := b"0000000000000000_0000000000000000_0010000011000100_1101101000001000"; -- 0.12800371834133112
	pesos_i(11000) := b"0000000000000000_0000000000000000_0000000011111101_1111111001100101"; -- 0.003875636738512213
	pesos_i(11001) := b"1111111111111111_1111111111111111_1101101110110101_0011011000011101"; -- -0.14176618375083627
	pesos_i(11002) := b"0000000000000000_0000000000000000_0000101110000011_0100001000010010"; -- 0.04497158952242628
	pesos_i(11003) := b"1111111111111111_1111111111111111_1110011011000000_1111101101000111"; -- -0.09861783515263729
	pesos_i(11004) := b"1111111111111111_1111111111111111_1110111110101110_1110100110000111"; -- -0.06373730135741414
	pesos_i(11005) := b"1111111111111111_1111111111111111_1111010000111101_1001100000100100"; -- -0.04593514548221267
	pesos_i(11006) := b"0000000000000000_0000000000000000_0010001110011101_1110000100101010"; -- 0.13912780075130424
	pesos_i(11007) := b"1111111111111111_1111111111111111_1111111100100110_0110111111001101"; -- -0.0033197521984920687
	pesos_i(11008) := b"1111111111111111_1111111111111111_1111001110010000_0101010111010010"; -- -0.048578869058225914
	pesos_i(11009) := b"1111111111111111_1111111111111111_1111011011101000_0000010011001011"; -- -0.03552217516275517
	pesos_i(11010) := b"0000000000000000_0000000000000000_0001101111100010_1101011010011110"; -- 0.10893002846270741
	pesos_i(11011) := b"0000000000000000_0000000000000000_0000001011110001_1101000011110000"; -- 0.011502321923186388
	pesos_i(11012) := b"1111111111111111_1111111111111111_1110000010011011_1001001101010001"; -- -0.1226261068480205
	pesos_i(11013) := b"1111111111111111_1111111111111111_1111001010110110_0010101100010001"; -- -0.05190783345747136
	pesos_i(11014) := b"1111111111111111_1111111111111111_1111000111111110_1010000011111010"; -- -0.05470842270829803
	pesos_i(11015) := b"1111111111111111_1111111111111111_1111001011000011_0011000101111010"; -- -0.05170908711119871
	pesos_i(11016) := b"0000000000000000_0000000000000000_0001011000000001_0011100111111101"; -- 0.08595621512624191
	pesos_i(11017) := b"1111111111111111_1111111111111111_1110100010011000_1000101001011000"; -- -0.09142241813701633
	pesos_i(11018) := b"0000000000000000_0000000000000000_0001111100110110_1000111011100110"; -- 0.12192624210810199
	pesos_i(11019) := b"0000000000000000_0000000000000000_0000111010111001_0101010011101101"; -- 0.05751543797382335
	pesos_i(11020) := b"1111111111111111_1111111111111111_1101101000000001_1010110010010110"; -- -0.14841195426386705
	pesos_i(11021) := b"1111111111111111_1111111111111111_1101011100011101_1110001000000011"; -- -0.15970027373885864
	pesos_i(11022) := b"1111111111111111_1111111111111111_1111001011101011_0111111000010101"; -- -0.05109416954655684
	pesos_i(11023) := b"1111111111111111_1111111111111111_1111111110101110_0000011010110100"; -- -0.0012508212691806164
	pesos_i(11024) := b"1111111111111111_1111111111111111_1101111010111001_0011101101100110"; -- -0.12998608368574335
	pesos_i(11025) := b"0000000000000000_0000000000000000_0001100110111010_1100101000011010"; -- 0.10050643091110237
	pesos_i(11026) := b"0000000000000000_0000000000000000_0000100011001010_0001001100000110"; -- 0.03433340915958508
	pesos_i(11027) := b"0000000000000000_0000000000000000_0000101010000110_1001000101001010"; -- 0.04111583761790295
	pesos_i(11028) := b"1111111111111111_1111111111111111_1110001010111111_0101010010100001"; -- -0.11426802698958971
	pesos_i(11029) := b"1111111111111111_1111111111111111_1111000101000011_0110010001011101"; -- -0.057565428943637385
	pesos_i(11030) := b"1111111111111111_1111111111111111_1111111100000011_1010101011110110"; -- -0.003850283472817592
	pesos_i(11031) := b"1111111111111111_1111111111111111_1110101000001111_0001100110111000"; -- -0.08570708523374508
	pesos_i(11032) := b"0000000000000000_0000000000000000_0000101111100001_1111001010111001"; -- 0.0464164450506504
	pesos_i(11033) := b"1111111111111111_1111111111111111_1101111111110011_1101010001111000"; -- -0.12518570006230273
	pesos_i(11034) := b"0000000000000000_0000000000000000_0000001111010100_1100110010100111"; -- 0.014965811580958886
	pesos_i(11035) := b"1111111111111111_1111111111111111_1111101111000111_0110001101010000"; -- -0.01648883145689252
	pesos_i(11036) := b"0000000000000000_0000000000000000_0001111100011011_0100001101000011"; -- 0.12150974635309157
	pesos_i(11037) := b"1111111111111111_1111111111111111_1111111101110111_1001010111011100"; -- -0.0020815218994056518
	pesos_i(11038) := b"0000000000000000_0000000000000000_0010001001011010_1111001000100010"; -- 0.1342002231757348
	pesos_i(11039) := b"1111111111111111_1111111111111111_1101011100011001_0001110110011001"; -- -0.1597730161797126
	pesos_i(11040) := b"1111111111111111_1111111111111111_1111000110000100_1111111011001110"; -- -0.056564402306161055
	pesos_i(11041) := b"1111111111111111_1111111111111111_1110111000000111_1100110000101111"; -- -0.07019351814747743
	pesos_i(11042) := b"0000000000000000_0000000000000000_0001001010110101_1101011011010001"; -- 0.07308714492739783
	pesos_i(11043) := b"0000000000000000_0000000000000000_0010100111111010_0101010010011100"; -- 0.16397599028897827
	pesos_i(11044) := b"0000000000000000_0000000000000000_0000101110011110_0010000000001011"; -- 0.04538154865301415
	pesos_i(11045) := b"1111111111111111_1111111111111111_1110111110100100_1111111111110110"; -- -0.06388855223170453
	pesos_i(11046) := b"0000000000000000_0000000000000000_0001001000011101_0111111111100110"; -- 0.0707626283004542
	pesos_i(11047) := b"0000000000000000_0000000000000000_0010010110000011_1011011011001000"; -- 0.14654104586769467
	pesos_i(11048) := b"0000000000000000_0000000000000000_0000000111011011_1011111000100001"; -- 0.00725925737671214
	pesos_i(11049) := b"1111111111111111_1111111111111111_1111011001101111_1011100111011010"; -- -0.037357696868694765
	pesos_i(11050) := b"0000000000000000_0000000000000000_0000101011001011_0101001011001001"; -- 0.04216496858725741
	pesos_i(11051) := b"0000000000000000_0000000000000000_0001011111011101_0000101010001111"; -- 0.0932165718016552
	pesos_i(11052) := b"0000000000000000_0000000000000000_0000110010000001_0010101100011001"; -- 0.0488459526653524
	pesos_i(11053) := b"1111111111111111_1111111111111111_1111011001100100_0110111000100111"; -- -0.03753005554507759
	pesos_i(11054) := b"0000000000000000_0000000000000000_0001010111011101_0100100111000110"; -- 0.08540783955612768
	pesos_i(11055) := b"0000000000000000_0000000000000000_0000110111000111_0000000110000010"; -- 0.053817838993860376
	pesos_i(11056) := b"1111111111111111_1111111111111111_1111010101100011_1111001011111111"; -- -0.0414436461498179
	pesos_i(11057) := b"1111111111111111_1111111111111111_1111010000100000_0111010111011010"; -- -0.046379694178851176
	pesos_i(11058) := b"0000000000000000_0000000000000000_0010001101011010_1010110000001001"; -- 0.1381022950477943
	pesos_i(11059) := b"0000000000000000_0000000000000000_0010001011100000_0011000101110101"; -- 0.13623341662333868
	pesos_i(11060) := b"1111111111111111_1111111111111111_1111010011101100_1100100111011111"; -- -0.043261893410246575
	pesos_i(11061) := b"1111111111111111_1111111111111111_1111000111110101_0011010000100010"; -- -0.05485223940986409
	pesos_i(11062) := b"0000000000000000_0000000000000000_0001100010101110_0100000101111001"; -- 0.0964089317659202
	pesos_i(11063) := b"1111111111111111_1111111111111111_1110000010111011_0011000101010101"; -- -0.12214366597832833
	pesos_i(11064) := b"1111111111111111_1111111111111111_1110110011110000_0111100110110000"; -- -0.07445563739741988
	pesos_i(11065) := b"0000000000000000_0000000000000000_0000010011001110_0110001100110000"; -- 0.018774222690030703
	pesos_i(11066) := b"0000000000000000_0000000000000000_0001101011010101_1110000010001100"; -- 0.10482600617655932
	pesos_i(11067) := b"1111111111111111_1111111111111111_1111011010010111_0011010001001001"; -- -0.03675530647949595
	pesos_i(11068) := b"0000000000000000_0000000000000000_0001001100111011_0000110110010110"; -- 0.07511982824868012
	pesos_i(11069) := b"0000000000000000_0000000000000000_0000110110101110_1101101101101100"; -- 0.05344935797144877
	pesos_i(11070) := b"0000000000000000_0000000000000000_0000000101101010_1101100101101110"; -- 0.005536641518596765
	pesos_i(11071) := b"1111111111111111_1111111111111111_1111111100010001_0101000011011011"; -- -0.003642031236667223
	pesos_i(11072) := b"1111111111111111_1111111111111111_1101100111011001_1111100011011010"; -- -0.14901776018005608
	pesos_i(11073) := b"0000000000000000_0000000000000000_0000000111000101_1111011000100101"; -- 0.006926902846738591
	pesos_i(11074) := b"0000000000000000_0000000000000000_0000100111111101_1011001111101110"; -- 0.039027448277604196
	pesos_i(11075) := b"1111111111111111_1111111111111111_1110101000100101_0001001001101011"; -- -0.08537182694369513
	pesos_i(11076) := b"1111111111111111_1111111111111111_1110001100001001_1010100110011111"; -- -0.11313381080514306
	pesos_i(11077) := b"1111111111111111_1111111111111111_1110111111010110_1101110011110101"; -- -0.06312769896510548
	pesos_i(11078) := b"0000000000000000_0000000000000000_0001001000010010_1110011011101100"; -- 0.07060092227085715
	pesos_i(11079) := b"1111111111111111_1111111111111111_1111001100101010_1000001010000101"; -- -0.05013260122004566
	pesos_i(11080) := b"0000000000000000_0000000000000000_0001100110010011_0100000111100010"; -- 0.09990321885005207
	pesos_i(11081) := b"1111111111111111_1111111111111111_1111010101101010_1101110000100110"; -- -0.04133819651952122
	pesos_i(11082) := b"1111111111111111_1111111111111111_1111111110110111_0001001101111011"; -- -0.0011127304964559503
	pesos_i(11083) := b"1111111111111111_1111111111111111_1111101000011100_1000110110111010"; -- -0.023001806287955052
	pesos_i(11084) := b"1111111111111111_1111111111111111_1111111101101100_1010110001011010"; -- -0.0022480278419423293
	pesos_i(11085) := b"0000000000000000_0000000000000000_0001111011111111_0111101011100000"; -- 0.12108581522011388
	pesos_i(11086) := b"0000000000000000_0000000000000000_0001101100110101_1000101000001110"; -- 0.10628569452040558
	pesos_i(11087) := b"0000000000000000_0000000000000000_0001101111011111_1101101101010011"; -- 0.10888453271543186
	pesos_i(11088) := b"0000000000000000_0000000000000000_0001010001001100_0011101110100110"; -- 0.07928822331321077
	pesos_i(11089) := b"1111111111111111_1111111111111111_1111101000100100_1010011111111110"; -- -0.022878170504729494
	pesos_i(11090) := b"0000000000000000_0000000000000000_0000001010000000_0101100101010101"; -- 0.009770949592821264
	pesos_i(11091) := b"1111111111111111_1111111111111111_1111010100001001_0100010111000101"; -- -0.04282726231710697
	pesos_i(11092) := b"1111111111111111_1111111111111111_1110011000010111_0100001101001011"; -- -0.1012075368660336
	pesos_i(11093) := b"0000000000000000_0000000000000000_0001110111010100_1101001111010001"; -- 0.11652873854183197
	pesos_i(11094) := b"0000000000000000_0000000000000000_0000100101011001_1010100111001000"; -- 0.036524401901649434
	pesos_i(11095) := b"0000000000000000_0000000000000000_0000110111001011_0000101110001010"; -- 0.05387947194952961
	pesos_i(11096) := b"1111111111111111_1111111111111111_1111111110011111_1110101010111001"; -- -0.0014661120234185033
	pesos_i(11097) := b"1111111111111111_1111111111111111_1111111011011110_0000100011111010"; -- -0.004424513674588798
	pesos_i(11098) := b"0000000000000000_0000000000000000_0001100111100010_0101111000000010"; -- 0.10111033958975886
	pesos_i(11099) := b"1111111111111111_1111111111111111_1110001110011110_1010101110100001"; -- -0.1108601315496149
	pesos_i(11100) := b"1111111111111111_1111111111111111_1110001010110100_0000010101111110"; -- -0.11444059069392053
	pesos_i(11101) := b"1111111111111111_1111111111111111_1111011000110001_0010110110100000"; -- -0.03831209989463959
	pesos_i(11102) := b"1111111111111111_1111111111111111_1111110110010000_1110001101000111"; -- -0.009507937671671095
	pesos_i(11103) := b"0000000000000000_0000000000000000_0001010101011101_1110000110100101"; -- 0.0834637669591704
	pesos_i(11104) := b"0000000000000000_0000000000000000_0001100001011110_0111011111100010"; -- 0.09519147174721786
	pesos_i(11105) := b"0000000000000000_0000000000000000_0001110011000000_1111110010011101"; -- 0.11231974452192148
	pesos_i(11106) := b"0000000000000000_0000000000000000_0010010010011101_0001111010100001"; -- 0.14302245545786318
	pesos_i(11107) := b"1111111111111111_1111111111111111_1101110011101011_0000010101101110"; -- -0.13703886097123158
	pesos_i(11108) := b"1111111111111111_1111111111111111_1110100101011001_0111011100101000"; -- -0.08847861550078978
	pesos_i(11109) := b"1111111111111111_1111111111111111_1101100110100011_0110111100101100"; -- -0.1498499409752928
	pesos_i(11110) := b"1111111111111111_1111111111111111_1101111001001001_0111111100001101"; -- -0.13169103558660844
	pesos_i(11111) := b"1111111111111111_1111111111111111_1110010101110101_1101110010010101"; -- -0.10367032396827063
	pesos_i(11112) := b"1111111111111111_1111111111111111_1110111011011000_1100000110111000"; -- -0.06700505502410889
	pesos_i(11113) := b"0000000000000000_0000000000000000_0000100111101000_1111101110001110"; -- 0.03871128298397454
	pesos_i(11114) := b"1111111111111111_1111111111111111_1111111101010101_1100011010111001"; -- -0.0025974081574195464
	pesos_i(11115) := b"1111111111111111_1111111111111111_1111111010011100_0001010101011111"; -- -0.005430855092682925
	pesos_i(11116) := b"1111111111111111_1111111111111111_1111101000010110_1110010010111111"; -- -0.023088172382889655
	pesos_i(11117) := b"1111111111111111_1111111111111111_1110000000100000_1000111011100100"; -- -0.1245032017326938
	pesos_i(11118) := b"1111111111111111_1111111111111111_1111001000010001_0011010110100010"; -- -0.05442490384370061
	pesos_i(11119) := b"1111111111111111_1111111111111111_1110100110011100_0100110011010001"; -- -0.0874588002527011
	pesos_i(11120) := b"1111111111111111_1111111111111111_1111011001110010_0000011010111001"; -- -0.03732259738522958
	pesos_i(11121) := b"1111111111111111_1111111111111111_1111010110111010_0100000100000011"; -- -0.04012674027212551
	pesos_i(11122) := b"1111111111111111_1111111111111111_1101100111001001_1001110110001010"; -- -0.14926734333904965
	pesos_i(11123) := b"0000000000000000_0000000000000000_0001011110000000_1011010101101101"; -- 0.09180768889261581
	pesos_i(11124) := b"0000000000000000_0000000000000000_0001010110010101_0011100110001110"; -- 0.08430824013790746
	pesos_i(11125) := b"1111111111111111_1111111111111111_1111111101011011_0010010110111101"; -- -0.0025154509237107115
	pesos_i(11126) := b"0000000000000000_0000000000000000_0001101000111110_0000100110000010"; -- 0.10250911167277905
	pesos_i(11127) := b"0000000000000000_0000000000000000_0001000000111110_1111100000010101"; -- 0.06346083186039937
	pesos_i(11128) := b"1111111111111111_1111111111111111_1110010010000000_1101110101111010"; -- -0.10740867388701188
	pesos_i(11129) := b"0000000000000000_0000000000000000_0000011111000101_0001000001110111"; -- 0.03035071283713986
	pesos_i(11130) := b"1111111111111111_1111111111111111_1111110000101000_1101000011100100"; -- -0.01500219767232268
	pesos_i(11131) := b"0000000000000000_0000000000000000_0000010001011010_1101100011010110"; -- 0.017011215418374408
	pesos_i(11132) := b"1111111111111111_1111111111111111_1110110100011101_1010001001000000"; -- -0.073766574288635
	pesos_i(11133) := b"0000000000000000_0000000000000000_0000010110010010_1001000011100110"; -- 0.02176766988650855
	pesos_i(11134) := b"1111111111111111_1111111111111111_1111100100011011_1111111011110011"; -- -0.026916566499588943
	pesos_i(11135) := b"1111111111111111_1111111111111111_1110100010100101_0000010001101100"; -- -0.09123203617497065
	pesos_i(11136) := b"1111111111111111_1111111111111111_1111000010110111_0001110000011111"; -- -0.059705965364888015
	pesos_i(11137) := b"1111111111111111_1111111111111111_1111001000011100_1010011001110001"; -- -0.05425033320506814
	pesos_i(11138) := b"0000000000000000_0000000000000000_0000011000110101_0101101001110100"; -- 0.02425160730262725
	pesos_i(11139) := b"1111111111111111_1111111111111111_1101110111011100_1100111111100011"; -- -0.13334942544509518
	pesos_i(11140) := b"0000000000000000_0000000000000000_0000111001011011_1100001101000111"; -- 0.05608768917324907
	pesos_i(11141) := b"0000000000000000_0000000000000000_0001110000010000_1011111011100010"; -- 0.10963051814439066
	pesos_i(11142) := b"1111111111111111_1111111111111111_1111000001101101_0001100011000011"; -- -0.06083531612204834
	pesos_i(11143) := b"1111111111111111_1111111111111111_1110110110011110_1011100011110101"; -- -0.07179683695880636
	pesos_i(11144) := b"1111111111111111_1111111111111111_1101110011101111_0010110111111101"; -- -0.1369754084052903
	pesos_i(11145) := b"1111111111111111_1111111111111111_1111110101001111_0001110011010001"; -- -0.010511588107998071
	pesos_i(11146) := b"1111111111111111_1111111111111111_1111000110110111_0111011010101010"; -- -0.055794318686390156
	pesos_i(11147) := b"0000000000000000_0000000000000000_0000000000101010_0000111110110010"; -- 0.0006418045877343484
	pesos_i(11148) := b"0000000000000000_0000000000000000_0010000011100111_0010011000100101"; -- 0.12852705387061192
	pesos_i(11149) := b"0000000000000000_0000000000000000_0001111001110100_0111010000101100"; -- 0.11896444380565785
	pesos_i(11150) := b"0000000000000000_0000000000000000_0001000101000111_0111010001000010"; -- 0.0674965534712548
	pesos_i(11151) := b"0000000000000000_0000000000000000_0000001100011101_1110101001011110"; -- 0.012175224285588232
	pesos_i(11152) := b"0000000000000000_0000000000000000_0010000000101010_1010000101011001"; -- 0.12565048626838232
	pesos_i(11153) := b"1111111111111111_1111111111111111_1111000111001101_0101010011010011"; -- -0.055460642396156584
	pesos_i(11154) := b"1111111111111111_1111111111111111_1111111000011000_1000000011000100"; -- -0.007438614040045841
	pesos_i(11155) := b"0000000000000000_0000000000000000_0001001101111111_0110000100101010"; -- 0.07616240772755707
	pesos_i(11156) := b"0000000000000000_0000000000000000_0001111011110110_1110011101110101"; -- 0.12095495802672514
	pesos_i(11157) := b"1111111111111111_1111111111111111_1110111010100110_1100100101100011"; -- -0.06776753745874992
	pesos_i(11158) := b"1111111111111111_1111111111111111_1110100000101100_1011110101111010"; -- -0.09306731971389097
	pesos_i(11159) := b"1111111111111111_1111111111111111_1111101100101111_1010000100001110"; -- -0.01880448736481529
	pesos_i(11160) := b"0000000000000000_0000000000000000_0010000011001111_1001100101111010"; -- 0.12816771727251114
	pesos_i(11161) := b"1111111111111111_1111111111111111_1111001100111111_1010110110110011"; -- -0.049809593006554444
	pesos_i(11162) := b"1111111111111111_1111111111111111_1110010001111000_1101101111011001"; -- -0.10753084140774301
	pesos_i(11163) := b"0000000000000000_0000000000000000_0001010110101001_0111101010100001"; -- 0.08461729462963861
	pesos_i(11164) := b"1111111111111111_1111111111111111_1111011000101100_0101001101010010"; -- -0.03838614697045492
	pesos_i(11165) := b"0000000000000000_0000000000000000_0000100011110100_1001000101111010"; -- 0.03498181551910495
	pesos_i(11166) := b"1111111111111111_1111111111111111_1111011101011101_0110001101001111"; -- -0.03373126338552771
	pesos_i(11167) := b"0000000000000000_0000000000000000_0000011100110001_1001010101111111"; -- 0.028100341342771652
	pesos_i(11168) := b"0000000000000000_0000000000000000_0001111010010100_1001011101000011"; -- 0.11945481677518625
	pesos_i(11169) := b"0000000000000000_0000000000000000_0001111110101100_1101010011100011"; -- 0.12373095074339638
	pesos_i(11170) := b"0000000000000000_0000000000000000_0001010010111100_1010111101010010"; -- 0.08100410221588732
	pesos_i(11171) := b"1111111111111111_1111111111111111_1110010010101111_1010011101001110"; -- -0.10669473967884062
	pesos_i(11172) := b"1111111111111111_1111111111111111_1110100110100011_0101111111001110"; -- -0.08735085707369991
	pesos_i(11173) := b"0000000000000000_0000000000000000_0000110101111010_0111100111011100"; -- 0.05265008567601061
	pesos_i(11174) := b"1111111111111111_1111111111111111_1111001101111001_0011001110101001"; -- -0.048931857336493016
	pesos_i(11175) := b"1111111111111111_1111111111111111_1110100100100010_1101011010001010"; -- -0.089312163534888
	pesos_i(11176) := b"0000000000000000_0000000000000000_0000010101111001_0110100011011010"; -- 0.021383813212606528
	pesos_i(11177) := b"0000000000000000_0000000000000000_0001000011010111_1000001001010100"; -- 0.06578840776835194
	pesos_i(11178) := b"0000000000000000_0000000000000000_0010000100011101_1110010000010111"; -- 0.12936235008362493
	pesos_i(11179) := b"0000000000000000_0000000000000000_0010001000110001_0110011011000100"; -- 0.13356630600923453
	pesos_i(11180) := b"0000000000000000_0000000000000000_0010000110111101_0111001100100000"; -- 0.1317970232168627
	pesos_i(11181) := b"0000000000000000_0000000000000000_0010000011100101_1111001000011001"; -- 0.12850869275721136
	pesos_i(11182) := b"1111111111111111_1111111111111111_1110001001010101_1101100111110001"; -- -0.11587751272081011
	pesos_i(11183) := b"0000000000000000_0000000000000000_0001011010100100_1010101001011101"; -- 0.08845009573629885
	pesos_i(11184) := b"1111111111111111_1111111111111111_1110110000101101_1101100010100000"; -- -0.07742544257891565
	pesos_i(11185) := b"1111111111111111_1111111111111111_1110110100111011_1000110100001101"; -- -0.07331007427221893
	pesos_i(11186) := b"1111111111111111_1111111111111111_1111010100001010_1110000001001000"; -- -0.04280279385082334
	pesos_i(11187) := b"0000000000000000_0000000000000000_0001111010000011_1100110100000100"; -- 0.11919862115655948
	pesos_i(11188) := b"1111111111111111_1111111111111111_1110011111111011_0011011000000110"; -- -0.09382307388533478
	pesos_i(11189) := b"1111111111111111_1111111111111111_1111011101111111_1011101100011011"; -- -0.03320723139364865
	pesos_i(11190) := b"0000000000000000_0000000000000000_0000000010100101_1011111000010001"; -- 0.0025290289746120855
	pesos_i(11191) := b"0000000000000000_0000000000000000_0001100101001100_0100011110101011"; -- 0.09882018964708848
	pesos_i(11192) := b"1111111111111111_1111111111111111_1110011001010001_1100000010000001"; -- -0.10031506394777978
	pesos_i(11193) := b"1111111111111111_1111111111111111_1111110101001000_1110000111001000"; -- -0.010606659626467379
	pesos_i(11194) := b"1111111111111111_1111111111111111_1111101110001101_0011101110100000"; -- -0.017376206929291146
	pesos_i(11195) := b"1111111111111111_1111111111111111_1110110010011001_0000101000011101"; -- -0.07578980238293713
	pesos_i(11196) := b"1111111111111111_1111111111111111_1110100001000101_1010110001101001"; -- -0.09268686700038077
	pesos_i(11197) := b"0000000000000000_0000000000000000_0001101101110010_1101100001010011"; -- 0.10722114578377363
	pesos_i(11198) := b"1111111111111111_1111111111111111_1110101100000110_1001101100001100"; -- -0.08193045573039731
	pesos_i(11199) := b"1111111111111111_1111111111111111_1110101110111100_0000000111011001"; -- -0.0791624874961602
	pesos_i(11200) := b"0000000000000000_0000000000000000_0000011001111010_0111011101001100"; -- 0.02530618287926157
	pesos_i(11201) := b"0000000000000000_0000000000000000_0001001001111000_0110001111000111"; -- 0.07214950192128196
	pesos_i(11202) := b"0000000000000000_0000000000000000_0000010001100001_0101011010001001"; -- 0.01711026053866747
	pesos_i(11203) := b"1111111111111111_1111111111111111_1110001001101100_0111100000101100"; -- -0.11553238790091584
	pesos_i(11204) := b"0000000000000000_0000000000000000_0000011110101001_0000010100011101"; -- 0.029922790084088782
	pesos_i(11205) := b"1111111111111111_1111111111111111_1110100001100010_1100101100100100"; -- -0.09224253055673082
	pesos_i(11206) := b"1111111111111111_1111111111111111_1101100110010010_1111011101110101"; -- -0.15010121719853745
	pesos_i(11207) := b"1111111111111111_1111111111111111_1111101011111111_1001001011010001"; -- -0.01953775780303556
	pesos_i(11208) := b"1111111111111111_1111111111111111_1110001110101110_1101110001100111"; -- -0.11061308373606533
	pesos_i(11209) := b"1111111111111111_1111111111111111_1110101100110100_1001000001101101"; -- -0.0812291845726571
	pesos_i(11210) := b"1111111111111111_1111111111111111_1101110111001010_0011011011101101"; -- -0.13363320072031534
	pesos_i(11211) := b"0000000000000000_0000000000000000_0000100000011110_0100100010111011"; -- 0.0317120986636623
	pesos_i(11212) := b"0000000000000000_0000000000000000_0010000010110010_0101110100101011"; -- 0.12772161758823683
	pesos_i(11213) := b"0000000000000000_0000000000000000_0001011010110000_0110011011010101"; -- 0.08862917610082618
	pesos_i(11214) := b"1111111111111111_1111111111111111_1110011011101010_1011100111111001"; -- -0.09798085857176694
	pesos_i(11215) := b"1111111111111111_1111111111111111_1111110101111100_0001101101010011"; -- -0.009825031411294203
	pesos_i(11216) := b"1111111111111111_1111111111111111_1110011001011010_1010011001111001"; -- -0.10017928644708983
	pesos_i(11217) := b"1111111111111111_1111111111111111_1111111110100001_0110101110001100"; -- -0.0014431746323975124
	pesos_i(11218) := b"1111111111111111_1111111111111111_1111001010110100_1110101010100110"; -- -0.05192693186354797
	pesos_i(11219) := b"0000000000000000_0000000000000000_0001110111001101_1110010000001010"; -- 0.11642289389363591
	pesos_i(11220) := b"0000000000000000_0000000000000000_0010010111010010_1110000010101101"; -- 0.14774898738897355
	pesos_i(11221) := b"0000000000000000_0000000000000000_0000000101100110_1000101011110110"; -- 0.005470929311326968
	pesos_i(11222) := b"1111111111111111_1111111111111111_1110011000011010_1000110011000101"; -- -0.10115738097285695
	pesos_i(11223) := b"0000000000000000_0000000000000000_0001000100010001_1011010111000001"; -- 0.06667648275033058
	pesos_i(11224) := b"1111111111111111_1111111111111111_1110111100001011_0010101111000000"; -- -0.06623579561874934
	pesos_i(11225) := b"1111111111111111_1111111111111111_1110000010100010_0110001101100010"; -- -0.12252215239854992
	pesos_i(11226) := b"1111111111111111_1111111111111111_1110100100100011_0110101011101001"; -- -0.08930332002637474
	pesos_i(11227) := b"0000000000000000_0000000000000000_0001101101010110_0011101110001101"; -- 0.10678455528317309
	pesos_i(11228) := b"1111111111111111_1111111111111111_1110000010000011_1010111101111101"; -- -0.12299063870140203
	pesos_i(11229) := b"0000000000000000_0000000000000000_0010000000100010_1111101110010010"; -- 0.12553379360698932
	pesos_i(11230) := b"1111111111111111_1111111111111111_1111101111101010_1111100110111001"; -- -0.015945808822945787
	pesos_i(11231) := b"0000000000000000_0000000000000000_0000110000101101_1010010010110101"; -- 0.047571462696146025
	pesos_i(11232) := b"0000000000000000_0000000000000000_0001101001010001_0110000011001100"; -- 0.10280423153511192
	pesos_i(11233) := b"1111111111111111_1111111111111111_1101110101000111_1101111010100011"; -- -0.13562210572691416
	pesos_i(11234) := b"0000000000000000_0000000000000000_0010010110011001_1100100101000011"; -- 0.1468778409430883
	pesos_i(11235) := b"1111111111111111_1111111111111111_1110101000011010_0000011110010101"; -- -0.08554031944542409
	pesos_i(11236) := b"0000000000000000_0000000000000000_0000010110010100_0000100011011110"; -- 0.02179007939125773
	pesos_i(11237) := b"0000000000000000_0000000000000000_0000001111111101_0010110011110101"; -- 0.015581903294448913
	pesos_i(11238) := b"1111111111111111_1111111111111111_1111001010110111_1100100110110101"; -- -0.051883118926741745
	pesos_i(11239) := b"0000000000000000_0000000000000000_0000110000010011_0000100101001100"; -- 0.04716547110306913
	pesos_i(11240) := b"1111111111111111_1111111111111111_1110111001111011_0000000011101110"; -- -0.06843561358264265
	pesos_i(11241) := b"1111111111111111_1111111111111111_1111111110001011_1001100001101111"; -- -0.001776192514333144
	pesos_i(11242) := b"0000000000000000_0000000000000000_0000110011001100_0111001101111000"; -- 0.049994675538491955
	pesos_i(11243) := b"0000000000000000_0000000000000000_0000111001100110_1001110101000001"; -- 0.05625326966298522
	pesos_i(11244) := b"0000000000000000_0000000000000000_0001000011011100_1100101101000100"; -- 0.06586904925497455
	pesos_i(11245) := b"1111111111111111_1111111111111111_1101101010000110_0101111001110110"; -- -0.1463871919924498
	pesos_i(11246) := b"0000000000000000_0000000000000000_0000100011110100_0110111010001101"; -- 0.03497973383416015
	pesos_i(11247) := b"0000000000000000_0000000000000000_0001010101110101_0111110010101111"; -- 0.08382395998932107
	pesos_i(11248) := b"1111111111111111_1111111111111111_1111100011011011_1110110101011110"; -- -0.02789417693963268
	pesos_i(11249) := b"1111111111111111_1111111111111111_1101110010011101_1001000100011001"; -- -0.1382207217224942
	pesos_i(11250) := b"1111111111111111_1111111111111111_1111110101000110_1101101111001100"; -- -0.010637533836220176
	pesos_i(11251) := b"1111111111111111_1111111111111111_1110000101101000_0010110110011110"; -- -0.11950411687901295
	pesos_i(11252) := b"1111111111111111_1111111111111111_1110010011110100_0110011010110010"; -- -0.10564573434610129
	pesos_i(11253) := b"0000000000000000_0000000000000000_0010010011000111_1110010101001101"; -- 0.14367516643135528
	pesos_i(11254) := b"1111111111111111_1111111111111111_1101100110001010_1110110000100010"; -- -0.15022396255439907
	pesos_i(11255) := b"0000000000000000_0000000000000000_0000000011000011_0100101110000100"; -- 0.0029799649400201254
	pesos_i(11256) := b"1111111111111111_1111111111111111_1110011010101010_1000110010001110"; -- -0.0989601280536735
	pesos_i(11257) := b"0000000000000000_0000000000000000_0010001101101100_0011111101001110"; -- 0.13837047254250537
	pesos_i(11258) := b"0000000000000000_0000000000000000_0000100011101000_1101010101001110"; -- 0.03480275304944734
	pesos_i(11259) := b"1111111111111111_1111111111111111_1110100101111100_1110001100010001"; -- -0.08793812592473796
	pesos_i(11260) := b"0000000000000000_0000000000000000_0001101111101001_1100110110110000"; -- 0.10903630771656994
	pesos_i(11261) := b"1111111111111111_1111111111111111_1110101101010100_0010110100011111"; -- -0.08074682225733182
	pesos_i(11262) := b"1111111111111111_1111111111111111_1111000101110100_1111011101110111"; -- -0.05680898051698728
	pesos_i(11263) := b"0000000000000000_0000000000000000_0000000101100000_0100001000010100"; -- 0.005375032408671707
	pesos_i(11264) := b"0000000000000000_0000000000000000_0000101010011100_1010001110110100"; -- 0.04145262860229979
	pesos_i(11265) := b"0000000000000000_0000000000000000_0001001011001000_1001000001100101"; -- 0.07337286429649813
	pesos_i(11266) := b"0000000000000000_0000000000000000_0000111011001000_1011111000000001"; -- 0.057750582826524545
	pesos_i(11267) := b"1111111111111111_1111111111111111_1111101111101101_1001101101011001"; -- -0.015905657570499655
	pesos_i(11268) := b"1111111111111111_1111111111111111_1110011010011101_0011111110111010"; -- -0.09916307168322774
	pesos_i(11269) := b"1111111111111111_1111111111111111_1110110111101010_1011101111111110"; -- -0.07063698810033313
	pesos_i(11270) := b"0000000000000000_0000000000000000_0010010100100000_1100111101110000"; -- 0.1450318954023304
	pesos_i(11271) := b"1111111111111111_1111111111111111_1111010101001111_1010001000101001"; -- -0.041753640194871655
	pesos_i(11272) := b"0000000000000000_0000000000000000_0000100001101010_1001001011100000"; -- 0.03287618616413344
	pesos_i(11273) := b"0000000000000000_0000000000000000_0001111111000001_1101100101101100"; -- 0.12405165569219356
	pesos_i(11274) := b"1111111111111111_1111111111111111_1110001011101011_0000111001010100"; -- -0.1136008305746661
	pesos_i(11275) := b"0000000000000000_0000000000000000_0000100110010111_1110100111001011"; -- 0.037474262330120134
	pesos_i(11276) := b"1111111111111111_1111111111111111_1110100110010010_0000001010001010"; -- -0.0876158154291193
	pesos_i(11277) := b"1111111111111111_1111111111111111_1111011100010100_1011000100110001"; -- -0.034840512858840815
	pesos_i(11278) := b"0000000000000000_0000000000000000_0001101110000111_0010001011100001"; -- 0.10753076543477504
	pesos_i(11279) := b"1111111111111111_1111111111111111_1101111001101010_0010100101001010"; -- -0.1311926074116067
	pesos_i(11280) := b"1111111111111111_1111111111111111_1110110111011100_1111110101010110"; -- -0.07084671641407703
	pesos_i(11281) := b"0000000000000000_0000000000000000_0001101100010101_0000110011011100"; -- 0.10578995095864636
	pesos_i(11282) := b"1111111111111111_1111111111111111_1101101101010100_0000101001011101"; -- -0.1432488941132658
	pesos_i(11283) := b"0000000000000000_0000000000000000_0000000110011100_1110110000110111"; -- 0.006300700497855059
	pesos_i(11284) := b"1111111111111111_1111111111111111_1111001111000000_0110010011110010"; -- -0.04784554563647424
	pesos_i(11285) := b"1111111111111111_1111111111111111_1101111010011111_1111010000110011"; -- -0.13037179712524521
	pesos_i(11286) := b"1111111111111111_1111111111111111_1110100110001000_0010000010111000"; -- -0.0877666045876589
	pesos_i(11287) := b"1111111111111111_1111111111111111_1111010001001111_0011110001111001"; -- -0.04566595130169952
	pesos_i(11288) := b"1111111111111111_1111111111111111_1110000000101010_0011100111101000"; -- -0.12435567935677964
	pesos_i(11289) := b"0000000000000000_0000000000000000_0010001010110010_0010111000010101"; -- 0.1355313111637311
	pesos_i(11290) := b"0000000000000000_0000000000000000_0001110000110010_0100100000100110"; -- 0.1101422397324461
	pesos_i(11291) := b"1111111111111111_1111111111111111_1110010010111010_0110101010001011"; -- -0.10653051487456808
	pesos_i(11292) := b"1111111111111111_1111111111111111_1111110110100101_1000100011000100"; -- -0.00919289790557389
	pesos_i(11293) := b"0000000000000000_0000000000000000_0000100111100111_0110000101111100"; -- 0.03868684071056225
	pesos_i(11294) := b"0000000000000000_0000000000000000_0010001100001000_1010001100001111"; -- 0.1368505392843833
	pesos_i(11295) := b"1111111111111111_1111111111111111_1110000111001111_0101101011101101"; -- -0.11792976103370077
	pesos_i(11296) := b"0000000000000000_0000000000000000_0010010111001010_0011111110111111"; -- 0.14761732487236284
	pesos_i(11297) := b"1111111111111111_1111111111111111_1101101100010100_0011010010110110"; -- -0.14422293247614104
	pesos_i(11298) := b"1111111111111111_1111111111111111_1110000010010000_1100000100100111"; -- -0.12279122162458202
	pesos_i(11299) := b"1111111111111111_1111111111111111_1101111101100100_1111001101010011"; -- -0.1273658679026926
	pesos_i(11300) := b"0000000000000000_0000000000000000_0010001011000011_0101101000000111"; -- 0.13579332985716566
	pesos_i(11301) := b"0000000000000000_0000000000000000_0001010011000100_0111110011010011"; -- 0.0811231626475759
	pesos_i(11302) := b"0000000000000000_0000000000000000_0010001100111011_1100000100101000"; -- 0.1376305315098774
	pesos_i(11303) := b"1111111111111111_1111111111111111_1110111001000010_1110000001100101"; -- -0.0692920449852018
	pesos_i(11304) := b"0000000000000000_0000000000000000_0001101111011111_1000111010101111"; -- 0.10887996462894227
	pesos_i(11305) := b"1111111111111111_1111111111111111_1111010111101101_0101101001011000"; -- -0.03934703212441146
	pesos_i(11306) := b"1111111111111111_1111111111111111_1111000000010110_1110010010100000"; -- -0.06215067952275029
	pesos_i(11307) := b"1111111111111111_1111111111111111_1110100100111001_1011111111010110"; -- -0.08896256471543643
	pesos_i(11308) := b"1111111111111111_1111111111111111_1110101111110111_0001110001001001"; -- -0.07826064314940569
	pesos_i(11309) := b"1111111111111111_1111111111111111_1110010010110010_0011000111001110"; -- -0.10665596700368568
	pesos_i(11310) := b"0000000000000000_0000000000000000_0001000000111111_0101111000010100"; -- 0.06346691109522759
	pesos_i(11311) := b"0000000000000000_0000000000000000_0000110111001100_1101101111111011"; -- 0.05390715492147877
	pesos_i(11312) := b"1111111111111111_1111111111111111_1110110001101000_1110101001100001"; -- -0.07652411588385048
	pesos_i(11313) := b"1111111111111111_1111111111111111_1101100000100110_0111001010100110"; -- -0.15566333238645344
	pesos_i(11314) := b"1111111111111111_1111111111111111_1110011101001110_0000010100111000"; -- -0.09646575330112156
	pesos_i(11315) := b"1111111111111111_1111111111111111_1101110001101111_1010100001010011"; -- -0.13892124161565272
	pesos_i(11316) := b"1111111111111111_1111111111111111_1111100010010110_1100010010110000"; -- -0.02894945809095646
	pesos_i(11317) := b"0000000000000000_0000000000000000_0000011110011010_0001000000111110"; -- 0.029694571527904497
	pesos_i(11318) := b"1111111111111111_1111111111111111_1101111010001001_1010010010100100"; -- -0.13071223261850293
	pesos_i(11319) := b"1111111111111111_1111111111111111_1110000100100000_0110010101001111"; -- -0.12059943023775513
	pesos_i(11320) := b"1111111111111111_1111111111111111_1110011110101111_1000001001010010"; -- -0.09497819427439122
	pesos_i(11321) := b"0000000000000000_0000000000000000_0010001110000111_1101101010000110"; -- 0.13879171142185745
	pesos_i(11322) := b"0000000000000000_0000000000000000_0001100101100000_0111001010100101"; -- 0.09912792708394355
	pesos_i(11323) := b"0000000000000000_0000000000000000_0000000110101010_0010011111000100"; -- 0.006502614267126988
	pesos_i(11324) := b"1111111111111111_1111111111111111_1111010101110001_0100010101010010"; -- -0.04124037507017389
	pesos_i(11325) := b"1111111111111111_1111111111111111_1111001011110001_0011101110010011"; -- -0.05100658084508249
	pesos_i(11326) := b"0000000000000000_0000000000000000_0001010010100001_1111010001100001"; -- 0.08059623113112523
	pesos_i(11327) := b"0000000000000000_0000000000000000_0001111110100001_1111100000010001"; -- 0.1235652009645964
	pesos_i(11328) := b"0000000000000000_0000000000000000_0000000111101000_1110011111010001"; -- 0.007460106302500083
	pesos_i(11329) := b"0000000000000000_0000000000000000_0000011110010000_0001001111011000"; -- 0.02954219841419978
	pesos_i(11330) := b"0000000000000000_0000000000000000_0000100011011001_0101011110111001"; -- 0.03456638583985343
	pesos_i(11331) := b"0000000000000000_0000000000000000_0000010011010110_1001100001100010"; -- 0.01889946369328379
	pesos_i(11332) := b"0000000000000000_0000000000000000_0001010110010000_1111000110011000"; -- 0.0842429157289467
	pesos_i(11333) := b"1111111111111111_1111111111111111_1101110011011000_1010001000101101"; -- -0.13731943519117035
	pesos_i(11334) := b"1111111111111111_1111111111111111_1101111100100011_1010100100110101"; -- -0.1283621069488708
	pesos_i(11335) := b"1111111111111111_1111111111111111_1111000101011001_1001001001010010"; -- -0.05722699646662873
	pesos_i(11336) := b"0000000000000000_0000000000000000_0001101011000111_1010100011101011"; -- 0.10460906722775572
	pesos_i(11337) := b"1111111111111111_1111111111111111_1111000011000000_0100110100001010"; -- -0.059565720723672784
	pesos_i(11338) := b"1111111111111111_1111111111111111_1111110011111110_0111100101000100"; -- -0.011742039558680336
	pesos_i(11339) := b"0000000000000000_0000000000000000_0000110111110100_1000010100011110"; -- 0.054512328834296554
	pesos_i(11340) := b"1111111111111111_1111111111111111_1101110101001110_0000001110000010"; -- -0.13552835540480518
	pesos_i(11341) := b"0000000000000000_0000000000000000_0000001111000010_0001010000111011"; -- 0.014680160859112496
	pesos_i(11342) := b"0000000000000000_0000000000000000_0000100100101011_0110111100010100"; -- 0.03581899871854652
	pesos_i(11343) := b"1111111111111111_1111111111111111_1110001111001100_0010000110110001"; -- -0.11016644898322252
	pesos_i(11344) := b"0000000000000000_0000000000000000_0001010011010101_0110110100011111"; -- 0.08138162626321772
	pesos_i(11345) := b"0000000000000000_0000000000000000_0000001111011010_0011001111111110"; -- 0.015048265015646111
	pesos_i(11346) := b"0000000000000000_0000000000000000_0010010011001001_0101000111010101"; -- 0.14369689422210152
	pesos_i(11347) := b"1111111111111111_1111111111111111_1110110100110110_0100010101011100"; -- -0.07339064115535604
	pesos_i(11348) := b"0000000000000000_0000000000000000_0000101111101001_1000010110001111"; -- 0.04653200863280581
	pesos_i(11349) := b"1111111111111111_1111111111111111_1111010101010001_0000111110001011"; -- -0.04173186170429775
	pesos_i(11350) := b"0000000000000000_0000000000000000_0001011111100001_0001001110001011"; -- 0.09327814245530013
	pesos_i(11351) := b"1111111111111111_1111111111111111_1111110100001111_0011001010111000"; -- -0.011486845050357733
	pesos_i(11352) := b"0000000000000000_0000000000000000_0000010000010010_0001100001100001"; -- 0.0159011113052094
	pesos_i(11353) := b"1111111111111111_1111111111111111_1110101111100101_1001011101101011"; -- -0.07852796198220631
	pesos_i(11354) := b"1111111111111111_1111111111111111_1111100100101010_1111110110010101"; -- -0.026687766118861915
	pesos_i(11355) := b"0000000000000000_0000000000000000_0010100010000010_0001100110010110"; -- 0.1582351676063534
	pesos_i(11356) := b"0000000000000000_0000000000000000_0001001110011011_1000110111000111"; -- 0.07659231286952674
	pesos_i(11357) := b"1111111111111111_1111111111111111_1101110110010110_1001110000011111"; -- -0.13442062616926323
	pesos_i(11358) := b"1111111111111111_1111111111111111_1111110011101001_1111111000101101"; -- -0.012054552133411592
	pesos_i(11359) := b"0000000000000000_0000000000000000_0001110110110001_1000111001101000"; -- 0.11599054366754423
	pesos_i(11360) := b"1111111111111111_1111111111111111_1111110100110100_0110010111101010"; -- -0.01091921835891824
	pesos_i(11361) := b"1111111111111111_1111111111111111_1101110101001110_1000010101111010"; -- -0.13552060859480633
	pesos_i(11362) := b"1111111111111111_1111111111111111_1101111011101101_0100101001011110"; -- -0.12919173435904371
	pesos_i(11363) := b"1111111111111111_1111111111111111_1111001110100101_1110101010100110"; -- -0.048249563682895874
	pesos_i(11364) := b"0000000000000000_0000000000000000_0000111100011011_0100110010011100"; -- 0.05901030349070943
	pesos_i(11365) := b"1111111111111111_1111111111111111_1110111110101011_0001011100100100"; -- -0.06379561789198933
	pesos_i(11366) := b"0000000000000000_0000000000000000_0000110010010011_1010000000011001"; -- 0.049127584616064854
	pesos_i(11367) := b"1111111111111111_1111111111111111_1110001100001010_1000001111010110"; -- -0.113120803976165
	pesos_i(11368) := b"0000000000000000_0000000000000000_0000001010101110_0000111001010100"; -- 0.01046838329535775
	pesos_i(11369) := b"1111111111111111_1111111111111111_1101111100011100_0001111111001101"; -- -0.1284771084016741
	pesos_i(11370) := b"0000000000000000_0000000000000000_0001100001100101_0010001100010011"; -- 0.09529322826651868
	pesos_i(11371) := b"1111111111111111_1111111111111111_1110000101100011_1011111100111100"; -- -0.11957173149298035
	pesos_i(11372) := b"1111111111111111_1111111111111111_1111011101101110_1000010100101111"; -- -0.033469844803146215
	pesos_i(11373) := b"0000000000000000_0000000000000000_0010000111110101_0111000101100001"; -- 0.13265141127882077
	pesos_i(11374) := b"0000000000000000_0000000000000000_0001100011001100_1001110011010100"; -- 0.09687214067534546
	pesos_i(11375) := b"1111111111111111_1111111111111111_1110110111010000_1011100001000101"; -- -0.07103393866234405
	pesos_i(11376) := b"0000000000000000_0000000000000000_0000000111100010_1011101101010111"; -- 0.007365902622684984
	pesos_i(11377) := b"0000000000000000_0000000000000000_0000011011001101_1000101100101101"; -- 0.0265738473807386
	pesos_i(11378) := b"0000000000000000_0000000000000000_0000110110100100_1000101010101100"; -- 0.05329195686619967
	pesos_i(11379) := b"0000000000000000_0000000000000000_0000001011110010_0110001100011010"; -- 0.011511033775631428
	pesos_i(11380) := b"1111111111111111_1111111111111111_1111010100000111_1111000000100010"; -- -0.042847625540604416
	pesos_i(11381) := b"1111111111111111_1111111111111111_1111000001001100_1000010100011011"; -- -0.061332398334407845
	pesos_i(11382) := b"0000000000000000_0000000000000000_0001101001011010_0001001010110001"; -- 0.10293690513190559
	pesos_i(11383) := b"1111111111111111_1111111111111111_1101101110010010_0110110110111010"; -- -0.14229692667618407
	pesos_i(11384) := b"1111111111111111_1111111111111111_1111001101011001_1100111110000100"; -- -0.04941084879031552
	pesos_i(11385) := b"0000000000000000_0000000000000000_0000000101110100_0011001111110110"; -- 0.005679366668285261
	pesos_i(11386) := b"1111111111111111_1111111111111111_1111111001100111_0110101111100001"; -- -0.006234414703625635
	pesos_i(11387) := b"1111111111111111_1111111111111111_1101101100110010_1101110101101111"; -- -0.143755112031711
	pesos_i(11388) := b"1111111111111111_1111111111111111_1111111000010101_0000011111001000"; -- -0.0074916017066812505
	pesos_i(11389) := b"0000000000000000_0000000000000000_0001110101010001_1001001000101110"; -- 0.11452592487386616
	pesos_i(11390) := b"1111111111111111_1111111111111111_1110010010001000_0111001110010111"; -- -0.10729291489465125
	pesos_i(11391) := b"1111111111111111_1111111111111111_1110110101010100_0000111110000001"; -- -0.07293608769582724
	pesos_i(11392) := b"1111111111111111_1111111111111111_1111110110101001_0101111101001111"; -- -0.009134333702066911
	pesos_i(11393) := b"1111111111111111_1111111111111111_1111001011011110_0101111100011010"; -- -0.05129438035776851
	pesos_i(11394) := b"0000000000000000_0000000000000000_0001110100010110_1001000101110001"; -- 0.11362561229180035
	pesos_i(11395) := b"1111111111111111_1111111111111111_1110000100111010_0110100010110000"; -- -0.12020250033916273
	pesos_i(11396) := b"1111111111111111_1111111111111111_1111011010111110_0011011001011001"; -- -0.03616009073773511
	pesos_i(11397) := b"0000000000000000_0000000000000000_0001011000111110_0110001010000111"; -- 0.08688941766843464
	pesos_i(11398) := b"0000000000000000_0000000000000000_0000110100110101_1001100000110001"; -- 0.051599037224328785
	pesos_i(11399) := b"0000000000000000_0000000000000000_0000111100000000_1010010110001100"; -- 0.05860361746114501
	pesos_i(11400) := b"1111111111111111_1111111111111111_1110011000000111_0010000110101101"; -- -0.10145368133361544
	pesos_i(11401) := b"1111111111111111_1111111111111111_1111001100010010_1111100111111110"; -- -0.050491691038754664
	pesos_i(11402) := b"1111111111111111_1111111111111111_1111110110010010_0101100000011010"; -- -0.009485715475502672
	pesos_i(11403) := b"1111111111111111_1111111111111111_1110110001010011_1110111110101110"; -- -0.07684423455423903
	pesos_i(11404) := b"1111111111111111_1111111111111111_1101101010100011_1110011101011101"; -- -0.1459365270722026
	pesos_i(11405) := b"0000000000000000_0000000000000000_0001001101010001_0101000010111111"; -- 0.07545952480484218
	pesos_i(11406) := b"0000000000000000_0000000000000000_0000001111001110_0000110010111000"; -- 0.014862818569293647
	pesos_i(11407) := b"0000000000000000_0000000000000000_0001111011110111_1101110110001000"; -- 0.12096962510049797
	pesos_i(11408) := b"1111111111111111_1111111111111111_1111110100000110_1011001001001111"; -- -0.011616569193504223
	pesos_i(11409) := b"0000000000000000_0000000000000000_0000010101000101_1110010000111001"; -- 0.020597709666015415
	pesos_i(11410) := b"0000000000000000_0000000000000000_0000001110110100_0100100000111111"; -- 0.014469638339603557
	pesos_i(11411) := b"0000000000000000_0000000000000000_0000100011011011_0001111011110110"; -- 0.034593520163814985
	pesos_i(11412) := b"0000000000000000_0000000000000000_0000000100001111_1000110010101000"; -- 0.004143515639164013
	pesos_i(11413) := b"1111111111111111_1111111111111111_1111000010010101_0001011011000010"; -- -0.06022508386078193
	pesos_i(11414) := b"0000000000000000_0000000000000000_0000010000100010_1100000000101010"; -- 0.016155252651025027
	pesos_i(11415) := b"0000000000000000_0000000000000000_0001101110111111_1101000000101000"; -- 0.1083955858530612
	pesos_i(11416) := b"1111111111111111_1111111111111111_1101111001111010_0111010000001100"; -- -0.13094401085015242
	pesos_i(11417) := b"0000000000000000_0000000000000000_0001011101110001_0000101000001001"; -- 0.0915685914138432
	pesos_i(11418) := b"1111111111111111_1111111111111111_1101111100110001_0011010010111010"; -- -0.1281554266901253
	pesos_i(11419) := b"1111111111111111_1111111111111111_1101100100110001_0011010111100011"; -- -0.1515928573803821
	pesos_i(11420) := b"0000000000000000_0000000000000000_0000101101101000_1111111110100110"; -- 0.04457090180250424
	pesos_i(11421) := b"1111111111111111_1111111111111111_1101111111111110_0111001111110110"; -- -0.12502360565961637
	pesos_i(11422) := b"0000000000000000_0000000000000000_0010010101101111_1100011100000110"; -- 0.14623683840822926
	pesos_i(11423) := b"0000000000000000_0000000000000000_0010000100111111_0111010101110100"; -- 0.12987455436250175
	pesos_i(11424) := b"1111111111111111_1111111111111111_1111110100111111_0010101110000100"; -- -0.010754852522983801
	pesos_i(11425) := b"0000000000000000_0000000000000000_0000001010011000_1010100001101100"; -- 0.010141874734124976
	pesos_i(11426) := b"1111111111111111_1111111111111111_1110111101001000_1001100100000000"; -- -0.06529849775472281
	pesos_i(11427) := b"0000000000000000_0000000000000000_0010001111011101_0101001001111101"; -- 0.14009585900194949
	pesos_i(11428) := b"1111111111111111_1111111111111111_1111001000010101_1101111110000101"; -- -0.05435374261789856
	pesos_i(11429) := b"1111111111111111_1111111111111111_1110111000111001_0110000100101011"; -- -0.06943695727540616
	pesos_i(11430) := b"0000000000000000_0000000000000000_0001001111010101_0111110010100100"; -- 0.07747630128554224
	pesos_i(11431) := b"1111111111111111_1111111111111111_1110111110110000_1101110101100100"; -- -0.06370750723278652
	pesos_i(11432) := b"0000000000000000_0000000000000000_0000001001001111_0110111000011111"; -- 0.009024508113557277
	pesos_i(11433) := b"0000000000000000_0000000000000000_0000101110011100_0100011100101110"; -- 0.045353363744837234
	pesos_i(11434) := b"0000000000000000_0000000000000000_0000010111001101_1000101011010010"; -- 0.022667576106016135
	pesos_i(11435) := b"0000000000000000_0000000000000000_0000100110001000_1011101110110100"; -- 0.03724263332652857
	pesos_i(11436) := b"0000000000000000_0000000000000000_0001101000011001_1010110011101000"; -- 0.10195427574850403
	pesos_i(11437) := b"0000000000000000_0000000000000000_0001011101100010_0110100101101011"; -- 0.09134539472437914
	pesos_i(11438) := b"0000000000000000_0000000000000000_0001101111110001_0100101100011011"; -- 0.10915059482350449
	pesos_i(11439) := b"1111111111111111_1111111111111111_1111111100110110_0010101101001010"; -- -0.0030796951563247794
	pesos_i(11440) := b"1111111111111111_1111111111111111_1111101011100000_0010100000110010"; -- -0.020017135336876185
	pesos_i(11441) := b"1111111111111111_1111111111111111_1111100111001000_0110000000110110"; -- -0.024286257532498398
	pesos_i(11442) := b"1111111111111111_1111111111111111_1111110000110000_0011111011111101"; -- -0.01488882384330017
	pesos_i(11443) := b"0000000000000000_0000000000000000_0000111011011100_1100111111100100"; -- 0.05805682495171606
	pesos_i(11444) := b"1111111111111111_1111111111111111_1110100100011001_1011000010010111"; -- -0.08945175467059766
	pesos_i(11445) := b"1111111111111111_1111111111111111_1101111100100100_0101111001010001"; -- -0.12835131193009072
	pesos_i(11446) := b"1111111111111111_1111111111111111_1110000001000100_1000101111001110"; -- -0.12395406930292875
	pesos_i(11447) := b"1111111111111111_1111111111111111_1111011001001111_1000010111010100"; -- -0.03784907889208557
	pesos_i(11448) := b"1111111111111111_1111111111111111_1111110010101111_1110000001011011"; -- -0.012941339296018093
	pesos_i(11449) := b"0000000000000000_0000000000000000_0000110101111100_0101000000100101"; -- 0.052678116775346985
	pesos_i(11450) := b"0000000000000000_0000000000000000_0001000011000110_1110000001100010"; -- 0.06553461452154412
	pesos_i(11451) := b"1111111111111111_1111111111111111_1111101101101010_0101011110001000"; -- -0.017908600993952913
	pesos_i(11452) := b"1111111111111111_1111111111111111_1110011001111011_0111111000110101"; -- -0.099678146381939
	pesos_i(11453) := b"1111111111111111_1111111111111111_1111011000000110_1000100001001111"; -- -0.038962822708991915
	pesos_i(11454) := b"1111111111111111_1111111111111111_1110100101001000_0001000010000000"; -- -0.08874413379917769
	pesos_i(11455) := b"0000000000000000_0000000000000000_0000001011110000_0010111001101111"; -- 0.011477377135782594
	pesos_i(11456) := b"1111111111111111_1111111111111111_1101101010001100_1001101011101000"; -- -0.1462920363295023
	pesos_i(11457) := b"1111111111111111_1111111111111111_1101110111100100_1110100100000100"; -- -0.1332258573341005
	pesos_i(11458) := b"1111111111111111_1111111111111111_1110111000110110_0000111010001101"; -- -0.06948765811642199
	pesos_i(11459) := b"1111111111111111_1111111111111111_1101100100011111_1100100100111000"; -- -0.1518587340031316
	pesos_i(11460) := b"0000000000000000_0000000000000000_0001111110001001_0000011000110000"; -- 0.12318457293491966
	pesos_i(11461) := b"0000000000000000_0000000000000000_0001011101110011_0100010111111000"; -- 0.09160268113019343
	pesos_i(11462) := b"1111111111111111_1111111111111111_1111101011010110_1101101011110101"; -- -0.020159068210349712
	pesos_i(11463) := b"0000000000000000_0000000000000000_0000111001010101_1100000100100101"; -- 0.05599600940993674
	pesos_i(11464) := b"0000000000000000_0000000000000000_0000010010111010_1001101111000010"; -- 0.018472418682650243
	pesos_i(11465) := b"1111111111111111_1111111111111111_1111001101101110_1100010011000110"; -- -0.04909105458493579
	pesos_i(11466) := b"0000000000000000_0000000000000000_0001111110010101_0010101001000000"; -- 0.12336982783771135
	pesos_i(11467) := b"1111111111111111_1111111111111111_1101101000111011_0000100111100001"; -- -0.14753664268057942
	pesos_i(11468) := b"0000000000000000_0000000000000000_0000000111111100_0000001111001000"; -- 0.007751690300585347
	pesos_i(11469) := b"0000000000000000_0000000000000000_0010000111011010_1010110111001001"; -- 0.1322430243484112
	pesos_i(11470) := b"0000000000000000_0000000000000000_0001111011000000_0000001000100111"; -- 0.12011731586163696
	pesos_i(11471) := b"1111111111111111_1111111111111111_1111111110100101_0101011001110001"; -- -0.0013833975204452034
	pesos_i(11472) := b"1111111111111111_1111111111111111_1110111100011001_0101111100110010"; -- -0.06601910610186175
	pesos_i(11473) := b"1111111111111111_1111111111111111_1110110000010010_0010001101010100"; -- -0.07784823616358999
	pesos_i(11474) := b"0000000000000000_0000000000000000_0010000110110111_0101011011010100"; -- 0.1317037838691458
	pesos_i(11475) := b"0000000000000000_0000000000000000_0010000010111011_1100000101010001"; -- 0.1278649161731405
	pesos_i(11476) := b"1111111111111111_1111111111111111_1111000010001010_0010011000000010"; -- -0.060392021555946133
	pesos_i(11477) := b"1111111111111111_1111111111111111_1101101111011011_1001000100011101"; -- -0.14118092568011872
	pesos_i(11478) := b"0000000000000000_0000000000000000_0001101110000111_1001000000111110"; -- 0.10753728406049806
	pesos_i(11479) := b"1111111111111111_1111111111111111_1101100001111100_1010000100001001"; -- -0.15434831161754176
	pesos_i(11480) := b"1111111111111111_1111111111111111_1110000000001101_0010000100001010"; -- -0.12479966638347086
	pesos_i(11481) := b"1111111111111111_1111111111111111_1110000111011011_1101100110000111"; -- -0.11773910956997743
	pesos_i(11482) := b"0000000000000000_0000000000000000_0001100100110000_0010101111000100"; -- 0.09839128056570876
	pesos_i(11483) := b"0000000000000000_0000000000000000_0010010111111111_1010011001101101"; -- 0.14843216102451046
	pesos_i(11484) := b"0000000000000000_0000000000000000_0000100011000101_1011011110100111"; -- 0.0342669280563002
	pesos_i(11485) := b"0000000000000000_0000000000000000_0001111111101111_1101000101100100"; -- 0.12475308113745363
	pesos_i(11486) := b"1111111111111111_1111111111111111_1101111000010110_0011001100110010"; -- -0.13247375523828334
	pesos_i(11487) := b"1111111111111111_1111111111111111_1101100111111010_0111000100011111"; -- -0.14852231012807893
	pesos_i(11488) := b"1111111111111111_1111111111111111_1101100101010010_0000001100111111"; -- -0.15109233592886406
	pesos_i(11489) := b"0000000000000000_0000000000000000_0000001101100110_0101000101000100"; -- 0.013279990353683937
	pesos_i(11490) := b"1111111111111111_1111111111111111_1111110110000000_1011001101011011"; -- -0.009754934644384441
	pesos_i(11491) := b"1111111111111111_1111111111111111_1111001110000111_1101111100110101"; -- -0.048708009255053086
	pesos_i(11492) := b"1111111111111111_1111111111111111_1111001101110101_0111000000110001"; -- -0.04898928458744468
	pesos_i(11493) := b"0000000000000000_0000000000000000_0000000000011100_1010100001000011"; -- 0.0004372751807108219
	pesos_i(11494) := b"0000000000000000_0000000000000000_0001001010000100_1011000011110110"; -- 0.0723372079465088
	pesos_i(11495) := b"1111111111111111_1111111111111111_1101110011010111_0111110001111001"; -- -0.13733694123162107
	pesos_i(11496) := b"0000000000000000_0000000000000000_0000000111000010_1010100011110111"; -- 0.006876526065112118
	pesos_i(11497) := b"0000000000000000_0000000000000000_0000010100111010_1100101110011011"; -- 0.02042839568783781
	pesos_i(11498) := b"1111111111111111_1111111111111111_1111100011000100_0111001000111111"; -- -0.028252467700336122
	pesos_i(11499) := b"0000000000000000_0000000000000000_0010101101100111_0100111101100101"; -- 0.16954513761794784
	pesos_i(11500) := b"0000000000000000_0000000000000000_0001001110000011_0011011111100110"; -- 0.07622098320307062
	pesos_i(11501) := b"1111111111111111_1111111111111111_1110101100101101_0001101110111100"; -- -0.08134295129008802
	pesos_i(11502) := b"1111111111111111_1111111111111111_1111111010010110_1101110100100001"; -- -0.005510501246994025
	pesos_i(11503) := b"1111111111111111_1111111111111111_1101111111010010_0000111001101001"; -- -0.1257010454123975
	pesos_i(11504) := b"0000000000000000_0000000000000000_0000111101110010_0111000111010001"; -- 0.060340035965036634
	pesos_i(11505) := b"0000000000000000_0000000000000000_0000110110011010_1110100111101010"; -- 0.05314504580326922
	pesos_i(11506) := b"0000000000000000_0000000000000000_0010000000011110_0100111010110100"; -- 0.12546245477830376
	pesos_i(11507) := b"0000000000000000_0000000000000000_0000101011110011_1011011111001001"; -- 0.04278134015655147
	pesos_i(11508) := b"1111111111111111_1111111111111111_1101111000001011_1010100110111110"; -- -0.1326345358214684
	pesos_i(11509) := b"1111111111111111_1111111111111111_1110110001001010_1010010000010011"; -- -0.07698607000048208
	pesos_i(11510) := b"1111111111111111_1111111111111111_1110001010101111_1111100100010110"; -- -0.11450236518440393
	pesos_i(11511) := b"1111111111111111_1111111111111111_1110010001101000_1100001011000100"; -- -0.10777647710254153
	pesos_i(11512) := b"0000000000000000_0000000000000000_0001101011001110_1101111000001011"; -- 0.10471904522827645
	pesos_i(11513) := b"1111111111111111_1111111111111111_1110101001110110_0111110010010101"; -- -0.08412953723770986
	pesos_i(11514) := b"1111111111111111_1111111111111111_1101110110111010_1100001011110001"; -- -0.13386899574657404
	pesos_i(11515) := b"0000000000000000_0000000000000000_0001110011111001_1000101100010110"; -- 0.11318272872295226
	pesos_i(11516) := b"1111111111111111_1111111111111111_1110101000011000_0111111001100111"; -- -0.0855637548252067
	pesos_i(11517) := b"1111111111111111_1111111111111111_1111111000001111_0000100110000110"; -- -0.007583050571846778
	pesos_i(11518) := b"0000000000000000_0000000000000000_0010000011111111_0000001001101100"; -- 0.12889113567218452
	pesos_i(11519) := b"0000000000000000_0000000000000000_0000011110011011_1000011110100110"; -- 0.029716947651971706
	pesos_i(11520) := b"0000000000000000_0000000000000000_0001111001101011_0001100101101010"; -- 0.11882170532559874
	pesos_i(11521) := b"1111111111111111_1111111111111111_1111100111000010_0101011110010110"; -- -0.02437832445476195
	pesos_i(11522) := b"0000000000000000_0000000000000000_0000111001100100_1001011001100101"; -- 0.056222343117493766
	pesos_i(11523) := b"0000000000000000_0000000000000000_0001101110101110_1010010011110101"; -- 0.10813361141258479
	pesos_i(11524) := b"1111111111111111_1111111111111111_1110110111100011_1100001000000011"; -- -0.07074344094801353
	pesos_i(11525) := b"0000000000000000_0000000000000000_0001110000000101_1110000001100110"; -- 0.10946466920085329
	pesos_i(11526) := b"1111111111111111_1111111111111111_1111110011000110_0111100110000101"; -- -0.01259651654335769
	pesos_i(11527) := b"1111111111111111_1111111111111111_1110011110001010_1010000010011001"; -- -0.09554096471088462
	pesos_i(11528) := b"1111111111111111_1111111111111111_1111100001000011_1000001101101101"; -- -0.03021982754741562
	pesos_i(11529) := b"0000000000000000_0000000000000000_0000010111110110_1001100111100010"; -- 0.02329408433910961
	pesos_i(11530) := b"0000000000000000_0000000000000000_0000000100001000_1100100011110001"; -- 0.0040402973087102405
	pesos_i(11531) := b"0000000000000000_0000000000000000_0000101101110000_0011100001001001"; -- 0.044681089193318674
	pesos_i(11532) := b"0000000000000000_0000000000000000_0000110100001000_1101100110000111"; -- 0.05091628594396874
	pesos_i(11533) := b"0000000000000000_0000000000000000_0010010101111011_1010010010001011"; -- 0.1464178885398134
	pesos_i(11534) := b"1111111111111111_1111111111111111_1111100100111001_0001001010110000"; -- -0.02647288516254062
	pesos_i(11535) := b"0000000000000000_0000000000000000_0001000010000011_1011001100000011"; -- 0.06450957128502588
	pesos_i(11536) := b"1111111111111111_1111111111111111_1110101101101110_0110100110000010"; -- -0.08034649455546869
	pesos_i(11537) := b"1111111111111111_1111111111111111_1111101010101000_0110100010011101"; -- -0.02086778794269218
	pesos_i(11538) := b"1111111111111111_1111111111111111_1110110110111110_0010011000101100"; -- -0.07131730480988009
	pesos_i(11539) := b"1111111111111111_1111111111111111_1101110001110100_1110101010110111"; -- -0.13884099044724954
	pesos_i(11540) := b"1111111111111111_1111111111111111_1111001101100000_1001000011011001"; -- -0.04930777264462511
	pesos_i(11541) := b"0000000000000000_0000000000000000_0001001101110100_0011001100010000"; -- 0.07599181305372159
	pesos_i(11542) := b"0000000000000000_0000000000000000_0000001011110110_0010011001100001"; -- 0.011568449753767269
	pesos_i(11543) := b"0000000000000000_0000000000000000_0001001111011111_1110100101011011"; -- 0.07763536896742738
	pesos_i(11544) := b"0000000000000000_0000000000000000_0000011010101000_0011100010110100"; -- 0.026004356328256192
	pesos_i(11545) := b"0000000000000000_0000000000000000_0001000000111000_0011010010010001"; -- 0.06335762545525755
	pesos_i(11546) := b"0000000000000000_0000000000000000_0001010110000110_0011010110100011"; -- 0.0840791247421937
	pesos_i(11547) := b"0000000000000000_0000000000000000_0001101100000111_0111000000010010"; -- 0.10558224150804842
	pesos_i(11548) := b"1111111111111111_1111111111111111_1111001110000011_1000111100011010"; -- -0.048773819129791
	pesos_i(11549) := b"1111111111111111_1111111111111111_1111111100100100_1011011100100110"; -- -0.0033460171493950768
	pesos_i(11550) := b"1111111111111111_1111111111111111_1111000111010001_1100111001011010"; -- -0.05539236348416545
	pesos_i(11551) := b"0000000000000000_0000000000000000_0001110001101011_1110010001100011"; -- 0.11102130324036338
	pesos_i(11552) := b"0000000000000000_0000000000000000_0000100101111111_1000001110011101"; -- 0.0371019610834145
	pesos_i(11553) := b"1111111111111111_1111111111111111_1111111111111100_1010011000101000"; -- -5.1131468074906216e-05
	pesos_i(11554) := b"1111111111111111_1111111111111111_1110101000100010_0010111100111101"; -- -0.08541588554065516
	pesos_i(11555) := b"1111111111111111_1111111111111111_1110111110100100_1011010110110001"; -- -0.06389297889127211
	pesos_i(11556) := b"0000000000000000_0000000000000000_0001010101100100_1101111100110011"; -- 0.08357043264425185
	pesos_i(11557) := b"1111111111111111_1111111111111111_1101100010100000_0100010010111100"; -- -0.15380449685522193
	pesos_i(11558) := b"0000000000000000_0000000000000000_0000000101100010_0100011101011000"; -- 0.005405863754366707
	pesos_i(11559) := b"0000000000000000_0000000000000000_0000111111111010_0101011100100011"; -- 0.06241364111856618
	pesos_i(11560) := b"1111111111111111_1111111111111111_1111011001100110_1011100110101011"; -- -0.037495036817204244
	pesos_i(11561) := b"1111111111111111_1111111111111111_1111100001101010_1110101000001000"; -- -0.02961861904355653
	pesos_i(11562) := b"0000000000000000_0000000000000000_0000111110010011_1000100000111000"; -- 0.06084491121856866
	pesos_i(11563) := b"0000000000000000_0000000000000000_0001000001001111_0001000101110110"; -- 0.06370648509624526
	pesos_i(11564) := b"0000000000000000_0000000000000000_0000000000010010_0101111000001100"; -- 0.00028026390417365505
	pesos_i(11565) := b"0000000000000000_0000000000000000_0010000110010010_0011110010101011"; -- 0.13113764925003
	pesos_i(11566) := b"0000000000000000_0000000000000000_0001001001100100_0111011001101010"; -- 0.0718454370459213
	pesos_i(11567) := b"0000000000000000_0000000000000000_0001100001010001_0000101010101001"; -- 0.09498659721578512
	pesos_i(11568) := b"1111111111111111_1111111111111111_1101101101010001_1101101101001100"; -- -0.14328221690699208
	pesos_i(11569) := b"0000000000000000_0000000000000000_0000001001100000_0110000100101110"; -- 0.009283136096765864
	pesos_i(11570) := b"1111111111111111_1111111111111111_1110000010111011_0110011001010100"; -- -0.12214050727594275
	pesos_i(11571) := b"1111111111111111_1111111111111111_1111001111100010_0111101111110001"; -- -0.047325376159766036
	pesos_i(11572) := b"1111111111111111_1111111111111111_1111001010011101_0011010100001101"; -- -0.05228870806595989
	pesos_i(11573) := b"0000000000000000_0000000000000000_0010001010001100_0011101000000110"; -- 0.1349521889482467
	pesos_i(11574) := b"0000000000000000_0000000000000000_0000111010000001_1101111001101110"; -- 0.056669141599584756
	pesos_i(11575) := b"1111111111111111_1111111111111111_1110111100101100_1110010101011010"; -- -0.06572119285845039
	pesos_i(11576) := b"1111111111111111_1111111111111111_1111110011110100_0000000010100101"; -- -0.01190181704932343
	pesos_i(11577) := b"1111111111111111_1111111111111111_1110001001001010_0010010111111111"; -- -0.11605608479066865
	pesos_i(11578) := b"0000000000000000_0000000000000000_0001111101010100_1111101110101101"; -- 0.12239048928365417
	pesos_i(11579) := b"1111111111111111_1111111111111111_1110101001000001_1011001101000100"; -- -0.08493499372446486
	pesos_i(11580) := b"1111111111111111_1111111111111111_1110001011100001_0011111001101101"; -- -0.11375055153567933
	pesos_i(11581) := b"0000000000000000_0000000000000000_0000001110010011_0101101000010100"; -- 0.013967161065179083
	pesos_i(11582) := b"1111111111111111_1111111111111111_1111110010011011_1011100110101000"; -- -0.013248821763422378
	pesos_i(11583) := b"0000000000000000_0000000000000000_0001101001011100_1000010111011110"; -- 0.10297428777003603
	pesos_i(11584) := b"1111111111111111_1111111111111111_1111100101101001_1100001000111000"; -- -0.02573000090663707
	pesos_i(11585) := b"1111111111111111_1111111111111111_1110100010000111_0001001001011011"; -- -0.0916889694590604
	pesos_i(11586) := b"1111111111111111_1111111111111111_1110110001101110_0011000110101001"; -- -0.07644357317241463
	pesos_i(11587) := b"1111111111111111_1111111111111111_1111111011001000_1001001000101000"; -- -0.004752030696975861
	pesos_i(11588) := b"0000000000000000_0000000000000000_0001101001101000_0101011111101110"; -- 0.1031546550462991
	pesos_i(11589) := b"0000000000000000_0000000000000000_0000010010100010_0011001111001001"; -- 0.01810001050794282
	pesos_i(11590) := b"1111111111111111_1111111111111111_1111000010010010_1010000010011010"; -- -0.06026264429305009
	pesos_i(11591) := b"0000000000000000_0000000000000000_0001010001000010_1010100100111000"; -- 0.07914216625915359
	pesos_i(11592) := b"0000000000000000_0000000000000000_0001010111100100_0110101011101011"; -- 0.08551662682298487
	pesos_i(11593) := b"1111111111111111_1111111111111111_1111011111101101_0110110111001110"; -- -0.03153337216319185
	pesos_i(11594) := b"1111111111111111_1111111111111111_1110000010110011_1010010101111101"; -- -0.12225881281949841
	pesos_i(11595) := b"1111111111111111_1111111111111111_1110100101010100_0111111110100001"; -- -0.08855440438641397
	pesos_i(11596) := b"1111111111111111_1111111111111111_1101110000010100_1101110000111101"; -- -0.14030669708011448
	pesos_i(11597) := b"1111111111111111_1111111111111111_1110110111111110_0011100000111010"; -- -0.07033966622629609
	pesos_i(11598) := b"1111111111111111_1111111111111111_1110111101000001_0011010000110011"; -- -0.06541131749208916
	pesos_i(11599) := b"1111111111111111_1111111111111111_1110101110010010_0010100011001110"; -- -0.07980103454985307
	pesos_i(11600) := b"0000000000000000_0000000000000000_0001101101111100_0010111001001010"; -- 0.10736359883445556
	pesos_i(11601) := b"0000000000000000_0000000000000000_0000011010101011_1110010010101010"; -- 0.026060382360803668
	pesos_i(11602) := b"1111111111111111_1111111111111111_1111010110010100_0101110001100001"; -- -0.04070494310560705
	pesos_i(11603) := b"1111111111111111_1111111111111111_1110001010010111_1111010010010111"; -- -0.11486884427635907
	pesos_i(11604) := b"1111111111111111_1111111111111111_1111001101000110_0110000110010010"; -- -0.04970731921986482
	pesos_i(11605) := b"1111111111111111_1111111111111111_1111101111000001_1100101111100111"; -- -0.016574150263066367
	pesos_i(11606) := b"1111111111111111_1111111111111111_1111100011011101_1011001001010101"; -- -0.02786717824488191
	pesos_i(11607) := b"1111111111111111_1111111111111111_1111001001000100_1010000010110010"; -- -0.05364032411717945
	pesos_i(11608) := b"1111111111111111_1111111111111111_1110001100011111_1100011001011110"; -- -0.11279640389632692
	pesos_i(11609) := b"0000000000000000_0000000000000000_0010011110100000_1011010111101000"; -- 0.1547959988190073
	pesos_i(11610) := b"0000000000000000_0000000000000000_0000111011001111_0001100000011010"; -- 0.05784750597823123
	pesos_i(11611) := b"1111111111111111_1111111111111111_1111000011011011_1010100111111001"; -- -0.05914819395795832
	pesos_i(11612) := b"1111111111111111_1111111111111111_1111001000111110_1001001001010001"; -- -0.05373273383269012
	pesos_i(11613) := b"1111111111111111_1111111111111111_1101111011011000_0000000111011110"; -- -0.1295164902477314
	pesos_i(11614) := b"0000000000000000_0000000000000000_0000000000101100_1001100011010111"; -- 0.0006804966912767431
	pesos_i(11615) := b"0000000000000000_0000000000000000_0010001000111011_0101011010011111"; -- 0.13371793166195284
	pesos_i(11616) := b"1111111111111111_1111111111111111_1111110111000010_0001100111001011"; -- -0.008757007448973054
	pesos_i(11617) := b"1111111111111111_1111111111111111_1111100111010110_1110010110111001"; -- -0.024064676495110897
	pesos_i(11618) := b"0000000000000000_0000000000000000_0001001111000011_0000001000111111"; -- 0.07719434775605524
	pesos_i(11619) := b"0000000000000000_0000000000000000_0000110100010010_1100000001110111"; -- 0.0510673800406812
	pesos_i(11620) := b"1111111111111111_1111111111111111_1111000011010011_0101001111001010"; -- -0.0592754013677721
	pesos_i(11621) := b"1111111111111111_1111111111111111_1111011010000000_1110011010101000"; -- -0.03709562676785753
	pesos_i(11622) := b"0000000000000000_0000000000000000_0000001110111100_1000100000110101"; -- 0.014595521030844332
	pesos_i(11623) := b"0000000000000000_0000000000000000_0001110010000010_0001000010110111"; -- 0.11135963880405618
	pesos_i(11624) := b"0000000000000000_0000000000000000_0001010101111111_1000011001101110"; -- 0.08397712875811614
	pesos_i(11625) := b"0000000000000000_0000000000000000_0000010001000011_0100010011101101"; -- 0.01665144719238954
	pesos_i(11626) := b"0000000000000000_0000000000000000_0001110000001101_1110010001100101"; -- 0.1095869775467445
	pesos_i(11627) := b"1111111111111111_1111111111111111_1101111000100001_1001011110111000"; -- -0.13229991674266464
	pesos_i(11628) := b"1111111111111111_1111111111111111_1110110000100111_1011011101101101"; -- -0.07751897420005893
	pesos_i(11629) := b"0000000000000000_0000000000000000_0000111010000111_1010111000010100"; -- 0.05675781230215912
	pesos_i(11630) := b"0000000000000000_0000000000000000_0000000010011101_0110000111010001"; -- 0.002401460148199912
	pesos_i(11631) := b"1111111111111111_1111111111111111_1111111111010111_0101111000001011"; -- -0.0006200048640872514
	pesos_i(11632) := b"0000000000000000_0000000000000000_0001101100101100_0100101000101110"; -- 0.10614455815711543
	pesos_i(11633) := b"1111111111111111_1111111111111111_1111110011001000_0111011100110110"; -- -0.01256613671688959
	pesos_i(11634) := b"0000000000000000_0000000000000000_0010000101001001_1110110011001010"; -- 0.13003425537273214
	pesos_i(11635) := b"1111111111111111_1111111111111111_1111000001101100_1011100100101001"; -- -0.060841014307480575
	pesos_i(11636) := b"1111111111111111_1111111111111111_1101111100010100_1010111010000100"; -- -0.12859067224225196
	pesos_i(11637) := b"1111111111111111_1111111111111111_1110010011011011_1001100010001011"; -- -0.10602423286322107
	pesos_i(11638) := b"1111111111111111_1111111111111111_1111110101110000_0011110011100110"; -- -0.010006135689436748
	pesos_i(11639) := b"1111111111111111_1111111111111111_1101101101011100_1100111011110110"; -- -0.14311510549018708
	pesos_i(11640) := b"0000000000000000_0000000000000000_0000101010101011_1101101111110101"; -- 0.04168486343119154
	pesos_i(11641) := b"1111111111111111_1111111111111111_1110100001101011_0001111111000000"; -- -0.09211541714510578
	pesos_i(11642) := b"0000000000000000_0000000000000000_0001010100111100_0000000001010110"; -- 0.0829467973134759
	pesos_i(11643) := b"1111111111111111_1111111111111111_1101111010100111_1011000111010011"; -- -0.13025368304070115
	pesos_i(11644) := b"0000000000000000_0000000000000000_0010011100000011_0011100111110100"; -- 0.1523929806585414
	pesos_i(11645) := b"0000000000000000_0000000000000000_0000010011001111_0100001111111000"; -- 0.0187876204823321
	pesos_i(11646) := b"1111111111111111_1111111111111111_1111010010100111_1000011110010000"; -- -0.044318702030092354
	pesos_i(11647) := b"1111111111111111_1111111111111111_1111110111000111_0001100001010110"; -- -0.008680800490298617
	pesos_i(11648) := b"1111111111111111_1111111111111111_1101101011001011_0011000100111100"; -- -0.14533703119131558
	pesos_i(11649) := b"0000000000000000_0000000000000000_0001000000110011_0000001110010000"; -- 0.06327841069999783
	pesos_i(11650) := b"1111111111111111_1111111111111111_1101110000000001_0011010101010010"; -- -0.1406065629626821
	pesos_i(11651) := b"0000000000000000_0000000000000000_0010100001111101_0000011011001000"; -- 0.1581577528088904
	pesos_i(11652) := b"0000000000000000_0000000000000000_0001110011000110_0110010010010101"; -- 0.11240223535781654
	pesos_i(11653) := b"0000000000000000_0000000000000000_0001011111110000_1110011111011110"; -- 0.09351967984184312
	pesos_i(11654) := b"0000000000000000_0000000000000000_0000110110111110_1101110111101011"; -- 0.053693647228532225
	pesos_i(11655) := b"1111111111111111_1111111111111111_1111010101111101_1101101010000111"; -- -0.04104837608758617
	pesos_i(11656) := b"1111111111111111_1111111111111111_1101100010000011_1000010101000110"; -- -0.15424315489859178
	pesos_i(11657) := b"0000000000000000_0000000000000000_0001100101000100_1101001111010110"; -- 0.09870647414040568
	pesos_i(11658) := b"0000000000000000_0000000000000000_0001101110001001_1000100010010010"; -- 0.10756734438837377
	pesos_i(11659) := b"0000000000000000_0000000000000000_0010001110011000_1010110100100001"; -- 0.13904840529580492
	pesos_i(11660) := b"0000000000000000_0000000000000000_0001111001110110_0001001101100100"; -- 0.11898919276938472
	pesos_i(11661) := b"0000000000000000_0000000000000000_0001000111101100_0111111111000101"; -- 0.07001493986903706
	pesos_i(11662) := b"1111111111111111_1111111111111111_1111010111111111_1001010100011101"; -- -0.03906887083687689
	pesos_i(11663) := b"1111111111111111_1111111111111111_1111101001110111_1010010101000001"; -- -0.021611854304208533
	pesos_i(11664) := b"1111111111111111_1111111111111111_1111101000000000_0000101011001001"; -- -0.0234368570453741
	pesos_i(11665) := b"0000000000000000_0000000000000000_0000110001000110_0011001000110010"; -- 0.04794610706407903
	pesos_i(11666) := b"1111111111111111_1111111111111111_1110111000111001_0010001001100011"; -- -0.06944069949068846
	pesos_i(11667) := b"1111111111111111_1111111111111111_1101111111011001_1010101100110110"; -- -0.12558488777236762
	pesos_i(11668) := b"1111111111111111_1111111111111111_1111011100101101_1110010100011100"; -- -0.03445594843928727
	pesos_i(11669) := b"0000000000000000_0000000000000000_0000100010100111_0010011101010111"; -- 0.03380056252072706
	pesos_i(11670) := b"0000000000000000_0000000000000000_0001101011100010_0110101100001101"; -- 0.10501736696713408
	pesos_i(11671) := b"1111111111111111_1111111111111111_1111011100100101_0010010101011001"; -- -0.03458944862851266
	pesos_i(11672) := b"1111111111111111_1111111111111111_1110000011011101_1100111001000110"; -- -0.12161551280342524
	pesos_i(11673) := b"0000000000000000_0000000000000000_0000110010010100_1111010000000000"; -- 0.04914784425908109
	pesos_i(11674) := b"0000000000000000_0000000000000000_0010011101111101_0010100011011101"; -- 0.15425353418564058
	pesos_i(11675) := b"0000000000000000_0000000000000000_0001010000111001_0111010101100110"; -- 0.07900174840652527
	pesos_i(11676) := b"1111111111111111_1111111111111111_1110110000110000_1001001100101001"; -- -0.07738380666968658
	pesos_i(11677) := b"1111111111111111_1111111111111111_1111100010010100_0111001001100010"; -- -0.028984881397329933
	pesos_i(11678) := b"0000000000000000_0000000000000000_0001000011111000_0010010101001111"; -- 0.066286403461401
	pesos_i(11679) := b"1111111111111111_1111111111111111_1111110011110100_0011001011111010"; -- -0.011898817136664947
	pesos_i(11680) := b"1111111111111111_1111111111111111_1111010010100100_1110010011111000"; -- -0.04435891107414471
	pesos_i(11681) := b"1111111111111111_1111111111111111_1101110101100000_1000100001111101"; -- -0.1352457709378754
	pesos_i(11682) := b"1111111111111111_1111111111111111_1110000000000011_0100011110100110"; -- -0.12494995315220818
	pesos_i(11683) := b"0000000000000000_0000000000000000_0001101110111111_0111111111100011"; -- 0.10839080123716406
	pesos_i(11684) := b"0000000000000000_0000000000000000_0010001010111110_1101000011000111"; -- 0.1357241139464708
	pesos_i(11685) := b"0000000000000000_0000000000000000_0010000101101110_0110100000111101"; -- 0.13059092997270427
	pesos_i(11686) := b"1111111111111111_1111111111111111_1101100110001111_0111010000000010"; -- -0.1501548286090247
	pesos_i(11687) := b"1111111111111111_1111111111111111_1101110101001101_0011000110000011"; -- -0.13554087204123672
	pesos_i(11688) := b"1111111111111111_1111111111111111_1111111101001101_0011011011110000"; -- -0.0027280486835342317
	pesos_i(11689) := b"1111111111111111_1111111111111111_1110010010001101_1001010100010011"; -- -0.10721462529921182
	pesos_i(11690) := b"0000000000000000_0000000000000000_0000110101010100_0000100100010101"; -- 0.05206352971734989
	pesos_i(11691) := b"0000000000000000_0000000000000000_0001000111000010_1000111101000101"; -- 0.06937499454840908
	pesos_i(11692) := b"0000000000000000_0000000000000000_0000111010001000_1010000110100100"; -- 0.0567723298619873
	pesos_i(11693) := b"0000000000000000_0000000000000000_0001010000010111_1010100100011101"; -- 0.07848603202577888
	pesos_i(11694) := b"0000000000000000_0000000000000000_0000101010000111_1000001011001010"; -- 0.041130232212980976
	pesos_i(11695) := b"1111111111111111_1111111111111111_1110010101101101_1001000110111101"; -- -0.10379685532948359
	pesos_i(11696) := b"0000000000000000_0000000000000000_0000110100010010_0111001011101100"; -- 0.05106275799554721
	pesos_i(11697) := b"0000000000000000_0000000000000000_0000101010101111_0000000100001101"; -- 0.041732850752436684
	pesos_i(11698) := b"0000000000000000_0000000000000000_0000110000010001_1110111110010111"; -- 0.04714868007464191
	pesos_i(11699) := b"0000000000000000_0000000000000000_0001101011100100_0001011010001111"; -- 0.10504284847243135
	pesos_i(11700) := b"0000000000000000_0000000000000000_0001010001011001_0111010000011111"; -- 0.07948995350262679
	pesos_i(11701) := b"1111111111111111_1111111111111111_1101111010100011_1100101111001001"; -- -0.13031317088027147
	pesos_i(11702) := b"0000000000000000_0000000000000000_0001011101000101_0001000110001111"; -- 0.09089765306599537
	pesos_i(11703) := b"0000000000000000_0000000000000000_0000001010111110_1100100001001001"; -- 0.010723607886369616
	pesos_i(11704) := b"1111111111111111_1111111111111111_1111110100001101_0110100010001100"; -- -0.011514154345845752
	pesos_i(11705) := b"0000000000000000_0000000000000000_0010001001101001_1100100001010100"; -- 0.13442661325902644
	pesos_i(11706) := b"0000000000000000_0000000000000000_0010001001110001_1000101111101101"; -- 0.13454508330328552
	pesos_i(11707) := b"0000000000000000_0000000000000000_0000100011100101_0110010001100101"; -- 0.03475024663333881
	pesos_i(11708) := b"0000000000000000_0000000000000000_0001100111010000_1110001011010011"; -- 0.10084359788459396
	pesos_i(11709) := b"1111111111111111_1111111111111111_1111111001011001_0011111101001101"; -- -0.006450694829335954
	pesos_i(11710) := b"1111111111111111_1111111111111111_1110010001011011_1111010111101001"; -- -0.10797179291774056
	pesos_i(11711) := b"1111111111111111_1111111111111111_1111010010110001_1101001101001001"; -- -0.04416160083664833
	pesos_i(11712) := b"1111111111111111_1111111111111111_1111000110000001_1000011000101101"; -- -0.0566173687538738
	pesos_i(11713) := b"0000000000000000_0000000000000000_0001111101101011_1011100111101101"; -- 0.12273752241150487
	pesos_i(11714) := b"1111111111111111_1111111111111111_1110110011011100_0111101100000000"; -- -0.07476073502246677
	pesos_i(11715) := b"0000000000000000_0000000000000000_0010010100000011_0000110001101010"; -- 0.1445777664080443
	pesos_i(11716) := b"0000000000000000_0000000000000000_0000111000101011_1011100111100101"; -- 0.05535470816081989
	pesos_i(11717) := b"0000000000000000_0000000000000000_0000100001101110_1111110010110001"; -- 0.0329435283809148
	pesos_i(11718) := b"0000000000000000_0000000000000000_0001001000000011_0111100111001011"; -- 0.07036553589402915
	pesos_i(11719) := b"1111111111111111_1111111111111111_1101101010100000_0100001110000111"; -- -0.14599206869800974
	pesos_i(11720) := b"0000000000000000_0000000000000000_0000111101111101_1011110111101110"; -- 0.06051241933276148
	pesos_i(11721) := b"1111111111111111_1111111111111111_1101110100000111_1000101110110000"; -- -0.13660361254415096
	pesos_i(11722) := b"1111111111111111_1111111111111111_1110010101110101_1110101001110000"; -- -0.10366949804058684
	pesos_i(11723) := b"0000000000000000_0000000000000000_0001000011110010_1011010010101000"; -- 0.06620339489052904
	pesos_i(11724) := b"0000000000000000_0000000000000000_0000001011010110_1010100001001101"; -- 0.011087912461464781
	pesos_i(11725) := b"1111111111111111_1111111111111111_1111100001110110_0110111000000001"; -- -0.029442906135953892
	pesos_i(11726) := b"0000000000000000_0000000000000000_0010010001101010_0100010010001010"; -- 0.14224651697516102
	pesos_i(11727) := b"1111111111111111_1111111111111111_1101101000011011_1011101111001011"; -- -0.14801431938046686
	pesos_i(11728) := b"0000000000000000_0000000000000000_0001101010101001_0101010100111001"; -- 0.10414631504133019
	pesos_i(11729) := b"1111111111111111_1111111111111111_1110101000101001_1111010011101011"; -- -0.08529729129361815
	pesos_i(11730) := b"1111111111111111_1111111111111111_1110110111010111_1011001010010101"; -- -0.07092746593433522
	pesos_i(11731) := b"0000000000000000_0000000000000000_0010000111110011_0101010010111011"; -- 0.1326191860686871
	pesos_i(11732) := b"0000000000000000_0000000000000000_0001110101110100_1101010011011101"; -- 0.1150639572774041
	pesos_i(11733) := b"1111111111111111_1111111111111111_1101110011011011_1000001101100110"; -- -0.1372754933417498
	pesos_i(11734) := b"0000000000000000_0000000000000000_0000100101010010_0011111011001100"; -- 0.03641121365727461
	pesos_i(11735) := b"0000000000000000_0000000000000000_0001011001101000_1111110111011110"; -- 0.0875395457536453
	pesos_i(11736) := b"1111111111111111_1111111111111111_1110100100011001_1010100111001100"; -- -0.0894521596405853
	pesos_i(11737) := b"0000000000000000_0000000000000000_0000001111001000_0010110111100101"; -- 0.014773243434179918
	pesos_i(11738) := b"1111111111111111_1111111111111111_1110001011011000_1000010110010101"; -- -0.1138836393974552
	pesos_i(11739) := b"1111111111111111_1111111111111111_1111011001010000_1011111011000110"; -- -0.03783042594611315
	pesos_i(11740) := b"0000000000000000_0000000000000000_0001101011110011_1110000011011110"; -- 0.10528378876002326
	pesos_i(11741) := b"1111111111111111_1111111111111111_1110001001000111_0110101000000000"; -- -0.11609780790837812
	pesos_i(11742) := b"0000000000000000_0000000000000000_0010110111101101_1011111000110100"; -- 0.17940891989158958
	pesos_i(11743) := b"0000000000000000_0000000000000000_0000100000001010_0101001001101111"; -- 0.03140750137128965
	pesos_i(11744) := b"0000000000000000_0000000000000000_0001010011010000_1101011001000011"; -- 0.08131159916315386
	pesos_i(11745) := b"0000000000000000_0000000000000000_0000011111101110_1010000011101110"; -- 0.030984933898544856
	pesos_i(11746) := b"1111111111111111_1111111111111111_1110011101100000_1010000100000100"; -- -0.09618180892887696
	pesos_i(11747) := b"1111111111111111_1111111111111111_1110010100000001_1101001010110000"; -- -0.10544093330038347
	pesos_i(11748) := b"0000000000000000_0000000000000000_0001111100000101_0000110010001101"; -- 0.12117079194014439
	pesos_i(11749) := b"0000000000000000_0000000000000000_0001000110000111_0000000000000100"; -- 0.06846618752009397
	pesos_i(11750) := b"0000000000000000_0000000000000000_0001000101001101_1100001010011011"; -- 0.06759277611443468
	pesos_i(11751) := b"0000000000000000_0000000000000000_0000001010001110_1110000010010111"; -- 0.00999263470634789
	pesos_i(11752) := b"0000000000000000_0000000000000000_0010000110101111_1010001000010101"; -- 0.13158619899776017
	pesos_i(11753) := b"0000000000000000_0000000000000000_0001011101010010_1011110011011001"; -- 0.09110622699565421
	pesos_i(11754) := b"1111111111111111_1111111111111111_1111110010110111_1010011000010111"; -- -0.012822741831821284
	pesos_i(11755) := b"1111111111111111_1111111111111111_1111110010010111_0010011111010101"; -- -0.013318548669453482
	pesos_i(11756) := b"1111111111111111_1111111111111111_1111011101101000_1000000101001010"; -- -0.033561629687417896
	pesos_i(11757) := b"1111111111111111_1111111111111111_1110001000101011_0111110001101011"; -- -0.11652395620644124
	pesos_i(11758) := b"1111111111111111_1111111111111111_1111110001101110_0111000101000001"; -- -0.01393978284931968
	pesos_i(11759) := b"1111111111111111_1111111111111111_1111111010101000_0000110100011001"; -- -0.005248242676977386
	pesos_i(11760) := b"1111111111111111_1111111111111111_1110000010000001_0111101111101001"; -- -0.12302423051160286
	pesos_i(11761) := b"0000000000000000_0000000000000000_0000001101100101_0010000101011111"; -- 0.013261876710432986
	pesos_i(11762) := b"1111111111111111_1111111111111111_1101110010011010_0100010100010100"; -- -0.13827102899393728
	pesos_i(11763) := b"0000000000000000_0000000000000000_0000000110000010_0110000000101101"; -- 0.005895625047235699
	pesos_i(11764) := b"0000000000000000_0000000000000000_0001100000101110_1110010001000101"; -- 0.09446551026218136
	pesos_i(11765) := b"1111111111111111_1111111111111111_1111110110000001_1000100110011100"; -- -0.009742164097404306
	pesos_i(11766) := b"1111111111111111_1111111111111111_1110101110010110_0111011110010001"; -- -0.07973530501489963
	pesos_i(11767) := b"1111111111111111_1111111111111111_1111100001001101_1001101100010110"; -- -0.030065829304869444
	pesos_i(11768) := b"0000000000000000_0000000000000000_0000100101110100_1111010011100110"; -- 0.0369408665236322
	pesos_i(11769) := b"0000000000000000_0000000000000000_0000110000001101_1100101001101100"; -- 0.04708542961185046
	pesos_i(11770) := b"1111111111111111_1111111111111111_1110011010010000_1010110111111111"; -- -0.09935486328743161
	pesos_i(11771) := b"1111111111111111_1111111111111111_1111100001101001_0010110011011111"; -- -0.029645152718971376
	pesos_i(11772) := b"0000000000000000_0000000000000000_0001101100010110_1101011001000110"; -- 0.1058172149470574
	pesos_i(11773) := b"1111111111111111_1111111111111111_1101110101011101_1000011010110110"; -- -0.13529165326420145
	pesos_i(11774) := b"1111111111111111_1111111111111111_1110000100100110_1010000101001100"; -- -0.12050430190873995
	pesos_i(11775) := b"0000000000000000_0000000000000000_0000000100100011_1011100011100100"; -- 0.0044513278464158494
	pesos_i(11776) := b"0000000000000000_0000000000000000_0000000111110101_1001110101001001"; -- 0.00765402824917872
	pesos_i(11777) := b"1111111111111111_1111111111111111_1101111111110010_1101100111001001"; -- -0.12520064194876337
	pesos_i(11778) := b"0000000000000000_0000000000000000_0010001010111001_1001000110001000"; -- 0.13564405034743282
	pesos_i(11779) := b"0000000000000000_0000000000000000_0001000111110010_1101110000100001"; -- 0.07011199772854217
	pesos_i(11780) := b"1111111111111111_1111111111111111_1110000110110010_0111001100011101"; -- -0.11837082428595415
	pesos_i(11781) := b"1111111111111111_1111111111111111_1111100000111111_0011101110001110"; -- -0.030285146511260564
	pesos_i(11782) := b"0000000000000000_0000000000000000_0001111110000011_1000111010111110"; -- 0.1231011595632608
	pesos_i(11783) := b"0000000000000000_0000000000000000_0000101111000000_1110100110011111"; -- 0.045912362323308226
	pesos_i(11784) := b"1111111111111111_1111111111111111_1111000100100001_0111110001100011"; -- -0.05808279604513611
	pesos_i(11785) := b"1111111111111111_1111111111111111_1111000110101000_0000010001001101"; -- -0.05603001702953926
	pesos_i(11786) := b"1111111111111111_1111111111111111_1111011010011011_1101100001000000"; -- -0.03668449827377395
	pesos_i(11787) := b"1111111111111111_1111111111111111_1110101010110111_0110111111111001"; -- -0.08313846745279388
	pesos_i(11788) := b"1111111111111111_1111111111111111_1110101001111001_0000010001111111"; -- -0.08409091849311356
	pesos_i(11789) := b"0000000000000000_0000000000000000_0010010101001010_0110110001100010"; -- 0.14566686054381126
	pesos_i(11790) := b"0000000000000000_0000000000000000_0001010101100011_0101011111111110"; -- 0.08354711487681053
	pesos_i(11791) := b"0000000000000000_0000000000000000_0000000110100110_0001101111010011"; -- 0.0064408674371105226
	pesos_i(11792) := b"1111111111111111_1111111111111111_1111110100110101_1111101100101110"; -- -0.010895062803946743
	pesos_i(11793) := b"1111111111111111_1111111111111111_1111001100000010_0100010000101111"; -- -0.05074666829491503
	pesos_i(11794) := b"1111111111111111_1111111111111111_1110111110001101_1110000000111111"; -- -0.06424139469597101
	pesos_i(11795) := b"1111111111111111_1111111111111111_1111011010010011_0101011010000001"; -- -0.03681430201159333
	pesos_i(11796) := b"0000000000000000_0000000000000000_0000010111110101_0101110110010100"; -- 0.023275231075445945
	pesos_i(11797) := b"1111111111111111_1111111111111111_1111010001111001_1110011000011000"; -- -0.045014971953697976
	pesos_i(11798) := b"0000000000000000_0000000000000000_0000100110001010_1110011100100001"; -- 0.03727573915164434
	pesos_i(11799) := b"1111111111111111_1111111111111111_1110001000101000_1001001101000000"; -- -0.11656837171413574
	pesos_i(11800) := b"1111111111111111_1111111111111111_1110111110111110_0000111100001101"; -- -0.06350618301725773
	pesos_i(11801) := b"1111111111111111_1111111111111111_1111011011111001_0011010001000000"; -- -0.03525994717157518
	pesos_i(11802) := b"0000000000000000_0000000000000000_0010001010111011_1101111110010110"; -- 0.13567922034360066
	pesos_i(11803) := b"0000000000000000_0000000000000000_0010000111000011_0110100001001010"; -- 0.13188792987310557
	pesos_i(11804) := b"1111111111111111_1111111111111111_1110100100010111_1001011101110001"; -- -0.08948377133610262
	pesos_i(11805) := b"1111111111111111_1111111111111111_1111011111100110_1000111001100110"; -- -0.03163824090767607
	pesos_i(11806) := b"1111111111111111_1111111111111111_1110100111110011_0101010010110101"; -- -0.08613081540884268
	pesos_i(11807) := b"1111111111111111_1111111111111111_1110010010110111_0111111000000111"; -- -0.10657512984233465
	pesos_i(11808) := b"0000000000000000_0000000000000000_0010001101100011_1011001000011100"; -- 0.13823998631168202
	pesos_i(11809) := b"1111111111111111_1111111111111111_1110110010000010_0111100100111001"; -- -0.07613413188549854
	pesos_i(11810) := b"0000000000000000_0000000000000000_0000001000110111_0011101101110110"; -- 0.008655277451247919
	pesos_i(11811) := b"1111111111111111_1111111111111111_1111100111100110_1011101101001110"; -- -0.023823064277477254
	pesos_i(11812) := b"1111111111111111_1111111111111111_1111000000001001_1111011010001001"; -- -0.06234797636932497
	pesos_i(11813) := b"1111111111111111_1111111111111111_1111100001101000_0100111010000111"; -- -0.02965840523689206
	pesos_i(11814) := b"0000000000000000_0000000000000000_0000110110011111_1101111111010001"; -- 0.053220737842696604
	pesos_i(11815) := b"1111111111111111_1111111111111111_1110111011101100_0000000101011111"; -- -0.06671134396748735
	pesos_i(11816) := b"0000000000000000_0000000000000000_0000010011101110_0101110000100110"; -- 0.01926208421491137
	pesos_i(11817) := b"0000000000000000_0000000000000000_0000110100111011_1101010011010101"; -- 0.05169420436635077
	pesos_i(11818) := b"0000000000000000_0000000000000000_0001000000111101_0100111100101100"; -- 0.06343550505042346
	pesos_i(11819) := b"1111111111111111_1111111111111111_1111110000001111_1000101011100010"; -- -0.015387840101803451
	pesos_i(11820) := b"1111111111111111_1111111111111111_1111001001010101_1100101100011110"; -- -0.05337839619219047
	pesos_i(11821) := b"1111111111111111_1111111111111111_1111011101110000_0110101111000110"; -- -0.033440841902585165
	pesos_i(11822) := b"1111111111111111_1111111111111111_1110101000001100_0101001000011000"; -- -0.0857495013958841
	pesos_i(11823) := b"0000000000000000_0000000000000000_0000110101110011_0010010000001010"; -- 0.05253815876815618
	pesos_i(11824) := b"1111111111111111_1111111111111111_1101110101011011_0110111110111101"; -- -0.1353235401424948
	pesos_i(11825) := b"1111111111111111_1111111111111111_1101111111101010_0011000100011110"; -- -0.12533276578523453
	pesos_i(11826) := b"0000000000000000_0000000000000000_0000101011110111_0001101001101011"; -- 0.04283299555071795
	pesos_i(11827) := b"1111111111111111_1111111111111111_1111001011100011_1111101010111111"; -- -0.051208809244877584
	pesos_i(11828) := b"0000000000000000_0000000000000000_0010000001100010_0001111101001000"; -- 0.12649722577135447
	pesos_i(11829) := b"0000000000000000_0000000000000000_0000110010010110_0000001101010110"; -- 0.04916401709606869
	pesos_i(11830) := b"0000000000000000_0000000000000000_0010011101100000_0011100101101000"; -- 0.1538120155381419
	pesos_i(11831) := b"0000000000000000_0000000000000000_0010001101110101_1100110010001001"; -- 0.13851621964041622
	pesos_i(11832) := b"0000000000000000_0000000000000000_0000001010110000_0111101110101000"; -- 0.010505417413267618
	pesos_i(11833) := b"0000000000000000_0000000000000000_0001100010001101_0110110110101100"; -- 0.0959080261307584
	pesos_i(11834) := b"1111111111111111_1111111111111111_1111010110010101_0110111011011110"; -- -0.04068858225733928
	pesos_i(11835) := b"0000000000000000_0000000000000000_0000111000011111_1101111111010100"; -- 0.05517386368520433
	pesos_i(11836) := b"1111111111111111_1111111111111111_1110110000001101_1000011100000011"; -- -0.07791858851385047
	pesos_i(11837) := b"0000000000000000_0000000000000000_0001010101111000_0010001000100001"; -- 0.08386433889730886
	pesos_i(11838) := b"1111111111111111_1111111111111111_1111110111011101_0011110001011001"; -- -0.008342960702130432
	pesos_i(11839) := b"0000000000000000_0000000000000000_0001110010011001_0011000010100100"; -- 0.11171249385577768
	pesos_i(11840) := b"1111111111111111_1111111111111111_1101110111010010_0110001000111110"; -- -0.13350854870642692
	pesos_i(11841) := b"1111111111111111_1111111111111111_1101111011111101_0010010010111001"; -- -0.1289498374644245
	pesos_i(11842) := b"0000000000000000_0000000000000000_0001111011011111_0111010101101100"; -- 0.12059720884333239
	pesos_i(11843) := b"1111111111111111_1111111111111111_1101110101101010_1100110101000111"; -- -0.13508908276477322
	pesos_i(11844) := b"0000000000000000_0000000000000000_0000101111111011_0000011011010010"; -- 0.046799112649893705
	pesos_i(11845) := b"0000000000000000_0000000000000000_0000000101000101_1001111011110011"; -- 0.004968580480196299
	pesos_i(11846) := b"1111111111111111_1111111111111111_1110111001100111_1001111111001011"; -- -0.06873132021517829
	pesos_i(11847) := b"1111111111111111_1111111111111111_1110001111100110_0011011001110001"; -- -0.10976848350275731
	pesos_i(11848) := b"0000000000000000_0000000000000000_0001010100001110_0101000101011100"; -- 0.08224972233496784
	pesos_i(11849) := b"1111111111111111_1111111111111111_1110111110000100_0000100101100011"; -- -0.0643915304281885
	pesos_i(11850) := b"1111111111111111_1111111111111111_1110011110000000_0101100011101000"; -- -0.09569782588950358
	pesos_i(11851) := b"0000000000000000_0000000000000000_0000110110010100_0011111010010110"; -- 0.05304328117683625
	pesos_i(11852) := b"1111111111111111_1111111111111111_1101110111100001_0111100101100001"; -- -0.13327828773930167
	pesos_i(11853) := b"1111111111111111_1111111111111111_1110001111110011_1101000010111011"; -- -0.1095609228438589
	pesos_i(11854) := b"1111111111111111_1111111111111111_1110111000101101_0111001110101100"; -- -0.06961895999667639
	pesos_i(11855) := b"0000000000000000_0000000000000000_0001111011000101_0111101101001010"; -- 0.12020083008385203
	pesos_i(11856) := b"1111111111111111_1111111111111111_1101111010001111_1010000100001101"; -- -0.13062089376680022
	pesos_i(11857) := b"1111111111111111_1111111111111111_1110010010101000_0110010110010011"; -- -0.10680546923050728
	pesos_i(11858) := b"0000000000000000_0000000000000000_0010000110011101_1000101001111010"; -- 0.13131013373390266
	pesos_i(11859) := b"1111111111111111_1111111111111111_1111111011110110_0010111110010100"; -- -0.004056002035133828
	pesos_i(11860) := b"0000000000000000_0000000000000000_0010010110100100_0100100110011100"; -- 0.1470380788738356
	pesos_i(11861) := b"0000000000000000_0000000000000000_0000001110111110_0100111011010110"; -- 0.014622618968293458
	pesos_i(11862) := b"1111111111111111_1111111111111111_1110100111011000_1100100011001111"; -- -0.08653588240239886
	pesos_i(11863) := b"0000000000000000_0000000000000000_0000111110011000_0011010111110001"; -- 0.06091630109743974
	pesos_i(11864) := b"0000000000000000_0000000000000000_0001000111000011_0101000111001010"; -- 0.069386588781436
	pesos_i(11865) := b"1111111111111111_1111111111111111_1110011111011000_1101010011111101"; -- -0.09434765645531333
	pesos_i(11866) := b"1111111111111111_1111111111111111_1111001111010111_0001100010100011"; -- -0.047499141821998214
	pesos_i(11867) := b"0000000000000000_0000000000000000_0001110000100110_0011010111001111"; -- 0.10995804127820584
	pesos_i(11868) := b"1111111111111111_1111111111111111_1111000110000010_1101100010111010"; -- -0.05659718949430683
	pesos_i(11869) := b"1111111111111111_1111111111111111_1111100101101011_1100100100000000"; -- -0.025699079075710583
	pesos_i(11870) := b"1111111111111111_1111111111111111_1101110001001001_0000101011010110"; -- -0.1395104625029493
	pesos_i(11871) := b"1111111111111111_1111111111111111_1101111001110001_0011011001000110"; -- -0.1310850218846391
	pesos_i(11872) := b"0000000000000000_0000000000000000_0001101110011000_1000101100110110"; -- 0.10779638356933906
	pesos_i(11873) := b"1111111111111111_1111111111111111_1111001100001000_0100000000101101"; -- -0.05065535440303977
	pesos_i(11874) := b"1111111111111111_1111111111111111_1110111100001110_0110100011000100"; -- -0.06618638239095595
	pesos_i(11875) := b"1111111111111111_1111111111111111_1101111000100100_1101100000111010"; -- -0.13225029552971246
	pesos_i(11876) := b"0000000000000000_0000000000000000_0001101011000111_1111001110011101"; -- 0.10461351949009086
	pesos_i(11877) := b"1111111111111111_1111111111111111_1110100101111101_0111011010001010"; -- -0.08792933586473094
	pesos_i(11878) := b"0000000000000000_0000000000000000_0001110001001011_0110110110101011"; -- 0.11052594579096803
	pesos_i(11879) := b"1111111111111111_1111111111111111_1111001011010000_0100111100011000"; -- -0.05150895757875578
	pesos_i(11880) := b"1111111111111111_1111111111111111_1110100101101111_0101111011101100"; -- -0.08814436654889604
	pesos_i(11881) := b"1111111111111111_1111111111111111_1110111011011010_0100111110111101"; -- -0.06698133118970358
	pesos_i(11882) := b"0000000000000000_0000000000000000_0001110001110110_1000011101101000"; -- 0.11118360802956491
	pesos_i(11883) := b"1111111111111111_1111111111111111_1111011010111101_1000101110010111"; -- -0.03617026860385329
	pesos_i(11884) := b"0000000000000000_0000000000000000_0001100111001101_0101100000011011"; -- 0.10078955317409884
	pesos_i(11885) := b"1111111111111111_1111111111111111_1111110001110111_1001101101000110"; -- -0.013799949129242388
	pesos_i(11886) := b"1111111111111111_1111111111111111_1111011110000110_1001110101100111"; -- -0.0331021902582508
	pesos_i(11887) := b"0000000000000000_0000000000000000_0001100000111011_1101100011001001"; -- 0.09466318998570548
	pesos_i(11888) := b"1111111111111111_1111111111111111_1111110101010101_1111010110100110"; -- -0.010407111058328403
	pesos_i(11889) := b"1111111111111111_1111111111111111_1110110010100100_0011010100000011"; -- -0.07561939885744107
	pesos_i(11890) := b"1111111111111111_1111111111111111_1101101110111101_0110101011001100"; -- -0.1416409731789745
	pesos_i(11891) := b"0000000000000000_0000000000000000_0000100111101011_1100110101000000"; -- 0.03875429920526068
	pesos_i(11892) := b"1111111111111111_1111111111111111_1110100000010000_0101011101110110"; -- -0.09350064631345671
	pesos_i(11893) := b"0000000000000000_0000000000000000_0000111111010011_0000101010000010"; -- 0.061813980908265835
	pesos_i(11894) := b"0000000000000000_0000000000000000_0010010000110111_1001010000000000"; -- 0.14147305484042594
	pesos_i(11895) := b"1111111111111111_1111111111111111_1110100011010001_1100101111111110"; -- -0.09054875426237245
	pesos_i(11896) := b"0000000000000000_0000000000000000_0001110110100010_1101011101100100"; -- 0.11576601201970972
	pesos_i(11897) := b"0000000000000000_0000000000000000_0001101101110110_0000001101101101"; -- 0.10726949138786236
	pesos_i(11898) := b"1111111111111111_1111111111111111_1101110000010011_1101100011011000"; -- -0.1403221582100063
	pesos_i(11899) := b"0000000000000000_0000000000000000_0000001010001000_0101011000100101"; -- 0.009892829892598494
	pesos_i(11900) := b"0000000000000000_0000000000000000_0001011010110110_1100101000101100"; -- 0.08872665008158771
	pesos_i(11901) := b"1111111111111111_1111111111111111_1111111111011110_1000011100000100"; -- -0.0005107511733925365
	pesos_i(11902) := b"1111111111111111_1111111111111111_1101011000011110_0110100000111010"; -- -0.163598524028427
	pesos_i(11903) := b"0000000000000000_0000000000000000_0000111001001111_1000110011000001"; -- 0.055901333909344465
	pesos_i(11904) := b"0000000000000000_0000000000000000_0000101011001010_1000111101001001"; -- 0.042153315840160126
	pesos_i(11905) := b"0000000000000000_0000000000000000_0001110110011011_1000100001001000"; -- 0.11565448528097426
	pesos_i(11906) := b"0000000000000000_0000000000000000_0001101100001010_1111110010011110"; -- 0.10563639503245438
	pesos_i(11907) := b"1111111111111111_1111111111111111_1110101011111101_0010111101000100"; -- -0.08207420915336285
	pesos_i(11908) := b"1111111111111111_1111111111111111_1111101101010111_0101100010010101"; -- -0.018198455441979382
	pesos_i(11909) := b"0000000000000000_0000000000000000_0010011001011011_1010101000001101"; -- 0.14983618569811585
	pesos_i(11910) := b"1111111111111111_1111111111111111_1111111010110010_0001101010110001"; -- -0.005094844657017936
	pesos_i(11911) := b"0000000000000000_0000000000000000_0001011010110001_1001100011101111"; -- 0.0886474211516082
	pesos_i(11912) := b"1111111111111111_1111111111111111_1111110101110001_1100100011001100"; -- -0.009982538503334032
	pesos_i(11913) := b"1111111111111111_1111111111111111_1111110011101000_1011110110011011"; -- -0.012073659654959028
	pesos_i(11914) := b"1111111111111111_1111111111111111_1111100101110011_1010100101101100"; -- -0.02557889094073678
	pesos_i(11915) := b"0000000000000000_0000000000000000_0000001111100011_0110111100010000"; -- 0.015189114950327584
	pesos_i(11916) := b"1111111111111111_1111111111111111_1110101100111001_1001010011101010"; -- -0.08115262297871106
	pesos_i(11917) := b"0000000000000000_0000000000000000_0010001100011111_0010000110001000"; -- 0.137193771104215
	pesos_i(11918) := b"0000000000000000_0000000000000000_0000000011100101_1010111100001101"; -- 0.0035046965058318264
	pesos_i(11919) := b"0000000000000000_0000000000000000_0000000101101011_0011000011010001"; -- 0.005541850013901753
	pesos_i(11920) := b"0000000000000000_0000000000000000_0001001111111100_0110010010110000"; -- 0.07806996639475207
	pesos_i(11921) := b"1111111111111111_1111111111111111_1110110110111101_0000000000010110"; -- -0.0713348336870017
	pesos_i(11922) := b"0000000000000000_0000000000000000_0001000001110100_0011001001011100"; -- 0.06427302125831794
	pesos_i(11923) := b"1111111111111111_1111111111111111_1101110111100100_0001101110001000"; -- -0.13323810509718265
	pesos_i(11924) := b"0000000000000000_0000000000000000_0001110110111100_0111101010011011"; -- 0.11615721012762602
	pesos_i(11925) := b"0000000000000000_0000000000000000_0000100101111110_0101111101100111"; -- 0.03708454394564848
	pesos_i(11926) := b"0000000000000000_0000000000000000_0000000110011100_0110100000000110"; -- 0.006292821464178824
	pesos_i(11927) := b"1111111111111111_1111111111111111_1110000101011111_0101101001101000"; -- -0.11963877630408774
	pesos_i(11928) := b"1111111111111111_1111111111111111_1101110011111110_1011110100011001"; -- -0.13673799655862576
	pesos_i(11929) := b"1111111111111111_1111111111111111_1110010111000010_0110010000110000"; -- -0.10250257325593579
	pesos_i(11930) := b"1111111111111111_1111111111111111_1101110110000011_1000111111011100"; -- -0.13471127397018223
	pesos_i(11931) := b"0000000000000000_0000000000000000_0001001010000101_0101100001001111"; -- 0.07234718246536584
	pesos_i(11932) := b"0000000000000000_0000000000000000_0000011111100101_0100111100111010"; -- 0.03084273492929536
	pesos_i(11933) := b"1111111111111111_1111111111111111_1111110001111111_0111000110000100"; -- -0.013680367629257284
	pesos_i(11934) := b"0000000000000000_0000000000000000_0001111101111010_1010101001001101"; -- 0.12296547303234454
	pesos_i(11935) := b"1111111111111111_1111111111111111_1111001010111011_0101110111111110"; -- -0.051828503996431165
	pesos_i(11936) := b"1111111111111111_1111111111111111_1111011000001100_0001110000110100"; -- -0.03887771341712513
	pesos_i(11937) := b"0000000000000000_0000000000000000_0001001110100011_0001100101001010"; -- 0.07670744000237015
	pesos_i(11938) := b"0000000000000000_0000000000000000_0000100010000000_0000101101010001"; -- 0.033203799550773745
	pesos_i(11939) := b"0000000000000000_0000000000000000_0000001110101100_1101001010000000"; -- 0.014355808449577017
	pesos_i(11940) := b"1111111111111111_1111111111111111_1110011110011011_0000011000011011"; -- -0.095290773723647
	pesos_i(11941) := b"0000000000000000_0000000000000000_0000110111000100_1101011111111000"; -- 0.05378484545442212
	pesos_i(11942) := b"0000000000000000_0000000000000000_0001001110100010_1111001111010011"; -- 0.07670520698839421
	pesos_i(11943) := b"1111111111111111_1111111111111111_1111001000010011_1101101001110011"; -- -0.05438456250889226
	pesos_i(11944) := b"0000000000000000_0000000000000000_0000110000101000_0011010100011100"; -- 0.04748851713918192
	pesos_i(11945) := b"0000000000000000_0000000000000000_0000110010101100_0010000010111111"; -- 0.04950146351348939
	pesos_i(11946) := b"1111111111111111_1111111111111111_1110100111100011_0000111111110110"; -- -0.08637905353075352
	pesos_i(11947) := b"1111111111111111_1111111111111111_1101111000011011_1010010111001010"; -- -0.13239063084902414
	pesos_i(11948) := b"1111111111111111_1111111111111111_1110111110000011_1100011010001100"; -- -0.06439551428311074
	pesos_i(11949) := b"0000000000000000_0000000000000000_0001100001000101_1010110011011011"; -- 0.0948131594477794
	pesos_i(11950) := b"1111111111111111_1111111111111111_1110101110110101_1011101010010101"; -- -0.07925828808787821
	pesos_i(11951) := b"1111111111111111_1111111111111111_1110111101011100_1111111111111101"; -- -0.06498718335110205
	pesos_i(11952) := b"0000000000000000_0000000000000000_0001110010111100_1000100100100000"; -- 0.11225182572707591
	pesos_i(11953) := b"1111111111111111_1111111111111111_1101111011010101_1100001011110111"; -- -0.12955075722207687
	pesos_i(11954) := b"0000000000000000_0000000000000000_0000101010111010_0101101000110111"; -- 0.04190601188911791
	pesos_i(11955) := b"0000000000000000_0000000000000000_0000101101100010_1101110011010010"; -- 0.044477273308250714
	pesos_i(11956) := b"1111111111111111_1111111111111111_1110010001000011_1010001100110011"; -- -0.10834293360913602
	pesos_i(11957) := b"0000000000000000_0000000000000000_0000110110001100_0011111010000111"; -- 0.052921207274977
	pesos_i(11958) := b"0000000000000000_0000000000000000_0001001110110011_0001101010011101"; -- 0.07695165960450472
	pesos_i(11959) := b"1111111111111111_1111111111111111_1111101010010110_0010110011010000"; -- -0.02114601068155408
	pesos_i(11960) := b"0000000000000000_0000000000000000_0000011111000010_0110100100101001"; -- 0.030310223217560273
	pesos_i(11961) := b"1111111111111111_1111111111111111_1111000101111010_1101101110111011"; -- -0.05671908087648016
	pesos_i(11962) := b"1111111111111111_1111111111111111_1111110000101100_1001111110100010"; -- -0.014944098440552635
	pesos_i(11963) := b"1111111111111111_1111111111111111_1110111101001011_0010011000000110"; -- -0.06525957440129324
	pesos_i(11964) := b"0000000000000000_0000000000000000_0001110101001000_1000111110000011"; -- 0.11438843675536714
	pesos_i(11965) := b"0000000000000000_0000000000000000_0001110100010111_0010101101010111"; -- 0.11363478550005925
	pesos_i(11966) := b"1111111111111111_1111111111111111_1111010111101110_1001110101111010"; -- -0.039327771913525
	pesos_i(11967) := b"1111111111111111_1111111111111111_1111110001111011_0101001000011101"; -- -0.01374327470408459
	pesos_i(11968) := b"0000000000000000_0000000000000000_0010010100010010_1011100010110111"; -- 0.14481691812344688
	pesos_i(11969) := b"0000000000000000_0000000000000000_0001011010111011_1100010001100100"; -- 0.08880259937853059
	pesos_i(11970) := b"0000000000000000_0000000000000000_0000101001011001_1001111110010000"; -- 0.04043004283948485
	pesos_i(11971) := b"1111111111111111_1111111111111111_1111101101100010_0111000100010100"; -- -0.018029148610998337
	pesos_i(11972) := b"0000000000000000_0000000000000000_0001011110010111_1011001011110100"; -- 0.09215849351082121
	pesos_i(11973) := b"0000000000000000_0000000000000000_0010100111010010_0011101110111010"; -- 0.16336415560010617
	pesos_i(11974) := b"0000000000000000_0000000000000000_0001001100101100_0111101000111100"; -- 0.07489742235822779
	pesos_i(11975) := b"1111111111111111_1111111111111111_1111100011000110_0101101100111000"; -- -0.02822332280208114
	pesos_i(11976) := b"0000000000000000_0000000000000000_0000110101011000_1110111101111100"; -- 0.05213829789923458
	pesos_i(11977) := b"1111111111111111_1111111111111111_1110001101100100_0000111110010100"; -- -0.1117544425493505
	pesos_i(11978) := b"1111111111111111_1111111111111111_1101110001101000_1000010101101110"; -- -0.13903013279450843
	pesos_i(11979) := b"1111111111111111_1111111111111111_1101110101101011_1001101000001111"; -- -0.13507687685406872
	pesos_i(11980) := b"0000000000000000_0000000000000000_0000011110001011_1000000000111010"; -- 0.029472364475342502
	pesos_i(11981) := b"1111111111111111_1111111111111111_1111101001101011_1111101000011000"; -- -0.02178990285861716
	pesos_i(11982) := b"0000000000000000_0000000000000000_0001101001100111_1000010110011101"; -- 0.10314211931558755
	pesos_i(11983) := b"0000000000000000_0000000000000000_0000110000001101_1000001101010010"; -- 0.04708119166672736
	pesos_i(11984) := b"0000000000000000_0000000000000000_0000011011011100_1100010110101011"; -- 0.02680621562630541
	pesos_i(11985) := b"1111111111111111_1111111111111111_1110011010110000_1100011100010110"; -- -0.0988650867255593
	pesos_i(11986) := b"1111111111111111_1111111111111111_1110100111101011_1010001110101101"; -- -0.0862481786834158
	pesos_i(11987) := b"1111111111111111_1111111111111111_1110110000110010_1000011011011101"; -- -0.07735402218445218
	pesos_i(11988) := b"0000000000000000_0000000000000000_0001101111000110_0001011111100100"; -- 0.10849141412677549
	pesos_i(11989) := b"1111111111111111_1111111111111111_1111000111010011_1110110101011000"; -- -0.055359998761621315
	pesos_i(11990) := b"0000000000000000_0000000000000000_0001100100111100_1100101110010101"; -- 0.09858391168166222
	pesos_i(11991) := b"0000000000000000_0000000000000000_0001100100000001_1000100001100111"; -- 0.09767963900414471
	pesos_i(11992) := b"1111111111111111_1111111111111111_1111111000010000_0100101100100111"; -- -0.007563879877347089
	pesos_i(11993) := b"0000000000000000_0000000000000000_0000100011000101_0010100101101000"; -- 0.03425844937229752
	pesos_i(11994) := b"1111111111111111_1111111111111111_1111010100110011_1001001101110001"; -- -0.04218176364426955
	pesos_i(11995) := b"1111111111111111_1111111111111111_1111111010001001_0011000111111000"; -- -0.005719067512948261
	pesos_i(11996) := b"0000000000000000_0000000000000000_0010001110001000_0100110100110100"; -- 0.13879854699279542
	pesos_i(11997) := b"1111111111111111_1111111111111111_1111001010110010_1001000010111000"; -- -0.051962809562189446
	pesos_i(11998) := b"0000000000000000_0000000000000000_0001111101110100_0000111001110000"; -- 0.12286463004406689
	pesos_i(11999) := b"1111111111111111_1111111111111111_1111011000001111_1001111010110011"; -- -0.03882415889954175
	pesos_i(12000) := b"1111111111111111_1111111111111111_1111110000110011_1011101001011000"; -- -0.014835694908201729
	pesos_i(12001) := b"1111111111111111_1111111111111111_1101100000101110_1110010101100101"; -- -0.15553442261347075
	pesos_i(12002) := b"0000000000000000_0000000000000000_0010011101000111_1100101111111111"; -- 0.1534392832502685
	pesos_i(12003) := b"1111111111111111_1111111111111111_1110111000110011_0011100100100010"; -- -0.06953089642548918
	pesos_i(12004) := b"1111111111111111_1111111111111111_1110010000000100_0100111010010010"; -- -0.1093092816589073
	pesos_i(12005) := b"0000000000000000_0000000000000000_0000011010011000_0111100010000010"; -- 0.025764018765304913
	pesos_i(12006) := b"0000000000000000_0000000000000000_0001111101100011_1010110001011101"; -- 0.12261464367227719
	pesos_i(12007) := b"0000000000000000_0000000000000000_0001110000011011_1001110000010110"; -- 0.10979629084798875
	pesos_i(12008) := b"1111111111111111_1111111111111111_1110000000110100_1111011101101100"; -- -0.12419179539796393
	pesos_i(12009) := b"1111111111111111_1111111111111111_1110000011001111_0001111101101010"; -- -0.12183955826307473
	pesos_i(12010) := b"1111111111111111_1111111111111111_1110100000000000_1001110101011110"; -- -0.09374062028521857
	pesos_i(12011) := b"1111111111111111_1111111111111111_1110001110110000_0100011011110111"; -- -0.11059147325850271
	pesos_i(12012) := b"0000000000000000_0000000000000000_0001011010111011_1110011001101011"; -- 0.08880462748571527
	pesos_i(12013) := b"1111111111111111_1111111111111111_1111101011010111_1111001011010011"; -- -0.020142386822158933
	pesos_i(12014) := b"1111111111111111_1111111111111111_1110101101110001_0111001000000001"; -- -0.08030021164436535
	pesos_i(12015) := b"1111111111111111_1111111111111111_1111110011101001_0010000111111011"; -- -0.012067676639505257
	pesos_i(12016) := b"1111111111111111_1111111111111111_1110101010001001_0001000110000101"; -- -0.08384600158437418
	pesos_i(12017) := b"1111111111111111_1111111111111111_1101101011100111_1100011101110100"; -- -0.1449008313702073
	pesos_i(12018) := b"0000000000000000_0000000000000000_0010010001111100_1000100011100101"; -- 0.14252524942569916
	pesos_i(12019) := b"0000000000000000_0000000000000000_0010000100011000_1011101101111011"; -- 0.12928363570583595
	pesos_i(12020) := b"1111111111111111_1111111111111111_1110001100111101_1110110011001111"; -- -0.11233634900092664
	pesos_i(12021) := b"0000000000000000_0000000000000000_0010011001011000_0111101101111011"; -- 0.14978763342913262
	pesos_i(12022) := b"1111111111111111_1111111111111111_1111001101000010_1000000001101011"; -- -0.049766515663245456
	pesos_i(12023) := b"0000000000000000_0000000000000000_0010001110100100_0111111110011100"; -- 0.13922879754068163
	pesos_i(12024) := b"1111111111111111_1111111111111111_1111101010001111_1100001010111001"; -- -0.021243886805241318
	pesos_i(12025) := b"1111111111111111_1111111111111111_1110010000110110_1100010101011100"; -- -0.10853926187450925
	pesos_i(12026) := b"1111111111111111_1111111111111111_1110001111010111_1100110001101101"; -- -0.10998842551466713
	pesos_i(12027) := b"0000000000000000_0000000000000000_0001101101111010_0101110010001111"; -- 0.10733583912810299
	pesos_i(12028) := b"1111111111111111_1111111111111111_1111000110101011_1111101000101101"; -- -0.055969585454267466
	pesos_i(12029) := b"0000000000000000_0000000000000000_0001001100110001_1000010101001101"; -- 0.07497437610197548
	pesos_i(12030) := b"0000000000000000_0000000000000000_0010000110011110_1010101101000000"; -- 0.13132734599650514
	pesos_i(12031) := b"1111111111111111_1111111111111111_1111000101001101_0010000100000110"; -- -0.057416854987628975
	pesos_i(12032) := b"1111111111111111_1111111111111111_1110000011000001_1110010010001111"; -- -0.122041430658916
	pesos_i(12033) := b"1111111111111111_1111111111111111_1101101000110111_1000110000100111"; -- -0.14758991278263273
	pesos_i(12034) := b"0000000000000000_0000000000000000_0000101111001000_0111110001010111"; -- 0.046027918994807106
	pesos_i(12035) := b"1111111111111111_1111111111111111_1110101011011100_1010010001110100"; -- -0.08257076429936897
	pesos_i(12036) := b"1111111111111111_1111111111111111_1110001111001101_1101110010011000"; -- -0.11014004981082047
	pesos_i(12037) := b"0000000000000000_0000000000000000_0001011100011101_0111101001001010"; -- 0.09029354386494022
	pesos_i(12038) := b"0000000000000000_0000000000000000_0001111111101000_1000011010000001"; -- 0.12464180621382089
	pesos_i(12039) := b"1111111111111111_1111111111111111_1111111101100101_1000010011000111"; -- -0.0023571981676787164
	pesos_i(12040) := b"1111111111111111_1111111111111111_1110100011110001_0000000100111000"; -- -0.09007255918128333
	pesos_i(12041) := b"0000000000000000_0000000000000000_0010000000111011_1001011100100110"; -- 0.12590927770703744
	pesos_i(12042) := b"1111111111111111_1111111111111111_1111011110111110_1100110000111000"; -- -0.03224490767242839
	pesos_i(12043) := b"1111111111111111_1111111111111111_1110100101001010_1011111010001101"; -- -0.08870324195904605
	pesos_i(12044) := b"1111111111111111_1111111111111111_1111001001111010_0101111111110100"; -- -0.0528202084043728
	pesos_i(12045) := b"1111111111111111_1111111111111111_1110101110000011_1100101001001001"; -- -0.08002029152271688
	pesos_i(12046) := b"0000000000000000_0000000000000000_0000010110011011_0111110100001101"; -- 0.02190381584642405
	pesos_i(12047) := b"1111111111111111_1111111111111111_1110011111010110_0110001101010011"; -- -0.094384948959624
	pesos_i(12048) := b"0000000000000000_0000000000000000_0000001110110110_0000000001010001"; -- 0.014495868547687158
	pesos_i(12049) := b"1111111111111111_1111111111111111_1111101001001000_0100000110000001"; -- -0.022334962920279033
	pesos_i(12050) := b"0000000000000000_0000000000000000_0000111110011100_0010000001000111"; -- 0.060976045012860094
	pesos_i(12051) := b"1111111111111111_1111111111111111_1111001111101010_0011101011111100"; -- -0.047207177714646026
	pesos_i(12052) := b"1111111111111111_1111111111111111_1111100110001100_1011010111110101"; -- -0.02519667407779944
	pesos_i(12053) := b"0000000000000000_0000000000000000_0010000101100111_1000000001001110"; -- 0.1304855527848565
	pesos_i(12054) := b"1111111111111111_1111111111111111_1110100111010000_1101010110010001"; -- -0.08665719241990558
	pesos_i(12055) := b"0000000000000000_0000000000000000_0000000101100000_1100001010101000"; -- 0.0053826960552669015
	pesos_i(12056) := b"0000000000000000_0000000000000000_0001110001100011_0101010000001010"; -- 0.11089062916140825
	pesos_i(12057) := b"0000000000000000_0000000000000000_0000110010010010_0000011010011100"; -- 0.049103177089253436
	pesos_i(12058) := b"1111111111111111_1111111111111111_1111110010100101_1110110111111011"; -- -0.013093115093581076
	pesos_i(12059) := b"0000000000000000_0000000000000000_0001011111100111_1100100001100010"; -- 0.09338047406620636
	pesos_i(12060) := b"0000000000000000_0000000000000000_0001000111000111_0100100000010001"; -- 0.06944704449733223
	pesos_i(12061) := b"0000000000000000_0000000000000000_0001101011001100_1101011101001010"; -- 0.10468812512284621
	pesos_i(12062) := b"1111111111111111_1111111111111111_1111000000101011_0011110000100101"; -- -0.06184028715194447
	pesos_i(12063) := b"0000000000000000_0000000000000000_0001010000101111_0111000000100001"; -- 0.07884884651803672
	pesos_i(12064) := b"0000000000000000_0000000000000000_0000011011100110_0010101010010011"; -- 0.026949559119185937
	pesos_i(12065) := b"1111111111111111_1111111111111111_1110100010010110_1001110110110111"; -- -0.09145178112449479
	pesos_i(12066) := b"1111111111111111_1111111111111111_1110100111100110_1110000110100001"; -- -0.08632078007773104
	pesos_i(12067) := b"0000000000000000_0000000000000000_0000010101111011_0100001110110101"; -- 0.021412116690409773
	pesos_i(12068) := b"0000000000000000_0000000000000000_0010000111000110_0010001101100111"; -- 0.13192960036557916
	pesos_i(12069) := b"1111111111111111_1111111111111111_1111100010110010_0101110000111001"; -- -0.028528438738019118
	pesos_i(12070) := b"1111111111111111_1111111111111111_1111110001000111_0110100101000001"; -- -0.01453535227121171
	pesos_i(12071) := b"0000000000000000_0000000000000000_0001111000111001_1000100110100111"; -- 0.11806545559106646
	pesos_i(12072) := b"1111111111111111_1111111111111111_1111000111001101_1000011000010101"; -- -0.05545770633249703
	pesos_i(12073) := b"0000000000000000_0000000000000000_0001011010001101_1100110100010111"; -- 0.0881012134658477
	pesos_i(12074) := b"0000000000000000_0000000000000000_0000110010011101_0010101100010001"; -- 0.04927319695518983
	pesos_i(12075) := b"0000000000000000_0000000000000000_0000111100110110_0011101001000000"; -- 0.05942119666945424
	pesos_i(12076) := b"0000000000000000_0000000000000000_0010000001110001_0100110011000001"; -- 0.12672881796786656
	pesos_i(12077) := b"1111111111111111_1111111111111111_1110111001000110_1001100100101000"; -- -0.06923525601619651
	pesos_i(12078) := b"0000000000000000_0000000000000000_0000011001111000_0110010000111000"; -- 0.02527452813426921
	pesos_i(12079) := b"1111111111111111_1111111111111111_1110010111000110_0010000011100111"; -- -0.1024455485712222
	pesos_i(12080) := b"0000000000000000_0000000000000000_0001101000110001_1001011100001100"; -- 0.10231918365885087
	pesos_i(12081) := b"0000000000000000_0000000000000000_0010001110110001_1101011111011011"; -- 0.13943242156792385
	pesos_i(12082) := b"1111111111111111_1111111111111111_1111010001110110_0010101110011110"; -- -0.045071863037298154
	pesos_i(12083) := b"0000000000000000_0000000000000000_0001110111100001_0000011000010001"; -- 0.11671483919934514
	pesos_i(12084) := b"1111111111111111_1111111111111111_1111011110100010_0010010011101011"; -- -0.03268212562834995
	pesos_i(12085) := b"1111111111111111_1111111111111111_1111101111100010_0000001100000011"; -- -0.016082584270097105
	pesos_i(12086) := b"1111111111111111_1111111111111111_1111001100011111_0000110011000100"; -- -0.05030746674059636
	pesos_i(12087) := b"1111111111111111_1111111111111111_1101100001010011_0111010000010011"; -- -0.15497660190469714
	pesos_i(12088) := b"1111111111111111_1111111111111111_1110001000111010_0101101100110101"; -- -0.11629705389861016
	pesos_i(12089) := b"1111111111111111_1111111111111111_1110001100100101_0101010111110010"; -- -0.11271155214188441
	pesos_i(12090) := b"0000000000000000_0000000000000000_0010001100000100_0000000111010110"; -- 0.13677989449394545
	pesos_i(12091) := b"0000000000000000_0000000000000000_0010000101011111_1110111111000011"; -- 0.13037012580402585
	pesos_i(12092) := b"1111111111111111_1111111111111111_1111111010110011_0110011010110011"; -- -0.005075055386859549
	pesos_i(12093) := b"0000000000000000_0000000000000000_0000110000100100_0111100111110111"; -- 0.04743158596727282
	pesos_i(12094) := b"0000000000000000_0000000000000000_0010011011011110_1110101000010111"; -- 0.15183890400550387
	pesos_i(12095) := b"0000000000000000_0000000000000000_0001101110000111_0001000001010001"; -- 0.10752965894615726
	pesos_i(12096) := b"1111111111111111_1111111111111111_1110011111011001_0001000111110011"; -- -0.09434402282890116
	pesos_i(12097) := b"0000000000000000_0000000000000000_0000110011001010_1011000100001101"; -- 0.049967828543916376
	pesos_i(12098) := b"1111111111111111_1111111111111111_1111110011011001_1111001011010111"; -- -0.012299368467566477
	pesos_i(12099) := b"0000000000000000_0000000000000000_0001000110101010_0110011111000110"; -- 0.06900642956794424
	pesos_i(12100) := b"1111111111111111_1111111111111111_1111111101000110_1110001000001100"; -- -0.002824661381396703
	pesos_i(12101) := b"0000000000000000_0000000000000000_0000100010111010_1111010101111010"; -- 0.034102766355131216
	pesos_i(12102) := b"0000000000000000_0000000000000000_0010010101011110_1100111010100111"; -- 0.14597789372730136
	pesos_i(12103) := b"1111111111111111_1111111111111111_1111000101000011_0110110101110000"; -- -0.057564888099608816
	pesos_i(12104) := b"1111111111111111_1111111111111111_1111111001010001_1101011101100001"; -- -0.006563700404501745
	pesos_i(12105) := b"1111111111111111_1111111111111111_1110000001110110_0111100111001101"; -- -0.12319220300140771
	pesos_i(12106) := b"0000000000000000_0000000000000000_0001010011101010_0001101010001101"; -- 0.08169713928506425
	pesos_i(12107) := b"1111111111111111_1111111111111111_1111110000101110_1010100000111111"; -- -0.014913067346990437
	pesos_i(12108) := b"1111111111111111_1111111111111111_1111000011000100_0111100010011101"; -- -0.05950208832152209
	pesos_i(12109) := b"1111111111111111_1111111111111111_1110110100000100_1111111111101101"; -- -0.07414246046948095
	pesos_i(12110) := b"0000000000000000_0000000000000000_0010001101110000_1000111100011010"; -- 0.13843626383483934
	pesos_i(12111) := b"1111111111111111_1111111111111111_1110110110101010_0111001000001011"; -- -0.07161795835869705
	pesos_i(12112) := b"1111111111111111_1111111111111111_1110001011101100_1001110000100001"; -- -0.11357711974323369
	pesos_i(12113) := b"0000000000000000_0000000000000000_0000110101010101_0010110000110110"; -- 0.05208088222512167
	pesos_i(12114) := b"1111111111111111_1111111111111111_1101011111010100_1101010111011010"; -- -0.1569086401503176
	pesos_i(12115) := b"1111111111111111_1111111111111111_1110010001000110_1010100001100101"; -- -0.10829684761555201
	pesos_i(12116) := b"1111111111111111_1111111111111111_1110100011010110_1001010100111010"; -- -0.09047572451749696
	pesos_i(12117) := b"1111111111111111_1111111111111111_1110011100111001_0000010100110101"; -- -0.09678618876745525
	pesos_i(12118) := b"1111111111111111_1111111111111111_1110010010011000_1111111100110011"; -- -0.10704045289589378
	pesos_i(12119) := b"0000000000000000_0000000000000000_0000001101110001_1000110011001111"; -- 0.013451386073491901
	pesos_i(12120) := b"1111111111111111_1111111111111111_1110111010011110_1110001001111001"; -- -0.06788811242241365
	pesos_i(12121) := b"1111111111111111_1111111111111111_1111001011001101_0010101000011110"; -- -0.051556937833538895
	pesos_i(12122) := b"0000000000000000_0000000000000000_0010010001100011_0100011111101110"; -- 0.14213990740287274
	pesos_i(12123) := b"0000000000000000_0000000000000000_0001001011001110_1100101011011011"; -- 0.0734679017045678
	pesos_i(12124) := b"0000000000000000_0000000000000000_0010010001111101_1100010110110101"; -- 0.1425441329592432
	pesos_i(12125) := b"1111111111111111_1111111111111111_1110110011010111_0000010111010001"; -- -0.07484401376480396
	pesos_i(12126) := b"1111111111111111_1111111111111111_1101111100100010_1110110010000001"; -- -0.1283733543498445
	pesos_i(12127) := b"0000000000000000_0000000000000000_0000010001111111_0111111001011001"; -- 0.01757039701777303
	pesos_i(12128) := b"0000000000000000_0000000000000000_0001110100010010_0000001011011000"; -- 0.11355607767347745
	pesos_i(12129) := b"0000000000000000_0000000000000000_0000001000000110_1011011101010110"; -- 0.007914980499410727
	pesos_i(12130) := b"1111111111111111_1111111111111111_1101110101111001_1001111011110110"; -- -0.13486296169884823
	pesos_i(12131) := b"1111111111111111_1111111111111111_1111100010101000_0011111001111110"; -- -0.028682798517529202
	pesos_i(12132) := b"1111111111111111_1111111111111111_1101101111100110_0111001101011110"; -- -0.14101485217690465
	pesos_i(12133) := b"0000000000000000_0000000000000000_0010011001000001_1000001100011010"; -- 0.14943713549604346
	pesos_i(12134) := b"1111111111111111_1111111111111111_1111100111101000_1111000011101000"; -- -0.023789351715649436
	pesos_i(12135) := b"1111111111111111_1111111111111111_1110001010110011_0100001111001010"; -- -0.11445213615051254
	pesos_i(12136) := b"1111111111111111_1111111111111111_1111100101011010_1010000011001011"; -- -0.025960875006913967
	pesos_i(12137) := b"1111111111111111_1111111111111111_1101110111110010_1001101010100001"; -- -0.13301690653996998
	pesos_i(12138) := b"1111111111111111_1111111111111111_1111110010111101_0001111101001100"; -- -0.012739223483213429
	pesos_i(12139) := b"1111111111111111_1111111111111111_1101101110111101_0001111110011101"; -- -0.1416454544895617
	pesos_i(12140) := b"0000000000000000_0000000000000000_0010001100001110_0100100000000110"; -- 0.13693666598795468
	pesos_i(12141) := b"1111111111111111_1111111111111111_1111110100111111_1000110100110101"; -- -0.0107490295854267
	pesos_i(12142) := b"1111111111111111_1111111111111111_1111101010111110_0101001110110111"; -- -0.02053334037569937
	pesos_i(12143) := b"0000000000000000_0000000000000000_0001100111000000_0111000010011000"; -- 0.10059264861629733
	pesos_i(12144) := b"0000000000000000_0000000000000000_0001001000010111_1100111001001111"; -- 0.07067574902334364
	pesos_i(12145) := b"1111111111111111_1111111111111111_1110110001000010_0111011100011101"; -- -0.0771108202878334
	pesos_i(12146) := b"0000000000000000_0000000000000000_0001101010100101_1110000010010011"; -- 0.10409358581867148
	pesos_i(12147) := b"0000000000000000_0000000000000000_0000101101110010_0001001111111100"; -- 0.04470944321563344
	pesos_i(12148) := b"1111111111111111_1111111111111111_1111011011100010_0100100111001010"; -- -0.03560961560439936
	pesos_i(12149) := b"1111111111111111_1111111111111111_1110111001011110_1111100110101010"; -- -0.0688632927768528
	pesos_i(12150) := b"0000000000000000_0000000000000000_0001011011100100_1101001011010110"; -- 0.0894290706057362
	pesos_i(12151) := b"1111111111111111_1111111111111111_1111101100110011_0100010001101111"; -- -0.01874897287424835
	pesos_i(12152) := b"0000000000000000_0000000000000000_0001010100101000_1000011011010111"; -- 0.08264963864445442
	pesos_i(12153) := b"0000000000000000_0000000000000000_0000001111100010_0110001111111001"; -- 0.015173195269527697
	pesos_i(12154) := b"0000000000000000_0000000000000000_0001001110011101_0111001101101011"; -- 0.07662125940823282
	pesos_i(12155) := b"1111111111111111_1111111111111111_1111010100000100_1010000000101001"; -- -0.04289816844293702
	pesos_i(12156) := b"1111111111111111_1111111111111111_1111110001110010_0111100000101111"; -- -0.01387833455224079
	pesos_i(12157) := b"0000000000000000_0000000000000000_0000011011111000_0100100101010100"; -- 0.027226050411207375
	pesos_i(12158) := b"1111111111111111_1111111111111111_1101101110100100_1011011001101101"; -- -0.14201793509873323
	pesos_i(12159) := b"0000000000000000_0000000000000000_0000010001101111_0100011001011000"; -- 0.01732291831098939
	pesos_i(12160) := b"1111111111111111_1111111111111111_1111100100000111_1011011101001110"; -- -0.027226012693538797
	pesos_i(12161) := b"1111111111111111_1111111111111111_1111001010001111_0010101010111010"; -- -0.052502946433691015
	pesos_i(12162) := b"1111111111111111_1111111111111111_1111101110000011_1100101100010000"; -- -0.017520245077104996
	pesos_i(12163) := b"0000000000000000_0000000000000000_0010011010111111_1100011001111010"; -- 0.15136375877239683
	pesos_i(12164) := b"1111111111111111_1111111111111111_1111000110110101_0011010110011000"; -- -0.055828714761527856
	pesos_i(12165) := b"1111111111111111_1111111111111111_1111010100011111_1111110000001011"; -- -0.04248070450361889
	pesos_i(12166) := b"0000000000000000_0000000000000000_0000110111000001_0111001010100000"; -- 0.05373302839118235
	pesos_i(12167) := b"1111111111111111_1111111111111111_1110000000110001_0100100100011010"; -- -0.12424796208216113
	pesos_i(12168) := b"1111111111111111_1111111111111111_1110000000110111_0011100011100000"; -- -0.12415737666207362
	pesos_i(12169) := b"1111111111111111_1111111111111111_1101110110111001_0011000010110101"; -- -0.1338929708318978
	pesos_i(12170) := b"0000000000000000_0000000000000000_0000101001110010_1000011110101001"; -- 0.040810087987176044
	pesos_i(12171) := b"0000000000000000_0000000000000000_0000101001110010_0001000111011010"; -- 0.04080306605421607
	pesos_i(12172) := b"0000000000000000_0000000000000000_0001000010010001_0001100111011101"; -- 0.06471406592131616
	pesos_i(12173) := b"0000000000000000_0000000000000000_0001111110011100_0000100000100110"; -- 0.12347460674697629
	pesos_i(12174) := b"1111111111111111_1111111111111111_1110101001110110_0100101010100001"; -- -0.08413251462549157
	pesos_i(12175) := b"0000000000000000_0000000000000000_0000101111101000_1000110000010011"; -- 0.04651713823205607
	pesos_i(12176) := b"0000000000000000_0000000000000000_0001011100110100_0011001111001100"; -- 0.09064029445653218
	pesos_i(12177) := b"1111111111111111_1111111111111111_1110100010001111_0010011001101011"; -- -0.09156570328071485
	pesos_i(12178) := b"1111111111111111_1111111111111111_1111101000011101_1101110000111111"; -- -0.02298186732185404
	pesos_i(12179) := b"0000000000000000_0000000000000000_0000011000010011_1011001101100001"; -- 0.02373810889459902
	pesos_i(12180) := b"0000000000000000_0000000000000000_0000010011010101_1000101001000010"; -- 0.018883362879624922
	pesos_i(12181) := b"1111111111111111_1111111111111111_1111011111100101_0101000100101101"; -- -0.0316571488166971
	pesos_i(12182) := b"1111111111111111_1111111111111111_1111101111100000_1100001001101111"; -- -0.016101692199168002
	pesos_i(12183) := b"0000000000000000_0000000000000000_0000001001110000_0110010101100111"; -- 0.009527528509115925
	pesos_i(12184) := b"0000000000000000_0000000000000000_0000100000101010_0100110111111010"; -- 0.03189551685694549
	pesos_i(12185) := b"0000000000000000_0000000000000000_0000111000011001_0100100110000011"; -- 0.05507335130432705
	pesos_i(12186) := b"0000000000000000_0000000000000000_0000111111001101_1110110010111110"; -- 0.06173591263308116
	pesos_i(12187) := b"1111111111111111_1111111111111111_1101110111111000_0001101010001001"; -- -0.13293298877550166
	pesos_i(12188) := b"1111111111111111_1111111111111111_1110000011110011_1111111001001010"; -- -0.12127695733670692
	pesos_i(12189) := b"0000000000000000_0000000000000000_0001011001010011_0010111000010001"; -- 0.08720672519278962
	pesos_i(12190) := b"0000000000000000_0000000000000000_0000010001011010_1011101101001110"; -- 0.017009455181140287
	pesos_i(12191) := b"0000000000000000_0000000000000000_0000010111001110_0111101001011111"; -- 0.02268185454733832
	pesos_i(12192) := b"1111111111111111_1111111111111111_1111000010010011_1101010110111011"; -- -0.06024421861574093
	pesos_i(12193) := b"1111111111111111_1111111111111111_1110110100111010_0100100001110011"; -- -0.0733294219393511
	pesos_i(12194) := b"1111111111111111_1111111111111111_1111000000000110_0000001011100011"; -- -0.062408275232296966
	pesos_i(12195) := b"0000000000000000_0000000000000000_0010000101111011_0011111111000110"; -- 0.13078688213240078
	pesos_i(12196) := b"1111111111111111_1111111111111111_1111000010100101_0111110101011100"; -- -0.05997482771547044
	pesos_i(12197) := b"1111111111111111_1111111111111111_1101110100001010_0010100110111000"; -- -0.13656367538428593
	pesos_i(12198) := b"0000000000000000_0000000000000000_0010010111101000_1011111110010111"; -- 0.1480827088227732
	pesos_i(12199) := b"0000000000000000_0000000000000000_0010001001010110_0110110011110110"; -- 0.13413125038786838
	pesos_i(12200) := b"1111111111111111_1111111111111111_1111110010010001_0100100001110100"; -- -0.013408157047759463
	pesos_i(12201) := b"0000000000000000_0000000000000000_0010010011001001_0001110110110011"; -- 0.14369378688256657
	pesos_i(12202) := b"0000000000000000_0000000000000000_0001000101100100_0101100110100111"; -- 0.06793747257571522
	pesos_i(12203) := b"1111111111111111_1111111111111111_1101100111001011_0100110001101100"; -- -0.14924166080932375
	pesos_i(12204) := b"1111111111111111_1111111111111111_1111111001010010_1111001101100000"; -- -0.006546772952528644
	pesos_i(12205) := b"0000000000000000_0000000000000000_0001110010000000_1001110100000110"; -- 0.11133748425370953
	pesos_i(12206) := b"1111111111111111_1111111111111111_1111000100111111_0001111111010110"; -- -0.05763054874331687
	pesos_i(12207) := b"1111111111111111_1111111111111111_1101110011101000_1001110110001001"; -- -0.13707557104696388
	pesos_i(12208) := b"1111111111111111_1111111111111111_1110001110100100_1000110011101000"; -- -0.1107704098215532
	pesos_i(12209) := b"1111111111111111_1111111111111111_1110111001111011_0111000100010001"; -- -0.06842892965446183
	pesos_i(12210) := b"1111111111111111_1111111111111111_1111111001011110_0101001110011010"; -- -0.0063731908113459695
	pesos_i(12211) := b"0000000000000000_0000000000000000_0001101110101111_1011000111001010"; -- 0.10814963513794237
	pesos_i(12212) := b"0000000000000000_0000000000000000_0000011110101001_1000111001010000"; -- 0.029930967788325873
	pesos_i(12213) := b"1111111111111111_1111111111111111_1111110111001110_1101111000010000"; -- -0.008562203464368751
	pesos_i(12214) := b"1111111111111111_1111111111111111_1111101101111011_1111100001001000"; -- -0.017639620208298595
	pesos_i(12215) := b"0000000000000000_0000000000000000_0000100100101100_0001010110010001"; -- 0.035828922155436524
	pesos_i(12216) := b"1111111111111111_1111111111111111_1111001100110100_0111001101010000"; -- -0.04998091974081276
	pesos_i(12217) := b"0000000000000000_0000000000000000_0001101000101001_0001111111111000"; -- 0.10219001592073315
	pesos_i(12218) := b"1111111111111111_1111111111111111_1110001100000101_0111100100110010"; -- -0.11319773227750114
	pesos_i(12219) := b"1111111111111111_1111111111111111_1111010011010101_1101110111010111"; -- -0.04361165518394148
	pesos_i(12220) := b"1111111111111111_1111111111111111_1111101010100011_0011110111000100"; -- -0.020946635980187776
	pesos_i(12221) := b"1111111111111111_1111111111111111_1111100101010110_0101110111010000"; -- -0.02602590252084646
	pesos_i(12222) := b"0000000000000000_0000000000000000_0010001101011101_1001111111110001"; -- 0.13814735073375128
	pesos_i(12223) := b"0000000000000000_0000000000000000_0000011111111111_1101110100111111"; -- 0.03124792840109534
	pesos_i(12224) := b"1111111111111111_1111111111111111_1110011110101010_1001111100100010"; -- -0.09505277074989177
	pesos_i(12225) := b"1111111111111111_1111111111111111_1101110010000100_0000010011101011"; -- -0.13861054675404802
	pesos_i(12226) := b"0000000000000000_0000000000000000_0001010111011101_0100011100010110"; -- 0.08540767939246768
	pesos_i(12227) := b"0000000000000000_0000000000000000_0001011011111001_1101110010011111"; -- 0.08975008856959313
	pesos_i(12228) := b"0000000000000000_0000000000000000_0001000011101000_1001101111001111"; -- 0.06604932609099493
	pesos_i(12229) := b"0000000000000000_0000000000000000_0000010110000011_0100001000100000"; -- 0.021534092688857583
	pesos_i(12230) := b"0000000000000000_0000000000000000_0010001001000100_0111110011111110"; -- 0.1338575477733071
	pesos_i(12231) := b"1111111111111111_1111111111111111_1111010100001010_1000101000000100"; -- -0.04280793564937506
	pesos_i(12232) := b"0000000000000000_0000000000000000_0001101011111110_1011010110101011"; -- 0.10544906074240598
	pesos_i(12233) := b"1111111111111111_1111111111111111_1110010001000110_1001101111100011"; -- -0.10829759312334952
	pesos_i(12234) := b"0000000000000000_0000000000000000_0000001010111000_1011101000111011"; -- 0.010631217322767625
	pesos_i(12235) := b"0000000000000000_0000000000000000_0010000101100001_0000011110111000"; -- 0.13038681267871935
	pesos_i(12236) := b"0000000000000000_0000000000000000_0001000001011111_1111101000110101"; -- 0.06396449840470281
	pesos_i(12237) := b"0000000000000000_0000000000000000_0001010000010011_0111011001000000"; -- 0.07842196528049339
	pesos_i(12238) := b"1111111111111111_1111111111111111_1111101011010010_1010111110011101"; -- -0.02022268691583633
	pesos_i(12239) := b"0000000000000000_0000000000000000_0000010010110010_1101001000101010"; -- 0.018353591179833317
	pesos_i(12240) := b"1111111111111111_1111111111111111_1110000100101001_0100101011101011"; -- -0.12046367427549456
	pesos_i(12241) := b"0000000000000000_0000000000000000_0000100100011110_0010000100101001"; -- 0.03561599021076017
	pesos_i(12242) := b"0000000000000000_0000000000000000_0001000101100100_0001111010110010"; -- 0.0679339585589529
	pesos_i(12243) := b"0000000000000000_0000000000000000_0000001011101101_0010000101101011"; -- 0.0114308247674996
	pesos_i(12244) := b"1111111111111111_1111111111111111_1111101100110011_1010100101101101"; -- -0.018742953182744607
	pesos_i(12245) := b"1111111111111111_1111111111111111_1110001110011101_1110000010111000"; -- -0.11087222585645595
	pesos_i(12246) := b"0000000000000000_0000000000000000_0000110111101111_1100001000011101"; -- 0.054439670705096393
	pesos_i(12247) := b"1111111111111111_1111111111111111_1110010001000011_1010011011101111"; -- -0.10834271114685728
	pesos_i(12248) := b"1111111111111111_1111111111111111_1101101101111000_1011010000001011"; -- -0.1426894638168547
	pesos_i(12249) := b"1111111111111111_1111111111111111_1111101011000011_0101011000110111"; -- -0.020456897246759177
	pesos_i(12250) := b"0000000000000000_0000000000000000_0000111111001010_1111101010100111"; -- 0.061690965414459724
	pesos_i(12251) := b"1111111111111111_1111111111111111_1111110110100000_0111000010111010"; -- -0.00927062480301349
	pesos_i(12252) := b"1111111111111111_1111111111111111_1110100110010111_1100110100101110"; -- -0.08752744323739912
	pesos_i(12253) := b"1111111111111111_1111111111111111_1110111100000110_0110011010010010"; -- -0.06630858355675068
	pesos_i(12254) := b"0000000000000000_0000000000000000_0000011010110001_1000100100110001"; -- 0.026146482845821294
	pesos_i(12255) := b"1111111111111111_1111111111111111_1111100110010001_1000000110110010"; -- -0.02512349512664853
	pesos_i(12256) := b"1111111111111111_1111111111111111_1111010001110111_0010100010100010"; -- -0.04505678214379859
	pesos_i(12257) := b"0000000000000000_0000000000000000_0000111111101010_1011110000101100"; -- 0.062175522667945925
	pesos_i(12258) := b"0000000000000000_0000000000000000_0000011001000011_0101111010000010"; -- 0.02446547206054522
	pesos_i(12259) := b"0000000000000000_0000000000000000_0001010001001001_1011001000101110"; -- 0.07924951202948724
	pesos_i(12260) := b"1111111111111111_1111111111111111_1110111101101001_0011011001110001"; -- -0.06480083218249519
	pesos_i(12261) := b"1111111111111111_1111111111111111_1110010010010110_0001010011101110"; -- -0.10708493421940894
	pesos_i(12262) := b"1111111111111111_1111111111111111_1110111001100100_1001000000100011"; -- -0.06877802976064734
	pesos_i(12263) := b"0000000000000000_0000000000000000_0000101000010110_0100110010011010"; -- 0.03940275918644908
	pesos_i(12264) := b"1111111111111111_1111111111111111_1101111101011001_1111111001010110"; -- -0.12753305823503927
	pesos_i(12265) := b"1111111111111111_1111111111111111_1111101101011101_1010110100100001"; -- -0.01810186342516411
	pesos_i(12266) := b"1111111111111111_1111111111111111_1111000110010010_1001101110001000"; -- -0.05635669650475051
	pesos_i(12267) := b"1111111111111111_1111111111111111_1111110011111010_1011011100110001"; -- -0.01179938355953927
	pesos_i(12268) := b"0000000000000000_0000000000000000_0000011010010100_0010101110111110"; -- 0.02569840793236651
	pesos_i(12269) := b"1111111111111111_1111111111111111_1111100111011011_0111010000011011"; -- -0.02399515477328019
	pesos_i(12270) := b"0000000000000000_0000000000000000_0001010010101001_1000000000111100"; -- 0.08071137878782245
	pesos_i(12271) := b"1111111111111111_1111111111111111_1110110010111110_1100111010110100"; -- -0.07521350956610376
	pesos_i(12272) := b"1111111111111111_1111111111111111_1101110101101010_1011101100100100"; -- -0.1350901640230864
	pesos_i(12273) := b"0000000000000000_0000000000000000_0000110111100001_1111111111011001"; -- 0.05422972726658426
	pesos_i(12274) := b"1111111111111111_1111111111111111_1111110100111101_0110101010000011"; -- -0.01078161524870571
	pesos_i(12275) := b"0000000000000000_0000000000000000_0001001100111001_1101000100111010"; -- 0.07510097188388683
	pesos_i(12276) := b"1111111111111111_1111111111111111_1111010010111011_1111010110011010"; -- -0.044006967506547784
	pesos_i(12277) := b"1111111111111111_1111111111111111_1101110101000111_1100000111001111"; -- -0.13562382400366577
	pesos_i(12278) := b"1111111111111111_1111111111111111_1110010001011101_1100000001110100"; -- -0.10794446148028784
	pesos_i(12279) := b"0000000000000000_0000000000000000_0001100101111101_1011011001111000"; -- 0.09957447472135209
	pesos_i(12280) := b"1111111111111111_1111111111111111_1111011100000100_0101000100011010"; -- -0.03509038081471578
	pesos_i(12281) := b"0000000000000000_0000000000000000_0001000111111000_1110101001101001"; -- 0.07020440171552013
	pesos_i(12282) := b"0000000000000000_0000000000000000_0001100010000010_1001101100000100"; -- 0.09574288226490293
	pesos_i(12283) := b"1111111111111111_1111111111111111_1111101000111001_1101110111001010"; -- -0.02255452940008365
	pesos_i(12284) := b"0000000000000000_0000000000000000_0001101100011001_1001001010100000"; -- 0.10585895922421183
	pesos_i(12285) := b"1111111111111111_1111111111111111_1111111000100011_1000111101010011"; -- -0.007269899565507412
	pesos_i(12286) := b"1111111111111111_1111111111111111_1101110110001010_0111110000111110"; -- -0.13460563174636458
	pesos_i(12287) := b"1111111111111111_1111111111111111_1110100010011000_0000011110001100"; -- -0.09143021431787668
	pesos_i(12288) := b"0000000000000000_0000000000000000_0010001111011101_1110111100000001"; -- 0.14010518811480804
	pesos_i(12289) := b"0000000000000000_0000000000000000_0000111100111001_1110111010110110"; -- 0.05947772919241856
	pesos_i(12290) := b"1111111111111111_1111111111111111_1110011110000001_0000011001100101"; -- -0.09568748495676123
	pesos_i(12291) := b"0000000000000000_0000000000000000_0010000010011110_0100111010001110"; -- 0.12741557095744682
	pesos_i(12292) := b"0000000000000000_0000000000000000_0000001011110101_0110000100011001"; -- 0.01155669084522869
	pesos_i(12293) := b"1111111111111111_1111111111111111_1110010001010000_0011111000001111"; -- -0.10815059778704943
	pesos_i(12294) := b"1111111111111111_1111111111111111_1110101011111011_1001100101100000"; -- -0.08209840206473137
	pesos_i(12295) := b"0000000000000000_0000000000000000_0001011110100110_0111101100101100"; -- 0.09238405052162121
	pesos_i(12296) := b"1111111111111111_1111111111111111_1110111101010110_0110100001000111"; -- -0.06508777883204327
	pesos_i(12297) := b"1111111111111111_1111111111111111_1110001010100100_1100110110010011"; -- -0.11467280546059687
	pesos_i(12298) := b"1111111111111111_1111111111111111_1110000110101000_0011111101101100"; -- -0.11852649326770671
	pesos_i(12299) := b"1111111111111111_1111111111111111_1110011000010000_0001101100001100"; -- -0.1013167472093986
	pesos_i(12300) := b"0000000000000000_0000000000000000_0000000001010011_1011001001100111"; -- 0.0012771130603472507
	pesos_i(12301) := b"0000000000000000_0000000000000000_0001011100110110_0101110101111010"; -- 0.09067329620222751
	pesos_i(12302) := b"1111111111111111_1111111111111111_1111100101011110_1011000010001011"; -- -0.02589890112066257
	pesos_i(12303) := b"1111111111111111_1111111111111111_1110111001110101_0100110000100110"; -- -0.06852268283578092
	pesos_i(12304) := b"1111111111111111_1111111111111111_1110100110000101_1100010000111010"; -- -0.0878026349767907
	pesos_i(12305) := b"1111111111111111_1111111111111111_1101110000001111_0110100011001101"; -- -0.14038987147452353
	pesos_i(12306) := b"0000000000000000_0000000000000000_0001011100000111_1110000010101101"; -- 0.08996395321829222
	pesos_i(12307) := b"1111111111111111_1111111111111111_1111101100101101_1101001101101111"; -- -0.018832002150160995
	pesos_i(12308) := b"0000000000000000_0000000000000000_0010001000011011_1001011110111010"; -- 0.13323353093884077
	pesos_i(12309) := b"0000000000000000_0000000000000000_0000000111101011_1001011101111110"; -- 0.007501095160945069
	pesos_i(12310) := b"0000000000000000_0000000000000000_0000000000010101_0010000100010000"; -- 0.00032240529697989266
	pesos_i(12311) := b"1111111111111111_1111111111111111_1110101101011001_1111010100001000"; -- -0.08065861286711047
	pesos_i(12312) := b"1111111111111111_1111111111111111_1110110001011011_1000111101011101"; -- -0.076727904983731
	pesos_i(12313) := b"0000000000000000_0000000000000000_0001110000110111_1100110100010101"; -- 0.11022645729060866
	pesos_i(12314) := b"0000000000000000_0000000000000000_0010001110110110_1011001100011000"; -- 0.13950652435973815
	pesos_i(12315) := b"0000000000000000_0000000000000000_0000011101110001_1010110010001100"; -- 0.029078277659082528
	pesos_i(12316) := b"0000000000000000_0000000000000000_0001000011010101_1011011111011100"; -- 0.06576108095298448
	pesos_i(12317) := b"1111111111111111_1111111111111111_1111010100001011_1111000111010101"; -- -0.042786488906827506
	pesos_i(12318) := b"0000000000000000_0000000000000000_0001000000000101_0000010001011110"; -- 0.06257655435882062
	pesos_i(12319) := b"1111111111111111_1111111111111111_1110100000011010_1000000100101011"; -- -0.09334557239847989
	pesos_i(12320) := b"1111111111111111_1111111111111111_1111010100000011_0100110011010110"; -- -0.04291839387182873
	pesos_i(12321) := b"0000000000000000_0000000000000000_0001001100000000_1000011101110111"; -- 0.07422682437350712
	pesos_i(12322) := b"1111111111111111_1111111111111111_1110010100000001_0001110011000110"; -- -0.10545177613332309
	pesos_i(12323) := b"1111111111111111_1111111111111111_1111000000000010_1111100101001100"; -- -0.06245462320285142
	pesos_i(12324) := b"0000000000000000_0000000000000000_0001110101011011_1101011101000000"; -- 0.11468262979832067
	pesos_i(12325) := b"0000000000000000_0000000000000000_0000011000000001_1001100001010000"; -- 0.02346183732016692
	pesos_i(12326) := b"0000000000000000_0000000000000000_0001101100001000_1101011101000111"; -- 0.10560365176921722
	pesos_i(12327) := b"0000000000000000_0000000000000000_0010000100100010_0100100011111011"; -- 0.12942939870880227
	pesos_i(12328) := b"0000000000000000_0000000000000000_0001000001111110_0111011110010111"; -- 0.06442973563671814
	pesos_i(12329) := b"0000000000000000_0000000000000000_0001101110011001_0000000000001110"; -- 0.10780334787325382
	pesos_i(12330) := b"1111111111111111_1111111111111111_1110010000011101_0000001010101011"; -- -0.10893233615576751
	pesos_i(12331) := b"0000000000000000_0000000000000000_0001000000110100_1010100110011100"; -- 0.06330356652246172
	pesos_i(12332) := b"1111111111111111_1111111111111111_1101110100010111_1101110110000001"; -- -0.1363545951187625
	pesos_i(12333) := b"1111111111111111_1111111111111111_1111110011110010_0101101100111110"; -- -0.011926934600690237
	pesos_i(12334) := b"0000000000000000_0000000000000000_0000101100101010_0000000100001110"; -- 0.043609681945827164
	pesos_i(12335) := b"1111111111111111_1111111111111111_1110010100001000_1000110100001110"; -- -0.10533827218908941
	pesos_i(12336) := b"0000000000000000_0000000000000000_0001000101111011_1001100110010100"; -- 0.06829223502849038
	pesos_i(12337) := b"0000000000000000_0000000000000000_0001101101001011_0110110000010110"; -- 0.10661960162549476
	pesos_i(12338) := b"0000000000000000_0000000000000000_0001010001100100_1100101010001110"; -- 0.07966295220259756
	pesos_i(12339) := b"0000000000000000_0000000000000000_0001100001101010_1000110000000001"; -- 0.09537577650972609
	pesos_i(12340) := b"1111111111111111_1111111111111111_1110010010000000_1010001111100000"; -- -0.10741210738957595
	pesos_i(12341) := b"0000000000000000_0000000000000000_0001111110010001_0111101011000100"; -- 0.12331359190858061
	pesos_i(12342) := b"0000000000000000_0000000000000000_0001100100000100_1011111100111001"; -- 0.09772868293078181
	pesos_i(12343) := b"1111111111111111_1111111111111111_1101011010111110_0100100100001010"; -- -0.16115897669560933
	pesos_i(12344) := b"0000000000000000_0000000000000000_0001010100011011_1111111010110101"; -- 0.08245841894653867
	pesos_i(12345) := b"0000000000000000_0000000000000000_0000101110110101_0111001001101100"; -- 0.04573741078429026
	pesos_i(12346) := b"0000000000000000_0000000000000000_0001010101010110_1101010110100011"; -- 0.08335623965769706
	pesos_i(12347) := b"1111111111111111_1111111111111111_1110101001110110_1010101101101110"; -- -0.08412674497042552
	pesos_i(12348) := b"0000000000000000_0000000000000000_0001101101001100_0000010101010111"; -- 0.1066287363487005
	pesos_i(12349) := b"0000000000000000_0000000000000000_0000111111101110_0011101000101101"; -- 0.062228809323369466
	pesos_i(12350) := b"0000000000000000_0000000000000000_0000010001000111_0001011111100100"; -- 0.016709797989123816
	pesos_i(12351) := b"1111111111111111_1111111111111111_1111011101111111_1111100000111110"; -- -0.033203587308983984
	pesos_i(12352) := b"0000000000000000_0000000000000000_0000111011111101_0101111000111111"; -- 0.05855359111107714
	pesos_i(12353) := b"0000000000000000_0000000000000000_0000101100101001_1011001001011001"; -- 0.04360499062873907
	pesos_i(12354) := b"1111111111111111_1111111111111111_1111111101110001_0001110100101000"; -- -0.002180269021546187
	pesos_i(12355) := b"0000000000000000_0000000000000000_0001111000110001_1110010000011100"; -- 0.11794877696746342
	pesos_i(12356) := b"0000000000000000_0000000000000000_0001101111110110_0011011001001100"; -- 0.10922564854093288
	pesos_i(12357) := b"0000000000000000_0000000000000000_0001011100000110_0111110010011101"; -- 0.08994273034008426
	pesos_i(12358) := b"0000000000000000_0000000000000000_0001000001100011_0001011011111001"; -- 0.06401198932165342
	pesos_i(12359) := b"1111111111111111_1111111111111111_1110100100000111_0010011111001001"; -- -0.08973456705343011
	pesos_i(12360) := b"0000000000000000_0000000000000000_0000110000100101_0101100010001010"; -- 0.04744485264462791
	pesos_i(12361) := b"1111111111111111_1111111111111111_1110101011000100_0000010100001000"; -- -0.08294647754706949
	pesos_i(12362) := b"1111111111111111_1111111111111111_1101101000000011_0000001111100101"; -- -0.1483914915564118
	pesos_i(12363) := b"0000000000000000_0000000000000000_0001000110000100_1011100111010001"; -- 0.0684314856740554
	pesos_i(12364) := b"0000000000000000_0000000000000000_0000101110101100_0001000111010100"; -- 0.045594324352502956
	pesos_i(12365) := b"0000000000000000_0000000000000000_0000011101100011_0111101000110010"; -- 0.028861653623428747
	pesos_i(12366) := b"0000000000000000_0000000000000000_0001001100110101_1010010111100010"; -- 0.07503735314298747
	pesos_i(12367) := b"0000000000000000_0000000000000000_0010010100001011_1100010110111100"; -- 0.1447108824606538
	pesos_i(12368) := b"0000000000000000_0000000000000000_0001000101000110_0010011011101101"; -- 0.06747668549003184
	pesos_i(12369) := b"1111111111111111_1111111111111111_1101111100110010_1010010000100000"; -- -0.1281335280284169
	pesos_i(12370) := b"1111111111111111_1111111111111111_1111010100011010_0010000100010001"; -- -0.04257005055769301
	pesos_i(12371) := b"1111111111111111_1111111111111111_1101101000111100_0010101101010001"; -- -0.1475193908050262
	pesos_i(12372) := b"1111111111111111_1111111111111111_1111111011000101_0000011010011011"; -- -0.004806124763542744
	pesos_i(12373) := b"0000000000000000_0000000000000000_0001101010100101_1101010100001001"; -- 0.10409289806107887
	pesos_i(12374) := b"0000000000000000_0000000000000000_0000011000111110_1000000001011111"; -- 0.024391196492158335
	pesos_i(12375) := b"1111111111111111_1111111111111111_1111110000011100_1000101110111111"; -- -0.015189424486465418
	pesos_i(12376) := b"0000000000000000_0000000000000000_0001001000100010_1100011111100010"; -- 0.07084321281195424
	pesos_i(12377) := b"1111111111111111_1111111111111111_1111110101000101_1010001000000110"; -- -0.01065623611123775
	pesos_i(12378) := b"1111111111111111_1111111111111111_1111100101101101_1101000010011101"; -- -0.025668107703706047
	pesos_i(12379) := b"0000000000000000_0000000000000000_0000001100000000_0110110010011110"; -- 0.01172522404158538
	pesos_i(12380) := b"1111111111111111_1111111111111111_1110000101011101_1111101111011010"; -- -0.11965967112748732
	pesos_i(12381) := b"0000000000000000_0000000000000000_0000001001110001_1010000010000111"; -- 0.00954631141993643
	pesos_i(12382) := b"1111111111111111_1111111111111111_1111000111011101_0011111101001010"; -- -0.05521778531319752
	pesos_i(12383) := b"1111111111111111_1111111111111111_1111100000011010_1000110110110011"; -- -0.030844825477861423
	pesos_i(12384) := b"0000000000000000_0000000000000000_0001101101110101_0101000011100110"; -- 0.10725885023096597
	pesos_i(12385) := b"1111111111111111_1111111111111111_1111111110011110_1010010111111111"; -- -0.001485467100835478
	pesos_i(12386) := b"1111111111111111_1111111111111111_1110111011000001_0100001011000011"; -- -0.06736357436131084
	pesos_i(12387) := b"1111111111111111_1111111111111111_1101110001111110_0111111011011000"; -- -0.13869483202694402
	pesos_i(12388) := b"0000000000000000_0000000000000000_0000100000101101_0000100100010010"; -- 0.03193718620906327
	pesos_i(12389) := b"0000000000000000_0000000000000000_0000000101101011_0100001101011010"; -- 0.005542954868803392
	pesos_i(12390) := b"0000000000000000_0000000000000000_0000010000110001_0010101100110110"; -- 0.016375256278737742
	pesos_i(12391) := b"1111111111111111_1111111111111111_1101110100110101_1101010100011001"; -- -0.1358973325259937
	pesos_i(12392) := b"0000000000000000_0000000000000000_0000011110000111_1010101101111000"; -- 0.02941390682090597
	pesos_i(12393) := b"1111111111111111_1111111111111111_1110000111000001_1011011011011110"; -- -0.11813790396983936
	pesos_i(12394) := b"1111111111111111_1111111111111111_1110110010000010_1001101100011111"; -- -0.07613211153916709
	pesos_i(12395) := b"1111111111111111_1111111111111111_1111110010111011_0000001000110110"; -- -0.012771474587954183
	pesos_i(12396) := b"1111111111111111_1111111111111111_1110101011100010_1010000100000100"; -- -0.0824794163843402
	pesos_i(12397) := b"1111111111111111_1111111111111111_1110101101101001_1101110010011010"; -- -0.08041592824246449
	pesos_i(12398) := b"0000000000000000_0000000000000000_0001100111000010_0100111110101101"; -- 0.10062120419317032
	pesos_i(12399) := b"0000000000000000_0000000000000000_0000100001010000_1110101001001011"; -- 0.03248466804465991
	pesos_i(12400) := b"0000000000000000_0000000000000000_0000000110110010_0000111100010100"; -- 0.006623213289001971
	pesos_i(12401) := b"0000000000000000_0000000000000000_0001101010001110_0110001110110100"; -- 0.10373519085119137
	pesos_i(12402) := b"0000000000000000_0000000000000000_0001000100000101_0100010011110110"; -- 0.06648665428369513
	pesos_i(12403) := b"1111111111111111_1111111111111111_1110000111011101_0010101110111110"; -- -0.11771895034885958
	pesos_i(12404) := b"1111111111111111_1111111111111111_1111111010010001_1010100010001010"; -- -0.005589929834370927
	pesos_i(12405) := b"0000000000000000_0000000000000000_0000111010110000_1111101000111110"; -- 0.05738796252643464
	pesos_i(12406) := b"0000000000000000_0000000000000000_0010011010001110_1101011111110000"; -- 0.15061711886993573
	pesos_i(12407) := b"0000000000000000_0000000000000000_0010000100101111_1001011100001010"; -- 0.12963241581945942
	pesos_i(12408) := b"0000000000000000_0000000000000000_0001111001111001_1110000010010010"; -- 0.11904719894256553
	pesos_i(12409) := b"1111111111111111_1111111111111111_1110110100110111_1101111010111010"; -- -0.07336624104454785
	pesos_i(12410) := b"0000000000000000_0000000000000000_0010001110100000_0111110101111001"; -- 0.13916763495366055
	pesos_i(12411) := b"1111111111111111_1111111111111111_1111000011010100_0101110101000010"; -- -0.05925957814773277
	pesos_i(12412) := b"1111111111111111_1111111111111111_1101101100110111_0111111011100010"; -- -0.14368445372362798
	pesos_i(12413) := b"1111111111111111_1111111111111111_1111001110011001_1100001101111001"; -- -0.048435004268819554
	pesos_i(12414) := b"0000000000000000_0000000000000000_0000110001011000_0011110101101100"; -- 0.04822143456644238
	pesos_i(12415) := b"0000000000000000_0000000000000000_0000100100000100_0101001000110001"; -- 0.035222184141850986
	pesos_i(12416) := b"1111111111111111_1111111111111111_1101111001001010_0010111001001000"; -- -0.13168059107228955
	pesos_i(12417) := b"1111111111111111_1111111111111111_1110011100110101_0100110110011010"; -- -0.09684290881355737
	pesos_i(12418) := b"1111111111111111_1111111111111111_1110110100111000_0100010101100000"; -- -0.07336012282298436
	pesos_i(12419) := b"0000000000000000_0000000000000000_0000001110111101_0110000110111011"; -- 0.014608486231060498
	pesos_i(12420) := b"1111111111111111_1111111111111111_1111011101000110_1110110100110000"; -- -0.034073997234184715
	pesos_i(12421) := b"0000000000000000_0000000000000000_0010101010110001_0011101100110011"; -- 0.16676683430618114
	pesos_i(12422) := b"0000000000000000_0000000000000000_0000101101010011_1000111110111000"; -- 0.044243795844966335
	pesos_i(12423) := b"1111111111111111_1111111111111111_1111000010101001_0111000100000101"; -- -0.0599145281644287
	pesos_i(12424) := b"1111111111111111_1111111111111111_1111111111010110_1110011000000001"; -- -0.0006271598853358244
	pesos_i(12425) := b"0000000000000000_0000000000000000_0001010101110101_1110001101000111"; -- 0.0838300751897399
	pesos_i(12426) := b"0000000000000000_0000000000000000_0001000010011101_0110110010000110"; -- 0.0649020983110794
	pesos_i(12427) := b"0000000000000000_0000000000000000_0001000000000111_0011101101100000"; -- 0.06261035048021768
	pesos_i(12428) := b"0000000000000000_0000000000000000_0001010111100010_1010011100111000"; -- 0.08548970335412187
	pesos_i(12429) := b"1111111111111111_1111111111111111_1110100111101011_0001001101011001"; -- -0.08625678142015927
	pesos_i(12430) := b"0000000000000000_0000000000000000_0001111101111001_1101110011011101"; -- 0.12295322797389004
	pesos_i(12431) := b"0000000000000000_0000000000000000_0001100001100111_1011010101100010"; -- 0.09533246661080966
	pesos_i(12432) := b"1111111111111111_1111111111111111_1101110100110001_1101101001001101"; -- -0.13595805757110235
	pesos_i(12433) := b"0000000000000000_0000000000000000_0001111101001000_0101000011000000"; -- 0.12219719597370884
	pesos_i(12434) := b"1111111111111111_1111111111111111_1110001000111101_0110010111011111"; -- -0.11625064185965633
	pesos_i(12435) := b"0000000000000000_0000000000000000_0001110110010101_0100000111110001"; -- 0.11555873993310177
	pesos_i(12436) := b"1111111111111111_1111111111111111_1110011011011010_1011111010010010"; -- -0.09822472510514978
	pesos_i(12437) := b"0000000000000000_0000000000000000_0000011101100111_1100110000010110"; -- 0.02892756971261322
	pesos_i(12438) := b"0000000000000000_0000000000000000_0000001100111110_1111010110001000"; -- 0.012679429797497399
	pesos_i(12439) := b"0000000000000000_0000000000000000_0001011010111110_0011100010011110"; -- 0.08884004466704407
	pesos_i(12440) := b"1111111111111111_1111111111111111_1110010111100110_1110001001101011"; -- -0.10194573288154679
	pesos_i(12441) := b"0000000000000000_0000000000000000_0001010110100010_0000101110110000"; -- 0.0845038704856801
	pesos_i(12442) := b"1111111111111111_1111111111111111_1110111110111100_1001011000011110"; -- -0.06352864994501191
	pesos_i(12443) := b"1111111111111111_1111111111111111_1111010001101101_0010011111111100"; -- -0.04520940881733222
	pesos_i(12444) := b"0000000000000000_0000000000000000_0000000110110101_0101001100110001"; -- 0.0066730493742326764
	pesos_i(12445) := b"0000000000000000_0000000000000000_0001101100001011_1101110111000000"; -- 0.10564981410326872
	pesos_i(12446) := b"0000000000000000_0000000000000000_0000000001011100_1010001010011010"; -- 0.0014135003042941032
	pesos_i(12447) := b"1111111111111111_1111111111111111_1111111110100100_1001011111010111"; -- -0.0013947582834029535
	pesos_i(12448) := b"1111111111111111_1111111111111111_1110010110111011_0101000111101101"; -- -0.10261047330384737
	pesos_i(12449) := b"1111111111111111_1111111111111111_1110000110101110_0110100011110100"; -- -0.11843246498393213
	pesos_i(12450) := b"1111111111111111_1111111111111111_1110000111100111_0001110001110000"; -- -0.11756727468957866
	pesos_i(12451) := b"0000000000000000_0000000000000000_0010101000000100_0101011100100001"; -- 0.16412872851240687
	pesos_i(12452) := b"0000000000000000_0000000000000000_0001111110000101_1101110010010111"; -- 0.12313631723435098
	pesos_i(12453) := b"1111111111111111_1111111111111111_1111101011011000_0111110110110011"; -- -0.02013410931817705
	pesos_i(12454) := b"1111111111111111_1111111111111111_1110111100110001_1011011000010101"; -- -0.06564771645940423
	pesos_i(12455) := b"0000000000000000_0000000000000000_0001001000001000_0101110100001100"; -- 0.07044011638930726
	pesos_i(12456) := b"0000000000000000_0000000000000000_0000011101000010_0110111101011011"; -- 0.02835746730907864
	pesos_i(12457) := b"1111111111111111_1111111111111111_1111111110101101_0011001111110101"; -- -0.0012633826188354744
	pesos_i(12458) := b"0000000000000000_0000000000000000_0000111000110011_1001110011011111"; -- 0.055475048376804004
	pesos_i(12459) := b"1111111111111111_1111111111111111_1111011100001011_1111000000111001"; -- -0.03497408495539864
	pesos_i(12460) := b"0000000000000000_0000000000000000_0001011100011001_0000001111011100"; -- 0.09022544977587985
	pesos_i(12461) := b"1111111111111111_1111111111111111_1111111011011110_1110110100010001"; -- -0.004410918492084963
	pesos_i(12462) := b"1111111111111111_1111111111111111_1110011100001101_1010010011100100"; -- -0.09744805743030362
	pesos_i(12463) := b"1111111111111111_1111111111111111_1111001111101001_1100011101001111"; -- -0.04721407250225152
	pesos_i(12464) := b"1111111111111111_1111111111111111_1110001001001010_0110000101001101"; -- -0.11605254996814587
	pesos_i(12465) := b"0000000000000000_0000000000000000_0010011000111111_1110110001010010"; -- 0.14941288952653736
	pesos_i(12466) := b"1111111111111111_1111111111111111_1101111010010001_1011110010011011"; -- -0.13058873389890183
	pesos_i(12467) := b"1111111111111111_1111111111111111_1101110100111001_0111011110001111"; -- -0.13584187273122758
	pesos_i(12468) := b"1111111111111111_1111111111111111_1110010110001000_0010011011110111"; -- -0.10339123209484308
	pesos_i(12469) := b"0000000000000000_0000000000000000_0010001010001001_0001000100010011"; -- 0.13490397180677882
	pesos_i(12470) := b"0000000000000000_0000000000000000_0001100000010010_1111010000100011"; -- 0.09403920990451069
	pesos_i(12471) := b"0000000000000000_0000000000000000_0000101010111110_1010111000010101"; -- 0.041972045985527326
	pesos_i(12472) := b"1111111111111111_1111111111111111_1110010111000011_0000100011101010"; -- -0.10249275486739735
	pesos_i(12473) := b"1111111111111111_1111111111111111_1110010101011010_1000011000100011"; -- -0.10408746390306602
	pesos_i(12474) := b"0000000000000000_0000000000000000_0000001001100111_0100101000010000"; -- 0.009388569800658596
	pesos_i(12475) := b"0000000000000000_0000000000000000_0001110101001100_1001001010101110"; -- 0.11444966085591786
	pesos_i(12476) := b"1111111111111111_1111111111111111_1111000001011011_0101110110110001"; -- -0.06110586575052013
	pesos_i(12477) := b"0000000000000000_0000000000000000_0000100001111010_0110110111100000"; -- 0.03311812124379627
	pesos_i(12478) := b"0000000000000000_0000000000000000_0000011110111110_0010110001110101"; -- 0.03024556979581314
	pesos_i(12479) := b"1111111111111111_1111111111111111_1101101001101100_1011100000101010"; -- -0.1467785738272748
	pesos_i(12480) := b"0000000000000000_0000000000000000_0000000110110101_0001000101010000"; -- 0.006669122746461741
	pesos_i(12481) := b"0000000000000000_0000000000000000_0001000110000100_1001010110111010"; -- 0.06842933446222085
	pesos_i(12482) := b"0000000000000000_0000000000000000_0001001010110100_0010110000100001"; -- 0.07306171224747378
	pesos_i(12483) := b"1111111111111111_1111111111111111_1110100110101100_0010010101101100"; -- -0.08721700765804022
	pesos_i(12484) := b"1111111111111111_1111111111111111_1110110000001011_1010100100011110"; -- -0.07794707303706672
	pesos_i(12485) := b"1111111111111111_1111111111111111_1111001101110111_1101001100001000"; -- -0.04895287569621213
	pesos_i(12486) := b"0000000000000000_0000000000000000_0000001011011011_0010000110111001"; -- 0.011156184773204347
	pesos_i(12487) := b"1111111111111111_1111111111111111_1101101100000011_0001111111000000"; -- -0.14448358111591225
	pesos_i(12488) := b"0000000000000000_0000000000000000_0010010100110001_0110101110101000"; -- 0.14528534759111747
	pesos_i(12489) := b"0000000000000000_0000000000000000_0010000101111110_0111101111010011"; -- 0.1308362379752511
	pesos_i(12490) := b"0000000000000000_0000000000000000_0000011101111100_1100011100011110"; -- 0.02924770822966666
	pesos_i(12491) := b"1111111111111111_1111111111111111_1101111110010000_1010110100101010"; -- -0.12669866292889845
	pesos_i(12492) := b"1111111111111111_1111111111111111_1101101110001011_1010111011010111"; -- -0.14239985695409435
	pesos_i(12493) := b"1111111111111111_1111111111111111_1111110001011100_0011000100000000"; -- -0.014218270688904987
	pesos_i(12494) := b"0000000000000000_0000000000000000_0000110011001001_1010101001111010"; -- 0.049952177690598246
	pesos_i(12495) := b"1111111111111111_1111111111111111_1101100111101000_1011111001100110"; -- -0.14879236227897855
	pesos_i(12496) := b"0000000000000000_0000000000000000_0000010110000100_1101001110100011"; -- 0.02155802478298285
	pesos_i(12497) := b"1111111111111111_1111111111111111_1110011110011000_0110010000101001"; -- -0.09533094412087935
	pesos_i(12498) := b"0000000000000000_0000000000000000_0001101100100011_0110010101101111"; -- 0.10600885346907864
	pesos_i(12499) := b"0000000000000000_0000000000000000_0000110010111110_1010111010101000"; -- 0.049784580188180605
	pesos_i(12500) := b"1111111111111111_1111111111111111_1110110110100011_0011010010100100"; -- -0.07172842969760417
	pesos_i(12501) := b"1111111111111111_1111111111111111_1111110110010010_0110001100111011"; -- -0.009485052246766816
	pesos_i(12502) := b"0000000000000000_0000000000000000_0001111000110010_0111111101011101"; -- 0.11795803086462349
	pesos_i(12503) := b"0000000000000000_0000000000000000_0010000111010010_0110110000010100"; -- 0.13211703772908098
	pesos_i(12504) := b"0000000000000000_0000000000000000_0000101101100111_1001100101001010"; -- 0.04454954202444463
	pesos_i(12505) := b"1111111111111111_1111111111111111_1111110100111000_1101110011010010"; -- -0.010851095871349598
	pesos_i(12506) := b"1111111111111111_1111111111111111_1110111101011111_1011111100110101"; -- -0.06494526819605777
	pesos_i(12507) := b"0000000000000000_0000000000000000_0000001110010111_0010110101110111"; -- 0.01402553702425218
	pesos_i(12508) := b"1111111111111111_1111111111111111_1111001000110011_0011100001100101"; -- -0.053905940484624534
	pesos_i(12509) := b"0000000000000000_0000000000000000_0001110011011111_1110010101001001"; -- 0.11279137631007836
	pesos_i(12510) := b"1111111111111111_1111111111111111_1110000110010101_1101100101100110"; -- -0.11880723239964847
	pesos_i(12511) := b"1111111111111111_1111111111111111_1111110110011000_1011011101001111"; -- -0.009388487921650122
	pesos_i(12512) := b"0000000000000000_0000000000000000_0001111011111111_0010100001011111"; -- 0.12108089741181187
	pesos_i(12513) := b"1111111111111111_1111111111111111_1101111011111000_0110010010100010"; -- -0.129022322156268
	pesos_i(12514) := b"1111111111111111_1111111111111111_1110001000100110_1010011110000101"; -- -0.11659768108983067
	pesos_i(12515) := b"1111111111111111_1111111111111111_1111011010100100_0111010010110011"; -- -0.03655310272284801
	pesos_i(12516) := b"1111111111111111_1111111111111111_1111101011110011_1000000110101101"; -- -0.01972188486424522
	pesos_i(12517) := b"0000000000000000_0000000000000000_0001001011100000_0101110100110111"; -- 0.07373602483443574
	pesos_i(12518) := b"1111111111111111_1111111111111111_1111011111010000_0011010001111110"; -- -0.031979293155921476
	pesos_i(12519) := b"1111111111111111_1111111111111111_1110000001100000_0110011100001001"; -- -0.12352901482501077
	pesos_i(12520) := b"1111111111111111_1111111111111111_1110111000010000_1001100110101000"; -- -0.07005920085024898
	pesos_i(12521) := b"1111111111111111_1111111111111111_1110101110000001_1000111110100111"; -- -0.0800543038887372
	pesos_i(12522) := b"1111111111111111_1111111111111111_1110110011010011_1101001011101000"; -- -0.07489282453608143
	pesos_i(12523) := b"1111111111111111_1111111111111111_1110010111101101_0111000101100110"; -- -0.10184565792319263
	pesos_i(12524) := b"1111111111111111_1111111111111111_1111110010111110_0110011001110000"; -- -0.012719724382817054
	pesos_i(12525) := b"1111111111111111_1111111111111111_1110110100011100_0111000000100001"; -- -0.07378482041262946
	pesos_i(12526) := b"1111111111111111_1111111111111111_1111010100010010_0000011100111000"; -- -0.04269366148597224
	pesos_i(12527) := b"1111111111111111_1111111111111111_1111110010100000_0100000101101000"; -- -0.013179695180873835
	pesos_i(12528) := b"1111111111111111_1111111111111111_1101111101001100_0111111000001101"; -- -0.12773906887615258
	pesos_i(12529) := b"1111111111111111_1111111111111111_1101111111011000_0100101011011000"; -- -0.12560589056891053
	pesos_i(12530) := b"1111111111111111_1111111111111111_1111011110011111_1110110011111100"; -- -0.03271597719005051
	pesos_i(12531) := b"1111111111111111_1111111111111111_1111000000000110_0101101001100101"; -- -0.06240305931800273
	pesos_i(12532) := b"1111111111111111_1111111111111111_1110000111010110_0100001011010011"; -- -0.11782438599641319
	pesos_i(12533) := b"1111111111111111_1111111111111111_1110001001101101_0111111110111101"; -- -0.11551667815344245
	pesos_i(12534) := b"1111111111111111_1111111111111111_1111110011100001_0000010010001110"; -- -0.012191500908530693
	pesos_i(12535) := b"1111111111111111_1111111111111111_1111110001100000_0111101000110000"; -- -0.014152873352494157
	pesos_i(12536) := b"0000000000000000_0000000000000000_0010010011100011_1001101011000110"; -- 0.1440979704340799
	pesos_i(12537) := b"0000000000000000_0000000000000000_0010010010111000_0101011000001010"; -- 0.1434377454860298
	pesos_i(12538) := b"0000000000000000_0000000000000000_0001100101111111_0110101100101101"; -- 0.0996005042943779
	pesos_i(12539) := b"1111111111111111_1111111111111111_1110001101001010_1111011011100011"; -- -0.11213738398653791
	pesos_i(12540) := b"1111111111111111_1111111111111111_1110101101011000_1001111001011010"; -- -0.0806790380281271
	pesos_i(12541) := b"1111111111111111_1111111111111111_1111010000110010_1110110010101000"; -- -0.0460979546854308
	pesos_i(12542) := b"0000000000000000_0000000000000000_0000111101101111_0101010110110010"; -- 0.06029258340434514
	pesos_i(12543) := b"1111111111111111_1111111111111111_1111110011010000_1010100011100001"; -- -0.012441105892066718
	pesos_i(12544) := b"1111111111111111_1111111111111111_1110111111100100_0101101110001110"; -- -0.06292178903800619
	pesos_i(12545) := b"1111111111111111_1111111111111111_1111010110100000_0110010010010110"; -- -0.04052134842299115
	pesos_i(12546) := b"1111111111111111_1111111111111111_1111000110101001_0111111001111010"; -- -0.056007476076460165
	pesos_i(12547) := b"0000000000000000_0000000000000000_0000010000001010_0011100101001111"; -- 0.015781003780793394
	pesos_i(12548) := b"1111111111111111_1111111111111111_1110010101000111_0001100011000010"; -- -0.10438390031029271
	pesos_i(12549) := b"1111111111111111_1111111111111111_1111110101111111_1000100000011011"; -- -0.00977277128343282
	pesos_i(12550) := b"1111111111111111_1111111111111111_1111001010110010_1101100000111111"; -- -0.05195854621823132
	pesos_i(12551) := b"1111111111111111_1111111111111111_1111110001111110_0011000000110010"; -- -0.01369951991373903
	pesos_i(12552) := b"1111111111111111_1111111111111111_1110000101001111_0010101001010100"; -- -0.11988578272123346
	pesos_i(12553) := b"0000000000000000_0000000000000000_0000001011011001_1111000011110011"; -- 0.011138018818704283
	pesos_i(12554) := b"0000000000000000_0000000000000000_0010001001101110_1110010000000010"; -- 0.13450455704508968
	pesos_i(12555) := b"0000000000000000_0000000000000000_0000001010111111_1100011101001101"; -- 0.010738808069105064
	pesos_i(12556) := b"1111111111111111_1111111111111111_1111011100110101_0100111010110100"; -- -0.0343428431976698
	pesos_i(12557) := b"0000000000000000_0000000000000000_0001011110001110_1110100010111001"; -- 0.09202436930960695
	pesos_i(12558) := b"1111111111111111_1111111111111111_1110110001011011_1100000100110011"; -- -0.07672493462417014
	pesos_i(12559) := b"1111111111111111_1111111111111111_1110001000011101_1111110010000001"; -- -0.11672994467465383
	pesos_i(12560) := b"1111111111111111_1111111111111111_1110100010001011_1010000010001010"; -- -0.09161945936263739
	pesos_i(12561) := b"0000000000000000_0000000000000000_0000111001001000_1000110100111000"; -- 0.05579455001027786
	pesos_i(12562) := b"0000000000000000_0000000000000000_0000111010100110_0111100110000110"; -- 0.057227702354054125
	pesos_i(12563) := b"1111111111111111_1111111111111111_1101110001110101_1011000110100100"; -- -0.13882913355722695
	pesos_i(12564) := b"0000000000000000_0000000000000000_0000111001111001_1100011001101111"; -- 0.05654564106500168
	pesos_i(12565) := b"1111111111111111_1111111111111111_1111010011000100_0111111100010100"; -- -0.043876702941989
	pesos_i(12566) := b"1111111111111111_1111111111111111_1101100010010010_0011110111010011"; -- -0.1540185318533208
	pesos_i(12567) := b"0000000000000000_0000000000000000_0001001100010101_0011101101110011"; -- 0.07454272791651947
	pesos_i(12568) := b"0000000000000000_0000000000000000_0001000111010110_0001111010100111"; -- 0.06967345782402133
	pesos_i(12569) := b"0000000000000000_0000000000000000_0000001010100010_1111001001100101"; -- 0.01029887177459446
	pesos_i(12570) := b"1111111111111111_1111111111111111_1110100110001100_0010001111011101"; -- -0.0877053818684376
	pesos_i(12571) := b"0000000000000000_0000000000000000_0010000001111010_0010010000100110"; -- 0.1268637267766025
	pesos_i(12572) := b"1111111111111111_1111111111111111_1111010010100000_1001011101011111"; -- -0.04442457144371421
	pesos_i(12573) := b"0000000000000000_0000000000000000_0000111110001111_0000000011101101"; -- 0.06077581208864725
	pesos_i(12574) := b"1111111111111111_1111111111111111_1111110001000010_0011001011010000"; -- -0.014614891301022784
	pesos_i(12575) := b"1111111111111111_1111111111111111_1110110101000100_0010011101111000"; -- -0.07317879992282322
	pesos_i(12576) := b"1111111111111111_1111111111111111_1110111011110100_0010001001001000"; -- -0.06658731221124418
	pesos_i(12577) := b"1111111111111111_1111111111111111_1111110111110011_1001010111001011"; -- -0.008001935911683973
	pesos_i(12578) := b"1111111111111111_1111111111111111_1111011010000101_1011010010111000"; -- -0.037022309369927044
	pesos_i(12579) := b"0000000000000000_0000000000000000_0001000110011001_1011010111001001"; -- 0.06875168005188313
	pesos_i(12580) := b"1111111111111111_1111111111111111_1110100101110001_0011110010010011"; -- -0.0881158964058235
	pesos_i(12581) := b"1111111111111111_1111111111111111_1101111000001000_1100010110001101"; -- -0.13267865467324946
	pesos_i(12582) := b"1111111111111111_1111111111111111_1111010011010100_1101010011111001"; -- -0.04362744255454411
	pesos_i(12583) := b"0000000000000000_0000000000000000_0001010111010110_0110001010001111"; -- 0.08530250537619996
	pesos_i(12584) := b"0000000000000000_0000000000000000_0010000001101110_0100010101000101"; -- 0.1266825955318626
	pesos_i(12585) := b"0000000000000000_0000000000000000_0000010110001101_0111111000000001"; -- 0.021690249675553375
	pesos_i(12586) := b"0000000000000000_0000000000000000_0000111100011010_1000000101010010"; -- 0.058998186602122624
	pesos_i(12587) := b"1111111111111111_1111111111111111_1110001010101100_1100110011110110"; -- -0.11455077157521211
	pesos_i(12588) := b"0000000000000000_0000000000000000_0000010110011111_1010110101101100"; -- 0.021967734171732003
	pesos_i(12589) := b"1111111111111111_1111111111111111_1101111001000101_1101010100111011"; -- -0.13174693410618277
	pesos_i(12590) := b"0000000000000000_0000000000000000_0001010111001010_1110110001000001"; -- 0.08512760716065482
	pesos_i(12591) := b"0000000000000000_0000000000000000_0001100110010101_0010000000101101"; -- 0.09993172748207556
	pesos_i(12592) := b"1111111111111111_1111111111111111_1111100101111101_1011110111000011"; -- -0.025425090700930787
	pesos_i(12593) := b"0000000000000000_0000000000000000_0010000111110000_0001111110000000"; -- 0.13257023695014972
	pesos_i(12594) := b"1111111111111111_1111111111111111_1110000110011010_1100010110110010"; -- -0.1187321128895754
	pesos_i(12595) := b"1111111111111111_1111111111111111_1110100101111011_1011011011000000"; -- -0.08795602625979275
	pesos_i(12596) := b"1111111111111111_1111111111111111_1110010010110001_0011011101010110"; -- -0.10667089614391738
	pesos_i(12597) := b"1111111111111111_1111111111111111_1110010000001111_1101110101000001"; -- -0.10913293038526811
	pesos_i(12598) := b"0000000000000000_0000000000000000_0001000111011101_0011010000010010"; -- 0.06978154611858063
	pesos_i(12599) := b"1111111111111111_1111111111111111_1110110111100101_0110111100110000"; -- -0.07071786009553545
	pesos_i(12600) := b"0000000000000000_0000000000000000_0000001001000010_0010001110101110"; -- 0.00882170675957132
	pesos_i(12601) := b"1111111111111111_1111111111111111_1110010001001010_0000111001001001"; -- -0.10824499813034309
	pesos_i(12602) := b"1111111111111111_1111111111111111_1111111110111111_0000111111101011"; -- -0.00099087253881772
	pesos_i(12603) := b"1111111111111111_1111111111111111_1110100010101001_0100011100111110"; -- -0.09116701834926973
	pesos_i(12604) := b"1111111111111111_1111111111111111_1111001110100100_1111011110100011"; -- -0.04826404824123269
	pesos_i(12605) := b"1111111111111111_1111111111111111_1110100010000001_0101111101000011"; -- -0.09177593816344476
	pesos_i(12606) := b"1111111111111111_1111111111111111_1111001111110001_1000101101110000"; -- -0.04709557078838042
	pesos_i(12607) := b"1111111111111111_1111111111111111_1111010101100111_0111010001111111"; -- -0.04139015111553849
	pesos_i(12608) := b"1111111111111111_1111111111111111_1110110101011111_1010110111011100"; -- -0.07275880226138624
	pesos_i(12609) := b"0000000000000000_0000000000000000_0000101100101100_0000011101100000"; -- 0.04364057619008702
	pesos_i(12610) := b"0000000000000000_0000000000000000_0001111000100100_1110001101101000"; -- 0.11775037090014746
	pesos_i(12611) := b"1111111111111111_1111111111111111_1111001010001111_0010000000101010"; -- -0.05250357602063883
	pesos_i(12612) := b"0000000000000000_0000000000000000_0000111011000010_1001000111101011"; -- 0.05765640237512153
	pesos_i(12613) := b"0000000000000000_0000000000000000_0001010010001110_1001001110001001"; -- 0.08030054190525897
	pesos_i(12614) := b"1111111111111111_1111111111111111_1111000110011000_0010010001010100"; -- -0.05627224883285858
	pesos_i(12615) := b"1111111111111111_1111111111111111_1101100110101111_0111011100011001"; -- -0.14966636324411944
	pesos_i(12616) := b"1111111111111111_1111111111111111_1110101110101001_0101001101111010"; -- -0.07944753903057135
	pesos_i(12617) := b"0000000000000000_0000000000000000_0010000000011011_1100110111111010"; -- 0.12542426435752174
	pesos_i(12618) := b"1111111111111111_1111111111111111_1110110010000001_0001100101110000"; -- -0.07615510001724647
	pesos_i(12619) := b"1111111111111111_1111111111111111_1111101010001010_1100110001101011"; -- -0.021319602829356483
	pesos_i(12620) := b"0000000000000000_0000000000000000_0001111110111100_1101101111111111"; -- 0.12397551523314404
	pesos_i(12621) := b"0000000000000000_0000000000000000_0000110110100111_1000011001111110"; -- 0.053337484118708596
	pesos_i(12622) := b"1111111111111111_1111111111111111_1101101010100110_0100101111101000"; -- -0.14590001661099106
	pesos_i(12623) := b"1111111111111111_1111111111111111_1110110101011110_0111000001110000"; -- -0.07277772195447019
	pesos_i(12624) := b"0000000000000000_0000000000000000_0000010101110111_0101111100110110"; -- 0.021352720877179588
	pesos_i(12625) := b"0000000000000000_0000000000000000_0010001010110111_0101001101010101"; -- 0.1356098253126453
	pesos_i(12626) := b"0000000000000000_0000000000000000_0010001101110110_1010110110111000"; -- 0.13852964161007444
	pesos_i(12627) := b"1111111111111111_1111111111111111_1101110101111001_0001110000000111"; -- -0.13487076596319056
	pesos_i(12628) := b"0000000000000000_0000000000000000_0000000100010001_0110100010001010"; -- 0.00417188034763679
	pesos_i(12629) := b"1111111111111111_1111111111111111_1111010000000011_1111101100111000"; -- -0.046814249900083274
	pesos_i(12630) := b"1111111111111111_1111111111111111_1111011001001101_0111011010000110"; -- -0.0378805086563001
	pesos_i(12631) := b"1111111111111111_1111111111111111_1101110000010011_0000111001010011"; -- -0.14033422918312727
	pesos_i(12632) := b"0000000000000000_0000000000000000_0001111110101110_1000001001111001"; -- 0.12375655618828181
	pesos_i(12633) := b"0000000000000000_0000000000000000_0010010111000000_1000001110111010"; -- 0.14746878910924482
	pesos_i(12634) := b"1111111111111111_1111111111111111_1101111000110000_1101000110110010"; -- -0.1320675792021562
	pesos_i(12635) := b"0000000000000000_0000000000000000_0000101000000111_1001101110110011"; -- 0.03917859187958258
	pesos_i(12636) := b"0000000000000000_0000000000000000_0010001010111101_1111111000001100"; -- 0.13571155340370922
	pesos_i(12637) := b"0000000000000000_0000000000000000_0001001110011101_0001110010000001"; -- 0.07661607878443966
	pesos_i(12638) := b"0000000000000000_0000000000000000_0000011101110011_0100111001000010"; -- 0.02910317538681229
	pesos_i(12639) := b"0000000000000000_0000000000000000_0001001111011011_0111111010101101"; -- 0.07756797537582455
	pesos_i(12640) := b"0000000000000000_0000000000000000_0010000001000010_0000110101101000"; -- 0.12600787918686088
	pesos_i(12641) := b"0000000000000000_0000000000000000_0001111000011000_0111111001111100"; -- 0.11756125000085607
	pesos_i(12642) := b"0000000000000000_0000000000000000_0001100110011011_1011101100010101"; -- 0.10003251323888616
	pesos_i(12643) := b"1111111111111111_1111111111111111_1110111111111000_0001100110010101"; -- -0.06262054551842537
	pesos_i(12644) := b"1111111111111111_1111111111111111_1111000110101100_1000011011111110"; -- -0.05596119202995491
	pesos_i(12645) := b"1111111111111111_1111111111111111_1101101110100011_1100101010100111"; -- -0.14203198846150678
	pesos_i(12646) := b"0000000000000000_0000000000000000_0010011110100101_1000110101111110"; -- 0.1548698836855503
	pesos_i(12647) := b"0000000000000000_0000000000000000_0000100000010001_0100111100010110"; -- 0.03151411330478663
	pesos_i(12648) := b"1111111111111111_1111111111111111_1101100110001001_0011000101111000"; -- -0.15025034733548565
	pesos_i(12649) := b"1111111111111111_1111111111111111_1111101011101010_0011110110001011"; -- -0.019863275050748114
	pesos_i(12650) := b"1111111111111111_1111111111111111_1101110100001001_1111011110111011"; -- -0.13656665499149526
	pesos_i(12651) := b"0000000000000000_0000000000000000_0000010010101001_0101010010101011"; -- 0.018208782015001417
	pesos_i(12652) := b"1111111111111111_1111111111111111_1111100110001110_1011010000011001"; -- -0.02516626737006096
	pesos_i(12653) := b"0000000000000000_0000000000000000_0000101000100000_0101011010111010"; -- 0.03955595045703303
	pesos_i(12654) := b"1111111111111111_1111111111111111_1110101110011001_0011111110011111"; -- -0.07969286319332461
	pesos_i(12655) := b"1111111111111111_1111111111111111_1111100000010101_0000010111010000"; -- -0.03092921903244501
	pesos_i(12656) := b"1111111111111111_1111111111111111_1101111101000000_1000101100101101"; -- -0.12792139197215344
	pesos_i(12657) := b"1111111111111111_1111111111111111_1111001001100100_0100101100001111"; -- -0.053157147280524376
	pesos_i(12658) := b"1111111111111111_1111111111111111_1110101111101011_1100111100000110"; -- -0.07843309500893145
	pesos_i(12659) := b"1111111111111111_1111111111111111_1111101011011100_1000000111101100"; -- -0.020072822544390433
	pesos_i(12660) := b"1111111111111111_1111111111111111_1111111101111100_1000010001100100"; -- -0.002006268974643785
	pesos_i(12661) := b"0000000000000000_0000000000000000_0001110001001010_1100101110101110"; -- 0.11051629057869274
	pesos_i(12662) := b"1111111111111111_1111111111111111_1111111011111010_1110000010010001"; -- -0.003984417567004351
	pesos_i(12663) := b"0000000000000000_0000000000000000_0010001011011110_1011111101100101"; -- 0.13621135927552014
	pesos_i(12664) := b"0000000000000000_0000000000000000_0010000100111000_0000011010011101"; -- 0.12976113626174002
	pesos_i(12665) := b"1111111111111111_1111111111111111_1111011110101100_0110010001111011"; -- -0.03252574912367738
	pesos_i(12666) := b"0000000000000000_0000000000000000_0010000111011101_0100010111000101"; -- 0.13228260101816808
	pesos_i(12667) := b"0000000000000000_0000000000000000_0000101010001110_0110000110010001"; -- 0.04123506355581273
	pesos_i(12668) := b"0000000000000000_0000000000000000_0000100100010100_0101010000000011"; -- 0.035466433385232
	pesos_i(12669) := b"0000000000000000_0000000000000000_0000111001111000_0000011000111101"; -- 0.05651892642777726
	pesos_i(12670) := b"0000000000000000_0000000000000000_0000100100000111_0001101110101011"; -- 0.03526471054738085
	pesos_i(12671) := b"1111111111111111_1111111111111111_1111100110010101_1010011101111000"; -- -0.025060208592838664
	pesos_i(12672) := b"1111111111111111_1111111111111111_1110111001111111_0111001011011111"; -- -0.06836778685289738
	pesos_i(12673) := b"0000000000000000_0000000000000000_0001101111101101_1111100000100011"; -- 0.10909987320288707
	pesos_i(12674) := b"1111111111111111_1111111111111111_1110101100011110_0011100000111111"; -- -0.08157013374973619
	pesos_i(12675) := b"1111111111111111_1111111111111111_1111001011000101_1110101111011101"; -- -0.0516674601163387
	pesos_i(12676) := b"1111111111111111_1111111111111111_1111010111011100_0011010110110110"; -- -0.03960861487580427
	pesos_i(12677) := b"0000000000000000_0000000000000000_0001000011001001_1010101001101110"; -- 0.06557717495441273
	pesos_i(12678) := b"0000000000000000_0000000000000000_0000011111000001_0001001001101000"; -- 0.030289793386583972
	pesos_i(12679) := b"1111111111111111_1111111111111111_1110000111010110_0110110101111000"; -- -0.11782184434016259
	pesos_i(12680) := b"0000000000000000_0000000000000000_0000001101011110_1010001100101000"; -- 0.013162801063992655
	pesos_i(12681) := b"0000000000000000_0000000000000000_0000100101001001_1101001101000110"; -- 0.03628273455323778
	pesos_i(12682) := b"1111111111111111_1111111111111111_1110111000101001_0110110001111010"; -- -0.06968042401299665
	pesos_i(12683) := b"0000000000000000_0000000000000000_0010000010110000_1000110010101100"; -- 0.1276939314608746
	pesos_i(12684) := b"1111111111111111_1111111111111111_1111010010101001_1001001010011111"; -- -0.04428752526837951
	pesos_i(12685) := b"0000000000000000_0000000000000000_0000000111111101_0110110011111101"; -- 0.0077732197906630225
	pesos_i(12686) := b"1111111111111111_1111111111111111_1110001111000110_1100101101010000"; -- -0.11024789142232361
	pesos_i(12687) := b"1111111111111111_1111111111111111_1110000001101101_0110101011011111"; -- -0.12333042194522399
	pesos_i(12688) := b"0000000000000000_0000000000000000_0010000111001111_1100110010000001"; -- 0.13207700883023668
	pesos_i(12689) := b"0000000000000000_0000000000000000_0001010111100101_0001110111110111"; -- 0.08552729870399707
	pesos_i(12690) := b"0000000000000000_0000000000000000_0000110010111110_0101110010101110"; -- 0.04977969415962086
	pesos_i(12691) := b"1111111111111111_1111111111111111_1110010010111011_0011100101011101"; -- -0.10651818727023464
	pesos_i(12692) := b"0000000000000000_0000000000000000_0001000100111111_0011000000001000"; -- 0.0673704165482085
	pesos_i(12693) := b"0000000000000000_0000000000000000_0001111010101010_1100101001001101"; -- 0.1197935521050599
	pesos_i(12694) := b"1111111111111111_1111111111111111_1111111111011100_1100110000010000"; -- -0.0005371533696649053
	pesos_i(12695) := b"0000000000000000_0000000000000000_0001101110010111_0101100110101110"; -- 0.10777817251316305
	pesos_i(12696) := b"1111111111111111_1111111111111111_1111001111110110_0100111011001111"; -- -0.04702289063844759
	pesos_i(12697) := b"0000000000000000_0000000000000000_0001000011010011_1001110100010000"; -- 0.06572896605281123
	pesos_i(12698) := b"0000000000000000_0000000000000000_0001110101100000_1000000110001001"; -- 0.11475381466121061
	pesos_i(12699) := b"0000000000000000_0000000000000000_0001101010001011_1111001110100101"; -- 0.10369799396652112
	pesos_i(12700) := b"1111111111111111_1111111111111111_1110111011011100_1011010011001010"; -- -0.06694479054678525
	pesos_i(12701) := b"1111111111111111_1111111111111111_1111111010101110_1111101111110011"; -- -0.005142453364590575
	pesos_i(12702) := b"0000000000000000_0000000000000000_0001010001101001_0000111011101111"; -- 0.0797280629658522
	pesos_i(12703) := b"0000000000000000_0000000000000000_0001110011101101_1001111010110001"; -- 0.1130007917675088
	pesos_i(12704) := b"1111111111111111_1111111111111111_1111011111111010_0110000011000000"; -- -0.03133578602000612
	pesos_i(12705) := b"1111111111111111_1111111111111111_1110010111111001_0000000110111010"; -- -0.10166920857520373
	pesos_i(12706) := b"1111111111111111_1111111111111111_1110001000111111_1111101110000011"; -- -0.1162112051281002
	pesos_i(12707) := b"0000000000000000_0000000000000000_0000001010010000_1100100000111110"; -- 0.010021701031817456
	pesos_i(12708) := b"1111111111111111_1111111111111111_1111000101001101_0001101110100111"; -- -0.05741717492560957
	pesos_i(12709) := b"0000000000000000_0000000000000000_0010010001111000_1001110110111110"; -- 0.14246545675845845
	pesos_i(12710) := b"1111111111111111_1111111111111111_1110011101100111_0001100010111001"; -- -0.09608312112796584
	pesos_i(12711) := b"0000000000000000_0000000000000000_0001101111000110_0111101001010000"; -- 0.10849728072006593
	pesos_i(12712) := b"1111111111111111_1111111111111111_1111001110000001_1100000010001010"; -- -0.04880139003601906
	pesos_i(12713) := b"1111111111111111_1111111111111111_1101111010100110_0001100101001100"; -- -0.1302780332271248
	pesos_i(12714) := b"0000000000000000_0000000000000000_0001110011111100_1000011000011011"; -- 0.11322820807757593
	pesos_i(12715) := b"0000000000000000_0000000000000000_0001010000110001_1100000010001011"; -- 0.07888415701531842
	pesos_i(12716) := b"0000000000000000_0000000000000000_0010010100101100_1110111110000001"; -- 0.14521691230683448
	pesos_i(12717) := b"1111111111111111_1111111111111111_1110001110101001_1110001000110000"; -- -0.11068903293517168
	pesos_i(12718) := b"1111111111111111_1111111111111111_1110001101000110_0010101010010111"; -- -0.11221059613686135
	pesos_i(12719) := b"1111111111111111_1111111111111111_1110111000110101_1110011110111100"; -- -0.0694899717944305
	pesos_i(12720) := b"0000000000000000_0000000000000000_0001011001101101_1110011110111101"; -- 0.08761452075581729
	pesos_i(12721) := b"1111111111111111_1111111111111111_1110111000001001_0010100100110000"; -- -0.07017271583937225
	pesos_i(12722) := b"0000000000000000_0000000000000000_0000101000011000_1001001000001111"; -- 0.0394374167195502
	pesos_i(12723) := b"0000000000000000_0000000000000000_0000111000010100_0101000110100010"; -- 0.05499754140276022
	pesos_i(12724) := b"0000000000000000_0000000000000000_0001101001100110_1001100111010100"; -- 0.10312806545704979
	pesos_i(12725) := b"1111111111111111_1111111111111111_1111011110111001_1001111010000000"; -- -0.032323926698279916
	pesos_i(12726) := b"0000000000000000_0000000000000000_0010000010110000_0000001101110010"; -- 0.12768575230820076
	pesos_i(12727) := b"1111111111111111_1111111111111111_1101111101100011_0010000101101100"; -- -0.1273936377228227
	pesos_i(12728) := b"1111111111111111_1111111111111111_1111100110111001_1101101010110010"; -- -0.024507838825613415
	pesos_i(12729) := b"0000000000000000_0000000000000000_0000011000100101_1111000111100101"; -- 0.024016493271585046
	pesos_i(12730) := b"1111111111111111_1111111111111111_1111011011100001_1100101010010110"; -- -0.03561719751200554
	pesos_i(12731) := b"0000000000000000_0000000000000000_0001010000111000_0111101000001111"; -- 0.07898676749825755
	pesos_i(12732) := b"1111111111111111_1111111111111111_1111101110011111_0111101001100010"; -- -0.017097808047684963
	pesos_i(12733) := b"0000000000000000_0000000000000000_0001011010001101_1100000110100101"; -- 0.08810053133546122
	pesos_i(12734) := b"1111111111111111_1111111111111111_1111011101110010_1111010110011101"; -- -0.03340210846346162
	pesos_i(12735) := b"0000000000000000_0000000000000000_0001111101100001_1110101001100010"; -- 0.12258782281439595
	pesos_i(12736) := b"0000000000000000_0000000000000000_0000111010110000_0011010011010110"; -- 0.057376196213870065
	pesos_i(12737) := b"1111111111111111_1111111111111111_1101111011000101_0000010110001110"; -- -0.1298061874509198
	pesos_i(12738) := b"0000000000000000_0000000000000000_0001110000011011_1111010000100100"; -- 0.10980153923422852
	pesos_i(12739) := b"0000000000000000_0000000000000000_0001000000001100_0011110010100111"; -- 0.06268672055365629
	pesos_i(12740) := b"0000000000000000_0000000000000000_0000110010101010_1100010000000001"; -- 0.04948067689576751
	pesos_i(12741) := b"0000000000000000_0000000000000000_0001000000001011_0010001010110000"; -- 0.06266991428845929
	pesos_i(12742) := b"1111111111111111_1111111111111111_1110011100011100_0110101101110111"; -- -0.0972225985083581
	pesos_i(12743) := b"1111111111111111_1111111111111111_1110010011011010_0011001111101011"; -- -0.10604548935618521
	pesos_i(12744) := b"0000000000000000_0000000000000000_0001110101100011_1010010011101111"; -- 0.1148017009676322
	pesos_i(12745) := b"0000000000000000_0000000000000000_0001011000011010_0101101111011001"; -- 0.08633970303380932
	pesos_i(12746) := b"1111111111111111_1111111111111111_1111110010000000_1110010011101011"; -- -0.01365823054004708
	pesos_i(12747) := b"0000000000000000_0000000000000000_0010001011101010_0111110111111010"; -- 0.1363905655339944
	pesos_i(12748) := b"0000000000000000_0000000000000000_0000010110100011_0000110000001100"; -- 0.02201915060386156
	pesos_i(12749) := b"1111111111111111_1111111111111111_1110111001110001_1000110000000110"; -- -0.06857991075891283
	pesos_i(12750) := b"1111111111111111_1111111111111111_1110001010000100_0100011101101001"; -- -0.11516908337331608
	pesos_i(12751) := b"1111111111111111_1111111111111111_1110010101111100_1101010101011011"; -- -0.10356394323494165
	pesos_i(12752) := b"0000000000000000_0000000000000000_0001110001000010_0100011011001110"; -- 0.11038630037443409
	pesos_i(12753) := b"1111111111111111_1111111111111111_1110111100100001_0100111000011111"; -- -0.0658980535741072
	pesos_i(12754) := b"1111111111111111_1111111111111111_1110010110001011_1100011010100100"; -- -0.1033359383437046
	pesos_i(12755) := b"0000000000000000_0000000000000000_0001100101100010_0000001000110001"; -- 0.09915174187577525
	pesos_i(12756) := b"1111111111111111_1111111111111111_1110001001001011_0001100110111100"; -- -0.11604155685926942
	pesos_i(12757) := b"1111111111111111_1111111111111111_1111011011100000_0000001100100100"; -- -0.035644344076028726
	pesos_i(12758) := b"0000000000000000_0000000000000000_0001100011110010_1101100111111110"; -- 0.09745562018489691
	pesos_i(12759) := b"1111111111111111_1111111111111111_1110101011101110_1011101011101000"; -- -0.08229476762851551
	pesos_i(12760) := b"0000000000000000_0000000000000000_0010001001101111_1110110111111101"; -- 0.13452041072132323
	pesos_i(12761) := b"0000000000000000_0000000000000000_0001101101010011_1111110010011101"; -- 0.10675028632061434
	pesos_i(12762) := b"0000000000000000_0000000000000000_0001000001101100_0110100010110000"; -- 0.06415418900942085
	pesos_i(12763) := b"0000000000000000_0000000000000000_0000011011001111_0111100100010111"; -- 0.026603286966820017
	pesos_i(12764) := b"0000000000000000_0000000000000000_0001110001111110_0101011101001011"; -- 0.11130281052945523
	pesos_i(12765) := b"1111111111111111_1111111111111111_1101110000111011_0110001010011000"; -- -0.13971885472584447
	pesos_i(12766) := b"0000000000000000_0000000000000000_0001001101110010_1011011011001000"; -- 0.07596914659110376
	pesos_i(12767) := b"1111111111111111_1111111111111111_1111101110000010_0001011111011011"; -- -0.01754618560963344
	pesos_i(12768) := b"1111111111111111_1111111111111111_1111111001010011_0011010110101011"; -- -0.006542821569099658
	pesos_i(12769) := b"1111111111111111_1111111111111111_1110001000100110_0011100000010001"; -- -0.11660432411530561
	pesos_i(12770) := b"1111111111111111_1111111111111111_1111010000101000_1111011100000110"; -- -0.046249924768392035
	pesos_i(12771) := b"1111111111111111_1111111111111111_1110011010101111_1011001001000001"; -- -0.09888158725317996
	pesos_i(12772) := b"0000000000000000_0000000000000000_0001011100001011_0000000100110111"; -- 0.09001166914940828
	pesos_i(12773) := b"0000000000000000_0000000000000000_0000101100100000_1011100100000011"; -- 0.043468058702765655
	pesos_i(12774) := b"1111111111111111_1111111111111111_1111101000110101_0011101101101000"; -- -0.02262524326326018
	pesos_i(12775) := b"1111111111111111_1111111111111111_1101111010101001_0100110010100111"; -- -0.1302291958956141
	pesos_i(12776) := b"0000000000000000_0000000000000000_0000010100011000_0111011100100110"; -- 0.019904562762471607
	pesos_i(12777) := b"0000000000000000_0000000000000000_0000001100001111_1100000000001011"; -- 0.011959078448052494
	pesos_i(12778) := b"0000000000000000_0000000000000000_0000101001000001_0111101000100001"; -- 0.04006160071718306
	pesos_i(12779) := b"1111111111111111_1111111111111111_1111111011011001_0000100110010000"; -- -0.004500772892656405
	pesos_i(12780) := b"1111111111111111_1111111111111111_1111010100000011_0111001001101111"; -- -0.0429161528986094
	pesos_i(12781) := b"1111111111111111_1111111111111111_1111111010100010_1110100001100000"; -- -0.005326725614432888
	pesos_i(12782) := b"1111111111111111_1111111111111111_1111000111011011_0111101011011000"; -- -0.055244753075316476
	pesos_i(12783) := b"0000000000000000_0000000000000000_0000011010110010_1010011101101011"; -- 0.026163543298312057
	pesos_i(12784) := b"0000000000000000_0000000000000000_0001100000101010_1000101000101101"; -- 0.09439910517221545
	pesos_i(12785) := b"0000000000000000_0000000000000000_0000010000110111_0101100000111000"; -- 0.016469491674073126
	pesos_i(12786) := b"1111111111111111_1111111111111111_1101111001000100_1110111100110001"; -- -0.13176064532676288
	pesos_i(12787) := b"0000000000000000_0000000000000000_0000110111011000_0011010001100101"; -- 0.05408027137369185
	pesos_i(12788) := b"0000000000000000_0000000000000000_0001110010111100_1001100010001110"; -- 0.11225274540082568
	pesos_i(12789) := b"0000000000000000_0000000000000000_0001100010011111_0011111101110111"; -- 0.0961799302101146
	pesos_i(12790) := b"0000000000000000_0000000000000000_0000100000111000_1011111101001001"; -- 0.032115893677130386
	pesos_i(12791) := b"0000000000000000_0000000000000000_0000111001001111_1011001011110110"; -- 0.05590361118918394
	pesos_i(12792) := b"1111111111111111_1111111111111111_1111000111111011_1000101101111100"; -- -0.054755479959910244
	pesos_i(12793) := b"0000000000000000_0000000000000000_0000101101000110_0101111010101011"; -- 0.044042507980250514
	pesos_i(12794) := b"0000000000000000_0000000000000000_0010010000001101_0110110000001000"; -- 0.1408298034073168
	pesos_i(12795) := b"0000000000000000_0000000000000000_0000001010110010_0101100101110010"; -- 0.0105338958516232
	pesos_i(12796) := b"0000000000000000_0000000000000000_0000101110101001_0011111110000110"; -- 0.04555127158453306
	pesos_i(12797) := b"0000000000000000_0000000000000000_0000011010011010_0011000000100010"; -- 0.025790222501200392
	pesos_i(12798) := b"1111111111111111_1111111111111111_1111000000101000_0111110110111100"; -- -0.06188215398763199
	pesos_i(12799) := b"0000000000000000_0000000000000000_0000101011010110_1110101011011110"; -- 0.042341880021565234
	pesos_i(12800) := b"0000000000000000_0000000000000000_0000111011111001_0110010100100101"; -- 0.05849296719664531
	pesos_i(12801) := b"0000000000000000_0000000000000000_0010000110110101_1001011101101011"; -- 0.13167711606469287
	pesos_i(12802) := b"1111111111111111_1111111111111111_1101100000101110_0110100011111000"; -- -0.15554183919318637
	pesos_i(12803) := b"0000000000000000_0000000000000000_0000111100100000_0101111000000000"; -- 0.05908763413047434
	pesos_i(12804) := b"1111111111111111_1111111111111111_1110001100011000_1110101000010010"; -- -0.11290108738230008
	pesos_i(12805) := b"1111111111111111_1111111111111111_1111000011000000_0010111110100011"; -- -0.05956747303652278
	pesos_i(12806) := b"1111111111111111_1111111111111111_1111011000110011_1011000101111010"; -- -0.038273723417289685
	pesos_i(12807) := b"1111111111111111_1111111111111111_1111011000100100_0100100001111000"; -- -0.038508864125363466
	pesos_i(12808) := b"0000000000000000_0000000000000000_0000001001100101_0010111100110110"; -- 0.009356451681747991
	pesos_i(12809) := b"0000000000000000_0000000000000000_0000001001110101_1000011110100001"; -- 0.009605862507814563
	pesos_i(12810) := b"1111111111111111_1111111111111111_1110101000111010_0111111001111111"; -- -0.0850449505130248
	pesos_i(12811) := b"1111111111111111_1111111111111111_1110100010011010_0011111111010101"; -- -0.09139634190565442
	pesos_i(12812) := b"0000000000000000_0000000000000000_0001101000010011_1110110111000011"; -- 0.1018665885786333
	pesos_i(12813) := b"0000000000000000_0000000000000000_0010000001101001_0110010111101010"; -- 0.12660824742420995
	pesos_i(12814) := b"1111111111111111_1111111111111111_1111100101011000_0111010000110001"; -- -0.025994050971674298
	pesos_i(12815) := b"1111111111111111_1111111111111111_1101011111101010_1100100100000101"; -- -0.15657371166917788
	pesos_i(12816) := b"1111111111111111_1111111111111111_1101101100101011_0010101001001001"; -- -0.14387260157878837
	pesos_i(12817) := b"1111111111111111_1111111111111111_1110010110110100_1111000000010110"; -- -0.10270785764688821
	pesos_i(12818) := b"0000000000000000_0000000000000000_0010000001000101_0101011101100100"; -- 0.12605806526651825
	pesos_i(12819) := b"0000000000000000_0000000000000000_0000111110100010_0011110011011110"; -- 0.06106930188205131
	pesos_i(12820) := b"0000000000000000_0000000000000000_0000110101001111_0010100010000111"; -- 0.05198911002316153
	pesos_i(12821) := b"1111111111111111_1111111111111111_1101110100001001_0011011011010111"; -- -0.13657815223480843
	pesos_i(12822) := b"0000000000000000_0000000000000000_0010101011011110_1011010011001000"; -- 0.16746072656348593
	pesos_i(12823) := b"1111111111111111_1111111111111111_1101111100101011_1101100001110100"; -- -0.12823722046244304
	pesos_i(12824) := b"0000000000000000_0000000000000000_0000100111111101_1011110110110101"; -- 0.03902803109343172
	pesos_i(12825) := b"1111111111111111_1111111111111111_1111010000110101_0011010000111001"; -- -0.046063171511113755
	pesos_i(12826) := b"0000000000000000_0000000000000000_0001110000011001_1111100101101101"; -- 0.10977133667434884
	pesos_i(12827) := b"0000000000000000_0000000000000000_0001100110100011_0011001000001101"; -- 0.10014641594356358
	pesos_i(12828) := b"0000000000000000_0000000000000000_0000100110000000_1111110011011011"; -- 0.03712444627087847
	pesos_i(12829) := b"0000000000000000_0000000000000000_0001000010111101_0010011010110100"; -- 0.06538621804806563
	pesos_i(12830) := b"1111111111111111_1111111111111111_1111111011011011_0000100110111000"; -- -0.004470245904884424
	pesos_i(12831) := b"0000000000000000_0000000000000000_0000011011110000_0011001010010010"; -- 0.02710262364795589
	pesos_i(12832) := b"0000000000000000_0000000000000000_0001000001111001_1001010101000111"; -- 0.06435521117107955
	pesos_i(12833) := b"1111111111111111_1111111111111111_1110011101010000_0010011100111010"; -- -0.09643320889564472
	pesos_i(12834) := b"0000000000000000_0000000000000000_0010010100010101_0001111001110011"; -- 0.14485349947210122
	pesos_i(12835) := b"1111111111111111_1111111111111111_1110110011010110_1100001010101111"; -- -0.0748480151390455
	pesos_i(12836) := b"0000000000000000_0000000000000000_0000100010111111_0101100011110010"; -- 0.034169730288849696
	pesos_i(12837) := b"1111111111111111_1111111111111111_1111001111001011_0111111011011011"; -- -0.047676154741772
	pesos_i(12838) := b"0000000000000000_0000000000000000_0000101001001001_0010110110000111"; -- 0.04017910528549373
	pesos_i(12839) := b"1111111111111111_1111111111111111_1111101100011111_0000110010000101"; -- -0.019057481419923725
	pesos_i(12840) := b"0000000000000000_0000000000000000_0000111001001110_0111110101111111"; -- 0.055885165790358834
	pesos_i(12841) := b"0000000000000000_0000000000000000_0000011011100101_1111011100010010"; -- 0.02694648929037016
	pesos_i(12842) := b"0000000000000000_0000000000000000_0001001010000011_1111101011111001"; -- 0.07232636059213175
	pesos_i(12843) := b"0000000000000000_0000000000000000_0000101100001101_0001101010011100"; -- 0.0431687003942535
	pesos_i(12844) := b"0000000000000000_0000000000000000_0001100100111010_0001110000011111"; -- 0.0985429359493156
	pesos_i(12845) := b"1111111111111111_1111111111111111_1110111000010101_0100010010000111"; -- -0.06998798095568669
	pesos_i(12846) := b"0000000000000000_0000000000000000_0001110111100011_0010110011110010"; -- 0.11674767416570966
	pesos_i(12847) := b"0000000000000000_0000000000000000_0010011100010110_0110110011000111"; -- 0.15268592691195207
	pesos_i(12848) := b"1111111111111111_1111111111111111_1110000110111010_0011001010101011"; -- -0.11825259516080434
	pesos_i(12849) := b"1111111111111111_1111111111111111_1110010100100000_0000110101011111"; -- -0.10497967185367571
	pesos_i(12850) := b"1111111111111111_1111111111111111_1111000111100000_0101100000101010"; -- -0.05517052623161917
	pesos_i(12851) := b"1111111111111111_1111111111111111_1110000011000010_1001110010101110"; -- -0.12203045615721174
	pesos_i(12852) := b"1111111111111111_1111111111111111_1101110111100110_0000110101101101"; -- -0.13320842838224087
	pesos_i(12853) := b"0000000000000000_0000000000000000_0001100100101111_0011101110101111"; -- 0.09837697041393922
	pesos_i(12854) := b"0000000000000000_0000000000000000_0001110100111100_1100000110110001"; -- 0.11420832220661695
	pesos_i(12855) := b"1111111111111111_1111111111111111_1110001011010001_1000001011000111"; -- -0.11399061819089336
	pesos_i(12856) := b"0000000000000000_0000000000000000_0001011110010111_1010111110011101"; -- 0.09215829457251311
	pesos_i(12857) := b"1111111111111111_1111111111111111_1111001010011100_1110010110110100"; -- -0.0522934374347788
	pesos_i(12858) := b"0000000000000000_0000000000000000_0001000100100011_1100000111110001"; -- 0.06695186735709009
	pesos_i(12859) := b"0000000000000000_0000000000000000_0000100011010110_0000001000001110"; -- 0.03451550343810574
	pesos_i(12860) := b"1111111111111111_1111111111111111_1110001100000010_1110001110010101"; -- -0.11323716749783627
	pesos_i(12861) := b"1111111111111111_1111111111111111_1111111011111011_0100111101000110"; -- -0.003977818795143632
	pesos_i(12862) := b"1111111111111111_1111111111111111_1110110110000000_0110101010011101"; -- -0.07225927037310731
	pesos_i(12863) := b"0000000000000000_0000000000000000_0001011001001011_0011011001011000"; -- 0.0870851483743514
	pesos_i(12864) := b"1111111111111111_1111111111111111_1111111100100011_1100000000100000"; -- -0.003360740883094351
	pesos_i(12865) := b"0000000000000000_0000000000000000_0000100100000101_0000011000101100"; -- 0.03523291171551689
	pesos_i(12866) := b"0000000000000000_0000000000000000_0000100111100010_0011111100000100"; -- 0.03860849234725682
	pesos_i(12867) := b"1111111111111111_1111111111111111_1111101000101011_1001111111111010"; -- -0.022771836767444296
	pesos_i(12868) := b"0000000000000000_0000000000000000_0000001000000101_1010110101100000"; -- 0.007899127963626395
	pesos_i(12869) := b"1111111111111111_1111111111111111_1110110001111111_1101100000010100"; -- -0.07617425443774051
	pesos_i(12870) := b"0000000000000000_0000000000000000_0000000001001100_0111000100101110"; -- 0.0011664140910401142
	pesos_i(12871) := b"1111111111111111_1111111111111111_1111111101010001_0000101101111100"; -- -0.0026696036766534247
	pesos_i(12872) := b"1111111111111111_1111111111111111_1110001000101001_0001111010111100"; -- -0.11656005762557363
	pesos_i(12873) := b"0000000000000000_0000000000000000_0000011011001001_0111100101000100"; -- 0.02651174453597552
	pesos_i(12874) := b"0000000000000000_0000000000000000_0001000100100010_0111010001011001"; -- 0.06693198377219998
	pesos_i(12875) := b"0000000000000000_0000000000000000_0001000000101010_0000011100100101"; -- 0.06314129495305243
	pesos_i(12876) := b"1111111111111111_1111111111111111_1110001001011111_0011110101011001"; -- -0.11573425850863159
	pesos_i(12877) := b"1111111111111111_1111111111111111_1111010011100100_0110001100100010"; -- -0.043390087297423274
	pesos_i(12878) := b"0000000000000000_0000000000000000_0010001101110001_0111000011100100"; -- 0.1384497219327634
	pesos_i(12879) := b"1111111111111111_1111111111111111_1111110110000110_1101000010101101"; -- -0.009661634217915575
	pesos_i(12880) := b"0000000000000000_0000000000000000_0000011010101100_0011111010110110"; -- 0.02606574965189168
	pesos_i(12881) := b"0000000000000000_0000000000000000_0000010000101001_1001001110010110"; -- 0.016259407133787943
	pesos_i(12882) := b"0000000000000000_0000000000000000_0001101100100100_0110000000001110"; -- 0.10602379159904379
	pesos_i(12883) := b"1111111111111111_1111111111111111_1111010101010101_0000110011011001"; -- -0.04167098716298188
	pesos_i(12884) := b"0000000000000000_0000000000000000_0000010011011000_0100011111101000"; -- 0.0189251844745939
	pesos_i(12885) := b"0000000000000000_0000000000000000_0001001001100001_0101010001100111"; -- 0.0717976333184207
	pesos_i(12886) := b"0000000000000000_0000000000000000_0000111100011000_1000111110001001"; -- 0.058968516353337094
	pesos_i(12887) := b"0000000000000000_0000000000000000_0010000001010100_1011001001001101"; -- 0.12629236592083054
	pesos_i(12888) := b"0000000000000000_0000000000000000_0000100010101110_0000010010000111"; -- 0.033905299177147394
	pesos_i(12889) := b"0000000000000000_0000000000000000_0000110111101111_0001111101101101"; -- 0.054429973733461194
	pesos_i(12890) := b"1111111111111111_1111111111111111_1111011101110100_0100010101011000"; -- -0.03338209737166693
	pesos_i(12891) := b"1111111111111111_1111111111111111_1111010100101010_0011111110100001"; -- -0.04232408818807519
	pesos_i(12892) := b"0000000000000000_0000000000000000_0001101001010101_1001000011001111"; -- 0.10286812844862236
	pesos_i(12893) := b"0000000000000000_0000000000000000_0001111011000001_0010111111000100"; -- 0.12013529343203709
	pesos_i(12894) := b"0000000000000000_0000000000000000_0000100101000000_0100101111110010"; -- 0.03613733916635621
	pesos_i(12895) := b"1111111111111111_1111111111111111_1111001110110110_1011101000011110"; -- -0.0479930568931806
	pesos_i(12896) := b"0000000000000000_0000000000000000_0001000000101011_1001011010100100"; -- 0.06316510670821214
	pesos_i(12897) := b"1111111111111111_1111111111111111_1110100010011101_0011010101111000"; -- -0.09135118313075262
	pesos_i(12898) := b"1111111111111111_1111111111111111_1110000100000011_0111011111110000"; -- -0.12104082476327338
	pesos_i(12899) := b"1111111111111111_1111111111111111_1111101100101100_1100000000001001"; -- -0.01884841704609668
	pesos_i(12900) := b"1111111111111111_1111111111111111_1101111101001110_1110010000010101"; -- -0.1277024696723007
	pesos_i(12901) := b"0000000000000000_0000000000000000_0010001011100101_1100001111010101"; -- 0.13631843514023237
	pesos_i(12902) := b"1111111111111111_1111111111111111_1110100110010110_1100001001101100"; -- -0.08754334313721926
	pesos_i(12903) := b"1111111111111111_1111111111111111_1111011011011001_1010110110110011"; -- -0.035740989607003074
	pesos_i(12904) := b"0000000000000000_0000000000000000_0010001101100110_0011110010101110"; -- 0.13827876336706552
	pesos_i(12905) := b"1111111111111111_1111111111111111_1110010100011101_1010011010100010"; -- -0.10501631313773727
	pesos_i(12906) := b"0000000000000000_0000000000000000_0001000111010011_1110101111011101"; -- 0.06963991297906487
	pesos_i(12907) := b"0000000000000000_0000000000000000_0001000011000101_1011001011000010"; -- 0.0655166362555771
	pesos_i(12908) := b"1111111111111111_1111111111111111_1111001110001010_1111111010001010"; -- -0.04866036551271551
	pesos_i(12909) := b"0000000000000000_0000000000000000_0000001110101000_1001001100111101"; -- 0.014291002639213183
	pesos_i(12910) := b"0000000000000000_0000000000000000_0000101110110001_1011011000101111"; -- 0.04568041464336472
	pesos_i(12911) := b"0000000000000000_0000000000000000_0010001010000110_1110111001010011"; -- 0.13487138284843256
	pesos_i(12912) := b"0000000000000000_0000000000000000_0001111011110101_0100110001000101"; -- 0.1209304493755426
	pesos_i(12913) := b"1111111111111111_1111111111111111_1110011100111110_0110110001110100"; -- -0.09670374065434703
	pesos_i(12914) := b"0000000000000000_0000000000000000_0000010001101001_1000010101000001"; -- 0.017235115461274132
	pesos_i(12915) := b"0000000000000000_0000000000000000_0010000111101010_0000001101100111"; -- 0.13247700946135807
	pesos_i(12916) := b"0000000000000000_0000000000000000_0001000000110110_0111100110101110"; -- 0.06333122733530609
	pesos_i(12917) := b"1111111111111111_1111111111111111_1110111111110100_0101000011101011"; -- -0.06267828242157192
	pesos_i(12918) := b"1111111111111111_1111111111111111_1111111011110011_1111111000010101"; -- -0.004089469832086165
	pesos_i(12919) := b"0000000000000000_0000000000000000_0001011110100010_0111001010111111"; -- 0.09232251327047034
	pesos_i(12920) := b"1111111111111111_1111111111111111_1110011000101101_0000010101010000"; -- -0.10087553787959415
	pesos_i(12921) := b"1111111111111111_1111111111111111_1110111011101100_1011001001110111"; -- -0.06670078844004053
	pesos_i(12922) := b"1111111111111111_1111111111111111_1111000101000010_1000100101010110"; -- -0.05757848407245958
	pesos_i(12923) := b"1111111111111111_1111111111111111_1111100010001010_1001111110001101"; -- -0.029134777161052873
	pesos_i(12924) := b"1111111111111111_1111111111111111_1111101010111010_0011001001011010"; -- -0.020596364082946895
	pesos_i(12925) := b"1111111111111111_1111111111111111_1110010010010000_0110110001011010"; -- -0.10717127604918983
	pesos_i(12926) := b"1111111111111111_1111111111111111_1110100110010110_0111100101011011"; -- -0.08754769830942827
	pesos_i(12927) := b"0000000000000000_0000000000000000_0010010010000011_0101101000001101"; -- 0.14262926871722162
	pesos_i(12928) := b"0000000000000000_0000000000000000_0010000010100001_0101100111010101"; -- 0.12746201950726133
	pesos_i(12929) := b"1111111111111111_1111111111111111_1101111101111100_1000000001001010"; -- -0.12700651350214126
	pesos_i(12930) := b"0000000000000000_0000000000000000_0000010011111100_0100100011110000"; -- 0.01947456228436625
	pesos_i(12931) := b"0000000000000000_0000000000000000_0001100010110101_1111101100111100"; -- 0.09652681563099223
	pesos_i(12932) := b"0000000000000000_0000000000000000_0000011000110100_0111000110010110"; -- 0.024237727217253768
	pesos_i(12933) := b"0000000000000000_0000000000000000_0001100101011101_1111011101000011"; -- 0.09909005527925129
	pesos_i(12934) := b"1111111111111111_1111111111111111_1110110000101111_1100011110110111"; -- -0.0773959330266722
	pesos_i(12935) := b"1111111111111111_1111111111111111_1101101010111001_1010111111100101"; -- -0.145604139837228
	pesos_i(12936) := b"1111111111111111_1111111111111111_1111111010110101_0110101001110001"; -- -0.00504431469633383
	pesos_i(12937) := b"0000000000000000_0000000000000000_0010001000000111_0101110111101011"; -- 0.13292490954772807
	pesos_i(12938) := b"1111111111111111_1111111111111111_1101011100000011_1100000011000111"; -- -0.1600989832687459
	pesos_i(12939) := b"1111111111111111_1111111111111111_1111100101001110_1110110011011111"; -- -0.026139445912985747
	pesos_i(12940) := b"0000000000000000_0000000000000000_0010010101000111_1100011000011000"; -- 0.14562643129667677
	pesos_i(12941) := b"1111111111111111_1111111111111111_1110110011111000_1001101110100010"; -- -0.07433154396588741
	pesos_i(12942) := b"1111111111111111_1111111111111111_1101111100110100_0100100111101110"; -- -0.1281083863793837
	pesos_i(12943) := b"1111111111111111_1111111111111111_1110110010001001_1100001100110101"; -- -0.07602291064073508
	pesos_i(12944) := b"0000000000000000_0000000000000000_0000010101111001_1001011101111101"; -- 0.0213865928692126
	pesos_i(12945) := b"1111111111111111_1111111111111111_1111001111111010_1011001111101111"; -- -0.04695582787710797
	pesos_i(12946) := b"0000000000000000_0000000000000000_0001011111000001_1110101000101101"; -- 0.0928026543041487
	pesos_i(12947) := b"1111111111111111_1111111111111111_1110000001001100_0101010100011001"; -- -0.12383525992543014
	pesos_i(12948) := b"1111111111111111_1111111111111111_1111101000011110_0101001010000010"; -- -0.022974818409840107
	pesos_i(12949) := b"1111111111111111_1111111111111111_1110000001010010_1001100101011101"; -- -0.12373963804382368
	pesos_i(12950) := b"1111111111111111_1111111111111111_1101010010100010_1001001011001111"; -- -0.16939432567610843
	pesos_i(12951) := b"1111111111111111_1111111111111111_1101101110100001_0100110010011010"; -- -0.14207001904592434
	pesos_i(12952) := b"1111111111111111_1111111111111111_1111101110110001_0111001001000111"; -- -0.016823632771259114
	pesos_i(12953) := b"0000000000000000_0000000000000000_0000011000100010_0101001110111011"; -- 0.023961289478857145
	pesos_i(12954) := b"0000000000000000_0000000000000000_0000111101110011_0110000100110001"; -- 0.060354303848061994
	pesos_i(12955) := b"1111111111111111_1111111111111111_1110100010011101_0101000000010111"; -- -0.09134959643475356
	pesos_i(12956) := b"1111111111111111_1111111111111111_1111010001100100_0111100100101001"; -- -0.045341899446823895
	pesos_i(12957) := b"0000000000000000_0000000000000000_0010001000110100_0101101110000101"; -- 0.13361141212734473
	pesos_i(12958) := b"1111111111111111_1111111111111111_1110001000001111_0001001111110011"; -- -0.11695742904762278
	pesos_i(12959) := b"0000000000000000_0000000000000000_0001001111111000_0111010101100100"; -- 0.0780099267393119
	pesos_i(12960) := b"1111111111111111_1111111111111111_1111100010100101_1000000000000001"; -- -0.02872467016419498
	pesos_i(12961) := b"0000000000000000_0000000000000000_0000001110110000_0101011110001111"; -- 0.014409515694465849
	pesos_i(12962) := b"1111111111111111_1111111111111111_1101110011111001_0111111011110001"; -- -0.1368179952226224
	pesos_i(12963) := b"0000000000000000_0000000000000000_0000100100101100_1100001101011100"; -- 0.03583928109539708
	pesos_i(12964) := b"1111111111111111_1111111111111111_1110001000100111_1001001100011110"; -- -0.11658363829282851
	pesos_i(12965) := b"1111111111111111_1111111111111111_1111010011100001_1000110010110110"; -- -0.04343338545122665
	pesos_i(12966) := b"0000000000000000_0000000000000000_0001010010101010_0011001100101001"; -- 0.0807220435779883
	pesos_i(12967) := b"0000000000000000_0000000000000000_0001111001101110_0100001001000000"; -- 0.11886991553673162
	pesos_i(12968) := b"0000000000000000_0000000000000000_0000101101100010_0000101111110010"; -- 0.0444648233999921
	pesos_i(12969) := b"1111111111111111_1111111111111111_1110001011010011_0110001011101111"; -- -0.1139619985446044
	pesos_i(12970) := b"1111111111111111_1111111111111111_1111001110101010_0101100000110011"; -- -0.04818199879283994
	pesos_i(12971) := b"0000000000000000_0000000000000000_0000010011000100_0000111011110011"; -- 0.018616613730070692
	pesos_i(12972) := b"0000000000000000_0000000000000000_0000110011011111_1000011001110010"; -- 0.050285723618494635
	pesos_i(12973) := b"0000000000000000_0000000000000000_0001101111010100_1000111100101011"; -- 0.10871214668748906
	pesos_i(12974) := b"1111111111111111_1111111111111111_1110001101011011_0100100000000001"; -- -0.11188840850760476
	pesos_i(12975) := b"1111111111111111_1111111111111111_1110111101011011_0001010111000000"; -- -0.06501640387261193
	pesos_i(12976) := b"0000000000000000_0000000000000000_0000111011100001_1100101101100001"; -- 0.058132849975213036
	pesos_i(12977) := b"0000000000000000_0000000000000000_0001010010100000_1110110110101110"; -- 0.08058057298789492
	pesos_i(12978) := b"1111111111111111_1111111111111111_1111001101110111_1011110000010111"; -- -0.04895424298539703
	pesos_i(12979) := b"1111111111111111_1111111111111111_1111100000010000_0110011000100111"; -- -0.030999770700092643
	pesos_i(12980) := b"1111111111111111_1111111111111111_1110011110001101_1101100100001100"; -- -0.09549182385120329
	pesos_i(12981) := b"1111111111111111_1111111111111111_1111011100110001_1100101100010101"; -- -0.03439646460141469
	pesos_i(12982) := b"1111111111111111_1111111111111111_1101110001101011_1100100010001110"; -- -0.13898035558722452
	pesos_i(12983) := b"0000000000000000_0000000000000000_0000000010011011_0101000000100010"; -- 0.002369888637757154
	pesos_i(12984) := b"1111111111111111_1111111111111111_1111000100111011_0000011110111000"; -- -0.05769302148726491
	pesos_i(12985) := b"1111111111111111_1111111111111111_1111011001000111_0111000110110100"; -- -0.03797234883676287
	pesos_i(12986) := b"0000000000000000_0000000000000000_0000111101101100_1110110000000001"; -- 0.06025576607099689
	pesos_i(12987) := b"0000000000000000_0000000000000000_0000001101100110_1011010100010111"; -- 0.01328594031527844
	pesos_i(12988) := b"0000000000000000_0000000000000000_0000111010001010_1100000010111101"; -- 0.05680470096382091
	pesos_i(12989) := b"1111111111111111_1111111111111111_1111000000100110_0010011000101101"; -- -0.061917890531956336
	pesos_i(12990) := b"0000000000000000_0000000000000000_0010000110101101_0101101110011001"; -- 0.13155148024265606
	pesos_i(12991) := b"0000000000000000_0000000000000000_0001011000110010_1001100010010010"; -- 0.08670953345596696
	pesos_i(12992) := b"1111111111111111_1111111111111111_1110001111101000_0010000100110000"; -- -0.10973923278719788
	pesos_i(12993) := b"0000000000000000_0000000000000000_0001110011100011_0100000110010100"; -- 0.11284265389616882
	pesos_i(12994) := b"0000000000000000_0000000000000000_0010001110101011_0111110100011111"; -- 0.13933546077114706
	pesos_i(12995) := b"0000000000000000_0000000000000000_0001111010110011_0011101110100001"; -- 0.11992237732223808
	pesos_i(12996) := b"0000000000000000_0000000000000000_0000000010010111_1001100110111101"; -- 0.0023132406641645075
	pesos_i(12997) := b"1111111111111111_1111111111111111_1111111001000101_0000111101001110"; -- -0.006758731404404717
	pesos_i(12998) := b"0000000000000000_0000000000000000_0000110011011110_0011011011100110"; -- 0.0502657234706088
	pesos_i(12999) := b"0000000000000000_0000000000000000_0000110000101010_1110111101110011"; -- 0.047530141411604526
	pesos_i(13000) := b"0000000000000000_0000000000000000_0001011101101010_1110110110010000"; -- 0.09147534144008491
	pesos_i(13001) := b"1111111111111111_1111111111111111_1111010000010110_0100101101011100"; -- -0.04653481486890552
	pesos_i(13002) := b"0000000000000000_0000000000000000_0000000011010010_1110001110101011"; -- 0.003217915747345288
	pesos_i(13003) := b"0000000000000000_0000000000000000_0001011100111001_1001100100001110"; -- 0.0907226238010489
	pesos_i(13004) := b"1111111111111111_1111111111111111_1110111110100011_1000010011111000"; -- -0.06391114177468789
	pesos_i(13005) := b"0000000000000000_0000000000000000_0000000000011010_0111000011111111"; -- 0.0004034636118229944
	pesos_i(13006) := b"0000000000000000_0000000000000000_0001000000100000_0010110111001000"; -- 0.06299100996336406
	pesos_i(13007) := b"0000000000000000_0000000000000000_0010011101001100_1111111000011011"; -- 0.15351856374452716
	pesos_i(13008) := b"0000000000000000_0000000000000000_0001100110000101_1011010000100101"; -- 0.099696406426595
	pesos_i(13009) := b"1111111111111111_1111111111111111_1110000111001010_1001010001011101"; -- -0.11800263146246086
	pesos_i(13010) := b"0000000000000000_0000000000000000_0000010000000001_0100101000000001"; -- 0.015644669804749198
	pesos_i(13011) := b"1111111111111111_1111111111111111_1111001100010101_0011010000110010"; -- -0.050457704292562654
	pesos_i(13012) := b"1111111111111111_1111111111111111_1101111100101100_1010001101110000"; -- -0.1282251216567398
	pesos_i(13013) := b"1111111111111111_1111111111111111_1110110010111001_0111110101011001"; -- -0.07529465266055041
	pesos_i(13014) := b"0000000000000000_0000000000000000_0001111011011111_0110011110001001"; -- 0.12059638112499003
	pesos_i(13015) := b"0000000000000000_0000000000000000_0001010101010100_0010000000001101"; -- 0.08331489855108483
	pesos_i(13016) := b"0000000000000000_0000000000000000_0000100110110010_0001110101011111"; -- 0.037874065033708305
	pesos_i(13017) := b"1111111111111111_1111111111111111_1111000010111111_1110011110101010"; -- -0.05957176303851701
	pesos_i(13018) := b"0000000000000000_0000000000000000_0010001011000000_0110010110110110"; -- 0.13574824988207146
	pesos_i(13019) := b"0000000000000000_0000000000000000_0000111110110010_0110110010111011"; -- 0.06131629533490797
	pesos_i(13020) := b"0000000000000000_0000000000000000_0001011111001011_1111111101100111"; -- 0.09295650738183202
	pesos_i(13021) := b"0000000000000000_0000000000000000_0000010000101000_1100000111110011"; -- 0.016246911756134734
	pesos_i(13022) := b"0000000000000000_0000000000000000_0001000010100100_0111111001100111"; -- 0.06500997555490805
	pesos_i(13023) := b"0000000000000000_0000000000000000_0001011000011000_0000011010001000"; -- 0.0863041003313726
	pesos_i(13024) := b"0000000000000000_0000000000000000_0000000111001001_1000011001101010"; -- 0.006981278205074879
	pesos_i(13025) := b"1111111111111111_1111111111111111_1110000000011011_1000000101000011"; -- -0.12458030804067753
	pesos_i(13026) := b"0000000000000000_0000000000000000_0000010011010001_1110100111000101"; -- 0.01882802076424292
	pesos_i(13027) := b"1111111111111111_1111111111111111_1110110110001010_1001001010101101"; -- -0.07210429451230697
	pesos_i(13028) := b"1111111111111111_1111111111111111_1110010100111110_1000111101010110"; -- -0.10451416160793958
	pesos_i(13029) := b"0000000000000000_0000000000000000_0001000111010101_1100100111110001"; -- 0.0696684087713046
	pesos_i(13030) := b"1111111111111111_1111111111111111_1111010111100010_1101011111100110"; -- -0.03950739503897016
	pesos_i(13031) := b"1111111111111111_1111111111111111_1101111011110010_0001101010100010"; -- -0.12911828559951571
	pesos_i(13032) := b"1111111111111111_1111111111111111_1111100111011111_1001000100001010"; -- -0.02393239498938427
	pesos_i(13033) := b"0000000000000000_0000000000000000_0001000111011100_1001100110111101"; -- 0.06977234701010669
	pesos_i(13034) := b"0000000000000000_0000000000000000_0000111000000001_1001110111100101"; -- 0.054712170099194636
	pesos_i(13035) := b"1111111111111111_1111111111111111_1111010111011111_0110101000111010"; -- -0.039559708487072284
	pesos_i(13036) := b"0000000000000000_0000000000000000_0001111111010111_1010001100111001"; -- 0.12438411850604425
	pesos_i(13037) := b"1111111111111111_1111111111111111_1110001110011001_0011100111000011"; -- -0.11094321232031726
	pesos_i(13038) := b"0000000000000000_0000000000000000_0001111111101110_1111011000100011"; -- 0.12474001263171383
	pesos_i(13039) := b"0000000000000000_0000000000000000_0000101001001000_1001111001111110"; -- 0.04017057962784503
	pesos_i(13040) := b"0000000000000000_0000000000000000_0000010100010001_0000100100010100"; -- 0.01979119059140302
	pesos_i(13041) := b"1111111111111111_1111111111111111_1110010111100110_0110001101110001"; -- -0.10195330130165955
	pesos_i(13042) := b"0000000000000000_0000000000000000_0000010011101010_1011001111110100"; -- 0.019206282760911724
	pesos_i(13043) := b"0000000000000000_0000000000000000_0010010010000110_1110100000111111"; -- 0.1426835207462939
	pesos_i(13044) := b"1111111111111111_1111111111111111_1111000101000000_0000010000111110"; -- -0.05761693462670657
	pesos_i(13045) := b"0000000000000000_0000000000000000_0000110111011010_0000000111001100"; -- 0.05410777316456094
	pesos_i(13046) := b"0000000000000000_0000000000000000_0001011110100100_0001000100000010"; -- 0.09234720515706397
	pesos_i(13047) := b"1111111111111111_1111111111111111_1110010001001100_0011100010010111"; -- -0.10821195905220393
	pesos_i(13048) := b"1111111111111111_1111111111111111_1110101011101100_0001100111111000"; -- -0.08233487801412143
	pesos_i(13049) := b"0000000000000000_0000000000000000_0000001000100011_1010011001001001"; -- 0.008356469076265909
	pesos_i(13050) := b"1111111111111111_1111111111111111_1110100001111001_1101111100010001"; -- -0.09189039071166809
	pesos_i(13051) := b"0000000000000000_0000000000000000_0000111100111001_0001110001000101"; -- 0.05946518589918185
	pesos_i(13052) := b"1111111111111111_1111111111111111_1110110001111011_0010111011111011"; -- -0.07624536860874628
	pesos_i(13053) := b"0000000000000000_0000000000000000_0001000011010000_1110011010111010"; -- 0.06568758061009276
	pesos_i(13054) := b"1111111111111111_1111111111111111_1111010000101001_0000010100000100"; -- -0.04624909077623901
	pesos_i(13055) := b"0000000000000000_0000000000000000_0010011001001001_1111011011010101"; -- 0.14956610388024535
	pesos_i(13056) := b"0000000000000000_0000000000000000_0001111101001001_1110100001110101"; -- 0.12222149707791953
	pesos_i(13057) := b"0000000000000000_0000000000000000_0000110101000100_0011001111011000"; -- 0.05182193770626356
	pesos_i(13058) := b"1111111111111111_1111111111111111_1101111111110011_1110010111110111"; -- -0.12518465732468623
	pesos_i(13059) := b"1111111111111111_1111111111111111_1111100010010000_1111100110110001"; -- -0.029037851706841068
	pesos_i(13060) := b"0000000000000000_0000000000000000_0000100010110110_0101010010000000"; -- 0.034032136206560565
	pesos_i(13061) := b"0000000000000000_0000000000000000_0001111001111010_0000110010011101"; -- 0.11904982401143537
	pesos_i(13062) := b"1111111111111111_1111111111111111_1111001001011101_1110111011100001"; -- -0.05325419426437027
	pesos_i(13063) := b"0000000000000000_0000000000000000_0010001101111000_0101010100000111"; -- 0.13855487268999067
	pesos_i(13064) := b"0000000000000000_0000000000000000_0001100010110010_1001110100111010"; -- 0.09647543578688964
	pesos_i(13065) := b"0000000000000000_0000000000000000_0001001110110011_0001011000100011"; -- 0.07695139275948802
	pesos_i(13066) := b"0000000000000000_0000000000000000_0001100111001000_0000011001011110"; -- 0.10070838722451347
	pesos_i(13067) := b"1111111111111111_1111111111111111_1111110001011100_0010000110100000"; -- -0.014219187256561365
	pesos_i(13068) := b"0000000000000000_0000000000000000_0010001011000110_1101111110011111"; -- 0.13584706906910493
	pesos_i(13069) := b"1111111111111111_1111111111111111_1111111011011000_0100001011111001"; -- -0.004512609750539709
	pesos_i(13070) := b"0000000000000000_0000000000000000_0001001010001001_1010110011010101"; -- 0.0724132555796931
	pesos_i(13071) := b"1111111111111111_1111111111111111_1110100101010010_0111000110011100"; -- -0.08858575760539113
	pesos_i(13072) := b"1111111111111111_1111111111111111_1110000001100100_1011011010010011"; -- -0.12346323877498047
	pesos_i(13073) := b"0000000000000000_0000000000000000_0000111111010001_1001110110001010"; -- 0.0617922269698216
	pesos_i(13074) := b"1111111111111111_1111111111111111_1111111010100010_0111101110011101"; -- -0.005333208155489971
	pesos_i(13075) := b"1111111111111111_1111111111111111_1101101001100110_0111110000111011"; -- -0.1468736988279905
	pesos_i(13076) := b"0000000000000000_0000000000000000_0000111110010110_1100101111100010"; -- 0.06089472062747545
	pesos_i(13077) := b"0000000000000000_0000000000000000_0010001110111100_1101010101010100"; -- 0.1396001176239184
	pesos_i(13078) := b"1111111111111111_1111111111111111_1111110010101001_0001010100011111"; -- -0.013045005789100578
	pesos_i(13079) := b"1111111111111111_1111111111111111_1110101100010111_0001100110110101"; -- -0.0816787656395158
	pesos_i(13080) := b"1111111111111111_1111111111111111_1110111001000001_0001011000001000"; -- -0.06931936558334419
	pesos_i(13081) := b"1111111111111111_1111111111111111_1101100101000011_1011010001100101"; -- -0.151310658754083
	pesos_i(13082) := b"1111111111111111_1111111111111111_1101101111110000_0010101101000100"; -- -0.14086656176097226
	pesos_i(13083) := b"0000000000000000_0000000000000000_0010010100100011_1110111110101110"; -- 0.1450795936393519
	pesos_i(13084) := b"0000000000000000_0000000000000000_0000010010101100_0111000100101100"; -- 0.018256257315791582
	pesos_i(13085) := b"1111111111111111_1111111111111111_1110110000100111_1011001001011000"; -- -0.07751927706610774
	pesos_i(13086) := b"1111111111111111_1111111111111111_1111011001010010_0111010100011011"; -- -0.03780429934030564
	pesos_i(13087) := b"0000000000000000_0000000000000000_0001011010101101_0001111101010110"; -- 0.08857913837928529
	pesos_i(13088) := b"1111111111111111_1111111111111111_1101110000001010_1010010011100111"; -- -0.14046258325832053
	pesos_i(13089) := b"1111111111111111_1111111111111111_1111000110111000_1101100100111100"; -- -0.05577318453725407
	pesos_i(13090) := b"1111111111111111_1111111111111111_1110100010111101_1000001010110101"; -- -0.09085829817557439
	pesos_i(13091) := b"1111111111111111_1111111111111111_1111101110111101_1101100001011000"; -- -0.0166344438597855
	pesos_i(13092) := b"0000000000000000_0000000000000000_0001101011110101_1001010100011111"; -- 0.10530979173776939
	pesos_i(13093) := b"0000000000000000_0000000000000000_0010000000001100_0111000010011011"; -- 0.12518981720185302
	pesos_i(13094) := b"0000000000000000_0000000000000000_0001101110101000_1000111010001011"; -- 0.10804072281420717
	pesos_i(13095) := b"1111111111111111_1111111111111111_1110001011111001_0111110100100001"; -- -0.11338060336600965
	pesos_i(13096) := b"0000000000000000_0000000000000000_0000111110101100_1011010010010011"; -- 0.061229024669835784
	pesos_i(13097) := b"0000000000000000_0000000000000000_0000000101010011_0011010001000000"; -- 0.005175843881879628
	pesos_i(13098) := b"0000000000000000_0000000000000000_0010110010101100_1111000100101110"; -- 0.17451388708000498
	pesos_i(13099) := b"1111111111111111_1111111111111111_1110111111011010_1111011110010110"; -- -0.06306507667414016
	pesos_i(13100) := b"0000000000000000_0000000000000000_0000101111100110_1010111101001110"; -- 0.04648872054197795
	pesos_i(13101) := b"1111111111111111_1111111111111111_1111100100111111_1001011110010011"; -- -0.026373411774868
	pesos_i(13102) := b"1111111111111111_1111111111111111_1110101000111101_0001101000110101"; -- -0.08500515175751286
	pesos_i(13103) := b"1111111111111111_1111111111111111_1110001100101011_1011111001100100"; -- -0.11261377395946098
	pesos_i(13104) := b"0000000000000000_0000000000000000_0010000010001001_1010111100011110"; -- 0.12710089187325835
	pesos_i(13105) := b"0000000000000000_0000000000000000_0010110010110000_0001010101011110"; -- 0.17456182039165147
	pesos_i(13106) := b"1111111111111111_1111111111111111_1101101001000010_1111111111000101"; -- -0.14741517483875705
	pesos_i(13107) := b"0000000000000000_0000000000000000_0001100110001011_0110011010010100"; -- 0.09978333584279059
	pesos_i(13108) := b"0000000000000000_0000000000000000_0000011010000011_0110101000110010"; -- 0.02544273113464393
	pesos_i(13109) := b"0000000000000000_0000000000000000_0000011110101011_0010111100100001"; -- 0.029955812003955296
	pesos_i(13110) := b"1111111111111111_1111111111111111_1110101001000010_1111000000110010"; -- -0.08491610323286373
	pesos_i(13111) := b"1111111111111111_1111111111111111_1111110111000100_0000100010101011"; -- -0.008727510646907393
	pesos_i(13112) := b"1111111111111111_1111111111111111_1110101100110100_1100110010010000"; -- -0.08122560002586468
	pesos_i(13113) := b"1111111111111111_1111111111111111_1110100011000011_0111101010101100"; -- -0.09076722425878782
	pesos_i(13114) := b"0000000000000000_0000000000000000_0000100101101100_0011010100101100"; -- 0.036807368578228736
	pesos_i(13115) := b"1111111111111111_1111111111111111_1110111000101110_1111110111010111"; -- -0.06959546574131227
	pesos_i(13116) := b"0000000000000000_0000000000000000_0001101000001101_1111001111101010"; -- 0.10177540265527593
	pesos_i(13117) := b"1111111111111111_1111111111111111_1111101001101010_1110100111100010"; -- -0.02180612789029217
	pesos_i(13118) := b"1111111111111111_1111111111111111_1111100101010011_1101011000100101"; -- -0.02606450651961599
	pesos_i(13119) := b"0000000000000000_0000000000000000_0000011101001110_1010001110100101"; -- 0.028543689618248755
	pesos_i(13120) := b"0000000000000000_0000000000000000_0000100001111110_1101101110101111"; -- 0.03318570168588103
	pesos_i(13121) := b"0000000000000000_0000000000000000_0000101011000010_1011010100010101"; -- 0.04203349846363309
	pesos_i(13122) := b"0000000000000000_0000000000000000_0010001100010111_0100101001100011"; -- 0.13707413603157906
	pesos_i(13123) := b"1111111111111111_1111111111111111_1110001001000000_1110001110010100"; -- -0.1161973727351349
	pesos_i(13124) := b"0000000000000000_0000000000000000_0000100001000111_0110100110010110"; -- 0.03233966734311619
	pesos_i(13125) := b"1111111111111111_1111111111111111_1101100001001100_1100000000011111"; -- -0.15507888073809722
	pesos_i(13126) := b"0000000000000000_0000000000000000_0001111111001111_0110001000111100"; -- 0.12425817467394405
	pesos_i(13127) := b"1111111111111111_1111111111111111_1110100010101101_1101101100110101"; -- -0.09109716368774629
	pesos_i(13128) := b"0000000000000000_0000000000000000_0001010111010000_0110100011100101"; -- 0.08521133027517869
	pesos_i(13129) := b"0000000000000000_0000000000000000_0000100100011001_1001011101101100"; -- 0.03554674506826003
	pesos_i(13130) := b"1111111111111111_1111111111111111_1110011010000110_0101001111110001"; -- -0.09951281886508137
	pesos_i(13131) := b"1111111111111111_1111111111111111_1110011101111011_0111001101110011"; -- -0.09577253757072873
	pesos_i(13132) := b"0000000000000000_0000000000000000_0010011101000111_0101000011011111"; -- 0.1534319443235286
	pesos_i(13133) := b"1111111111111111_1111111111111111_1111000011001001_0100101010101110"; -- -0.059428532065124925
	pesos_i(13134) := b"0000000000000000_0000000000000000_0000101100010010_1111001111000001"; -- 0.04325793713446086
	pesos_i(13135) := b"1111111111111111_1111111111111111_1101010010110010_1110101010011010"; -- -0.16914495231785345
	pesos_i(13136) := b"1111111111111111_1111111111111111_1110111000011010_0111110111001110"; -- -0.06990827290506799
	pesos_i(13137) := b"1111111111111111_1111111111111111_1110011111101011_0111100111101111"; -- -0.09406316672534167
	pesos_i(13138) := b"1111111111111111_1111111111111111_1110100000001110_1001010110101100"; -- -0.09352745582712853
	pesos_i(13139) := b"0000000000000000_0000000000000000_0001110101000001_0011010000101011"; -- 0.11427618076358383
	pesos_i(13140) := b"1111111111111111_1111111111111111_1101101011000000_0100001000110111"; -- -0.14550386576641278
	pesos_i(13141) := b"1111111111111111_1111111111111111_1101110000010001_0110000000101111"; -- -0.14035986765152225
	pesos_i(13142) := b"0000000000000000_0000000000000000_0001000111010100_1110000101110010"; -- 0.06965455095149072
	pesos_i(13143) := b"1111111111111111_1111111111111111_1110011101100101_0110110001110000"; -- -0.09610864887769287
	pesos_i(13144) := b"1111111111111111_1111111111111111_1110001011111001_0001101111111001"; -- -0.11338639429996356
	pesos_i(13145) := b"0000000000000000_0000000000000000_0001101011010100_0011011000110011"; -- 0.10480059371598623
	pesos_i(13146) := b"1111111111111111_1111111111111111_1110000100101001_0101011101100100"; -- -0.12046293067912806
	pesos_i(13147) := b"1111111111111111_1111111111111111_1111001011000011_0001100011110001"; -- -0.051710549439636405
	pesos_i(13148) := b"0000000000000000_0000000000000000_0001001000101101_0011010001010000"; -- 0.0710022636672688
	pesos_i(13149) := b"0000000000000000_0000000000000000_0001101111100110_0100000100000000"; -- 0.10898214570952822
	pesos_i(13150) := b"0000000000000000_0000000000000000_0001100110010010_1001101000000010"; -- 0.09989321279728594
	pesos_i(13151) := b"0000000000000000_0000000000000000_0000111010000010_1010110000001010"; -- 0.05668139692970138
	pesos_i(13152) := b"1111111111111111_1111111111111111_1110011000110100_1111011110110011"; -- -0.10075427899060467
	pesos_i(13153) := b"1111111111111111_1111111111111111_1101111100100110_1010010110000101"; -- -0.12831655035997064
	pesos_i(13154) := b"1111111111111111_1111111111111111_1110111010101101_0011001110001010"; -- -0.06766965748135181
	pesos_i(13155) := b"0000000000000000_0000000000000000_0000001110000011_0001000010011100"; -- 0.013718641278067253
	pesos_i(13156) := b"1111111111111111_1111111111111111_1111000001011101_1110100100010111"; -- -0.06106703932901992
	pesos_i(13157) := b"0000000000000000_0000000000000000_0000101111101101_0100000000110100"; -- 0.04658890969924786
	pesos_i(13158) := b"0000000000000000_0000000000000000_0001110010001111_0110000101001010"; -- 0.11156280567199621
	pesos_i(13159) := b"0000000000000000_0000000000000000_0000010110100110_1011010111010001"; -- 0.022075046172843803
	pesos_i(13160) := b"0000000000000000_0000000000000000_0001011001010000_0110010001001011"; -- 0.08716418114162638
	pesos_i(13161) := b"1111111111111111_1111111111111111_1110110001001100_0011001001000110"; -- -0.07696233554525708
	pesos_i(13162) := b"0000000000000000_0000000000000000_0010100001011110_0010100110111111"; -- 0.15768681445595584
	pesos_i(13163) := b"0000000000000000_0000000000000000_0001110000101111_1111101001010111"; -- 0.11010708458280628
	pesos_i(13164) := b"1111111111111111_1111111111111111_1110001110011001_1100011111000110"; -- -0.11093474774855157
	pesos_i(13165) := b"0000000000000000_0000000000000000_0001000010101101_1111000101101110"; -- 0.0651541607544984
	pesos_i(13166) := b"1111111111111111_1111111111111111_1111101101000101_0010000110101010"; -- -0.01847638699694702
	pesos_i(13167) := b"1111111111111111_1111111111111111_1110101001001001_0011000111001110"; -- -0.08482063986612606
	pesos_i(13168) := b"0000000000000000_0000000000000000_0001101000010101_1111101100100000"; -- 0.10189790286683356
	pesos_i(13169) := b"0000000000000000_0000000000000000_0000110001101011_0101000101000001"; -- 0.0485125335663238
	pesos_i(13170) := b"1111111111111111_1111111111111111_1110001010000010_1000000010110010"; -- -0.11519618648728713
	pesos_i(13171) := b"0000000000000000_0000000000000000_0001011110100011_1001000010110101"; -- 0.0923395579003347
	pesos_i(13172) := b"1111111111111111_1111111111111111_1110011100010101_0100101010000010"; -- -0.09733137441736907
	pesos_i(13173) := b"0000000000000000_0000000000000000_0000100111010101_0100110000110111"; -- 0.03841091472969775
	pesos_i(13174) := b"0000000000000000_0000000000000000_0000000000010010_1110001100101110"; -- 0.0002881991040821143
	pesos_i(13175) := b"0000000000000000_0000000000000000_0010000000011110_0111011010111100"; -- 0.12546484080811832
	pesos_i(13176) := b"1111111111111111_1111111111111111_1110011111110110_1101011110001111"; -- -0.09388973960070186
	pesos_i(13177) := b"1111111111111111_1111111111111111_1110011010000011_0110100011101011"; -- -0.09955734507888432
	pesos_i(13178) := b"1111111111111111_1111111111111111_1101101000100101_1000101000011000"; -- -0.14786469384633416
	pesos_i(13179) := b"0000000000000000_0000000000000000_0001001010001011_1010011110111011"; -- 0.0724434691280562
	pesos_i(13180) := b"0000000000000000_0000000000000000_0000011000000000_0011110101011001"; -- 0.02344115661254393
	pesos_i(13181) := b"1111111111111111_1111111111111111_1111111010010111_1001101011000010"; -- -0.005499198586876231
	pesos_i(13182) := b"0000000000000000_0000000000000000_0000100000010111_0001011100111010"; -- 0.03160233654852285
	pesos_i(13183) := b"1111111111111111_1111111111111111_1110111000111100_1100000111000111"; -- -0.06938542269973409
	pesos_i(13184) := b"1111111111111111_1111111111111111_1110111001100000_1001100111110111"; -- -0.06883847915033903
	pesos_i(13185) := b"0000000000000000_0000000000000000_0000011100101111_1101000101111100"; -- 0.02807339942344058
	pesos_i(13186) := b"0000000000000000_0000000000000000_0001110001110111_0001011010010101"; -- 0.11119214185617665
	pesos_i(13187) := b"1111111111111111_1111111111111111_1111101010001000_0101101000101011"; -- -0.021356930253665432
	pesos_i(13188) := b"0000000000000000_0000000000000000_0001110101101010_1111010011100001"; -- 0.11491327755812782
	pesos_i(13189) := b"0000000000000000_0000000000000000_0001111101110011_1100110100011011"; -- 0.1228607360287277
	pesos_i(13190) := b"0000000000000000_0000000000000000_0010000010111000_0000100100110011"; -- 0.12780816544940526
	pesos_i(13191) := b"0000000000000000_0000000000000000_0001010011101101_0101101110100010"; -- 0.08174679476929247
	pesos_i(13192) := b"1111111111111111_1111111111111111_1110011010000000_0000011001010101"; -- -0.09960899749423824
	pesos_i(13193) := b"1111111111111111_1111111111111111_1111101000000100_1011110111011101"; -- -0.023365148111929433
	pesos_i(13194) := b"0000000000000000_0000000000000000_0000110101101110_0010110001110111"; -- 0.05246236722155359
	pesos_i(13195) := b"1111111111111111_1111111111111111_1111101011111011_1001100010000100"; -- -0.019598453259858345
	pesos_i(13196) := b"0000000000000000_0000000000000000_0000111011000111_0011010011100110"; -- 0.05772715197841394
	pesos_i(13197) := b"0000000000000000_0000000000000000_0000000110011100_0111000001010100"; -- 0.006293316343001885
	pesos_i(13198) := b"1111111111111111_1111111111111111_1110000111101010_1101000111000000"; -- -0.11751069131133238
	pesos_i(13199) := b"1111111111111111_1111111111111111_1111011011011111_1011101000000111"; -- -0.03564870182921901
	pesos_i(13200) := b"0000000000000000_0000000000000000_0001001001110000_0101110100010100"; -- 0.07202703226351033
	pesos_i(13201) := b"1111111111111111_1111111111111111_1111111010110001_0011101000110100"; -- -0.0051082251205149054
	pesos_i(13202) := b"0000000000000000_0000000000000000_0001101011111100_0101101011101011"; -- 0.10541313392868235
	pesos_i(13203) := b"1111111111111111_1111111111111111_1110110101110111_0010000011111100"; -- -0.07240098800650983
	pesos_i(13204) := b"0000000000000000_0000000000000000_0001010001111101_1101101110010100"; -- 0.08004543642282007
	pesos_i(13205) := b"0000000000000000_0000000000000000_0010010100011010_0011100011110110"; -- 0.1449313735812335
	pesos_i(13206) := b"1111111111111111_1111111111111111_1101011001010001_0010011000100100"; -- -0.16282426478254328
	pesos_i(13207) := b"1111111111111111_1111111111111111_1111011100101011_0110100011001010"; -- -0.03449387624250671
	pesos_i(13208) := b"0000000000000000_0000000000000000_0010000101110010_1111111001010111"; -- 0.13066091168160182
	pesos_i(13209) := b"0000000000000000_0000000000000000_0010001001101110_0101010100011001"; -- 0.1344960389601222
	pesos_i(13210) := b"0000000000000000_0000000000000000_0000000101000011_0001011111010000"; -- 0.004930008185008231
	pesos_i(13211) := b"1111111111111111_1111111111111111_1110101001011100_1111000110011000"; -- -0.08451929120041621
	pesos_i(13212) := b"0000000000000000_0000000000000000_0001010001101101_0111011010000001"; -- 0.07979527129505729
	pesos_i(13213) := b"1111111111111111_1111111111111111_1111100110100001_0001000000011010"; -- -0.024886125297808148
	pesos_i(13214) := b"1111111111111111_1111111111111111_1111101110000100_0101001011000101"; -- -0.01751215645841514
	pesos_i(13215) := b"1111111111111111_1111111111111111_1111101110101100_0111100011010000"; -- -0.01689953735540136
	pesos_i(13216) := b"1111111111111111_1111111111111111_1111101000100111_0101000111100111"; -- -0.02283752546262889
	pesos_i(13217) := b"0000000000000000_0000000000000000_0000011000010101_1101000001100111"; -- 0.023770356241242286
	pesos_i(13218) := b"0000000000000000_0000000000000000_0001100100010000_1110110011010011"; -- 0.09791450638157204
	pesos_i(13219) := b"0000000000000000_0000000000000000_0001010001110100_1010000101110001"; -- 0.07990464210820825
	pesos_i(13220) := b"0000000000000000_0000000000000000_0001101111101011_0010110010110011"; -- 0.10905722978680676
	pesos_i(13221) := b"1111111111111111_1111111111111111_1110101101011111_1101110001110010"; -- -0.08056852541652766
	pesos_i(13222) := b"0000000000000000_0000000000000000_0001110101111110_0101111010111110"; -- 0.11520950461228346
	pesos_i(13223) := b"0000000000000000_0000000000000000_0001110010001010_1101111100100000"; -- 0.11149401214583674
	pesos_i(13224) := b"1111111111111111_1111111111111111_1101110001001111_1100000111101101"; -- -0.13940799682591412
	pesos_i(13225) := b"0000000000000000_0000000000000000_0001001100001000_0111101101001110"; -- 0.07434816989708071
	pesos_i(13226) := b"1111111111111111_1111111111111111_1101110011001011_0001111100110011"; -- -0.1375256063126623
	pesos_i(13227) := b"1111111111111111_1111111111111111_1110101111010110_1101111111111101"; -- -0.07875251828775953
	pesos_i(13228) := b"1111111111111111_1111111111111111_1111101000011011_0010000001000110"; -- -0.023023588981425137
	pesos_i(13229) := b"0000000000000000_0000000000000000_0000111001100010_0110100001111101"; -- 0.056189089361257154
	pesos_i(13230) := b"0000000000000000_0000000000000000_0000000111001100_0000110110101111"; -- 0.007019858552227013
	pesos_i(13231) := b"0000000000000000_0000000000000000_0001101111110011_0110000111110111"; -- 0.1091824749241478
	pesos_i(13232) := b"1111111111111111_1111111111111111_1111100110110010_0110011000100101"; -- -0.024621597242610285
	pesos_i(13233) := b"0000000000000000_0000000000000000_0000011111111110_0111100011110110"; -- 0.03122669220826253
	pesos_i(13234) := b"0000000000000000_0000000000000000_0000000110101100_1011000000110011"; -- 0.006541264040578339
	pesos_i(13235) := b"1111111111111111_1111111111111111_1110100001101010_1010110110101010"; -- -0.09212221719709257
	pesos_i(13236) := b"0000000000000000_0000000000000000_0000001111100100_0011100010111110"; -- 0.015201136031869133
	pesos_i(13237) := b"0000000000000000_0000000000000000_0001100100111110_1001000001001111"; -- 0.09861089646367371
	pesos_i(13238) := b"1111111111111111_1111111111111111_1110011100011001_1011001101010110"; -- -0.09726409091256585
	pesos_i(13239) := b"1111111111111111_1111111111111111_1110111001010101_1101110101111010"; -- -0.0690023018670084
	pesos_i(13240) := b"0000000000000000_0000000000000000_0010000101011011_0101011101100001"; -- 0.13030000809448802
	pesos_i(13241) := b"0000000000000000_0000000000000000_0000000101011110_1111010010111101"; -- 0.005355163622320924
	pesos_i(13242) := b"0000000000000000_0000000000000000_0001000100000110_1000100110001110"; -- 0.06650600156482749
	pesos_i(13243) := b"0000000000000000_0000000000000000_0001001001000101_0111001101110101"; -- 0.07137223830189723
	pesos_i(13244) := b"1111111111111111_1111111111111111_1110000001110000_1000101111011101"; -- -0.12328267919287292
	pesos_i(13245) := b"0000000000000000_0000000000000000_0000001001101110_0001111111101001"; -- 0.009492868886206748
	pesos_i(13246) := b"0000000000000000_0000000000000000_0000010111001111_0000001101100010"; -- 0.022690020871893722
	pesos_i(13247) := b"1111111111111111_1111111111111111_1110101010000100_0100100001000100"; -- -0.08391903247650631
	pesos_i(13248) := b"0000000000000000_0000000000000000_0001010110101010_1010001110100101"; -- 0.08463499820975122
	pesos_i(13249) := b"1111111111111111_1111111111111111_1110001010111101_0000000101100100"; -- -0.1143035060658169
	pesos_i(13250) := b"0000000000000000_0000000000000000_0000111001000110_1110100110001111"; -- 0.05576953629629466
	pesos_i(13251) := b"0000000000000000_0000000000000000_0001001110110011_0101001010110001"; -- 0.0769550019364856
	pesos_i(13252) := b"1111111111111111_1111111111111111_1110110010111011_1010111101110011"; -- -0.07526114890779602
	pesos_i(13253) := b"0000000000000000_0000000000000000_0001000001000010_0000000111100111"; -- 0.06350719338893944
	pesos_i(13254) := b"0000000000000000_0000000000000000_0000000011000111_0001111100001001"; -- 0.0030383487481284916
	pesos_i(13255) := b"0000000000000000_0000000000000000_0000000011011100_1001011001011100"; -- 0.00336589567402313
	pesos_i(13256) := b"0000000000000000_0000000000000000_0001110000101110_0010111001011000"; -- 0.11007966655302992
	pesos_i(13257) := b"0000000000000000_0000000000000000_0010001010011000_0010100001000000"; -- 0.13513423490961626
	pesos_i(13258) := b"1111111111111111_1111111111111111_1110000101010100_0000100000101100"; -- -0.11981152464616089
	pesos_i(13259) := b"0000000000000000_0000000000000000_0001001011000000_1001001000100001"; -- 0.07325089737840797
	pesos_i(13260) := b"1111111111111111_1111111111111111_1111011010011101_0101111000010001"; -- -0.03666126334079538
	pesos_i(13261) := b"1111111111111111_1111111111111111_1110011100110110_1000101001010000"; -- -0.0968240313801637
	pesos_i(13262) := b"0000000000000000_0000000000000000_0000111100101110_0011011010011010"; -- 0.05929890869027312
	pesos_i(13263) := b"0000000000000000_0000000000000000_0000110101010011_0110101011101101"; -- 0.05205410287652862
	pesos_i(13264) := b"1111111111111111_1111111111111111_1110100011011010_0001010100001001"; -- -0.09042233019438548
	pesos_i(13265) := b"0000000000000000_0000000000000000_0010001100000111_0101100100011011"; -- 0.13683087267577482
	pesos_i(13266) := b"0000000000000000_0000000000000000_0000111111110001_0001100110100110"; -- 0.062272646898319
	pesos_i(13267) := b"1111111111111111_1111111111111111_1101110000110001_0000100010001001"; -- -0.1398768105737162
	pesos_i(13268) := b"0000000000000000_0000000000000000_0001101110010000_1100001001111100"; -- 0.10767760777878518
	pesos_i(13269) := b"0000000000000000_0000000000000000_0010000110111101_1110010101010111"; -- 0.13180383083907565
	pesos_i(13270) := b"1111111111111111_1111111111111111_1110110001011000_1110111010011000"; -- -0.07676800535262839
	pesos_i(13271) := b"1111111111111111_1111111111111111_1101111001110011_0111100001111110"; -- -0.13105055746603878
	pesos_i(13272) := b"1111111111111111_1111111111111111_1110111101011111_0111101100101010"; -- -0.06494932381850103
	pesos_i(13273) := b"0000000000000000_0000000000000000_0001001000100011_0000001111010001"; -- 0.0708467851773189
	pesos_i(13274) := b"1111111111111111_1111111111111111_1110000100110011_1101011100100101"; -- -0.12030272810968648
	pesos_i(13275) := b"0000000000000000_0000000000000000_0010001111110100_0110110110011001"; -- 0.14044842705743008
	pesos_i(13276) := b"1111111111111111_1111111111111111_1101100101101000_1100011000010100"; -- -0.15074502954828925
	pesos_i(13277) := b"0000000000000000_0000000000000000_0001110000111010_1110101000111111"; -- 0.11027397198527383
	pesos_i(13278) := b"0000000000000000_0000000000000000_0000010110000101_0111001111101111"; -- 0.021567579107917643
	pesos_i(13279) := b"1111111111111111_1111111111111111_1111110100011110_1010111000010100"; -- -0.011250610557187467
	pesos_i(13280) := b"1111111111111111_1111111111111111_1110100000001000_0100011010000000"; -- -0.09362372765807585
	pesos_i(13281) := b"0000000000000000_0000000000000000_0000101001101100_1111101011111001"; -- 0.040725408377542495
	pesos_i(13282) := b"1111111111111111_1111111111111111_1110101110110111_0010100100110100"; -- -0.07923643574045694
	pesos_i(13283) := b"1111111111111111_1111111111111111_1101110000101101_0010111011110001"; -- -0.1399355565234818
	pesos_i(13284) := b"1111111111111111_1111111111111111_1111100001101010_1110011100011110"; -- -0.02961879273840623
	pesos_i(13285) := b"1111111111111111_1111111111111111_1110100100000100_0101000100000110"; -- -0.08977788555287539
	pesos_i(13286) := b"1111111111111111_1111111111111111_1111111101101000_0100010111101010"; -- -0.002315168817575298
	pesos_i(13287) := b"0000000000000000_0000000000000000_0001101110100001_0010100110001101"; -- 0.1079278917739646
	pesos_i(13288) := b"1111111111111111_1111111111111111_1111001110100100_0011010100110100"; -- -0.04827563733009984
	pesos_i(13289) := b"1111111111111111_1111111111111111_1111110001010100_1111101000011110"; -- -0.014328353510247017
	pesos_i(13290) := b"1111111111111111_1111111111111111_1101101001111010_0001000010110110"; -- -0.14657493167706484
	pesos_i(13291) := b"0000000000000000_0000000000000000_0001110001111100_1101001100110110"; -- 0.11127967906062852
	pesos_i(13292) := b"0000000000000000_0000000000000000_0000111000110110_0011110101101110"; -- 0.0555151361449066
	pesos_i(13293) := b"1111111111111111_1111111111111111_1111001011001011_0010111100110001"; -- -0.05158715310010361
	pesos_i(13294) := b"1111111111111111_1111111111111111_1111000010101001_1111101001000011"; -- -0.05990634792313335
	pesos_i(13295) := b"0000000000000000_0000000000000000_0001110110101101_0101101110101000"; -- 0.11592648356753951
	pesos_i(13296) := b"0000000000000000_0000000000000000_0000111100100111_1100000111011110"; -- 0.05920039811143189
	pesos_i(13297) := b"0000000000000000_0000000000000000_0000111000010000_0111011011111011"; -- 0.054938732353945655
	pesos_i(13298) := b"1111111111111111_1111111111111111_1111100100011001_0011011111010010"; -- -0.026958953233988364
	pesos_i(13299) := b"0000000000000000_0000000000000000_0001100101001101_0110111010110111"; -- 0.09883777593944278
	pesos_i(13300) := b"0000000000000000_0000000000000000_0010001010100010_0001011001101011"; -- 0.13528576009153484
	pesos_i(13301) := b"1111111111111111_1111111111111111_1111101111101001_0101111011100101"; -- -0.01597029598714495
	pesos_i(13302) := b"1111111111111111_1111111111111111_1111100101101000_1011000100111111"; -- -0.025746271257116222
	pesos_i(13303) := b"1111111111111111_1111111111111111_1111111110100101_0001101101010011"; -- -0.0013869211533409768
	pesos_i(13304) := b"0000000000000000_0000000000000000_0000010111010011_0011110011010010"; -- 0.022754479741173214
	pesos_i(13305) := b"0000000000000000_0000000000000000_0001000110011011_0101110101001000"; -- 0.06877692234791971
	pesos_i(13306) := b"1111111111111111_1111111111111111_1101100101010101_0110001111010101"; -- -0.1510408023798428
	pesos_i(13307) := b"0000000000000000_0000000000000000_0000100101001011_0001100011100001"; -- 0.03630214201589473
	pesos_i(13308) := b"0000000000000000_0000000000000000_0001011000101110_1011000000000010"; -- 0.08664989522046855
	pesos_i(13309) := b"1111111111111111_1111111111111111_1101111001000011_1101011111011101"; -- -0.13177729469590851
	pesos_i(13310) := b"1111111111111111_1111111111111111_1111101100011000_1100111100100100"; -- -0.019152692599690272
	pesos_i(13311) := b"0000000000000000_0000000000000000_0000110011110101_1000101011110100"; -- 0.05062168554351779
	pesos_i(13312) := b"0000000000000000_0000000000000000_0010001110000010_0011111100100111"; -- 0.1387061567276578
	pesos_i(13313) := b"1111111111111111_1111111111111111_1111010011010010_1100101001111000"; -- -0.04365858625690243
	pesos_i(13314) := b"1111111111111111_1111111111111111_1111000101010000_0100110011010001"; -- -0.05736846825706001
	pesos_i(13315) := b"1111111111111111_1111111111111111_1111001001110110_0101100101010101"; -- -0.052881638277210576
	pesos_i(13316) := b"1111111111111111_1111111111111111_1110010110101000_1100101101100111"; -- -0.10289314973438614
	pesos_i(13317) := b"1111111111111111_1111111111111111_1111111100101011_0011011100110110"; -- -0.0032468313566323516
	pesos_i(13318) := b"0000000000000000_0000000000000000_0000000000011101_1100000111010000"; -- 0.00045405691820674874
	pesos_i(13319) := b"0000000000000000_0000000000000000_0010000011110000_1011010100100110"; -- 0.12867290657454813
	pesos_i(13320) := b"0000000000000000_0000000000000000_0001000010001100_1111010100101100"; -- 0.06465084374502854
	pesos_i(13321) := b"0000000000000000_0000000000000000_0001101110000000_1101101010111011"; -- 0.10743491246461308
	pesos_i(13322) := b"0000000000000000_0000000000000000_0000100010001100_0010110100000110"; -- 0.033388914100117725
	pesos_i(13323) := b"0000000000000000_0000000000000000_0001110001110000_0001000101011101"; -- 0.11108501940934579
	pesos_i(13324) := b"1111111111111111_1111111111111111_1111110100000011_1001111001100100"; -- -0.011663532805714999
	pesos_i(13325) := b"1111111111111111_1111111111111111_1111011001111001_1100000111101101"; -- -0.03720462762281311
	pesos_i(13326) := b"1111111111111111_1111111111111111_1110001000110000_0001000011100011"; -- -0.11645407152951427
	pesos_i(13327) := b"1111111111111111_1111111111111111_1110110011001000_0000011101100000"; -- -0.07507280266472044
	pesos_i(13328) := b"1111111111111111_1111111111111111_1110011001101111_0001111101111001"; -- -0.09986689838190915
	pesos_i(13329) := b"0000000000000000_0000000000000000_0000011100001000_0001111110011000"; -- 0.027467703379618274
	pesos_i(13330) := b"1111111111111111_1111111111111111_1101111111000000_1001100100111101"; -- -0.12596742877550213
	pesos_i(13331) := b"0000000000000000_0000000000000000_0001010101100010_1110010000001111"; -- 0.08354020461383992
	pesos_i(13332) := b"0000000000000000_0000000000000000_0000100100100001_1101110100010001"; -- 0.03567296654554933
	pesos_i(13333) := b"0000000000000000_0000000000000000_0000111000100011_0010100000001111"; -- 0.055223945310242356
	pesos_i(13334) := b"1111111111111111_1111111111111111_1111111111010011_1010100000000010"; -- -0.0006766313721675876
	pesos_i(13335) := b"0000000000000000_0000000000000000_0000001001010001_0100101110010110"; -- 0.009052967178134818
	pesos_i(13336) := b"1111111111111111_1111111111111111_1110001101010111_1001010101011110"; -- -0.1119448323157929
	pesos_i(13337) := b"0000000000000000_0000000000000000_0000110110110011_0110011110001010"; -- 0.0535187447386225
	pesos_i(13338) := b"0000000000000000_0000000000000000_0001011001001011_0110111100101000"; -- 0.08708853456269505
	pesos_i(13339) := b"0000000000000000_0000000000000000_0001101011101010_1101110111101010"; -- 0.1051462837350034
	pesos_i(13340) := b"0000000000000000_0000000000000000_0000110101001010_0001110100011101"; -- 0.051912135746352485
	pesos_i(13341) := b"1111111111111111_1111111111111111_1110000010101110_0000011110100001"; -- -0.12234451590136991
	pesos_i(13342) := b"1111111111111111_1111111111111111_1110011010011101_0101111100100110"; -- -0.09916119894425449
	pesos_i(13343) := b"0000000000000000_0000000000000000_0001011100001101_1011100010100000"; -- 0.09005311878814817
	pesos_i(13344) := b"0000000000000000_0000000000000000_0001000110010110_0110101111010110"; -- 0.06870149583511481
	pesos_i(13345) := b"0000000000000000_0000000000000000_0001101010101111_1110100110100100"; -- 0.10424671409636783
	pesos_i(13346) := b"1111111111111111_1111111111111111_1110000111010110_1101001000011001"; -- -0.11781584637930284
	pesos_i(13347) := b"1111111111111111_1111111111111111_1111100010010110_1111111001101110"; -- -0.028946016397795975
	pesos_i(13348) := b"1111111111111111_1111111111111111_1111010101111000_1001010000110111"; -- -0.041128861111143764
	pesos_i(13349) := b"0000000000000000_0000000000000000_0000100111010010_0110000110110101"; -- 0.03836641957756913
	pesos_i(13350) := b"0000000000000000_0000000000000000_0000011100011011_1010110000011111"; -- 0.027765996421113014
	pesos_i(13351) := b"1111111111111111_1111111111111111_1111010011110000_1101010101010111"; -- -0.043200174672684624
	pesos_i(13352) := b"0000000000000000_0000000000000000_0000000010110100_0010010001001100"; -- 0.0027487455775216945
	pesos_i(13353) := b"1111111111111111_1111111111111111_1110000110111100_0111001111100001"; -- -0.11821819070945722
	pesos_i(13354) := b"0000000000000000_0000000000000000_0010000010111000_1110011000111010"; -- 0.12782133972529278
	pesos_i(13355) := b"0000000000000000_0000000000000000_0001001001110101_1011001001110110"; -- 0.07210841549040625
	pesos_i(13356) := b"1111111111111111_1111111111111111_1111011100110110_1000100010110111"; -- -0.03432412665931281
	pesos_i(13357) := b"1111111111111111_1111111111111111_1101110011111101_1011100000110001"; -- -0.13675354774397466
	pesos_i(13358) := b"0000000000000000_0000000000000000_0001010111110101_0111001010010100"; -- 0.08577648280602614
	pesos_i(13359) := b"1111111111111111_1111111111111111_1110001111101001_1110000110100110"; -- -0.1097125024553323
	pesos_i(13360) := b"0000000000000000_0000000000000000_0001011100011110_1010011000100101"; -- 0.09031141668028789
	pesos_i(13361) := b"0000000000000000_0000000000000000_0000110001011110_1010001100101101"; -- 0.048319052097788744
	pesos_i(13362) := b"0000000000000000_0000000000000000_0010000111100010_0000111111011101"; -- 0.13235568196627887
	pesos_i(13363) := b"1111111111111111_1111111111111111_1111010110001010_1111001010101100"; -- -0.04084857265151332
	pesos_i(13364) := b"0000000000000000_0000000000000000_0000111111101011_0010010110011110"; -- 0.0621818076838518
	pesos_i(13365) := b"0000000000000000_0000000000000000_0001011110010111_0101100011011000"; -- 0.09215312271181846
	pesos_i(13366) := b"1111111111111111_1111111111111111_1110101100011110_1111001000001111"; -- -0.0815590584865239
	pesos_i(13367) := b"0000000000000000_0000000000000000_0001011000011101_1001110010110010"; -- 0.0863893446874113
	pesos_i(13368) := b"1111111111111111_1111111111111111_1101110000100000_0100001110101111"; -- -0.14013268441710347
	pesos_i(13369) := b"1111111111111111_1111111111111111_1110001001001010_0110011000101111"; -- -0.1160522589402671
	pesos_i(13370) := b"0000000000000000_0000000000000000_0001101010101111_1000100000100101"; -- 0.1042409028670796
	pesos_i(13371) := b"0000000000000000_0000000000000000_0010001101100001_1101101100001101"; -- 0.13821190889310392
	pesos_i(13372) := b"1111111111111111_1111111111111111_1101111000010000_1111001101100111"; -- -0.1325538514048824
	pesos_i(13373) := b"0000000000000000_0000000000000000_0001001101111110_0010100000000011"; -- 0.0761437423992783
	pesos_i(13374) := b"0000000000000000_0000000000000000_0001011000111100_1110111000000000"; -- 0.08686721325728024
	pesos_i(13375) := b"1111111111111111_1111111111111111_1111100111101010_0111001101111011"; -- -0.023766310236143354
	pesos_i(13376) := b"0000000000000000_0000000000000000_0000101100110010_0000010010111000"; -- 0.0437319707851911
	pesos_i(13377) := b"0000000000000000_0000000000000000_0000011101010011_1111011011101011"; -- 0.028624947033471727
	pesos_i(13378) := b"0000000000000000_0000000000000000_0000100101010010_0000101011000100"; -- 0.036408112413317234
	pesos_i(13379) := b"1111111111111111_1111111111111111_1110101100111100_1001101110100111"; -- -0.081106444988006
	pesos_i(13380) := b"0000000000000000_0000000000000000_0001111011100001_1111110110100100"; -- 0.12063584559076952
	pesos_i(13381) := b"0000000000000000_0000000000000000_0001010001010100_0001000110001101"; -- 0.07940778443890813
	pesos_i(13382) := b"0000000000000000_0000000000000000_0001110000001110_0100000010010000"; -- 0.10959247119101118
	pesos_i(13383) := b"1111111111111111_1111111111111111_1111100101100001_0011101110101011"; -- -0.025860090925677436
	pesos_i(13384) := b"0000000000000000_0000000000000000_0001001001011000_0101111001111111"; -- 0.07166090576195372
	pesos_i(13385) := b"0000000000000000_0000000000000000_0000110010101010_1011010110111100"; -- 0.049479826348883815
	pesos_i(13386) := b"1111111111111111_1111111111111111_1110010100110010_0101100001110110"; -- -0.10470053787017021
	pesos_i(13387) := b"1111111111111111_1111111111111111_1111010110000110_0001011010000001"; -- -0.04092273095575649
	pesos_i(13388) := b"1111111111111111_1111111111111111_1111111001110111_0010000101000101"; -- -0.005994721175590387
	pesos_i(13389) := b"0000000000000000_0000000000000000_0001100100111111_1011100011011010"; -- 0.09862857166459242
	pesos_i(13390) := b"1111111111111111_1111111111111111_1110111011111001_0101000101001110"; -- -0.06650821535888168
	pesos_i(13391) := b"0000000000000000_0000000000000000_0000100100100100_0100010111100111"; -- 0.035709732988469786
	pesos_i(13392) := b"0000000000000000_0000000000000000_0000000001011010_1010011011111100"; -- 0.0013832440471730884
	pesos_i(13393) := b"0000000000000000_0000000000000000_0001111100101110_1000011001100010"; -- 0.12180366422600904
	pesos_i(13394) := b"1111111111111111_1111111111111111_1110101011001010_0011100111110011"; -- -0.08285177046281823
	pesos_i(13395) := b"0000000000000000_0000000000000000_0000101101111110_1110101001110010"; -- 0.04490533147172265
	pesos_i(13396) := b"1111111111111111_1111111111111111_1111000000001001_0011011011111101"; -- -0.062359393269325776
	pesos_i(13397) := b"1111111111111111_1111111111111111_1110011010101011_1100001101000110"; -- -0.09894160775685018
	pesos_i(13398) := b"0000000000000000_0000000000000000_0001101001010000_0010111011000111"; -- 0.1027859913092225
	pesos_i(13399) := b"0000000000000000_0000000000000000_0010000001100101_1011111110010000"; -- 0.12655255582566463
	pesos_i(13400) := b"1111111111111111_1111111111111111_1110101010001010_0111011111010100"; -- -0.08382464485747605
	pesos_i(13401) := b"1111111111111111_1111111111111111_1110101100011011_1010110100110011"; -- -0.08160893919122296
	pesos_i(13402) := b"0000000000000000_0000000000000000_0000000110111101_0010001010011001"; -- 0.006792223237822337
	pesos_i(13403) := b"0000000000000000_0000000000000000_0000100110111110_0011101001010100"; -- 0.038058896568403396
	pesos_i(13404) := b"1111111111111111_1111111111111111_1101111001001011_1100110110101110"; -- -0.13165583142606302
	pesos_i(13405) := b"0000000000000000_0000000000000000_0001000000100110_0100101111010000"; -- 0.06308435269289486
	pesos_i(13406) := b"0000000000000000_0000000000000000_0001011011100010_0000101010011001"; -- 0.0893866179014836
	pesos_i(13407) := b"0000000000000000_0000000000000000_0001111100111100_1111100100011111"; -- 0.12202412605197178
	pesos_i(13408) := b"1111111111111111_1111111111111111_1101100101101101_1101111101110011"; -- -0.15066722326587767
	pesos_i(13409) := b"0000000000000000_0000000000000000_0000100111001000_1011101010010001"; -- 0.038219128096547095
	pesos_i(13410) := b"1111111111111111_1111111111111111_1110111010110110_1110001100111101"; -- -0.06752185582401478
	pesos_i(13411) := b"1111111111111111_1111111111111111_1110110010000101_1010001101000110"; -- -0.07608584917321073
	pesos_i(13412) := b"0000000000000000_0000000000000000_0001001011001010_0111111100001101"; -- 0.07340234822649322
	pesos_i(13413) := b"1111111111111111_1111111111111111_1110101011100011_1000111111110110"; -- -0.08246517416633449
	pesos_i(13414) := b"0000000000000000_0000000000000000_0001000011110111_0000100101111001"; -- 0.06626948558971497
	pesos_i(13415) := b"0000000000000000_0000000000000000_0000101111011111_1000111000011101"; -- 0.046379930539545464
	pesos_i(13416) := b"1111111111111111_1111111111111111_1101101111100110_1011000110110100"; -- -0.1410111366625153
	pesos_i(13417) := b"0000000000000000_0000000000000000_0001110101001101_0110101110100110"; -- 0.11446259312964667
	pesos_i(13418) := b"1111111111111111_1111111111111111_1101101000101010_1011011011101001"; -- -0.1477857285119593
	pesos_i(13419) := b"1111111111111111_1111111111111111_1110000101011000_1010010000111111"; -- -0.11974118671363275
	pesos_i(13420) := b"0000000000000000_0000000000000000_0010001010000010_1111000000101000"; -- 0.13481045706637462
	pesos_i(13421) := b"1111111111111111_1111111111111111_1110010010000101_0110100011110110"; -- -0.1073393249189236
	pesos_i(13422) := b"0000000000000000_0000000000000000_0010001111110110_0111011010010001"; -- 0.14047947914350975
	pesos_i(13423) := b"0000000000000000_0000000000000000_0001100001001101_0000000001111010"; -- 0.09492495516530972
	pesos_i(13424) := b"0000000000000000_0000000000000000_0010010111010110_1001111101111011"; -- 0.1478061367101554
	pesos_i(13425) := b"0000000000000000_0000000000000000_0000011100010101_0001010100011011"; -- 0.027665442635267344
	pesos_i(13426) := b"0000000000000000_0000000000000000_0010011011011110_1111110011101101"; -- 0.15184002664427754
	pesos_i(13427) := b"0000000000000000_0000000000000000_0010001010101100_1100100000001100"; -- 0.13544893534331282
	pesos_i(13428) := b"0000000000000000_0000000000000000_0001101000110100_0100110100001110"; -- 0.1023605499372558
	pesos_i(13429) := b"1111111111111111_1111111111111111_1111100010011001_0110011000001011"; -- -0.0289093229355265
	pesos_i(13430) := b"1111111111111111_1111111111111111_1111011010010110_1111110000111011"; -- -0.03675864747866518
	pesos_i(13431) := b"1111111111111111_1111111111111111_1111100010010000_1111011100000000"; -- -0.029038012037682737
	pesos_i(13432) := b"1111111111111111_1111111111111111_1110110110011010_1010101010111011"; -- -0.07185872021605771
	pesos_i(13433) := b"1111111111111111_1111111111111111_1111010011111010_1111001111100111"; -- -0.04304576500595988
	pesos_i(13434) := b"0000000000000000_0000000000000000_0001100101101000_0010110000011001"; -- 0.09924579245737068
	pesos_i(13435) := b"1111111111111111_1111111111111111_1110000111001010_1111100001010000"; -- -0.11799667394795983
	pesos_i(13436) := b"1111111111111111_1111111111111111_1111100111001101_0101011101001101"; -- -0.02421049472336303
	pesos_i(13437) := b"0000000000000000_0000000000000000_0001110101101101_1011010110110110"; -- 0.11495528883362907
	pesos_i(13438) := b"1111111111111111_1111111111111111_1111111100000001_0011000111101001"; -- -0.003888016262075474
	pesos_i(13439) := b"1111111111111111_1111111111111111_1110100111001110_0111111011100010"; -- -0.08669287662429327
	pesos_i(13440) := b"0000000000000000_0000000000000000_0001100100000010_0110011111011110"; -- 0.09769295850225686
	pesos_i(13441) := b"1111111111111111_1111111111111111_1110110001101111_0011110001000010"; -- -0.07642768270357247
	pesos_i(13442) := b"0000000000000000_0000000000000000_0001111111001111_0011111100000001"; -- 0.12425607467131142
	pesos_i(13443) := b"0000000000000000_0000000000000000_0000010101111001_1001100100000011"; -- 0.021386683690403387
	pesos_i(13444) := b"1111111111111111_1111111111111111_1110111100010100_0111110101111011"; -- -0.0660935950381285
	pesos_i(13445) := b"1111111111111111_1111111111111111_1111010100110110_1001001010010010"; -- -0.04213603905309445
	pesos_i(13446) := b"1111111111111111_1111111111111111_1110001001111010_0100011100111001"; -- -0.1153216825628964
	pesos_i(13447) := b"1111111111111111_1111111111111111_1111010011011100_0000100101001010"; -- -0.04351751265159534
	pesos_i(13448) := b"1111111111111111_1111111111111111_1110011110101001_0011111111101000"; -- -0.09507370548953886
	pesos_i(13449) := b"1111111111111111_1111111111111111_1101101110010110_1011111010111101"; -- -0.14223106267809657
	pesos_i(13450) := b"0000000000000000_0000000000000000_0010001000000001_0001010001001011"; -- 0.13282896837550903
	pesos_i(13451) := b"0000000000000000_0000000000000000_0000001000001101_0100000111000011"; -- 0.008014783991432144
	pesos_i(13452) := b"0000000000000000_0000000000000000_0000000101001101_1011000110011101"; -- 0.0050917634119159215
	pesos_i(13453) := b"0000000000000000_0000000000000000_0001011111110111_1111101011010100"; -- 0.09362762135182323
	pesos_i(13454) := b"1111111111111111_1111111111111111_1111000100011010_0100111111010000"; -- -0.05819226429206041
	pesos_i(13455) := b"1111111111111111_1111111111111111_1110110101101100_1101000111000100"; -- -0.07255829770462001
	pesos_i(13456) := b"1111111111111111_1111111111111111_1111101100100110_0010011010111010"; -- -0.018949107712407955
	pesos_i(13457) := b"0000000000000000_0000000000000000_0001110001000111_0011100101101110"; -- 0.1104617970446314
	pesos_i(13458) := b"0000000000000000_0000000000000000_0010000011000010_1111100101011010"; -- 0.12797506764087396
	pesos_i(13459) := b"1111111111111111_1111111111111111_1110011000101011_1101000101010111"; -- -0.10089389445288047
	pesos_i(13460) := b"1111111111111111_1111111111111111_1110100110001101_0100101101100110"; -- -0.08768776664823173
	pesos_i(13461) := b"0000000000000000_0000000000000000_0001100001101111_0000111000010011"; -- 0.09544456456581621
	pesos_i(13462) := b"0000000000000000_0000000000000000_0000001110111100_0110101110101011"; -- 0.014593819858255069
	pesos_i(13463) := b"0000000000000000_0000000000000000_0001110101101011_0001010000101110"; -- 0.11491514326757496
	pesos_i(13464) := b"1111111111111111_1111111111111111_1111011000001001_0001101011000100"; -- -0.038923575478712155
	pesos_i(13465) := b"0000000000000000_0000000000000000_0000011011001010_1111111100000100"; -- 0.026534975503359395
	pesos_i(13466) := b"1111111111111111_1111111111111111_1110111100011000_1100111111001110"; -- -0.06602765298480862
	pesos_i(13467) := b"1111111111111111_1111111111111111_1111001011001000_0111100011001101"; -- -0.051628541920071575
	pesos_i(13468) := b"0000000000000000_0000000000000000_0000110001010110_1100111101011010"; -- 0.04819961498420921
	pesos_i(13469) := b"1111111111111111_1111111111111111_1111101110001010_1101001001111001"; -- -0.017412991907947952
	pesos_i(13470) := b"0000000000000000_0000000000000000_0000110110010101_0100110000101011"; -- 0.05305934964913322
	pesos_i(13471) := b"0000000000000000_0000000000000000_0010001010001100_0110001101101101"; -- 0.13495465659778755
	pesos_i(13472) := b"0000000000000000_0000000000000000_0001011110000001_1000011011001111"; -- 0.09182016901793921
	pesos_i(13473) := b"0000000000000000_0000000000000000_0000001100111001_0101101001101111"; -- 0.012593891273661893
	pesos_i(13474) := b"1111111111111111_1111111111111111_1111011001110111_0111100110001100"; -- -0.03723945942569025
	pesos_i(13475) := b"0000000000000000_0000000000000000_0001000010011110_1110111010111110"; -- 0.06492511884999712
	pesos_i(13476) := b"0000000000000000_0000000000000000_0001111110010101_1110110111100011"; -- 0.12338148880923185
	pesos_i(13477) := b"1111111111111111_1111111111111111_1110011110001110_1111110100111001"; -- -0.09547440864282457
	pesos_i(13478) := b"0000000000000000_0000000000000000_0000110101010011_0011010110111010"; -- 0.052050931857222205
	pesos_i(13479) := b"0000000000000000_0000000000000000_0001111011111111_0111101100000010"; -- 0.12108582310395778
	pesos_i(13480) := b"1111111111111111_1111111111111111_1110011110010000_0000110001010000"; -- -0.09545825046819342
	pesos_i(13481) := b"0000000000000000_0000000000000000_0000010011100000_0101010011100110"; -- 0.019048029194455706
	pesos_i(13482) := b"1111111111111111_1111111111111111_1111001101110001_1010110001001111"; -- -0.04904673634245298
	pesos_i(13483) := b"1111111111111111_1111111111111111_1111000111010101_1000000000110110"; -- -0.055335985920175704
	pesos_i(13484) := b"1111111111111111_1111111111111111_1110100110110011_0010010110010010"; -- -0.08711018733488936
	pesos_i(13485) := b"1111111111111111_1111111111111111_1111101011111000_1001000001011111"; -- -0.019644715125158363
	pesos_i(13486) := b"0000000000000000_0000000000000000_0001101100011100_0101100110100100"; -- 0.10590133918638296
	pesos_i(13487) := b"1111111111111111_1111111111111111_1111001101010111_0111101101000110"; -- -0.04944638762316269
	pesos_i(13488) := b"0000000000000000_0000000000000000_0010001101010101_0011001011100000"; -- 0.13801877952948907
	pesos_i(13489) := b"1111111111111111_1111111111111111_1110010101110011_1100001010111010"; -- -0.10370238269784308
	pesos_i(13490) := b"0000000000000000_0000000000000000_0001001000010010_1001110001111101"; -- 0.07059648574345673
	pesos_i(13491) := b"0000000000000000_0000000000000000_0000111100001010_0000000001001110"; -- 0.05874635602096877
	pesos_i(13492) := b"1111111111111111_1111111111111111_1110100100001010_0100011101000011"; -- -0.08968691446598318
	pesos_i(13493) := b"0000000000000000_0000000000000000_0010010000101110_1001001010001110"; -- 0.14133563961084714
	pesos_i(13494) := b"1111111111111111_1111111111111111_1111101011100100_1101010100011000"; -- -0.019945794828485165
	pesos_i(13495) := b"0000000000000000_0000000000000000_0001111100100001_0011001101010001"; -- 0.12160034872265506
	pesos_i(13496) := b"1111111111111111_1111111111111111_1101110000111110_1110000110110011"; -- -0.13966550245280748
	pesos_i(13497) := b"0000000000000000_0000000000000000_0010001011110010_1000011101010100"; -- 0.1365131931147877
	pesos_i(13498) := b"0000000000000000_0000000000000000_0000000100110001_1100110100110010"; -- 0.004666161310465375
	pesos_i(13499) := b"0000000000000000_0000000000000000_0001010011010101_0100001110110100"; -- 0.08137915746419146
	pesos_i(13500) := b"1111111111111111_1111111111111111_1111101101011010_0110101101110111"; -- -0.01815155367417317
	pesos_i(13501) := b"0000000000000000_0000000000000000_0000010011001000_1110100111110100"; -- 0.018690702551084733
	pesos_i(13502) := b"0000000000000000_0000000000000000_0000011111010111_0111000000000001"; -- 0.03063106559621257
	pesos_i(13503) := b"0000000000000000_0000000000000000_0001000101011110_0100010001100010"; -- 0.06784465202066044
	pesos_i(13504) := b"0000000000000000_0000000000000000_0000110000000100_0011011110000001"; -- 0.046939343457002285
	pesos_i(13505) := b"1111111111111111_1111111111111111_1110011111000100_0101110100101011"; -- -0.09465997404526175
	pesos_i(13506) := b"1111111111111111_1111111111111111_1111110101100011_1001001100111110"; -- -0.010199353615187035
	pesos_i(13507) := b"1111111111111111_1111111111111111_1110100010011111_1110001110000110"; -- -0.0913102909800747
	pesos_i(13508) := b"1111111111111111_1111111111111111_1111110011010101_1101000100110100"; -- -0.012362408394243941
	pesos_i(13509) := b"0000000000000000_0000000000000000_0000100100011010_1100001111110110"; -- 0.03556465880832137
	pesos_i(13510) := b"0000000000000000_0000000000000000_0000101111111100_1001100110000010"; -- 0.04682311458285205
	pesos_i(13511) := b"1111111111111111_1111111111111111_1111101110011111_1110101010011111"; -- -0.0170911181250193
	pesos_i(13512) := b"0000000000000000_0000000000000000_0001111110111111_1011000011001010"; -- 0.124018716161187
	pesos_i(13513) := b"0000000000000000_0000000000000000_0001011001001011_1111001100101010"; -- 0.08709640289002815
	pesos_i(13514) := b"0000000000000000_0000000000000000_0001010111111011_1010000001101011"; -- 0.08587076773678431
	pesos_i(13515) := b"1111111111111111_1111111111111111_1111110111100111_0100010111000101"; -- -0.008189811160722654
	pesos_i(13516) := b"1111111111111111_1111111111111111_1111000100110000_0001110100110011"; -- -0.05785958773005501
	pesos_i(13517) := b"0000000000000000_0000000000000000_0000100100000110_1111011111110001"; -- 0.03526258124944047
	pesos_i(13518) := b"0000000000000000_0000000000000000_0001111101011100_1101101000100100"; -- 0.12251056082068364
	pesos_i(13519) := b"0000000000000000_0000000000000000_0001111101001011_1011110100111010"; -- 0.12224943797712955
	pesos_i(13520) := b"1111111111111111_1111111111111111_1110011001100001_1101101101111100"; -- -0.10006931522828197
	pesos_i(13521) := b"1111111111111111_1111111111111111_1110010111010100_1111011011100010"; -- -0.10221917133529118
	pesos_i(13522) := b"0000000000000000_0000000000000000_0000001101001110_1111010100111111"; -- 0.012923553420983055
	pesos_i(13523) := b"0000000000000000_0000000000000000_0000001010100111_1010010101011100"; -- 0.01037057390542882
	pesos_i(13524) := b"0000000000000000_0000000000000000_0001001101100100_0111111000010010"; -- 0.0757521431969646
	pesos_i(13525) := b"1111111111111111_1111111111111111_1111000101110101_0101110011100111"; -- -0.05680293435269159
	pesos_i(13526) := b"1111111111111111_1111111111111111_1111010111111100_1100001100110010"; -- -0.0391119005199021
	pesos_i(13527) := b"0000000000000000_0000000000000000_0001110100100001_0011001111111000"; -- 0.11378788761113139
	pesos_i(13528) := b"1111111111111111_1111111111111111_1110101010110010_1010011111011101"; -- -0.0832114301590139
	pesos_i(13529) := b"1111111111111111_1111111111111111_1110001101100111_1100111001111011"; -- -0.11169728744099708
	pesos_i(13530) := b"0000000000000000_0000000000000000_0001000001010010_0100101000010011"; -- 0.06375563576437562
	pesos_i(13531) := b"1111111111111111_1111111111111111_1110000110110110_1001111001110100"; -- -0.11830720573908271
	pesos_i(13532) := b"0000000000000000_0000000000000000_0000000000001000_0001001111001100"; -- 0.00012325030838714616
	pesos_i(13533) := b"1111111111111111_1111111111111111_1110010010100111_0110101100100000"; -- -0.10682039704957896
	pesos_i(13534) := b"0000000000000000_0000000000000000_0001000001101100_1010101000100111"; -- 0.0641580910308392
	pesos_i(13535) := b"0000000000000000_0000000000000000_0000011010011110_0110111111101100"; -- 0.02585505978523497
	pesos_i(13536) := b"0000000000000000_0000000000000000_0001001111011011_0000110011010001"; -- 0.07756118872718823
	pesos_i(13537) := b"0000000000000000_0000000000000000_0001001011001111_1000111000011000"; -- 0.0734795388651699
	pesos_i(13538) := b"0000000000000000_0000000000000000_0010001100110101_1001000101110110"; -- 0.1375361358819789
	pesos_i(13539) := b"1111111111111111_1111111111111111_1110010100110111_1010101110010001"; -- -0.10461929051410054
	pesos_i(13540) := b"0000000000000000_0000000000000000_0001100001101010_1011101000111000"; -- 0.09537853114627352
	pesos_i(13541) := b"1111111111111111_1111111111111111_1110010110001101_0101111111000011"; -- -0.10331155293357326
	pesos_i(13542) := b"0000000000000000_0000000000000000_0010011001011101_1100110101011110"; -- 0.14986880817852027
	pesos_i(13543) := b"0000000000000000_0000000000000000_0010000011000001_0001011110100100"; -- 0.1279463552638547
	pesos_i(13544) := b"1111111111111111_1111111111111111_1111100001001000_0000000100111100"; -- -0.030151293655186675
	pesos_i(13545) := b"1111111111111111_1111111111111111_1111110111000111_0010001011000111"; -- -0.00868017802216194
	pesos_i(13546) := b"1111111111111111_1111111111111111_1110111011110001_1110110000001101"; -- -0.06662106206215715
	pesos_i(13547) := b"0000000000000000_0000000000000000_0001100101110101_0011000111101000"; -- 0.09944450295186695
	pesos_i(13548) := b"1111111111111111_1111111111111111_1111111001100100_1011111010111111"; -- -0.006275251846503721
	pesos_i(13549) := b"0000000000000000_0000000000000000_0001010000111110_0010000010110100"; -- 0.07907299425710791
	pesos_i(13550) := b"1111111111111111_1111111111111111_1111001101001001_1100110100101010"; -- -0.049655129704020674
	pesos_i(13551) := b"1111111111111111_1111111111111111_1110101110110100_1111100100010010"; -- -0.0792698222262394
	pesos_i(13552) := b"1111111111111111_1111111111111111_1111010111000100_1101010011111011"; -- -0.03996533277963225
	pesos_i(13553) := b"0000000000000000_0000000000000000_0000000011110100_0111101101100110"; -- 0.003730499566144359
	pesos_i(13554) := b"1111111111111111_1111111111111111_1111010000010110_1100010101101000"; -- -0.04652754024345225
	pesos_i(13555) := b"1111111111111111_1111111111111111_1110000101110101_1110101001010011"; -- -0.11929450476933506
	pesos_i(13556) := b"1111111111111111_1111111111111111_1110100101100101_0001011111110111"; -- -0.08830118377564113
	pesos_i(13557) := b"1111111111111111_1111111111111111_1111110000011100_1011011111111100"; -- -0.015186787663801327
	pesos_i(13558) := b"0000000000000000_0000000000000000_0001111001000001_0000010111001111"; -- 0.11817966761048254
	pesos_i(13559) := b"0000000000000000_0000000000000000_0000011101000101_1100111010000011"; -- 0.028408915544444403
	pesos_i(13560) := b"1111111111111111_1111111111111111_1111000101111101_0010010001111111"; -- -0.056684226036116406
	pesos_i(13561) := b"1111111111111111_1111111111111111_1110100111111010_1011000100101010"; -- -0.08601849299902511
	pesos_i(13562) := b"1111111111111111_1111111111111111_1111001110101100_1101001101111001"; -- -0.04814413351895566
	pesos_i(13563) := b"1111111111111111_1111111111111111_1110001011101100_1111010101101101"; -- -0.11357179722728773
	pesos_i(13564) := b"1111111111111111_1111111111111111_1111011010100100_0000101100000000"; -- -0.03655940291090474
	pesos_i(13565) := b"0000000000000000_0000000000000000_0000000100111110_1101110110010101"; -- 0.00486550221897143
	pesos_i(13566) := b"0000000000000000_0000000000000000_0001010000000111_1110111001010010"; -- 0.0782460166260681
	pesos_i(13567) := b"0000000000000000_0000000000000000_0001011101111001_0110110001101101"; -- 0.09169652626593663
	pesos_i(13568) := b"0000000000000000_0000000000000000_0010100110001100_1100010000111010"; -- 0.16230417639070163
	pesos_i(13569) := b"1111111111111111_1111111111111111_1110001011010010_1110100101011000"; -- -0.11396924581148489
	pesos_i(13570) := b"1111111111111111_1111111111111111_1110000111001000_1100000010000101"; -- -0.11803051705491104
	pesos_i(13571) := b"0000000000000000_0000000000000000_0001011110101100_1111011000001100"; -- 0.09248292720406939
	pesos_i(13572) := b"0000000000000000_0000000000000000_0001011101001101_0010000111110010"; -- 0.09102069995371409
	pesos_i(13573) := b"1111111111111111_1111111111111111_1101100001010000_0000110001001011"; -- -0.15502856407189664
	pesos_i(13574) := b"0000000000000000_0000000000000000_0000010010000001_0111010011101001"; -- 0.017600352158546124
	pesos_i(13575) := b"1111111111111111_1111111111111111_1111100011001101_0101010011011100"; -- -0.028116890315029983
	pesos_i(13576) := b"0000000000000000_0000000000000000_0010001101001011_0101010010001011"; -- 0.13786819830429117
	pesos_i(13577) := b"1111111111111111_1111111111111111_1111001011111110_0110111111101001"; -- -0.05080509722975839
	pesos_i(13578) := b"1111111111111111_1111111111111111_1110111000010111_0010001011001100"; -- -0.06995947370549305
	pesos_i(13579) := b"0000000000000000_0000000000000000_0000111001011010_0000100011100011"; -- 0.056061320685818136
	pesos_i(13580) := b"1111111111111111_1111111111111111_1110000111000001_0101111001011011"; -- -0.1181431797697398
	pesos_i(13581) := b"0000000000000000_0000000000000000_0010000101111001_1100101001011011"; -- 0.1307646247942245
	pesos_i(13582) := b"0000000000000000_0000000000000000_0001110000001001_0010101101110000"; -- 0.10951491811983474
	pesos_i(13583) := b"1111111111111111_1111111111111111_1111011111101001_1100110011101110"; -- -0.03158873740733868
	pesos_i(13584) := b"1111111111111111_1111111111111111_1110100001000101_1101011101001111"; -- -0.09268431012195136
	pesos_i(13585) := b"0000000000000000_0000000000000000_0001000110010110_1100111010110010"; -- 0.06870738835246834
	pesos_i(13586) := b"1111111111111111_1111111111111111_1111100110000000_1000010011011111"; -- -0.02538270516971716
	pesos_i(13587) := b"0000000000000000_0000000000000000_0000010111010111_1011111100001100"; -- 0.02282327694324552
	pesos_i(13588) := b"1111111111111111_1111111111111111_1101101110000101_1001111010011010"; -- -0.14249237757546235
	pesos_i(13589) := b"1111111111111111_1111111111111111_1111111010001111_0111100010010111"; -- -0.005623305416236737
	pesos_i(13590) := b"0000000000000000_0000000000000000_0001100111000010_1011000011111110"; -- 0.10062700473888964
	pesos_i(13591) := b"0000000000000000_0000000000000000_0000011001011110_1110011110010110"; -- 0.024885629753451183
	pesos_i(13592) := b"1111111111111111_1111111111111111_1111001011110101_0101110000000001"; -- -0.05094361293525018
	pesos_i(13593) := b"1111111111111111_1111111111111111_1110111001101110_0101011111001101"; -- -0.06862879989210238
	pesos_i(13594) := b"1111111111111111_1111111111111111_1111111010100100_1100000011110100"; -- -0.005298557663633499
	pesos_i(13595) := b"0000000000000000_0000000000000000_0010001100110010_0100010000100011"; -- 0.1374857507180645
	pesos_i(13596) := b"0000000000000000_0000000000000000_0001000001010000_1000111000001111"; -- 0.06372917036721426
	pesos_i(13597) := b"0000000000000000_0000000000000000_0001111100011101_0100010101001011"; -- 0.12154038506015945
	pesos_i(13598) := b"1111111111111111_1111111111111111_1111011000001011_1000011010111001"; -- -0.038886623306551606
	pesos_i(13599) := b"0000000000000000_0000000000000000_0010001111101011_1011000011010101"; -- 0.1403151054791773
	pesos_i(13600) := b"0000000000000000_0000000000000000_0000000111111010_0000000111101000"; -- 0.0077210608705153136
	pesos_i(13601) := b"1111111111111111_1111111111111111_1101100111101010_0010010100000110"; -- -0.148770986566793
	pesos_i(13602) := b"0000000000000000_0000000000000000_0001011111010010_0010001110000101"; -- 0.09305021272161162
	pesos_i(13603) := b"0000000000000000_0000000000000000_0010010110101011_0001100101111100"; -- 0.1471420218511582
	pesos_i(13604) := b"0000000000000000_0000000000000000_0000111101101111_1100001011001010"; -- 0.0602990858785975
	pesos_i(13605) := b"1111111111111111_1111111111111111_1110000010011110_0101110001000101"; -- -0.12258361168681571
	pesos_i(13606) := b"1111111111111111_1111111111111111_1111000001100010_1010000000010110"; -- -0.0609950967227682
	pesos_i(13607) := b"1111111111111111_1111111111111111_1111100101001101_0010101110001111"; -- -0.02616622690012129
	pesos_i(13608) := b"0000000000000000_0000000000000000_0000011011010001_0011000001110100"; -- 0.026629474945928495
	pesos_i(13609) := b"0000000000000000_0000000000000000_0001111001010100_0011011010111100"; -- 0.11847250060708153
	pesos_i(13610) := b"0000000000000000_0000000000000000_0001011110100100_0101010100111101"; -- 0.09235127190489312
	pesos_i(13611) := b"1111111111111111_1111111111111111_1111010000110000_1101101010100101"; -- -0.046129545941360844
	pesos_i(13612) := b"0000000000000000_0000000000000000_0000010101011101_1010001000100100"; -- 0.020959981648792467
	pesos_i(13613) := b"1111111111111111_1111111111111111_1111011010110110_1010011100000000"; -- -0.03627544638694793
	pesos_i(13614) := b"1111111111111111_1111111111111111_1111110100011001_0111110000100000"; -- -0.01132988183874002
	pesos_i(13615) := b"1111111111111111_1111111111111111_1110000000110101_1010110101101110"; -- -0.12418094693765544
	pesos_i(13616) := b"0000000000000000_0000000000000000_0001111011101100_0111001011001000"; -- 0.12079541574820292
	pesos_i(13617) := b"1111111111111111_1111111111111111_1111000101110001_0001101011101010"; -- -0.05686790274610461
	pesos_i(13618) := b"1111111111111111_1111111111111111_1111110011111010_0101010101100101"; -- -0.011805212845432803
	pesos_i(13619) := b"0000000000000000_0000000000000000_0000011000010010_1111100011000000"; -- 0.023726984843419844
	pesos_i(13620) := b"0000000000000000_0000000000000000_0000110000001100_1011001101111100"; -- 0.047068803552886805
	pesos_i(13621) := b"0000000000000000_0000000000000000_0010000100111001_1000000000101011"; -- 0.12978364046972507
	pesos_i(13622) := b"1111111111111111_1111111111111111_1111111010001001_0101010110010000"; -- -0.0057169458705776475
	pesos_i(13623) := b"0000000000000000_0000000000000000_0001000000011101_0101011011101000"; -- 0.06294768490616341
	pesos_i(13624) := b"1111111111111111_1111111111111111_1111011110111111_0110101100011101"; -- -0.03223543695066723
	pesos_i(13625) := b"0000000000000000_0000000000000000_0001110011000111_1010110010011101"; -- 0.11242178766688661
	pesos_i(13626) := b"1111111111111111_1111111111111111_1101101101010010_1001100110111001"; -- -0.14327086662714095
	pesos_i(13627) := b"1111111111111111_1111111111111111_1110001111101101_0000010011000000"; -- -0.10966463395430781
	pesos_i(13628) := b"1111111111111111_1111111111111111_1110111001101010_1011001001000101"; -- -0.06868444274935402
	pesos_i(13629) := b"0000000000000000_0000000000000000_0000010101011001_0011110011010001"; -- 0.02089290714245432
	pesos_i(13630) := b"1111111111111111_1111111111111111_1111100110010110_1011100000100110"; -- -0.02504395553656249
	pesos_i(13631) := b"1111111111111111_1111111111111111_1110110011001010_1000111010010100"; -- -0.07503422629116102
	pesos_i(13632) := b"1111111111111111_1111111111111111_1111000010011100_1000101110100110"; -- -0.06011130530656842
	pesos_i(13633) := b"1111111111111111_1111111111111111_1110100011010010_1001000011011011"; -- -0.09053702032196423
	pesos_i(13634) := b"1111111111111111_1111111111111111_1110000100101000_1000010010111010"; -- -0.12047548731528455
	pesos_i(13635) := b"0000000000000000_0000000000000000_0000011101010110_1010010101011001"; -- 0.028665861384845774
	pesos_i(13636) := b"0000000000000000_0000000000000000_0010001101010101_0001111101000101"; -- 0.13801761076467453
	pesos_i(13637) := b"0000000000000000_0000000000000000_0000101101010111_1001111110011101"; -- 0.04430577844173227
	pesos_i(13638) := b"0000000000000000_0000000000000000_0000101000111011_0110011001101011"; -- 0.039968873186310344
	pesos_i(13639) := b"0000000000000000_0000000000000000_0000011110100101_1000111110100000"; -- 0.02987001084504815
	pesos_i(13640) := b"0000000000000000_0000000000000000_0000110001111101_1110011011101111"; -- 0.048796113448804315
	pesos_i(13641) := b"1111111111111111_1111111111111111_1110001010100010_0010001011111000"; -- -0.11471349195689576
	pesos_i(13642) := b"1111111111111111_1111111111111111_1110000011010100_0110001100000000"; -- -0.12175923578901336
	pesos_i(13643) := b"0000000000000000_0000000000000000_0000001010010000_0111011010000011"; -- 0.010016829561585157
	pesos_i(13644) := b"0000000000000000_0000000000000000_0001110011000011_1010010011011100"; -- 0.11236029021022169
	pesos_i(13645) := b"0000000000000000_0000000000000000_0001010000011000_1111110001100101"; -- 0.07850625482364718
	pesos_i(13646) := b"1111111111111111_1111111111111111_1111010000111101_1110010111010011"; -- -0.045930515214659844
	pesos_i(13647) := b"0000000000000000_0000000000000000_0001000001010010_0101010011111110"; -- 0.0637562866555301
	pesos_i(13648) := b"0000000000000000_0000000000000000_0000000111100101_1100111100010101"; -- 0.007412855773247506
	pesos_i(13649) := b"0000000000000000_0000000000000000_0000001101101001_0001000111110101"; -- 0.013321993221142145
	pesos_i(13650) := b"1111111111111111_1111111111111111_1110100101101011_1000110000000011"; -- -0.08820271425874592
	pesos_i(13651) := b"0000000000000000_0000000000000000_0001101001111110_1111101100001011"; -- 0.10350007073715273
	pesos_i(13652) := b"1111111111111111_1111111111111111_1111100100011011_1110000101011011"; -- -0.026918330432836816
	pesos_i(13653) := b"1111111111111111_1111111111111111_1111011001000000_0110000100111111"; -- -0.03808014124241319
	pesos_i(13654) := b"0000000000000000_0000000000000000_0010001010100111_0101001000111000"; -- 0.13536561849704729
	pesos_i(13655) := b"1111111111111111_1111111111111111_1110001010010110_0001011010110100"; -- -0.11489732849984133
	pesos_i(13656) := b"1111111111111111_1111111111111111_1111110000011111_1111101010010111"; -- -0.01513704129498936
	pesos_i(13657) := b"1111111111111111_1111111111111111_1101111000101001_1100111111101100"; -- -0.13217449645257864
	pesos_i(13658) := b"0000000000000000_0000000000000000_0000010111111111_1100010101101100"; -- 0.02343400840998964
	pesos_i(13659) := b"1111111111111111_1111111111111111_1110000100101110_0100010011000010"; -- -0.1203877474959652
	pesos_i(13660) := b"1111111111111111_1111111111111111_1111001010111010_0010101101111101"; -- -0.05184677318669279
	pesos_i(13661) := b"0000000000000000_0000000000000000_0000110110111010_0100001100000011"; -- 0.053623378973279
	pesos_i(13662) := b"1111111111111111_1111111111111111_1101111100110010_0110110001111101"; -- -0.12813684417750007
	pesos_i(13663) := b"0000000000000000_0000000000000000_0001001110101010_1110010000101000"; -- 0.07682634333024403
	pesos_i(13664) := b"1111111111111111_1111111111111111_1111010100011110_0001111100011011"; -- -0.04250913222167889
	pesos_i(13665) := b"1111111111111111_1111111111111111_1110001011110011_1000000101101100"; -- -0.11347190009446173
	pesos_i(13666) := b"1111111111111111_1111111111111111_1110111111000001_0010000100001000"; -- -0.0634593348461233
	pesos_i(13667) := b"0000000000000000_0000000000000000_0001100001001011_1011000010010101"; -- 0.0949049343398382
	pesos_i(13668) := b"1111111111111111_1111111111111111_1111000111000000_0100100000110000"; -- -0.055659759852207495
	pesos_i(13669) := b"0000000000000000_0000000000000000_0000110010000100_1100010110001111"; -- 0.04890093565018036
	pesos_i(13670) := b"1111111111111111_1111111111111111_1110001010000110_0001000110010000"; -- -0.11514177546161843
	pesos_i(13671) := b"0000000000000000_0000000000000000_0000110001111111_1101101001101110"; -- 0.04882588557529348
	pesos_i(13672) := b"0000000000000000_0000000000000000_0000011110101110_1100000110011101"; -- 0.030010319438492274
	pesos_i(13673) := b"1111111111111111_1111111111111111_1101110010111100_0101000100000101"; -- -0.1377515184139865
	pesos_i(13674) := b"0000000000000000_0000000000000000_0000000000001100_0100000111111011"; -- 0.00018703818061689383
	pesos_i(13675) := b"0000000000000000_0000000000000000_0000111001111011_0001111010110111"; -- 0.056566161875348284
	pesos_i(13676) := b"1111111111111111_1111111111111111_1110111011110110_0110100001101110"; -- -0.0665526134760633
	pesos_i(13677) := b"1111111111111111_1111111111111111_1110001100100010_1000110111111100"; -- -0.112753988358309
	pesos_i(13678) := b"0000000000000000_0000000000000000_0001000001111010_0000100111111000"; -- 0.0643621665126604
	pesos_i(13679) := b"0000000000000000_0000000000000000_0010000010010110_1100110110101010"; -- 0.1273010768237202
	pesos_i(13680) := b"0000000000000000_0000000000000000_0001000011110000_1101011001001010"; -- 0.0661748820131563
	pesos_i(13681) := b"1111111111111111_1111111111111111_1101110111000000_0011000100100101"; -- -0.13378613326753827
	pesos_i(13682) := b"0000000000000000_0000000000000000_0000101100010000_1010010000110001"; -- 0.04322267725133423
	pesos_i(13683) := b"1111111111111111_1111111111111111_1111110111011111_0101111101101000"; -- -0.008310353377468167
	pesos_i(13684) := b"1111111111111111_1111111111111111_1111011000011110_0000001101101110"; -- -0.03860453179180427
	pesos_i(13685) := b"1111111111111111_1111111111111111_1101101110100101_1111000110101011"; -- -0.14199914532719704
	pesos_i(13686) := b"0000000000000000_0000000000000000_0000101000000001_0111101000101000"; -- 0.03908503987167745
	pesos_i(13687) := b"1111111111111111_1111111111111111_1110010111001100_1001011010001111"; -- -0.10234698298168848
	pesos_i(13688) := b"0000000000000000_0000000000000000_0000001100110000_0001111111001001"; -- 0.012453066329933562
	pesos_i(13689) := b"1111111111111111_1111111111111111_1110000010100011_0001001111111001"; -- -0.12251162696759443
	pesos_i(13690) := b"1111111111111111_1111111111111111_1110111001000011_0100101001111010"; -- -0.06928572209345209
	pesos_i(13691) := b"1111111111111111_1111111111111111_1111000011010011_1001100011100000"; -- -0.05927128353541661
	pesos_i(13692) := b"1111111111111111_1111111111111111_1101110010100101_0010000010010100"; -- -0.13810535790047135
	pesos_i(13693) := b"1111111111111111_1111111111111111_1101101010001100_0111001110000000"; -- -0.14629438508922965
	pesos_i(13694) := b"0000000000000000_0000000000000000_0000011011100110_1011001001100010"; -- 0.026957654037948805
	pesos_i(13695) := b"1111111111111111_1111111111111111_1111010011001100_0111010000111101"; -- -0.04375527872753025
	pesos_i(13696) := b"1111111111111111_1111111111111111_1111011100001000_0110101111011101"; -- -0.03502775047078328
	pesos_i(13697) := b"1111111111111111_1111111111111111_1110001101110001_1101011011000101"; -- -0.11154420555817503
	pesos_i(13698) := b"0000000000000000_0000000000000000_0000011010010100_1101110110000000"; -- 0.02570900315033978
	pesos_i(13699) := b"0000000000000000_0000000000000000_0001101101000101_0000010111010011"; -- 0.1065219535869721
	pesos_i(13700) := b"0000000000000000_0000000000000000_0001001101000101_1101110011010111"; -- 0.075284769523838
	pesos_i(13701) := b"1111111111111111_1111111111111111_1111111101111101_1000110000100101"; -- -0.0019905481627107563
	pesos_i(13702) := b"0000000000000000_0000000000000000_0010000011000001_0010000011111100"; -- 0.1279469123874257
	pesos_i(13703) := b"1111111111111111_1111111111111111_1101111101010110_0100000110011010"; -- -0.1275900838707107
	pesos_i(13704) := b"1111111111111111_1111111111111111_1111110010101101_0101001111111111"; -- -0.012980222883149335
	pesos_i(13705) := b"1111111111111111_1111111111111111_1111100000000000_0101001000100110"; -- -0.031245103637016353
	pesos_i(13706) := b"1111111111111111_1111111111111111_1110100111000110_0001101011000101"; -- -0.08682091427043262
	pesos_i(13707) := b"0000000000000000_0000000000000000_0000000101000100_0101100111000011"; -- 0.004949197834451649
	pesos_i(13708) := b"1111111111111111_1111111111111111_1110101001011110_1001110011001110"; -- -0.0844938275689256
	pesos_i(13709) := b"1111111111111111_1111111111111111_1111111100010011_0110011011000001"; -- -0.0036102083642445496
	pesos_i(13710) := b"1111111111111111_1111111111111111_1111011110100101_1001110001100101"; -- -0.032629228057490606
	pesos_i(13711) := b"0000000000000000_0000000000000000_0001100111001000_0001111011000110"; -- 0.10070984202132773
	pesos_i(13712) := b"0000000000000000_0000000000000000_0000010111111101_0011001110111101"; -- 0.02339480740275189
	pesos_i(13713) := b"1111111111111111_1111111111111111_1110011010100100_0000100000001111"; -- -0.09905957830821738
	pesos_i(13714) := b"0000000000000000_0000000000000000_0000001110011100_0111001100011001"; -- 0.014105981453221282
	pesos_i(13715) := b"1111111111111111_1111111111111111_1111000000010110_1001011110100000"; -- -0.06215526919916097
	pesos_i(13716) := b"1111111111111111_1111111111111111_1110010110110010_0001001011100001"; -- -0.10275156038865475
	pesos_i(13717) := b"1111111111111111_1111111111111111_1111010111000101_0110100110100101"; -- -0.03995647171325675
	pesos_i(13718) := b"0000000000000000_0000000000000000_0001100111110011_0001110111011101"; -- 0.10136591575078874
	pesos_i(13719) := b"1111111111111111_1111111111111111_1110000010111001_1010010101100100"; -- -0.12216726586097792
	pesos_i(13720) := b"0000000000000000_0000000000000000_0001101101100000_0011001001111001"; -- 0.1069366021075131
	pesos_i(13721) := b"1111111111111111_1111111111111111_1101101110001101_0010010000101111"; -- -0.1423776039285669
	pesos_i(13722) := b"0000000000000000_0000000000000000_0000111001010001_0100011000110111"; -- 0.055927646997966325
	pesos_i(13723) := b"0000000000000000_0000000000000000_0001011000010100_1100000110110001"; -- 0.08625422068946494
	pesos_i(13724) := b"0000000000000000_0000000000000000_0001001110111000_0101101111111100"; -- 0.07703184978618774
	pesos_i(13725) := b"0000000000000000_0000000000000000_0000110110101110_1010110011010001"; -- 0.05344658001874331
	pesos_i(13726) := b"1111111111111111_1111111111111111_1111111110010101_1001101010001000"; -- -0.001623479703403421
	pesos_i(13727) := b"1111111111111111_1111111111111111_1111110010111110_0110001010101011"; -- -0.012719948934028263
	pesos_i(13728) := b"0000000000000000_0000000000000000_0000100011010001_1111000110010111"; -- 0.034453486763610534
	pesos_i(13729) := b"1111111111111111_1111111111111111_1110100000110100_1010000001101100"; -- -0.09294698117272505
	pesos_i(13730) := b"1111111111111111_1111111111111111_1110111001111110_1000001010000010"; -- -0.0683821137515226
	pesos_i(13731) := b"0000000000000000_0000000000000000_0001011010110000_0000100011111110"; -- 0.08862358276836439
	pesos_i(13732) := b"0000000000000000_0000000000000000_0010010010011010_1100010000110101"; -- 0.142986548474864
	pesos_i(13733) := b"1111111111111111_1111111111111111_1111100101010100_1110111110011011"; -- -0.026047730113011175
	pesos_i(13734) := b"0000000000000000_0000000000000000_0010000110101001_0110000011101000"; -- 0.13149076144352762
	pesos_i(13735) := b"1111111111111111_1111111111111111_1110100001010100_0000100001010000"; -- -0.09246776622168598
	pesos_i(13736) := b"1111111111111111_1111111111111111_1111001000100101_1100101100001101"; -- -0.054110822054957125
	pesos_i(13737) := b"1111111111111111_1111111111111111_1110100101111010_1001111000000000"; -- -0.08797276016572647
	pesos_i(13738) := b"1111111111111111_1111111111111111_1110011000111011_1010110110111011"; -- -0.10065187624946292
	pesos_i(13739) := b"0000000000000000_0000000000000000_0001011010000100_1111110011101101"; -- 0.08796673581420482
	pesos_i(13740) := b"1111111111111111_1111111111111111_1110000111001011_0111110110101100"; -- -0.11798872517680525
	pesos_i(13741) := b"0000000000000000_0000000000000000_0000111111110100_0001111010001111"; -- 0.062318716048418474
	pesos_i(13742) := b"0000000000000000_0000000000000000_0001001001100001_1011000100000000"; -- 0.07180315260787701
	pesos_i(13743) := b"0000000000000000_0000000000000000_0000000011010000_1001000011000011"; -- 0.0031824565949219587
	pesos_i(13744) := b"1111111111111111_1111111111111111_1111110110101011_1111111010111100"; -- -0.00909431361125465
	pesos_i(13745) := b"0000000000000000_0000000000000000_0000010010101100_0011011010001000"; -- 0.01825276198140938
	pesos_i(13746) := b"1111111111111111_1111111111111111_1110001011101011_0110110100001100"; -- -0.11359518497180705
	pesos_i(13747) := b"0000000000000000_0000000000000000_0000101001111100_0101001110100100"; -- 0.040959575249035825
	pesos_i(13748) := b"1111111111111111_1111111111111111_1111100110000100_1001000000001101"; -- -0.025321003787162583
	pesos_i(13749) := b"0000000000000000_0000000000000000_0010001011010100_0011010001000010"; -- 0.13605047803513304
	pesos_i(13750) := b"1111111111111111_1111111111111111_1110010101111000_1101011010101111"; -- -0.1036248991368028
	pesos_i(13751) := b"1111111111111111_1111111111111111_1111010000000011_1110101100010110"; -- -0.04681521145207713
	pesos_i(13752) := b"0000000000000000_0000000000000000_0000010010111000_0010000111001111"; -- 0.01843463236071433
	pesos_i(13753) := b"0000000000000000_0000000000000000_0000001001011101_0100101100011111"; -- 0.009236045031067506
	pesos_i(13754) := b"0000000000000000_0000000000000000_0001101000110101_0110010011111111"; -- 0.10237723559144912
	pesos_i(13755) := b"0000000000000000_0000000000000000_0001000001101011_1010101110000101"; -- 0.06414291388426133
	pesos_i(13756) := b"0000000000000000_0000000000000000_0000011010011011_0010110110101001"; -- 0.02580533379233881
	pesos_i(13757) := b"0000000000000000_0000000000000000_0000110001110110_1110010010000000"; -- 0.048689156730317394
	pesos_i(13758) := b"1111111111111111_1111111111111111_1110111111110010_1011000011010011"; -- -0.06270308353968873
	pesos_i(13759) := b"0000000000000000_0000000000000000_0001011100101011_1000100001110100"; -- 0.09050801126344614
	pesos_i(13760) := b"1111111111111111_1111111111111111_1110101010100111_0000100111110011"; -- -0.08338868917740583
	pesos_i(13761) := b"1111111111111111_1111111111111111_1101011011000001_1110011000001110"; -- -0.16110384134272676
	pesos_i(13762) := b"1111111111111111_1111111111111111_1111000101010110_1001110110001000"; -- -0.05727210444105317
	pesos_i(13763) := b"1111111111111111_1111111111111111_1110111110110011_0000110100100011"; -- -0.06367414380558516
	pesos_i(13764) := b"0000000000000000_0000000000000000_0001101100001010_0110101001100001"; -- 0.10562767862295783
	pesos_i(13765) := b"1111111111111111_1111111111111111_1111001000010100_1101011010100010"; -- -0.054369531147613656
	pesos_i(13766) := b"1111111111111111_1111111111111111_1110111011001000_1001000001000011"; -- -0.06725214361411297
	pesos_i(13767) := b"0000000000000000_0000000000000000_0000101100101001_0010110101110000"; -- 0.04359706854155313
	pesos_i(13768) := b"1111111111111111_1111111111111111_1110111001010101_1011001011111110"; -- -0.06900483418937095
	pesos_i(13769) := b"0000000000000000_0000000000000000_0001000010111000_0001010001110110"; -- 0.06530883675168449
	pesos_i(13770) := b"0000000000000000_0000000000000000_0000111100111000_1001100110100110"; -- 0.05945740043392687
	pesos_i(13771) := b"0000000000000000_0000000000000000_0000010000001111_0101000110101010"; -- 0.015858749352566724
	pesos_i(13772) := b"1111111111111111_1111111111111111_1110010011100010_0001100110000001"; -- -0.1059249936217082
	pesos_i(13773) := b"1111111111111111_1111111111111111_1111110001111001_0011000100110011"; -- -0.013775753992842085
	pesos_i(13774) := b"0000000000000000_0000000000000000_0000010010001111_1001001100000001"; -- 0.01781576892469797
	pesos_i(13775) := b"1111111111111111_1111111111111111_1110100110110111_0111010111000111"; -- -0.0870443714484173
	pesos_i(13776) := b"0000000000000000_0000000000000000_0001011001001101_1011000010001001"; -- 0.08712294903580504
	pesos_i(13777) := b"1111111111111111_1111111111111111_1110000111100010_0001111010100011"; -- -0.11764343758404157
	pesos_i(13778) := b"1111111111111111_1111111111111111_1110110000011011_1110100000101100"; -- -0.0776991742461452
	pesos_i(13779) := b"0000000000000000_0000000000000000_0000110111110111_0001010111011001"; -- 0.054551473123878334
	pesos_i(13780) := b"0000000000000000_0000000000000000_0000000000101011_1110011100010110"; -- 0.0006699017957035725
	pesos_i(13781) := b"0000000000000000_0000000000000000_0000110110111000_1100001010111110"; -- 0.053600474715717966
	pesos_i(13782) := b"0000000000000000_0000000000000000_0010010001101100_1110000101000000"; -- 0.14228637523294357
	pesos_i(13783) := b"0000000000000000_0000000000000000_0001001010110011_0010111011100001"; -- 0.07304661735733817
	pesos_i(13784) := b"0000000000000000_0000000000000000_0001100011011001_0010111010000111"; -- 0.0970639305347534
	pesos_i(13785) := b"1111111111111111_1111111111111111_1111100100110000_1000011000001111"; -- -0.026603337597923674
	pesos_i(13786) := b"0000000000000000_0000000000000000_0001000111010001_0000100100001110"; -- 0.06959587663651397
	pesos_i(13787) := b"0000000000000000_0000000000000000_0010011010000000_1111011110100001"; -- 0.1504053847445051
	pesos_i(13788) := b"0000000000000000_0000000000000000_0001111010000001_1001101001001001"; -- 0.11916507993982395
	pesos_i(13789) := b"1111111111111111_1111111111111111_1111001010110000_0000011101010010"; -- -0.05200151683046355
	pesos_i(13790) := b"0000000000000000_0000000000000000_0000000101000110_1110001100011101"; -- 0.004987902347162797
	pesos_i(13791) := b"0000000000000000_0000000000000000_0000001101111010_1110010110001100"; -- 0.013594004425166494
	pesos_i(13792) := b"0000000000000000_0000000000000000_0010001000110000_0110000000111000"; -- 0.13355065684538248
	pesos_i(13793) := b"0000000000000000_0000000000000000_0001011001001000_0001011001111000"; -- 0.08703747200845449
	pesos_i(13794) := b"1111111111111111_1111111111111111_1101101010010101_1100011011101101"; -- -0.14615208361137558
	pesos_i(13795) := b"0000000000000000_0000000000000000_0010011010010111_0110100110000110"; -- 0.15074786684412958
	pesos_i(13796) := b"0000000000000000_0000000000000000_0000010111101010_1110011011001101"; -- 0.023115563516280344
	pesos_i(13797) := b"1111111111111111_1111111111111111_1111100110111110_0101100100010100"; -- -0.02443927064552779
	pesos_i(13798) := b"1111111111111111_1111111111111111_1101111011001100_0000100110001100"; -- -0.12969913809100142
	pesos_i(13799) := b"0000000000000000_0000000000000000_0001111101011000_1111001001100010"; -- 0.12245097067220509
	pesos_i(13800) := b"0000000000000000_0000000000000000_0000100101110010_0101111111010110"; -- 0.03690146412852396
	pesos_i(13801) := b"0000000000000000_0000000000000000_0000001010101011_0000000010111010"; -- 0.010421796127557923
	pesos_i(13802) := b"1111111111111111_1111111111111111_1111001000100100_1011001111111000"; -- -0.054127456627492625
	pesos_i(13803) := b"1111111111111111_1111111111111111_1111011100111101_1011110000000110"; -- -0.034214256759636706
	pesos_i(13804) := b"0000000000000000_0000000000000000_0001000110111101_1101010000111000"; -- 0.06930281041735095
	pesos_i(13805) := b"0000000000000000_0000000000000000_0000010101000011_1000011110011001"; -- 0.020561671196416158
	pesos_i(13806) := b"0000000000000000_0000000000000000_0001000111110010_1000011011011001"; -- 0.07010691458853116
	pesos_i(13807) := b"0000000000000000_0000000000000000_0010000010110000_0011011000101110"; -- 0.12768877613725782
	pesos_i(13808) := b"1111111111111111_1111111111111111_1110101110101011_1010101110001001"; -- -0.07941177270495596
	pesos_i(13809) := b"1111111111111111_1111111111111111_1111101101100111_0100000101110000"; -- -0.017955694435361668
	pesos_i(13810) := b"0000000000000000_0000000000000000_0010010000111100_0101110101001110"; -- 0.14154608882074757
	pesos_i(13811) := b"1111111111111111_1111111111111111_1111011011000100_0110111000000101"; -- -0.036065219566725586
	pesos_i(13812) := b"0000000000000000_0000000000000000_0001100011100111_0011010101011100"; -- 0.09727796073645514
	pesos_i(13813) := b"1111111111111111_1111111111111111_1110010011010011_1000100000000101"; -- -0.10614728803679978
	pesos_i(13814) := b"0000000000000000_0000000000000000_0010010000010101_0001011001000010"; -- 0.14094676132597433
	pesos_i(13815) := b"0000000000000000_0000000000000000_0000001001100101_1101100011111011"; -- 0.009366570644049655
	pesos_i(13816) := b"0000000000000000_0000000000000000_0000110010101100_1100010111000111"; -- 0.04951130019908627
	pesos_i(13817) := b"0000000000000000_0000000000000000_0001100000101100_1001101100011100"; -- 0.09443063195784218
	pesos_i(13818) := b"0000000000000000_0000000000000000_0010011001001011_0101100100111111"; -- 0.14958722857666695
	pesos_i(13819) := b"1111111111111111_1111111111111111_1101110001000111_1000011100001110"; -- -0.13953357599684962
	pesos_i(13820) := b"0000000000000000_0000000000000000_0010000110111011_1010011100111011"; -- 0.13176961115713456
	pesos_i(13821) := b"1111111111111111_1111111111111111_1111110100010101_0111000010010110"; -- -0.011391604670924201
	pesos_i(13822) := b"0000000000000000_0000000000000000_0001010100110001_1011010000110101"; -- 0.08278967189741072
	pesos_i(13823) := b"1111111111111111_1111111111111111_1110001101000010_0010101101110111"; -- -0.11227157927693474
	pesos_i(13824) := b"0000000000000000_0000000000000000_0001100100011100_0011110100111000"; -- 0.09808714509259096
	pesos_i(13825) := b"0000000000000000_0000000000000000_0000011011100110_1100101100101110"; -- 0.026959131859846223
	pesos_i(13826) := b"1111111111111111_1111111111111111_1110001011001111_0111000101100001"; -- -0.11402217282209097
	pesos_i(13827) := b"0000000000000000_0000000000000000_0000000010001100_1100101101100100"; -- 0.0021483535753019194
	pesos_i(13828) := b"0000000000000000_0000000000000000_0001000100110111_0001111000011110"; -- 0.06724727856549745
	pesos_i(13829) := b"1111111111111111_1111111111111111_1111101101001101_0001000110110110"; -- -0.018355267565282572
	pesos_i(13830) := b"0000000000000000_0000000000000000_0010011010101111_1000000011010101"; -- 0.15111546715084392
	pesos_i(13831) := b"0000000000000000_0000000000000000_0010001111101111_1011001110101011"; -- 0.1403763095404574
	pesos_i(13832) := b"0000000000000000_0000000000000000_0000011100100011_0111101000010100"; -- 0.02788508400511063
	pesos_i(13833) := b"0000000000000000_0000000000000000_0010001110000000_0101100000011100"; -- 0.13867712662814094
	pesos_i(13834) := b"1111111111111111_1111111111111111_1111110011011001_1101100010110010"; -- -0.012300926681833269
	pesos_i(13835) := b"1111111111111111_1111111111111111_1111010001100110_0011001101110000"; -- -0.04531553758012429
	pesos_i(13836) := b"0000000000000000_0000000000000000_0001010101011101_1010011100000111"; -- 0.08346027294474033
	pesos_i(13837) := b"0000000000000000_0000000000000000_0010001101101100_0011000101111101"; -- 0.13836964895483608
	pesos_i(13838) := b"0000000000000000_0000000000000000_0001101000001011_0101001101110100"; -- 0.10173532088841883
	pesos_i(13839) := b"0000000000000000_0000000000000000_0000111110100011_1100001111100010"; -- 0.0610926081929966
	pesos_i(13840) := b"1111111111111111_1111111111111111_1110101110101001_1000010100101100"; -- -0.07944457709741887
	pesos_i(13841) := b"1111111111111111_1111111111111111_1101111001111111_0001100100110101"; -- -0.13087313131743283
	pesos_i(13842) := b"1111111111111111_1111111111111111_1111110111001000_1000110001010111"; -- -0.008658627203389106
	pesos_i(13843) := b"1111111111111111_1111111111111111_1111101000010011_0010101111110010"; -- -0.02314496357890534
	pesos_i(13844) := b"0000000000000000_0000000000000000_0001100011111001_1101011011001011"; -- 0.09756224104475476
	pesos_i(13845) := b"1111111111111111_1111111111111111_1110100001001011_0101010011000010"; -- -0.09260053875433773
	pesos_i(13846) := b"1111111111111111_1111111111111111_1110011000101010_0010001111110101"; -- -0.10091948754651331
	pesos_i(13847) := b"0000000000000000_0000000000000000_0000110100001100_1111111010000000"; -- 0.05097952492529349
	pesos_i(13848) := b"0000000000000000_0000000000000000_0010011011100000_0000101011111000"; -- 0.1518561224584457
	pesos_i(13849) := b"1111111111111111_1111111111111111_1110110101101011_1101101011001001"; -- -0.07257301897045698
	pesos_i(13850) := b"0000000000000000_0000000000000000_0001100000010100_0110110000100001"; -- 0.09406162084766624
	pesos_i(13851) := b"1111111111111111_1111111111111111_1110010000001101_1111110010101001"; -- -0.1091615759570535
	pesos_i(13852) := b"1111111111111111_1111111111111111_1101111001010000_0100001100010101"; -- -0.13158779844746507
	pesos_i(13853) := b"1111111111111111_1111111111111111_1110001010011110_0111000011011101"; -- -0.1147698841751187
	pesos_i(13854) := b"1111111111111111_1111111111111111_1111001111110111_1100100111111111"; -- -0.04700028927846873
	pesos_i(13855) := b"1111111111111111_1111111111111111_1111100011111101_1001110111110100"; -- -0.027380111684626496
	pesos_i(13856) := b"1111111111111111_1111111111111111_1101111100010100_1101011100011110"; -- -0.12858825214406083
	pesos_i(13857) := b"0000000000000000_0000000000000000_0010000100101110_0111000000111010"; -- 0.12961484360423287
	pesos_i(13858) := b"1111111111111111_1111111111111111_1111011110000111_0111001000010010"; -- -0.03308951433302263
	pesos_i(13859) := b"1111111111111111_1111111111111111_1111110000101110_1000110101101001"; -- -0.014914667093243256
	pesos_i(13860) := b"1111111111111111_1111111111111111_1110111011000110_0110110101001010"; -- -0.06728474565917451
	pesos_i(13861) := b"1111111111111111_1111111111111111_1111110011011101_1100001001100000"; -- -0.012241222025060538
	pesos_i(13862) := b"0000000000000000_0000000000000000_0000101001101111_1110110111101111"; -- 0.040770407430339925
	pesos_i(13863) := b"1111111111111111_1111111111111111_1111000000110001_0100111001101010"; -- -0.061747645598999354
	pesos_i(13864) := b"1111111111111111_1111111111111111_1111111000011001_0011100111110100"; -- -0.007427575932994702
	pesos_i(13865) := b"0000000000000000_0000000000000000_0010001001010100_0101000001101111"; -- 0.13409903240518853
	pesos_i(13866) := b"0000000000000000_0000000000000000_0001000101001000_1111111100000010"; -- 0.06752008252546204
	pesos_i(13867) := b"1111111111111111_1111111111111111_1101111011000011_0001010001010010"; -- -0.1298358250166745
	pesos_i(13868) := b"0000000000000000_0000000000000000_0001011001100111_1010011001100001"; -- 0.08751907212349214
	pesos_i(13869) := b"1111111111111111_1111111111111111_1111011011010110_0100101001101001"; -- -0.035792683926843254
	pesos_i(13870) := b"0000000000000000_0000000000000000_0001011111001001_0101101101001100"; -- 0.09291620824350721
	pesos_i(13871) := b"0000000000000000_0000000000000000_0000001100111111_1111100011110100"; -- 0.012694892480559966
	pesos_i(13872) := b"0000000000000000_0000000000000000_0010011110110100_0100110111010100"; -- 0.15509497088516133
	pesos_i(13873) := b"1111111111111111_1111111111111111_1110100110011110_0000111111011111"; -- -0.08743191535262636
	pesos_i(13874) := b"0000000000000000_0000000000000000_0001111011110000_1001011001001010"; -- 0.12085856740419545
	pesos_i(13875) := b"1111111111111111_1111111111111111_1111011101111110_0011010011111101"; -- -0.03323048421528183
	pesos_i(13876) := b"1111111111111111_1111111111111111_1111011001101011_1111000111000011"; -- -0.03741539933898768
	pesos_i(13877) := b"0000000000000000_0000000000000000_0001010010001101_0101111010111110"; -- 0.08028213644406118
	pesos_i(13878) := b"0000000000000000_0000000000000000_0001010101110110_0000110100010011"; -- 0.08383256641582018
	pesos_i(13879) := b"1111111111111111_1111111111111111_1110100010000001_1101111111111001"; -- -0.09176826646990122
	pesos_i(13880) := b"1111111111111111_1111111111111111_1101110011111010_0010100011000110"; -- -0.13680787246171278
	pesos_i(13881) := b"1111111111111111_1111111111111111_1110111001000100_1000000101111111"; -- -0.06926718387375315
	pesos_i(13882) := b"0000000000000000_0000000000000000_0000111111100111_0001001111000100"; -- 0.062119708384727974
	pesos_i(13883) := b"1111111111111111_1111111111111111_1111111001000111_1011110000000011"; -- -0.0067179195366125115
	pesos_i(13884) := b"0000000000000000_0000000000000000_0001000001000000_0110001110010101"; -- 0.06348249797816183
	pesos_i(13885) := b"1111111111111111_1111111111111111_1111111000010001_1111100100111110"; -- -0.007538244700948085
	pesos_i(13886) := b"1111111111111111_1111111111111111_1111110000010000_0110101001111100"; -- -0.01537451245224816
	pesos_i(13887) := b"0000000000000000_0000000000000000_0010010001000101_0011011001100101"; -- 0.14168109872807932
	pesos_i(13888) := b"0000000000000000_0000000000000000_0001001110100001_0101111010011100"; -- 0.07668105426875578
	pesos_i(13889) := b"0000000000000000_0000000000000000_0000100010100001_1011000011011100"; -- 0.0337172067680917
	pesos_i(13890) := b"0000000000000000_0000000000000000_0000110001000011_1010000010010101"; -- 0.04790691034309948
	pesos_i(13891) := b"1111111111111111_1111111111111111_1110000111111010_1011110001110110"; -- -0.11726781961241947
	pesos_i(13892) := b"1111111111111111_1111111111111111_1110100010110101_1101111000011010"; -- -0.09097492087123339
	pesos_i(13893) := b"0000000000000000_0000000000000000_0001101101111000_1000010111110001"; -- 0.10730778830799727
	pesos_i(13894) := b"1111111111111111_1111111111111111_1101000101011111_1000110110111001"; -- -0.18213571769585826
	pesos_i(13895) := b"1111111111111111_1111111111111111_1110001000010100_0000010100000100"; -- -0.11688202533439669
	pesos_i(13896) := b"1111111111111111_1111111111111111_1110100100010011_0001110001011010"; -- -0.08955214321160422
	pesos_i(13897) := b"1111111111111111_1111111111111111_1110010110111010_1110001011110001"; -- -0.1026170884910577
	pesos_i(13898) := b"1111111111111111_1111111111111111_1111110111000000_1011001010011100"; -- -0.0087784165839228
	pesos_i(13899) := b"0000000000000000_0000000000000000_0010001101110110_0110100110111110"; -- 0.13852558987607544
	pesos_i(13900) := b"1111111111111111_1111111111111111_1110100010001111_0101100100101111"; -- -0.09156267748796545
	pesos_i(13901) := b"1111111111111111_1111111111111111_1110110011111010_1100100011110111"; -- -0.07429832435142686
	pesos_i(13902) := b"1111111111111111_1111111111111111_1101101011010101_0010011001010100"; -- -0.145185093461198
	pesos_i(13903) := b"1111111111111111_1111111111111111_1110010010110011_1001111111011000"; -- -0.10663414922791113
	pesos_i(13904) := b"1111111111111111_1111111111111111_1111110001100000_0101101100111011"; -- -0.014154718518358894
	pesos_i(13905) := b"0000000000000000_0000000000000000_0010011101010100_0100110100001100"; -- 0.15363008053699717
	pesos_i(13906) := b"1111111111111111_1111111111111111_1111110101011011_0101111101000011"; -- -0.01032452212446073
	pesos_i(13907) := b"1111111111111111_1111111111111111_1101111001011011_1001010111001001"; -- -0.13141502233354874
	pesos_i(13908) := b"1111111111111111_1111111111111111_1101111110100111_1110110110100010"; -- -0.1263438682038786
	pesos_i(13909) := b"0000000000000000_0000000000000000_0000111001100111_1100101111111001"; -- 0.056271313023150665
	pesos_i(13910) := b"0000000000000000_0000000000000000_0000110110011010_1111001100100010"; -- 0.05314559539360975
	pesos_i(13911) := b"1111111111111111_1111111111111111_1101110110101100_1110010010110010"; -- -0.13408060698614618
	pesos_i(13912) := b"1111111111111111_1111111111111111_1111111010111101_0101101010111110"; -- -0.004923180118636118
	pesos_i(13913) := b"0000000000000000_0000000000000000_0000111011111100_1110010011000011"; -- 0.058546350167547966
	pesos_i(13914) := b"0000000000000000_0000000000000000_0000011011000011_1101110110111100"; -- 0.02642618017879569
	pesos_i(13915) := b"1111111111111111_1111111111111111_1110000111101010_1011001000001010"; -- -0.11751258135654635
	pesos_i(13916) := b"1111111111111111_1111111111111111_1110101101010101_1011100100111101"; -- -0.08072321190816421
	pesos_i(13917) := b"0000000000000000_0000000000000000_0000101110011000_0101011101011001"; -- 0.04529329230072903
	pesos_i(13918) := b"0000000000000000_0000000000000000_0001000010110111_1111100111001010"; -- 0.06530724690620707
	pesos_i(13919) := b"1111111111111111_1111111111111111_1101111111101111_1010000001110100"; -- -0.12524983577059662
	pesos_i(13920) := b"0000000000000000_0000000000000000_0001000101000101_1110100111111010"; -- 0.06747305257667595
	pesos_i(13921) := b"0000000000000000_0000000000000000_0001101110110101_0110001011011010"; -- 0.10823648278112886
	pesos_i(13922) := b"0000000000000000_0000000000000000_0000110111101000_1010101111110101"; -- 0.05433153849888838
	pesos_i(13923) := b"0000000000000000_0000000000000000_0000111001111110_0100000000001111"; -- 0.056613925611685184
	pesos_i(13924) := b"0000000000000000_0000000000000000_0001100101000111_1110010100101000"; -- 0.09875328275434199
	pesos_i(13925) := b"1111111111111111_1111111111111111_1111101100111010_0000111001010111"; -- -0.01864538558880732
	pesos_i(13926) := b"0000000000000000_0000000000000000_0000101001001011_0011010000101110"; -- 0.04021001925341065
	pesos_i(13927) := b"0000000000000000_0000000000000000_0001010101011011_0101100101100110"; -- 0.08342512845198678
	pesos_i(13928) := b"0000000000000000_0000000000000000_0001111010000010_0111000111110011"; -- 0.11917793443272764
	pesos_i(13929) := b"1111111111111111_1111111111111111_1111111010101001_1110000100000000"; -- -0.005220353594345984
	pesos_i(13930) := b"1111111111111111_1111111111111111_1101101101011111_1111001010011110"; -- -0.14306720400306738
	pesos_i(13931) := b"0000000000000000_0000000000000000_0001110110111100_0001000111011100"; -- 0.116150966810188
	pesos_i(13932) := b"0000000000000000_0000000000000000_0000000010101101_1101010111000010"; -- 0.0026525114602819746
	pesos_i(13933) := b"1111111111111111_1111111111111111_1101110111011001_0000101101011000"; -- -0.13340691665256083
	pesos_i(13934) := b"0000000000000000_0000000000000000_0010011000010100_1010000110000110"; -- 0.14875230342381857
	pesos_i(13935) := b"0000000000000000_0000000000000000_0000011010010100_0111001001110101"; -- 0.025702623062728976
	pesos_i(13936) := b"1111111111111111_1111111111111111_1110001000001010_0011100001000111"; -- -0.11703155774502398
	pesos_i(13937) := b"1111111111111111_1111111111111111_1101101000110011_0011110000000111"; -- -0.14765572392428775
	pesos_i(13938) := b"1111111111111111_1111111111111111_1110100000001010_1110110001011011"; -- -0.09358332425191843
	pesos_i(13939) := b"0000000000000000_0000000000000000_0000000011010101_0110011111010111"; -- 0.0032563114957152293
	pesos_i(13940) := b"0000000000000000_0000000000000000_0001001111101110_1010101111011111"; -- 0.07786058612058944
	pesos_i(13941) := b"1111111111111111_1111111111111111_1110000101010010_1010011100101101"; -- -0.11983256480415935
	pesos_i(13942) := b"1111111111111111_1111111111111111_1111000101010110_0001110010101011"; -- -0.057279785507386084
	pesos_i(13943) := b"0000000000000000_0000000000000000_0001010010011000_0001010000001111"; -- 0.08044553159916075
	pesos_i(13944) := b"1111111111111111_1111111111111111_1110010000111011_1001010000100111"; -- -0.10846590098440623
	pesos_i(13945) := b"0000000000000000_0000000000000000_0000000011100111_0111110110000001"; -- 0.0035322608899036553
	pesos_i(13946) := b"0000000000000000_0000000000000000_0010010110100011_1010010010101001"; -- 0.14702824722945976
	pesos_i(13947) := b"1111111111111111_1111111111111111_1111110111110100_1111010001011011"; -- -0.007981040736885275
	pesos_i(13948) := b"0000000000000000_0000000000000000_0001001011010000_1101111100000110"; -- 0.073499621277809
	pesos_i(13949) := b"0000000000000000_0000000000000000_0010001000100101_1010100111001111"; -- 0.13338719664503976
	pesos_i(13950) := b"1111111111111111_1111111111111111_1110011100100101_0001000100110110"; -- -0.09709064888759197
	pesos_i(13951) := b"1111111111111111_1111111111111111_1110000100011111_1101101110011100"; -- -0.12060763785804345
	pesos_i(13952) := b"0000000000000000_0000000000000000_0001101000101110_0111001010010111"; -- 0.10227123449062073
	pesos_i(13953) := b"1111111111111111_1111111111111111_1101101001001101_1000011110010100"; -- -0.1472544922535862
	pesos_i(13954) := b"1111111111111111_1111111111111111_1110111100100011_0110010000010010"; -- -0.06586622762515808
	pesos_i(13955) := b"0000000000000000_0000000000000000_0010010010111101_1001010100110101"; -- 0.14351780447803952
	pesos_i(13956) := b"1111111111111111_1111111111111111_1111001010100011_0101011101100111"; -- -0.052195107697408726
	pesos_i(13957) := b"0000000000000000_0000000000000000_0001111011110010_0110110000101001"; -- 0.120886573908111
	pesos_i(13958) := b"0000000000000000_0000000000000000_0001000111010000_1111001101000001"; -- 0.0695945771695958
	pesos_i(13959) := b"1111111111111111_1111111111111111_1111101000001000_1101001011000111"; -- -0.02330286646966768
	pesos_i(13960) := b"1111111111111111_1111111111111111_1110010011010001_0101010011001010"; -- -0.1061808591993189
	pesos_i(13961) := b"0000000000000000_0000000000000000_0000000100001110_0011110111000011"; -- 0.004123554271627171
	pesos_i(13962) := b"0000000000000000_0000000000000000_0001111111011111_0100100001011101"; -- 0.12450077322691015
	pesos_i(13963) := b"0000000000000000_0000000000000000_0000111000101000_0010110111101010"; -- 0.05530058825884648
	pesos_i(13964) := b"0000000000000000_0000000000000000_0001011111001100_0101010100101110"; -- 0.09296161997808891
	pesos_i(13965) := b"1111111111111111_1111111111111111_1110011101101011_0001011010000110"; -- -0.09602221696268792
	pesos_i(13966) := b"1111111111111111_1111111111111111_1111001010110000_1011101101110001"; -- -0.05199078064659833
	pesos_i(13967) := b"1111111111111111_1111111111111111_1111011011001011_0011011010101011"; -- -0.03596170730596103
	pesos_i(13968) := b"0000000000000000_0000000000000000_0000111001110010_1101001010010000"; -- 0.05643955234896559
	pesos_i(13969) := b"1111111111111111_1111111111111111_1101101110101000_1111100000011001"; -- -0.14195298577074872
	pesos_i(13970) := b"0000000000000000_0000000000000000_0000100001010101_1000010010100011"; -- 0.03255490293077774
	pesos_i(13971) := b"1111111111111111_1111111111111111_1111111011010101_0000010111000011"; -- -0.00456203441477633
	pesos_i(13972) := b"1111111111111111_1111111111111111_1110001101100011_1010011010110000"; -- -0.11176069450730393
	pesos_i(13973) := b"1111111111111111_1111111111111111_1110111011111111_1010000110101000"; -- -0.06641187330984637
	pesos_i(13974) := b"1111111111111111_1111111111111111_1111010000000010_0000001101000110"; -- -0.046844287303866305
	pesos_i(13975) := b"0000000000000000_0000000000000000_0010011000001100_0000111110111111"; -- 0.14862154390701843
	pesos_i(13976) := b"1111111111111111_1111111111111111_1101110110010100_0100110011011001"; -- -0.13445586873284876
	pesos_i(13977) := b"1111111111111111_1111111111111111_1110111101000110_0100110111111001"; -- -0.06533348720136269
	pesos_i(13978) := b"1111111111111111_1111111111111111_1110111010011110_1100001010001001"; -- -0.06789001620215111
	pesos_i(13979) := b"1111111111111111_1111111111111111_1101101011110011_0101010110111100"; -- -0.1447245040420632
	pesos_i(13980) := b"1111111111111111_1111111111111111_1110101001000000_0111110100101100"; -- -0.08495347660316839
	pesos_i(13981) := b"0000000000000000_0000000000000000_0000001101101100_1001010110101010"; -- 0.013375619897713985
	pesos_i(13982) := b"0000000000000000_0000000000000000_0001100101011011_0011010100110000"; -- 0.09904796992723844
	pesos_i(13983) := b"0000000000000000_0000000000000000_0000100111101100_1111000101011100"; -- 0.03877171028658879
	pesos_i(13984) := b"1111111111111111_1111111111111111_1111100010100101_1100111100011100"; -- -0.028719955186965233
	pesos_i(13985) := b"1111111111111111_1111111111111111_1101101111001110_0011110110000000"; -- -0.14138427370659137
	pesos_i(13986) := b"0000000000000000_0000000000000000_0010001011110010_0100001001010010"; -- 0.13650907991355035
	pesos_i(13987) := b"1111111111111111_1111111111111111_1111001101011000_1000110100010101"; -- -0.04943006732609874
	pesos_i(13988) := b"1111111111111111_1111111111111111_1110110010101100_0100101001001101"; -- -0.07549605972174833
	pesos_i(13989) := b"1111111111111111_1111111111111111_1101110001011000_0001100001011101"; -- -0.1392807745044831
	pesos_i(13990) := b"0000000000000000_0000000000000000_0000100010001001_1110101010011110"; -- 0.033354438332830284
	pesos_i(13991) := b"1111111111111111_1111111111111111_1101111010011110_0110111100111110"; -- -0.13039498075845385
	pesos_i(13992) := b"1111111111111111_1111111111111111_1110000010111001_1000100111010111"; -- -0.12216890811693987
	pesos_i(13993) := b"1111111111111111_1111111111111111_1110111010011101_0111101001001011"; -- -0.06790958097381375
	pesos_i(13994) := b"0000000000000000_0000000000000000_0000100110010101_0101000100110101"; -- 0.0374346499616606
	pesos_i(13995) := b"0000000000000000_0000000000000000_0001110101001110_1101011101001110"; -- 0.11448426876814835
	pesos_i(13996) := b"1111111111111111_1111111111111111_1111000000010101_0001001000011001"; -- -0.06217848671893035
	pesos_i(13997) := b"1111111111111111_1111111111111111_1111111101000101_0010110010101111"; -- -0.002850730179028372
	pesos_i(13998) := b"1111111111111111_1111111111111111_1110000110010101_1100101000110101"; -- -0.1188081378534019
	pesos_i(13999) := b"0000000000000000_0000000000000000_0010000000101000_0101111110001010"; -- 0.12561604621013045
	pesos_i(14000) := b"1111111111111111_1111111111111111_1101110101000101_1011010100000101"; -- -0.13565510388269614
	pesos_i(14001) := b"0000000000000000_0000000000000000_0000011000010110_1100110111101000"; -- 0.023785466314347806
	pesos_i(14002) := b"1111111111111111_1111111111111111_1110001111000101_1110011110110001"; -- -0.11026145862431333
	pesos_i(14003) := b"0000000000000000_0000000000000000_0001111101110011_0011111001001111"; -- 0.12285222469429538
	pesos_i(14004) := b"1111111111111111_1111111111111111_1111011111000110_0101000011101110"; -- -0.03213018608238272
	pesos_i(14005) := b"1111111111111111_1111111111111111_1101101111001011_0111001010000000"; -- -0.14142689097266187
	pesos_i(14006) := b"0000000000000000_0000000000000000_0001110101111001_1100101110010000"; -- 0.11513969674905881
	pesos_i(14007) := b"0000000000000000_0000000000000000_0010011111111111_1001111110111000"; -- 0.15624426128140198
	pesos_i(14008) := b"0000000000000000_0000000000000000_0001011100001110_0111000100001101"; -- 0.09006411134053821
	pesos_i(14009) := b"0000000000000000_0000000000000000_0001011010110010_1100011100100111"; -- 0.0886654349587529
	pesos_i(14010) := b"0000000000000000_0000000000000000_0001110101010110_1101100110001111"; -- 0.1146064733220116
	pesos_i(14011) := b"1111111111111111_1111111111111111_1110001100100001_0111010010010100"; -- -0.1127707612749452
	pesos_i(14012) := b"1111111111111111_1111111111111111_1111011110010101_0001011100111100"; -- -0.032881305563535454
	pesos_i(14013) := b"1111111111111111_1111111111111111_1111011000110101_1011000000110110"; -- -0.03824328114768278
	pesos_i(14014) := b"0000000000000000_0000000000000000_0001111101010110_1110110010000001"; -- 0.12242010255394858
	pesos_i(14015) := b"0000000000000000_0000000000000000_0000111111110101_1000100111100101"; -- 0.06234037236076487
	pesos_i(14016) := b"1111111111111111_1111111111111111_1111000100100010_1001101010010010"; -- -0.05806573810296969
	pesos_i(14017) := b"1111111111111111_1111111111111111_1111001001001010_0101101011010010"; -- -0.05355293622746208
	pesos_i(14018) := b"1111111111111111_1111111111111111_1110110100001011_1010101101101101"; -- -0.07404068555572922
	pesos_i(14019) := b"1111111111111111_1111111111111111_1111100010011111_0001111111111101"; -- -0.028821945922720138
	pesos_i(14020) := b"1111111111111111_1111111111111111_1111111111001000_1000111101000001"; -- -0.000845953499848188
	pesos_i(14021) := b"1111111111111111_1111111111111111_1110011011001011_0111111110101010"; -- -0.0984573563504596
	pesos_i(14022) := b"1111111111111111_1111111111111111_1110000011001000_0110000110000111"; -- -0.12194242906101063
	pesos_i(14023) := b"1111111111111111_1111111111111111_1111011111100101_0100000001110010"; -- -0.031658145951628615
	pesos_i(14024) := b"1111111111111111_1111111111111111_1111111111010101_1111111010100100"; -- -0.0006409500535271433
	pesos_i(14025) := b"1111111111111111_1111111111111111_1111010101011110_1000010100100010"; -- -0.04152648844225876
	pesos_i(14026) := b"0000000000000000_0000000000000000_0010000101110011_0011000011101111"; -- 0.1306639274786345
	pesos_i(14027) := b"1111111111111111_1111111111111111_1110010010001001_1110001001000100"; -- -0.10727105933590798
	pesos_i(14028) := b"1111111111111111_1111111111111111_1111101001001110_1100101101111010"; -- -0.022235186196920158
	pesos_i(14029) := b"0000000000000000_0000000000000000_0000000100100010_0001011001101011"; -- 0.00442638494568956
	pesos_i(14030) := b"1111111111111111_1111111111111111_1110011000101100_0001001100101001"; -- -0.10088997122674427
	pesos_i(14031) := b"1111111111111111_1111111111111111_1110001000000000_1111111001011010"; -- -0.11717233948139986
	pesos_i(14032) := b"1111111111111111_1111111111111111_1101111111110101_1100100000101010"; -- -0.1251559160601992
	pesos_i(14033) := b"1111111111111111_1111111111111111_1110000000101100_1011000010101000"; -- -0.12431808367492556
	pesos_i(14034) := b"0000000000000000_0000000000000000_0001110110010001_0000010011101101"; -- 0.11549406801478414
	pesos_i(14035) := b"1111111111111111_1111111111111111_1101111111000111_1001111001100001"; -- -0.12586031077866788
	pesos_i(14036) := b"1111111111111111_1111111111111111_1111110011011010_1111111001110001"; -- -0.012283418184525446
	pesos_i(14037) := b"1111111111111111_1111111111111111_1111001011101111_1011000000001000"; -- -0.05103015722392654
	pesos_i(14038) := b"1111111111111111_1111111111111111_1110011001011111_1011100010110110"; -- -0.10010190534000045
	pesos_i(14039) := b"1111111111111111_1111111111111111_1111011011100011_0101011011100111"; -- -0.03559357518391087
	pesos_i(14040) := b"0000000000000000_0000000000000000_0010001110000100_1101010100000011"; -- 0.13874560672844558
	pesos_i(14041) := b"1111111111111111_1111111111111111_1111111001100000_1110011101001110"; -- -0.006333869309761921
	pesos_i(14042) := b"1111111111111111_1111111111111111_1110000100001110_1110000111011100"; -- -0.12086666462982458
	pesos_i(14043) := b"1111111111111111_1111111111111111_1111110111101011_0010010111000011"; -- -0.008130683772084986
	pesos_i(14044) := b"1111111111111111_1111111111111111_1111111010111101_0011010100111110"; -- -0.004925415367705474
	pesos_i(14045) := b"0000000000000000_0000000000000000_0000001100000011_0001110010110100"; -- 0.011766237245548386
	pesos_i(14046) := b"1111111111111111_1111111111111111_1110111111001111_0001011100100100"; -- -0.06324630136089981
	pesos_i(14047) := b"0000000000000000_0000000000000000_0000111010001111_1000100010010011"; -- 0.056877647258440675
	pesos_i(14048) := b"0000000000000000_0000000000000000_0000010000100111_0011111101100110"; -- 0.016223871537705926
	pesos_i(14049) := b"0000000000000000_0000000000000000_0001111111110011_1011010110110010"; -- 0.12481246557564761
	pesos_i(14050) := b"1111111111111111_1111111111111111_1110111101111101_1101010101001110"; -- -0.06448618732741104
	pesos_i(14051) := b"1111111111111111_1111111111111111_1111001010110000_0011000100100111"; -- -0.05199902333704698
	pesos_i(14052) := b"0000000000000000_0000000000000000_0010011100100011_1101100010100111"; -- 0.15289072103640305
	pesos_i(14053) := b"0000000000000000_0000000000000000_0010001011001001_1111110011000111"; -- 0.13589458331995735
	pesos_i(14054) := b"0000000000000000_0000000000000000_0001000111000010_1011000110101101"; -- 0.06937704544370621
	pesos_i(14055) := b"0000000000000000_0000000000000000_0001001100111010_1011111101010110"; -- 0.07511516434055103
	pesos_i(14056) := b"0000000000000000_0000000000000000_0001111011111100_1111110110100011"; -- 0.12104783284478139
	pesos_i(14057) := b"0000000000000000_0000000000000000_0010011101001000_0101100011100000"; -- 0.15344768025321998
	pesos_i(14058) := b"0000000000000000_0000000000000000_0001110001110011_0000100000001001"; -- 0.11113023961923457
	pesos_i(14059) := b"1111111111111111_1111111111111111_1110010000001100_0000100100100000"; -- -0.10919135060598584
	pesos_i(14060) := b"1111111111111111_1111111111111111_1110110110110001_1011100100011010"; -- -0.07150691141246632
	pesos_i(14061) := b"1111111111111111_1111111111111111_1111001000101000_0111110010001010"; -- -0.054069725375999286
	pesos_i(14062) := b"1111111111111111_1111111111111111_1110111000000101_1110010111110011"; -- -0.07022250001233155
	pesos_i(14063) := b"1111111111111111_1111111111111111_1111100110000110_1010100100010101"; -- -0.02528899412272758
	pesos_i(14064) := b"1111111111111111_1111111111111111_1111000000110010_0111101100000011"; -- -0.06172972854340566
	pesos_i(14065) := b"1111111111111111_1111111111111111_1110101011001001_0101001110001101"; -- -0.0828655034034412
	pesos_i(14066) := b"1111111111111111_1111111111111111_1111101011010010_0111111111101111"; -- -0.02022552894658494
	pesos_i(14067) := b"1111111111111111_1111111111111111_1110010010101010_0011011011101001"; -- -0.10677773289936385
	pesos_i(14068) := b"1111111111111111_1111111111111111_1110000111111011_1000111111010011"; -- -0.1172552213009578
	pesos_i(14069) := b"1111111111111111_1111111111111111_1110100111001100_1001001000110011"; -- -0.08672224283599078
	pesos_i(14070) := b"1111111111111111_1111111111111111_1111001110001000_0010001011111110"; -- -0.04870396887845128
	pesos_i(14071) := b"1111111111111111_1111111111111111_1111110110010101_0011110111111100"; -- -0.009441495945973714
	pesos_i(14072) := b"0000000000000000_0000000000000000_0001000110110010_0001101101010110"; -- 0.06912394372557353
	pesos_i(14073) := b"1111111111111111_1111111111111111_1101101111111100_1000100110100011"; -- -0.14067783134460124
	pesos_i(14074) := b"1111111111111111_1111111111111111_1110011011000000_0001111001101011"; -- -0.09863099954476093
	pesos_i(14075) := b"0000000000000000_0000000000000000_0010100101100101_1110011100101101"; -- 0.16171116687067114
	pesos_i(14076) := b"1111111111111111_1111111111111111_1110111111000100_0001001111000010"; -- -0.06341434964412766
	pesos_i(14077) := b"0000000000000000_0000000000000000_0000010001010101_1001000111101001"; -- 0.016930694048858212
	pesos_i(14078) := b"0000000000000000_0000000000000000_0001100010100111_0000001001110100"; -- 0.09629836390236808
	pesos_i(14079) := b"0000000000000000_0000000000000000_0001000011111111_0011011101000111"; -- 0.06639428600402156
	pesos_i(14080) := b"0000000000000000_0000000000000000_0000011011001101_1100001110010111"; -- 0.026577209743407524
	pesos_i(14081) := b"1111111111111111_1111111111111111_1111110101000000_1110110000000100"; -- -0.010728119778610972
	pesos_i(14082) := b"1111111111111111_1111111111111111_1111111011100100_1010110001011100"; -- -0.0043232227808442025
	pesos_i(14083) := b"1111111111111111_1111111111111111_1110110011111100_1001101000101001"; -- -0.07427059654976596
	pesos_i(14084) := b"1111111111111111_1111111111111111_1110110100100111_0111101010010110"; -- -0.07361635050639603
	pesos_i(14085) := b"0000000000000000_0000000000000000_0001000001100000_0010011110111000"; -- 0.0639672111085125
	pesos_i(14086) := b"0000000000000000_0000000000000000_0010001101011101_1000000011100010"; -- 0.1381454993327933
	pesos_i(14087) := b"0000000000000000_0000000000000000_0001101100101010_1001001101000000"; -- 0.10611839600111228
	pesos_i(14088) := b"0000000000000000_0000000000000000_0001001110110001_0101011110000001"; -- 0.07692477120233877
	pesos_i(14089) := b"0000000000000000_0000000000000000_0010100000111001_1111011100100111"; -- 0.15713448250621742
	pesos_i(14090) := b"0000000000000000_0000000000000000_0000101010101000_1010101101000011"; -- 0.041636184508059323
	pesos_i(14091) := b"0000000000000000_0000000000000000_0010011001000100_1000110111011111"; -- 0.14948355387575632
	pesos_i(14092) := b"1111111111111111_1111111111111111_1111100111011101_1101111100101110"; -- -0.023958255048928796
	pesos_i(14093) := b"1111111111111111_1111111111111111_1110011010100110_1001101001010101"; -- -0.09902034199938191
	pesos_i(14094) := b"0000000000000000_0000000000000000_0001010101111101_0000000010101011"; -- 0.08393863855736095
	pesos_i(14095) := b"0000000000000000_0000000000000000_0001111111011101_0101001110100011"; -- 0.12447092747358943
	pesos_i(14096) := b"0000000000000000_0000000000000000_0010010011010011_0100101001111010"; -- 0.1438490435772437
	pesos_i(14097) := b"1111111111111111_1111111111111111_1111111000000101_1000101111000100"; -- -0.007727875429156258
	pesos_i(14098) := b"1111111111111111_1111111111111111_1110011100010010_0111010000000001"; -- -0.09737467750932613
	pesos_i(14099) := b"0000000000000000_0000000000000000_0001000001011111_0110100111001000"; -- 0.06395589009802978
	pesos_i(14100) := b"0000000000000000_0000000000000000_0001000111101100_1000011010001011"; -- 0.07001534365317001
	pesos_i(14101) := b"0000000000000000_0000000000000000_0001011011010000_1000110100111011"; -- 0.0891197460781368
	pesos_i(14102) := b"1111111111111111_1111111111111111_1101000011110000_1111010111001100"; -- -0.1838232399799788
	pesos_i(14103) := b"0000000000000000_0000000000000000_0001100000101011_0110110110111010"; -- 0.09441266809690835
	pesos_i(14104) := b"1111111111111111_1111111111111111_1111011010010110_1111110010111010"; -- -0.036758618016509426
	pesos_i(14105) := b"1111111111111111_1111111111111111_1111001001011110_0010111111110100"; -- -0.05325031566873973
	pesos_i(14106) := b"0000000000000000_0000000000000000_0000000100100001_1111000001001000"; -- 0.004424111997441232
	pesos_i(14107) := b"1111111111111111_1111111111111111_1101110011100000_1000000110001111"; -- -0.13719930891421667
	pesos_i(14108) := b"0000000000000000_0000000000000000_0000110111011000_1001111111001111"; -- 0.05408667380072193
	pesos_i(14109) := b"1111111111111111_1111111111111111_1110011101100010_0000000001001110"; -- -0.09616087059122007
	pesos_i(14110) := b"0000000000000000_0000000000000000_0001111100010110_1101100111111101"; -- 0.12144243654121877
	pesos_i(14111) := b"1111111111111111_1111111111111111_1110110010111100_0001101000111110"; -- -0.07525478352259854
	pesos_i(14112) := b"1111111111111111_1111111111111111_1110010010110011_0000011001110101"; -- -0.10664329193913424
	pesos_i(14113) := b"1111111111111111_1111111111111111_1101111100111100_0100000010011101"; -- -0.12798687145329343
	pesos_i(14114) := b"1111111111111111_1111111111111111_1111001111101110_0111101011100101"; -- -0.047142333082923746
	pesos_i(14115) := b"1111111111111111_1111111111111111_1110001001001011_1011010101110000"; -- -0.11603227632168073
	pesos_i(14116) := b"1111111111111111_1111111111111111_1111111000011110_1000101011111111"; -- -0.007346451590860064
	pesos_i(14117) := b"0000000000000000_0000000000000000_0010100000110000_1110011011110010"; -- 0.1569961872583494
	pesos_i(14118) := b"1111111111111111_1111111111111111_1110001000001000_1111100101110111"; -- -0.11705056037155459
	pesos_i(14119) := b"0000000000000000_0000000000000000_0001011000001101_1101001011110110"; -- 0.08614843848513619
	pesos_i(14120) := b"1111111111111111_1111111111111111_1111101110011111_1110111111001011"; -- -0.01709080970521319
	pesos_i(14121) := b"1111111111111111_1111111111111111_1110110100101111_0010010000100110"; -- -0.07349943226885831
	pesos_i(14122) := b"1111111111111111_1111111111111111_1110111101000101_0011110110101101"; -- -0.06534971736018806
	pesos_i(14123) := b"0000000000000000_0000000000000000_0010000011011000_1111100101101101"; -- 0.12831076531170718
	pesos_i(14124) := b"1111111111111111_1111111111111111_1101011111011000_1011010111001110"; -- -0.15684951510404546
	pesos_i(14125) := b"0000000000000000_0000000000000000_0010001001001101_1101001100001001"; -- 0.13400000537071172
	pesos_i(14126) := b"0000000000000000_0000000000000000_0010001010010010_0101000100001011"; -- 0.1350451136525648
	pesos_i(14127) := b"0000000000000000_0000000000000000_0010001000010011_0110011001100111"; -- 0.13310852066514456
	pesos_i(14128) := b"1111111111111111_1111111111111111_1111000100000010_1101010001110011"; -- -0.05855056957560502
	pesos_i(14129) := b"1111111111111111_1111111111111111_1110100111101011_0010100001111100"; -- -0.08625552151033673
	pesos_i(14130) := b"1111111111111111_1111111111111111_1101101110110100_1000010001011011"; -- -0.14177677890998608
	pesos_i(14131) := b"0000000000000000_0000000000000000_0001101011111111_1101000010001011"; -- 0.10546592132557159
	pesos_i(14132) := b"0000000000000000_0000000000000000_0001011011110101_1000001001101111"; -- 0.08968367774049138
	pesos_i(14133) := b"0000000000000000_0000000000000000_0010001111010110_1001001000011100"; -- 0.13999283964426096
	pesos_i(14134) := b"1111111111111111_1111111111111111_1110110011000011_0111110011100111"; -- -0.07514209130114637
	pesos_i(14135) := b"1111111111111111_1111111111111111_1111010011100010_0000000011110001"; -- -0.0434264574978261
	pesos_i(14136) := b"1111111111111111_1111111111111111_1110000001100111_0010110100110101"; -- -0.1234256501651316
	pesos_i(14137) := b"1111111111111111_1111111111111111_1110001100011111_0110111101001111"; -- -0.11280159299864327
	pesos_i(14138) := b"0000000000000000_0000000000000000_0010010110011111_0000100010110001"; -- 0.14695791552392298
	pesos_i(14139) := b"1111111111111111_1111111111111111_1111011110101101_0010011010100111"; -- -0.03251417568613016
	pesos_i(14140) := b"0000000000000000_0000000000000000_0000010010010001_1011111110001010"; -- 0.017848941077987898
	pesos_i(14141) := b"1111111111111111_1111111111111111_1101111001011010_1111010111001111"; -- -0.13142455767838326
	pesos_i(14142) := b"1111111111111111_1111111111111111_1111111011110101_1100110010010010"; -- -0.004061903406912469
	pesos_i(14143) := b"1111111111111111_1111111111111111_1111101111110111_0111000011001001"; -- -0.015755606557815376
	pesos_i(14144) := b"1111111111111111_1111111111111111_1111000111110100_1111001100111110"; -- -0.054856107027872934
	pesos_i(14145) := b"0000000000000000_0000000000000000_0000010101000110_0001010101001101"; -- 0.02060063486526854
	pesos_i(14146) := b"1111111111111111_1111111111111111_1111110111100010_0111100100010110"; -- -0.008263046287494021
	pesos_i(14147) := b"1111111111111111_1111111111111111_1111011100010011_1100010101011000"; -- -0.03485457051871183
	pesos_i(14148) := b"1111111111111111_1111111111111111_1111001010000100_0010011111101111"; -- -0.05267095965321838
	pesos_i(14149) := b"1111111111111111_1111111111111111_1111001000001100_1100000100101100"; -- -0.05449288052786027
	pesos_i(14150) := b"0000000000000000_0000000000000000_0000010011000001_1011000100101010"; -- 0.018580506190590724
	pesos_i(14151) := b"0000000000000000_0000000000000000_0000110101000000_1011011001111011"; -- 0.05176868928718867
	pesos_i(14152) := b"0000000000000000_0000000000000000_0000000001111111_0111010101110000"; -- 0.0019448660969860429
	pesos_i(14153) := b"0000000000000000_0000000000000000_0001001100011001_1001000100111111"; -- 0.07460887700671304
	pesos_i(14154) := b"0000000000000000_0000000000000000_0010010100111011_0111000011110011"; -- 0.14543825074565314
	pesos_i(14155) := b"0000000000000000_0000000000000000_0001100101011101_0010010000000001"; -- 0.09907746344112353
	pesos_i(14156) := b"1111111111111111_1111111111111111_1110110000100011_1100101110101000"; -- -0.07757880357631802
	pesos_i(14157) := b"0000000000000000_0000000000000000_0010000000011111_0001011100110100"; -- 0.12547440553733238
	pesos_i(14158) := b"0000000000000000_0000000000000000_0000011100001101_0110110001101010"; -- 0.027548576275032013
	pesos_i(14159) := b"1111111111111111_1111111111111111_1111110111001010_1010010011101000"; -- -0.008626645499936289
	pesos_i(14160) := b"0000000000000000_0000000000000000_0001100011111011_0010110001011110"; -- 0.09758260051268386
	pesos_i(14161) := b"0000000000000000_0000000000000000_0001010011111101_0000110001001010"; -- 0.08198620614892867
	pesos_i(14162) := b"0000000000000000_0000000000000000_0000001111011100_1000001100100110"; -- 0.015083500619998365
	pesos_i(14163) := b"1111111111111111_1111111111111111_1110100100011010_1010000001001100"; -- -0.08943746697734015
	pesos_i(14164) := b"0000000000000000_0000000000000000_0000001001110000_1100111001000001"; -- 0.0095337780129147
	pesos_i(14165) := b"1111111111111111_1111111111111111_1111010111111100_0110111011100111"; -- -0.03911692493873075
	pesos_i(14166) := b"0000000000000000_0000000000000000_0010001000101010_0101001001001001"; -- 0.13345827364566265
	pesos_i(14167) := b"1111111111111111_1111111111111111_1101101001010000_0110010100111000"; -- -0.14721076385828424
	pesos_i(14168) := b"0000000000000000_0000000000000000_0000001110110111_1001010001100010"; -- 0.014519952737490663
	pesos_i(14169) := b"0000000000000000_0000000000000000_0010000100010000_1001110011010010"; -- 0.1291597379329309
	pesos_i(14170) := b"1111111111111111_1111111111111111_1110111110110000_0001000111111100"; -- -0.06371963121937038
	pesos_i(14171) := b"1111111111111111_1111111111111111_1111111101110101_1111101010101001"; -- -0.0021060312729042825
	pesos_i(14172) := b"0000000000000000_0000000000000000_0001100000111100_0000111110111110"; -- 0.09466646575806609
	pesos_i(14173) := b"1111111111111111_1111111111111111_1111001001011101_0111111000101100"; -- -0.053260912193646356
	pesos_i(14174) := b"0000000000000000_0000000000000000_0001110110010111_1000110000001000"; -- 0.11559367365405296
	pesos_i(14175) := b"1111111111111111_1111111111111111_1111010100110101_1011110110100011"; -- -0.04214873091431081
	pesos_i(14176) := b"0000000000000000_0000000000000000_0010000100001011_1010101100100111"; -- 0.1290842981946425
	pesos_i(14177) := b"0000000000000000_0000000000000000_0000001111010111_1010011110001110"; -- 0.015009376687453085
	pesos_i(14178) := b"0000000000000000_0000000000000000_0010010101011000_1010000100101100"; -- 0.14588363005161437
	pesos_i(14179) := b"0000000000000000_0000000000000000_0000100110111101_0100111000111101"; -- 0.03804482453972443
	pesos_i(14180) := b"0000000000000000_0000000000000000_0001011010010100_0111111001101011"; -- 0.08820333596669877
	pesos_i(14181) := b"1111111111111111_1111111111111111_1101110010110110_1111111010100010"; -- -0.13783272314601192
	pesos_i(14182) := b"0000000000000000_0000000000000000_0001011011010011_0100010100001111"; -- 0.08916122061808396
	pesos_i(14183) := b"0000000000000000_0000000000000000_0000000101010101_0001000011010011"; -- 0.005204249805037083
	pesos_i(14184) := b"0000000000000000_0000000000000000_0001110001001101_1100001010010111"; -- 0.11056152528200132
	pesos_i(14185) := b"0000000000000000_0000000000000000_0010000011100010_1011101110110000"; -- 0.12845967328510563
	pesos_i(14186) := b"0000000000000000_0000000000000000_0001010111010110_1010100110110010"; -- 0.0853067454298791
	pesos_i(14187) := b"0000000000000000_0000000000000000_0000000000101001_1101110111100011"; -- 0.0006388357287287669
	pesos_i(14188) := b"0000000000000000_0000000000000000_0010000001000001_1100100101110110"; -- 0.1260038294067683
	pesos_i(14189) := b"1111111111111111_1111111111111111_1110111111100100_1101010001101000"; -- -0.06291458568023249
	pesos_i(14190) := b"0000000000000000_0000000000000000_0001000111110001_0101010011100101"; -- 0.07008867815846842
	pesos_i(14191) := b"0000000000000000_0000000000000000_0001101010010011_1100100101001010"; -- 0.10381753969766268
	pesos_i(14192) := b"0000000000000000_0000000000000000_0000010001011010_1110010101110100"; -- 0.01701196749531165
	pesos_i(14193) := b"0000000000000000_0000000000000000_0000001100100000_0101110011110000"; -- 0.012212570696548363
	pesos_i(14194) := b"1111111111111111_1111111111111111_1110100010001001_1110100110011011"; -- -0.09164562191867853
	pesos_i(14195) := b"1111111111111111_1111111111111111_1111001010001000_1011000010110010"; -- -0.05260177277137778
	pesos_i(14196) := b"0000000000000000_0000000000000000_0001001110111000_1111111100100011"; -- 0.0770415745132655
	pesos_i(14197) := b"1111111111111111_1111111111111111_1111001101000010_0000010010110100"; -- -0.04977388949815158
	pesos_i(14198) := b"0000000000000000_0000000000000000_0001101110001010_1101100111010000"; -- 0.10758744541459962
	pesos_i(14199) := b"1111111111111111_1111111111111111_1111011101111000_1101111001011011"; -- -0.033311941851070434
	pesos_i(14200) := b"0000000000000000_0000000000000000_0001000001011100_0100010001000011"; -- 0.0639078772830682
	pesos_i(14201) := b"1111111111111111_1111111111111111_1101110001111001_1001011000001100"; -- -0.13876974300024006
	pesos_i(14202) := b"0000000000000000_0000000000000000_0000101111010101_0001110100110110"; -- 0.04622061313563223
	pesos_i(14203) := b"1111111111111111_1111111111111111_1111111011000011_1000011011000010"; -- -0.004829003847069905
	pesos_i(14204) := b"0000000000000000_0000000000000000_0000001011101110_0010010011000011"; -- 0.011446283002487836
	pesos_i(14205) := b"0000000000000000_0000000000000000_0000111000010000_1111010110011010"; -- 0.05494627962952428
	pesos_i(14206) := b"0000000000000000_0000000000000000_0010001010100000_1000100010111011"; -- 0.1352620559062307
	pesos_i(14207) := b"1111111111111111_1111111111111111_1110100011001001_1101101011110110"; -- -0.0906699322042407
	pesos_i(14208) := b"1111111111111111_1111111111111111_1111001010000011_1101010010000100"; -- -0.05267593168107421
	pesos_i(14209) := b"1111111111111111_1111111111111111_1111011100111101_0001110110100111"; -- -0.03422369643102002
	pesos_i(14210) := b"0000000000000000_0000000000000000_0000010111011110_0011010110111101"; -- 0.022921904306422988
	pesos_i(14211) := b"1111111111111111_1111111111111111_1101111110000001_1000100001100101"; -- -0.12692973647667818
	pesos_i(14212) := b"1111111111111111_1111111111111111_1111001100000010_1011110111100001"; -- -0.05073941474850112
	pesos_i(14213) := b"1111111111111111_1111111111111111_1111100110101001_1100010010010001"; -- -0.024753298307961535
	pesos_i(14214) := b"0000000000000000_0000000000000000_0010000011101011_0100111001001011"; -- 0.12859048212531365
	pesos_i(14215) := b"1111111111111111_1111111111111111_1111101000101001_1110100110011110"; -- -0.022797964964319614
	pesos_i(14216) := b"0000000000000000_0000000000000000_0010010001100011_1111101000010001"; -- 0.14215052513234006
	pesos_i(14217) := b"1111111111111111_1111111111111111_1101111110100011_1101110100000110"; -- -0.12640589337166544
	pesos_i(14218) := b"0000000000000000_0000000000000000_0000000111110011_0000000011100010"; -- 0.007614188306289857
	pesos_i(14219) := b"1111111111111111_1111111111111111_1101111010110011_0110011100100001"; -- -0.1300750298477502
	pesos_i(14220) := b"1111111111111111_1111111111111111_1111000110011011_0100100001010100"; -- -0.05622432667012645
	pesos_i(14221) := b"0000000000000000_0000000000000000_0010010000100011_0011111001111110"; -- 0.14116278248108854
	pesos_i(14222) := b"1111111111111111_1111111111111111_1110110110000011_0001101111110110"; -- -0.07221818196447057
	pesos_i(14223) := b"1111111111111111_1111111111111111_1111110111000011_1101101011011000"; -- -0.008730242092821187
	pesos_i(14224) := b"1111111111111111_1111111111111111_1111110010101100_1001111011111111"; -- -0.012991011266667426
	pesos_i(14225) := b"0000000000000000_0000000000000000_0001010011001110_1001011110000101"; -- 0.0812773418474226
	pesos_i(14226) := b"0000000000000000_0000000000000000_0000010110011001_0010100010011010"; -- 0.021868264679560344
	pesos_i(14227) := b"0000000000000000_0000000000000000_0001100001011010_1000111001110110"; -- 0.0951317822717745
	pesos_i(14228) := b"0000000000000000_0000000000000000_0000010010010001_1101001010101010"; -- 0.01785008098443618
	pesos_i(14229) := b"0000000000000000_0000000000000000_0001100000000111_0001010111001111"; -- 0.09385811142415863
	pesos_i(14230) := b"0000000000000000_0000000000000000_0001111110001000_1100010000100101"; -- 0.12318063650398481
	pesos_i(14231) := b"1111111111111111_1111111111111111_1101110100101101_0010110100000011"; -- -0.13602942169417148
	pesos_i(14232) := b"0000000000000000_0000000000000000_0010001011111011_1101000100100011"; -- 0.13665492148137776
	pesos_i(14233) := b"0000000000000000_0000000000000000_0001100110111011_0001110001110001"; -- 0.10051133876911798
	pesos_i(14234) := b"0000000000000000_0000000000000000_0001111100100010_0101101001111101"; -- 0.12161794224090289
	pesos_i(14235) := b"1111111111111111_1111111111111111_1111000111101000_1000101000111111"; -- -0.0550454708796368
	pesos_i(14236) := b"0000000000000000_0000000000000000_0001000110010100_1001011010011010"; -- 0.06867352732021605
	pesos_i(14237) := b"1111111111111111_1111111111111111_1110000100100110_1111110011010010"; -- -0.12049884667134822
	pesos_i(14238) := b"0000000000000000_0000000000000000_0000111001111101_1011000000111011"; -- 0.05660535271536183
	pesos_i(14239) := b"0000000000000000_0000000000000000_0010100110010101_1110110000100000"; -- 0.16244388374526014
	pesos_i(14240) := b"0000000000000000_0000000000000000_0001011010000110_1001111111001111"; -- 0.08799170302385256
	pesos_i(14241) := b"1111111111111111_1111111111111111_1110100010000001_1111000110101100"; -- -0.09176721140914762
	pesos_i(14242) := b"1111111111111111_1111111111111111_1101110011000111_0101111111110001"; -- -0.1375827824432688
	pesos_i(14243) := b"1111111111111111_1111111111111111_1110001111101000_1101111000111011"; -- -0.10972796497581937
	pesos_i(14244) := b"0000000000000000_0000000000000000_0000110011001000_0011110010000111"; -- 0.049930365620219505
	pesos_i(14245) := b"0000000000000000_0000000000000000_0000100100101010_0101100000110110"; -- 0.03580237684880453
	pesos_i(14246) := b"1111111111111111_1111111111111111_1101110001101011_1100110011011101"; -- -0.13898009874247272
	pesos_i(14247) := b"1111111111111111_1111111111111111_1110101111100001_0101110110000110"; -- -0.07859244812281134
	pesos_i(14248) := b"1111111111111111_1111111111111111_1111000110110111_0001110001101010"; -- -0.05579969799908188
	pesos_i(14249) := b"1111111111111111_1111111111111111_1111001100000011_1110100100000010"; -- -0.05072158523907008
	pesos_i(14250) := b"1111111111111111_1111111111111111_1111110110101011_0011010000011010"; -- -0.009106391604095761
	pesos_i(14251) := b"1111111111111111_1111111111111111_1110111111010101_1110111011000010"; -- -0.06314189680487584
	pesos_i(14252) := b"0000000000000000_0000000000000000_0001101011111111_0100111001000001"; -- 0.10545815550109025
	pesos_i(14253) := b"1111111111111111_1111111111111111_1111000100111011_1111111010101001"; -- -0.057678302502683444
	pesos_i(14254) := b"1111111111111111_1111111111111111_1110010000000111_0001100100000111"; -- -0.10926669679518014
	pesos_i(14255) := b"1111111111111111_1111111111111111_1111000111010101_0000100111011101"; -- -0.05534303997763355
	pesos_i(14256) := b"0000000000000000_0000000000000000_0001011000011100_1001001010110001"; -- 0.08637348953175536
	pesos_i(14257) := b"0000000000000000_0000000000000000_0001011100111110_1010010000110010"; -- 0.09079958167085336
	pesos_i(14258) := b"1111111111111111_1111111111111111_1111101110101011_0101110100101101"; -- -0.016916443386559517
	pesos_i(14259) := b"0000000000000000_0000000000000000_0000010010000111_0010011010010000"; -- 0.017687234934804896
	pesos_i(14260) := b"0000000000000000_0000000000000000_0010010000000000_1110001111001111"; -- 0.1406385784275559
	pesos_i(14261) := b"0000000000000000_0000000000000000_0001110000011011_0001110111101110"; -- 0.109788771159047
	pesos_i(14262) := b"0000000000000000_0000000000000000_0001100100110001_1001011011110011"; -- 0.09841292802464201
	pesos_i(14263) := b"1111111111111111_1111111111111111_1110101001000010_0001010011101110"; -- -0.08492917242225832
	pesos_i(14264) := b"1111111111111111_1111111111111111_1111001001111111_1010111100001011"; -- -0.052739200341604016
	pesos_i(14265) := b"1111111111111111_1111111111111111_1110101110101100_1101010110010000"; -- -0.0793940090163427
	pesos_i(14266) := b"0000000000000000_0000000000000000_0000111101110100_1000101111001100"; -- 0.06037210200465223
	pesos_i(14267) := b"0000000000000000_0000000000000000_0001100110001111_0001100101001110"; -- 0.099839765051126
	pesos_i(14268) := b"0000000000000000_0000000000000000_0001110100100111_0001100001100100"; -- 0.11387779654932925
	pesos_i(14269) := b"0000000000000000_0000000000000000_0000111011011010_1000011011001110"; -- 0.058021951025171624
	pesos_i(14270) := b"1111111111111111_1111111111111111_1110100001101000_0000101000110111"; -- -0.09216247706984745
	pesos_i(14271) := b"1111111111111111_1111111111111111_1111100110100111_1000011101001000"; -- -0.024787468845069115
	pesos_i(14272) := b"0000000000000000_0000000000000000_0001000011100110_1110001010111010"; -- 0.06602303552338157
	pesos_i(14273) := b"1111111111111111_1111111111111111_1111110011100010_0110011001101010"; -- -0.012170409245961763
	pesos_i(14274) := b"1111111111111111_1111111111111111_1110111000101011_0000101010111110"; -- -0.06965573188489661
	pesos_i(14275) := b"1111111111111111_1111111111111111_1101011110110111_0111111010100011"; -- -0.1573563434178917
	pesos_i(14276) := b"1111111111111111_1111111111111111_1111011010010100_0001000100011111"; -- -0.036803178624987644
	pesos_i(14277) := b"1111111111111111_1111111111111111_1110001110001010_1101101111000111"; -- -0.11116243732025523
	pesos_i(14278) := b"1111111111111111_1111111111111111_1110001000001110_1100001110010101"; -- -0.11696221934032108
	pesos_i(14279) := b"1111111111111111_1111111111111111_1110010101110001_1000101000101001"; -- -0.10373627182989013
	pesos_i(14280) := b"0000000000000000_0000000000000000_0000111000000100_1111110010111011"; -- 0.05476359906711035
	pesos_i(14281) := b"0000000000000000_0000000000000000_0010010000110111_1001100011111101"; -- 0.1414733522654414
	pesos_i(14282) := b"0000000000000000_0000000000000000_0000101111010100_0110001110100001"; -- 0.04620955168712261
	pesos_i(14283) := b"1111111111111111_1111111111111111_1111111000110001_0010000001010110"; -- -0.007062891915609016
	pesos_i(14284) := b"0000000000000000_0000000000000000_0000010101001000_0101011010000111"; -- 0.020635040294715662
	pesos_i(14285) := b"1111111111111111_1111111111111111_1110011101101010_0101111110001011"; -- -0.09603312364401696
	pesos_i(14286) := b"1111111111111111_1111111111111111_1111010111011000_0100011100100000"; -- -0.039668612171394384
	pesos_i(14287) := b"1111111111111111_1111111111111111_1110010111111010_0111100001000000"; -- -0.10164688520478675
	pesos_i(14288) := b"1111111111111111_1111111111111111_1110011010000001_1001111101001111"; -- -0.09958462069725188
	pesos_i(14289) := b"1111111111111111_1111111111111111_1101100000100110_1000011101000100"; -- -0.1556621035993623
	pesos_i(14290) := b"0000000000000000_0000000000000000_0000100000000101_0101100000001111"; -- 0.03133154271997338
	pesos_i(14291) := b"0000000000000000_0000000000000000_0000111000110101_1000110010100111"; -- 0.055504599277035244
	pesos_i(14292) := b"1111111111111111_1111111111111111_1111100101010001_0100110111100110"; -- -0.026103144882046198
	pesos_i(14293) := b"1111111111111111_1111111111111111_1111110010010010_1001110011010011"; -- -0.013387869360239803
	pesos_i(14294) := b"1111111111111111_1111111111111111_1111110101010101_1000001110111010"; -- -0.010413901474442813
	pesos_i(14295) := b"0000000000000000_0000000000000000_0000001100111100_0000100101110011"; -- 0.012634840641911171
	pesos_i(14296) := b"0000000000000000_0000000000000000_0001001000110111_0101011110100110"; -- 0.07115695775434655
	pesos_i(14297) := b"0000000000000000_0000000000000000_0001010111000001_0101110011100011"; -- 0.0849817327120742
	pesos_i(14298) := b"0000000000000000_0000000000000000_0000110101101100_1001111100000001"; -- 0.05243867652561402
	pesos_i(14299) := b"1111111111111111_1111111111111111_1110111010010111_0011010100100110"; -- -0.0680052550134594
	pesos_i(14300) := b"0000000000000000_0000000000000000_0001000010101001_0101100001101010"; -- 0.06508400530859329
	pesos_i(14301) := b"1111111111111111_1111111111111111_1111101000011011_0100001101100110"; -- -0.02302149551016725
	pesos_i(14302) := b"1111111111111111_1111111111111111_1110000010010010_0000000100000011"; -- -0.12277215643774607
	pesos_i(14303) := b"0000000000000000_0000000000000000_0001011010011111_1110110101100010"; -- 0.08837779659167154
	pesos_i(14304) := b"0000000000000000_0000000000000000_0001100110111110_0010010110100000"; -- 0.10055766252323275
	pesos_i(14305) := b"1111111111111111_1111111111111111_1111101101111001_0100001111001011"; -- -0.017680895694616477
	pesos_i(14306) := b"1111111111111111_1111111111111111_1110000000011001_1100111111111010"; -- -0.12460613387919076
	pesos_i(14307) := b"1111111111111111_1111111111111111_1110010111011110_0000101100111010"; -- -0.1020806295939952
	pesos_i(14308) := b"1111111111111111_1111111111111111_1111001100100111_1011010011110101"; -- -0.050175371386562986
	pesos_i(14309) := b"1111111111111111_1111111111111111_1111110101001100_1011100001001011"; -- -0.010548097222744936
	pesos_i(14310) := b"1111111111111111_1111111111111111_1111100110111010_1110100111000110"; -- -0.024491681311427368
	pesos_i(14311) := b"0000000000000000_0000000000000000_0001111111111010_0111000010101001"; -- 0.12491516236671624
	pesos_i(14312) := b"0000000000000000_0000000000000000_0001101100001101_0110110000100011"; -- 0.10567355959915245
	pesos_i(14313) := b"1111111111111111_1111111111111111_1110011010110101_1001110111101010"; -- -0.09879124682513332
	pesos_i(14314) := b"1111111111111111_1111111111111111_1111001100000001_0100011110001100"; -- -0.05076172674920871
	pesos_i(14315) := b"0000000000000000_0000000000000000_0001101010001011_1110100100000010"; -- 0.10369736009243134
	pesos_i(14316) := b"1111111111111111_1111111111111111_1110110101101111_1000111010100100"; -- -0.07251652229370992
	pesos_i(14317) := b"1111111111111111_1111111111111111_1110010011000001_0110010000000000"; -- -0.10642409315121096
	pesos_i(14318) := b"1111111111111111_1111111111111111_1110110100100111_0001010000111111"; -- -0.07362245055625362
	pesos_i(14319) := b"1111111111111111_1111111111111111_1110010010011001_1010000100011011"; -- -0.10703080262338746
	pesos_i(14320) := b"1111111111111111_1111111111111111_1111000101010100_0010100110011101"; -- -0.05730953126233948
	pesos_i(14321) := b"1111111111111111_1111111111111111_1111010000000000_1011110010000011"; -- -0.04686376375417348
	pesos_i(14322) := b"1111111111111111_1111111111111111_1111111110101000_1111110010001001"; -- -0.0013277210884821092
	pesos_i(14323) := b"0000000000000000_0000000000000000_0001101001100101_0001001000110111"; -- 0.10310472332779082
	pesos_i(14324) := b"0000000000000000_0000000000000000_0001111011010110_0100100111010111"; -- 0.12045728196308957
	pesos_i(14325) := b"1111111111111111_1111111111111111_1111011010100011_1011010000000000"; -- -0.03656458843858236
	pesos_i(14326) := b"0000000000000000_0000000000000000_0010000001010011_0011001001010111"; -- 0.1262694799033492
	pesos_i(14327) := b"0000000000000000_0000000000000000_0001000111110110_1100111010010111"; -- 0.07017222590211439
	pesos_i(14328) := b"1111111111111111_1111111111111111_1111001101101100_1101000110110100"; -- -0.04912080139311167
	pesos_i(14329) := b"1111111111111111_1111111111111111_1111011000000110_0011011010010011"; -- -0.038967694502767006
	pesos_i(14330) := b"1111111111111111_1111111111111111_1110100110010011_1001000100111111"; -- -0.08759205062086658
	pesos_i(14331) := b"1111111111111111_1111111111111111_1101011101110100_0011000100110011"; -- -0.15838329801499743
	pesos_i(14332) := b"0000000000000000_0000000000000000_0001011101000110_1100001101111001"; -- 0.09092351633210047
	pesos_i(14333) := b"0000000000000000_0000000000000000_0000100010011000_0010111001001111"; -- 0.03357209621435732
	pesos_i(14334) := b"1111111111111111_1111111111111111_1110000011000101_0110101000001111"; -- -0.12198769692459797
	pesos_i(14335) := b"0000000000000000_0000000000000000_0001101110111011_1011100110000010"; -- 0.10833320065994106
	pesos_i(14336) := b"0000000000000000_0000000000000000_0001100001110000_0101111110010010"; -- 0.09546468091896233
	pesos_i(14337) := b"0000000000000000_0000000000000000_0001111001110001_0010101001100010"; -- 0.1189142693945019
	pesos_i(14338) := b"1111111111111111_1111111111111111_1110001110111000_0010010111000100"; -- -0.11047138178570101
	pesos_i(14339) := b"1111111111111111_1111111111111111_1110100011110001_0001101010011111"; -- -0.09007104511414646
	pesos_i(14340) := b"0000000000000000_0000000000000000_0001110110101011_0110101011100101"; -- 0.11589687444672903
	pesos_i(14341) := b"0000000000000000_0000000000000000_0001010000101011_1011101001101011"; -- 0.0787922392825439
	pesos_i(14342) := b"1111111111111111_1111111111111111_1111100010011010_1111100100100011"; -- -0.02888529681502934
	pesos_i(14343) := b"1111111111111111_1111111111111111_1111001110011110_0100011101010110"; -- -0.04836610935010778
	pesos_i(14344) := b"0000000000000000_0000000000000000_0000110101111111_1001100011001101"; -- 0.05272822386888849
	pesos_i(14345) := b"1111111111111111_1111111111111111_1110010110110000_0100010011111111"; -- -0.102779090612429
	pesos_i(14346) := b"1111111111111111_1111111111111111_1111101011111010_1001110011100111"; -- -0.01961345059544574
	pesos_i(14347) := b"0000000000000000_0000000000000000_0010011100000000_0101100110011110"; -- 0.15234909158771548
	pesos_i(14348) := b"1111111111111111_1111111111111111_1110000011011101_0100101111100110"; -- -0.12162328376554055
	pesos_i(14349) := b"0000000000000000_0000000000000000_0001010001010100_1010101111100000"; -- 0.07941698288380596
	pesos_i(14350) := b"0000000000000000_0000000000000000_0001101000111000_1110011011010000"; -- 0.1024307496226588
	pesos_i(14351) := b"1111111111111111_1111111111111111_1111001001000110_1110010001011011"; -- -0.05360577367069472
	pesos_i(14352) := b"0000000000000000_0000000000000000_0001011110010000_0110011100100111"; -- 0.09204716403873885
	pesos_i(14353) := b"1111111111111111_1111111111111111_1101110110010101_1101110011111101"; -- -0.13443201842143368
	pesos_i(14354) := b"0000000000000000_0000000000000000_0001110111010000_1010110101101010"; -- 0.11646541440842825
	pesos_i(14355) := b"1111111111111111_1111111111111111_1101111011010101_0011101100011001"; -- -0.1295588554955135
	pesos_i(14356) := b"0000000000000000_0000000000000000_0000011110111101_1010111011001000"; -- 0.030238078792669574
	pesos_i(14357) := b"1111111111111111_1111111111111111_1110011101100011_0100101110100001"; -- -0.09614112211275377
	pesos_i(14358) := b"0000000000000000_0000000000000000_0000001100011000_1111000001000010"; -- 0.012099281528810481
	pesos_i(14359) := b"0000000000000000_0000000000000000_0000100111011000_0111000011010100"; -- 0.038458873474249464
	pesos_i(14360) := b"0000000000000000_0000000000000000_0001111111000111_0111001010100111"; -- 0.12413708278084247
	pesos_i(14361) := b"1111111111111111_1111111111111111_1101110001010011_0110011010000110"; -- -0.1393524096644678
	pesos_i(14362) := b"1111111111111111_1111111111111111_1101101110101011_0110100000011111"; -- -0.1419157908875615
	pesos_i(14363) := b"1111111111111111_1111111111111111_1111111110010111_0001111100100001"; -- -0.0016003174141715185
	pesos_i(14364) := b"0000000000000000_0000000000000000_0001000000101010_0000111011111011"; -- 0.06314176194997548
	pesos_i(14365) := b"0000000000000000_0000000000000000_0000101011100010_0111000111111111"; -- 0.04251778094428836
	pesos_i(14366) := b"0000000000000000_0000000000000000_0010011011101101_0001001001001001"; -- 0.15205492279683003
	pesos_i(14367) := b"0000000000000000_0000000000000000_0001100101010101_0100110001000111"; -- 0.09895779357178132
	pesos_i(14368) := b"0000000000000000_0000000000000000_0010001010110011_0000100101111010"; -- 0.13554438817491815
	pesos_i(14369) := b"0000000000000000_0000000000000000_0000010101011111_1011111000101001"; -- 0.020992169429893553
	pesos_i(14370) := b"1111111111111111_1111111111111111_1101100101100000_1010001100011001"; -- -0.15086918489809503
	pesos_i(14371) := b"1111111111111111_1111111111111111_1111100110000100_1101001011100111"; -- -0.025317019091304235
	pesos_i(14372) := b"1111111111111111_1111111111111111_1110000110111110_1000001000010111"; -- -0.11818682617819326
	pesos_i(14373) := b"1111111111111111_1111111111111111_1101101110101001_0000100111111001"; -- -0.14195192013987365
	pesos_i(14374) := b"0000000000000000_0000000000000000_0001000110000100_1001110000011100"; -- 0.06842971511468078
	pesos_i(14375) := b"0000000000000000_0000000000000000_0001010011011010_0010111001001110"; -- 0.08145417588719026
	pesos_i(14376) := b"1111111111111111_1111111111111111_1111001110000010_1111011001100011"; -- -0.048782921623209734
	pesos_i(14377) := b"1111111111111111_1111111111111111_1111001101100001_0010111010100000"; -- -0.04929836836808173
	pesos_i(14378) := b"1111111111111111_1111111111111111_1111011101100110_0001101010001110"; -- -0.03359827073087034
	pesos_i(14379) := b"1111111111111111_1111111111111111_1110010000011001_0011001111111000"; -- -0.10899043273766286
	pesos_i(14380) := b"1111111111111111_1111111111111111_1110101010000001_1111100011100111"; -- -0.08395428043518774
	pesos_i(14381) := b"1111111111111111_1111111111111111_1101110101111100_1111100000000001"; -- -0.1348118779282342
	pesos_i(14382) := b"0000000000000000_0000000000000000_0000110011111010_1100101110101010"; -- 0.0507018366541534
	pesos_i(14383) := b"0000000000000000_0000000000000000_0001011100001100_1100100001000010"; -- 0.0900387918788946
	pesos_i(14384) := b"0000000000000000_0000000000000000_0001101101010111_0010100110100010"; -- 0.10679874611040448
	pesos_i(14385) := b"1111111111111111_1111111111111111_1101011000111011_0011101100110100"; -- -0.16315870255832782
	pesos_i(14386) := b"0000000000000000_0000000000000000_0000111010010001_1101111001101001"; -- 0.056913281047844884
	pesos_i(14387) := b"0000000000000000_0000000000000000_0001001000000011_1100001011110011"; -- 0.07036989635156124
	pesos_i(14388) := b"0000000000000000_0000000000000000_0001011001110011_0010011111101101"; -- 0.08769464057743499
	pesos_i(14389) := b"1111111111111111_1111111111111111_1101111101000111_0110101111110000"; -- -0.12781644251146068
	pesos_i(14390) := b"1111111111111111_1111111111111111_1111110011100010_0010001001110110"; -- -0.012174459570063832
	pesos_i(14391) := b"1111111111111111_1111111111111111_1110010011001100_0101010110101010"; -- -0.10625710093940388
	pesos_i(14392) := b"0000000000000000_0000000000000000_0010000001001111_0000100001110111"; -- 0.12620594891802892
	pesos_i(14393) := b"1111111111111111_1111111111111111_1110101111000001_0001011110001101"; -- -0.07908489999666214
	pesos_i(14394) := b"0000000000000000_0000000000000000_0000010010100101_1100000111101111"; -- 0.01815425953879617
	pesos_i(14395) := b"0000000000000000_0000000000000000_0010001100000000_0010110010111010"; -- 0.13672141601805185
	pesos_i(14396) := b"1111111111111111_1111111111111111_1111110101001111_0100100111000100"; -- -0.01050890891924052
	pesos_i(14397) := b"0000000000000000_0000000000000000_0000000010010010_1110001100000010"; -- 0.002241313854510505
	pesos_i(14398) := b"1111111111111111_1111111111111111_1111100001010111_0010001010101000"; -- -0.02992041977047181
	pesos_i(14399) := b"1111111111111111_1111111111111111_1111000000000000_0011000101011100"; -- -0.06249705804801939
	pesos_i(14400) := b"0000000000000000_0000000000000000_0001011100001100_0010001101010111"; -- 0.09002896180227683
	pesos_i(14401) := b"1111111111111111_1111111111111111_1101001011010110_0101110000000101"; -- -0.17641663440197233
	pesos_i(14402) := b"0000000000000000_0000000000000000_0010000110111110_0111001100111001"; -- 0.1318122876746408
	pesos_i(14403) := b"0000000000000000_0000000000000000_0010010011101100_1110101000011100"; -- 0.14424002818893003
	pesos_i(14404) := b"0000000000000000_0000000000000000_0010011010000100_1111010110001011"; -- 0.1504662955553311
	pesos_i(14405) := b"0000000000000000_0000000000000000_0000001001110100_1101011011000001"; -- 0.0095953199468509
	pesos_i(14406) := b"1111111111111111_1111111111111111_1110111101011111_0111010000101001"; -- -0.06494974136974008
	pesos_i(14407) := b"0000000000000000_0000000000000000_0001011010110000_1011111001100110"; -- 0.08863439539319896
	pesos_i(14408) := b"0000000000000000_0000000000000000_0001011000111010_1111001101101010"; -- 0.08683701833546645
	pesos_i(14409) := b"1111111111111111_1111111111111111_1111001111001100_1010000101001111"; -- -0.04765884218047568
	pesos_i(14410) := b"1111111111111111_1111111111111111_1110101100001110_0010111010010000"; -- -0.08181485150711001
	pesos_i(14411) := b"1111111111111111_1111111111111111_1101110111101100_0110100101111101"; -- -0.13311138819673426
	pesos_i(14412) := b"1111111111111111_1111111111111111_1110111011101001_0000111010000101"; -- -0.06675633681477529
	pesos_i(14413) := b"0000000000000000_0000000000000000_0010010101111010_0010011000110000"; -- 0.1463950983344307
	pesos_i(14414) := b"0000000000000000_0000000000000000_0010100000101100_0010110000101101"; -- 0.1569240197612126
	pesos_i(14415) := b"1111111111111111_1111111111111111_1110011110001111_0110101100111010"; -- -0.09546785201634075
	pesos_i(14416) := b"1111111111111111_1111111111111111_1110111110011010_0000000011011101"; -- -0.06405634502029438
	pesos_i(14417) := b"1111111111111111_1111111111111111_1111001001101100_1111111111110101"; -- -0.05302429452838342
	pesos_i(14418) := b"0000000000000000_0000000000000000_0010000001110001_0001100001111110"; -- 0.12672570299390268
	pesos_i(14419) := b"0000000000000000_0000000000000000_0001011010100101_0101111101011001"; -- 0.08846088325621315
	pesos_i(14420) := b"0000000000000000_0000000000000000_0000111110100110_0111001111001111"; -- 0.06113361179298966
	pesos_i(14421) := b"0000000000000000_0000000000000000_0001001000110011_1110110100100010"; -- 0.07110483250170128
	pesos_i(14422) := b"1111111111111111_1111111111111111_1111011101000011_1111010001011001"; -- -0.034119346898883664
	pesos_i(14423) := b"1111111111111111_1111111111111111_1101010110010001_1001100101011111"; -- -0.1657470840434537
	pesos_i(14424) := b"0000000000000000_0000000000000000_0000110101011000_0011000000111100"; -- 0.05212689847693558
	pesos_i(14425) := b"1111111111111111_1111111111111111_1110111110001111_1101110001011111"; -- -0.06421110797742817
	pesos_i(14426) := b"1111111111111111_1111111111111111_1111100110011110_0100111100101100"; -- -0.024928142247458488
	pesos_i(14427) := b"0000000000000000_0000000000000000_0000110010111001_1111110000111110"; -- 0.049712910728833014
	pesos_i(14428) := b"1111111111111111_1111111111111111_1110101100100101_1000001101110000"; -- -0.08145884051789097
	pesos_i(14429) := b"1111111111111111_1111111111111111_1110100000111000_1010111000110000"; -- -0.0928851253740793
	pesos_i(14430) := b"0000000000000000_0000000000000000_0001001000101011_0010010011011000"; -- 0.0709708238923897
	pesos_i(14431) := b"0000000000000000_0000000000000000_0001111000101010_0000010000100101"; -- 0.11782861609778336
	pesos_i(14432) := b"1111111111111111_1111111111111111_1110001010011110_1001101011001001"; -- -0.11476738531879213
	pesos_i(14433) := b"1111111111111111_1111111111111111_1110101111111101_1011010010010011"; -- -0.07816001327027648
	pesos_i(14434) := b"0000000000000000_0000000000000000_0000011100100011_1100010110101101"; -- 0.027889589919482826
	pesos_i(14435) := b"0000000000000000_0000000000000000_0010000000011101_0110100111111111"; -- 0.12544882285651607
	pesos_i(14436) := b"1111111111111111_1111111111111111_1101111000101010_0000010101100101"; -- -0.13217130937510935
	pesos_i(14437) := b"0000000000000000_0000000000000000_0001010011110111_1000011100110100"; -- 0.08190197961304525
	pesos_i(14438) := b"0000000000000000_0000000000000000_0000101101001000_0101000100110010"; -- 0.044072222449082946
	pesos_i(14439) := b"1111111111111111_1111111111111111_1111101011101000_1101110001001011"; -- -0.019884330433292654
	pesos_i(14440) := b"1111111111111111_1111111111111111_1111010000100111_1111101011011010"; -- -0.046264955305838046
	pesos_i(14441) := b"1111111111111111_1111111111111111_1101101000100010_1001111000010101"; -- -0.14790927872840448
	pesos_i(14442) := b"0000000000000000_0000000000000000_0000100010010010_0001000110110100"; -- 0.033478838490374405
	pesos_i(14443) := b"1111111111111111_1111111111111111_1110011000000101_0111110011100001"; -- -0.1014787626636297
	pesos_i(14444) := b"1111111111111111_1111111111111111_1101011101001010_1111101001110011"; -- -0.1590121716702264
	pesos_i(14445) := b"0000000000000000_0000000000000000_0001001101110111_0100110111010110"; -- 0.07603918533628601
	pesos_i(14446) := b"1111111111111111_1111111111111111_1110011111000110_0110101101100100"; -- -0.09462860871331617
	pesos_i(14447) := b"0000000000000000_0000000000000000_0001000100111011_0001001001011111"; -- 0.06730761360230568
	pesos_i(14448) := b"1111111111111111_1111111111111111_1101011010000110_1001010011000001"; -- -0.16200895582411765
	pesos_i(14449) := b"1111111111111111_1111111111111111_1110111111000010_0001011010100111"; -- -0.06344469472527284
	pesos_i(14450) := b"1111111111111111_1111111111111111_1101111111100001_0101011110000011"; -- -0.1254678064408401
	pesos_i(14451) := b"1111111111111111_1111111111111111_1110101010111101_0100110011110011"; -- -0.08304900236625513
	pesos_i(14452) := b"1111111111111111_1111111111111111_1111111001000001_1100100000001100"; -- -0.006808754910056439
	pesos_i(14453) := b"0000000000000000_0000000000000000_0001111001011101_1001100010011111"; -- 0.1186156643944563
	pesos_i(14454) := b"1111111111111111_1111111111111111_1110010001110101_0101001001100111"; -- -0.10758481006868789
	pesos_i(14455) := b"1111111111111111_1111111111111111_1101111000100101_0101001011000011"; -- -0.13224299191670794
	pesos_i(14456) := b"0000000000000000_0000000000000000_0001010000011001_0000110001010110"; -- 0.07850720490255861
	pesos_i(14457) := b"0000000000000000_0000000000000000_0001101000001110_0100110101110000"; -- 0.10178073862006082
	pesos_i(14458) := b"0000000000000000_0000000000000000_0001111100100001_1001101100101101"; -- 0.12160653913136774
	pesos_i(14459) := b"0000000000000000_0000000000000000_0001110000000001_0010000000001110"; -- 0.10939216947137627
	pesos_i(14460) := b"0000000000000000_0000000000000000_0001110000011000_0010110110100111"; -- 0.10974393204370396
	pesos_i(14461) := b"1111111111111111_1111111111111111_1101111111101101_1010100001101010"; -- -0.12527987861995274
	pesos_i(14462) := b"1111111111111111_1111111111111111_1110010001011000_0100110100111000"; -- -0.10802762406299816
	pesos_i(14463) := b"1111111111111111_1111111111111111_1110001110100001_1111000101101110"; -- -0.11081019462558178
	pesos_i(14464) := b"0000000000000000_0000000000000000_0000100110010110_0011100001110111"; -- 0.03744843397440167
	pesos_i(14465) := b"1111111111111111_1111111111111111_1110001111011111_1010011011010000"; -- -0.10986859731743442
	pesos_i(14466) := b"1111111111111111_1111111111111111_1111011110010110_0111010010001000"; -- -0.03286048591169776
	pesos_i(14467) := b"1111111111111111_1111111111111111_1111101110011000_1011111010001101"; -- -0.017200556288042727
	pesos_i(14468) := b"0000000000000000_0000000000000000_0001011111111111_1011101000001001"; -- 0.09374582976038376
	pesos_i(14469) := b"1111111111111111_1111111111111111_1111010100000111_1000100101100011"; -- -0.0428537495483791
	pesos_i(14470) := b"1111111111111111_1111111111111111_1111101111000010_0011110111000011"; -- -0.01656736361026203
	pesos_i(14471) := b"1111111111111111_1111111111111111_1110110010110111_0011000001000001"; -- -0.07532976554834227
	pesos_i(14472) := b"0000000000000000_0000000000000000_0001110100111101_0000111101010001"; -- 0.11421294905266766
	pesos_i(14473) := b"1111111111111111_1111111111111111_1111011111010010_1101101101110100"; -- -0.031938823844585296
	pesos_i(14474) := b"0000000000000000_0000000000000000_0000011110000011_1010010001110011"; -- 0.029352453192264177
	pesos_i(14475) := b"0000000000000000_0000000000000000_0001000111110010_1011000110100100"; -- 0.07010946518486691
	pesos_i(14476) := b"1111111111111111_1111111111111111_1101101010000100_0110101011000001"; -- -0.14641697685240676
	pesos_i(14477) := b"1111111111111111_1111111111111111_1101101000001011_0001111101011110"; -- -0.1482677837356926
	pesos_i(14478) := b"1111111111111111_1111111111111111_1110001110011011_1001100000100001"; -- -0.11090707017777061
	pesos_i(14479) := b"0000000000000000_0000000000000000_0001000010101010_1000101000101100"; -- 0.06510222974576547
	pesos_i(14480) := b"1111111111111111_1111111111111111_1101100100100111_1111110100100000"; -- -0.15173356972089502
	pesos_i(14481) := b"0000000000000000_0000000000000000_0000111111011101_1001010011010111"; -- 0.06197481390123376
	pesos_i(14482) := b"1111111111111111_1111111111111111_1111110111010101_1100111100100010"; -- -0.008456281894483478
	pesos_i(14483) := b"0000000000000000_0000000000000000_0010000001011101_0110111100000000"; -- 0.12642568351402186
	pesos_i(14484) := b"0000000000000000_0000000000000000_0001010001111110_0101001001000101"; -- 0.08005251101174397
	pesos_i(14485) := b"1111111111111111_1111111111111111_1110100011010111_1100101000011110"; -- -0.09045731332960724
	pesos_i(14486) := b"0000000000000000_0000000000000000_0000100100000010_0011010101011110"; -- 0.03518994862065684
	pesos_i(14487) := b"1111111111111111_1111111111111111_1101101101100110_1001101000111101"; -- -0.1429656601998063
	pesos_i(14488) := b"0000000000000000_0000000000000000_0000001110100110_1111001101111101"; -- 0.014266222122519705
	pesos_i(14489) := b"1111111111111111_1111111111111111_1111100100001010_1000010100000100"; -- -0.027183233815287082
	pesos_i(14490) := b"0000000000000000_0000000000000000_0001100101101100_1110100101101011"; -- 0.09931811209557667
	pesos_i(14491) := b"0000000000000000_0000000000000000_0010010100111011_0100110001100000"; -- 0.14543607083777374
	pesos_i(14492) := b"1111111111111111_1111111111111111_1111011011110011_1000110011011011"; -- -0.03534621864939259
	pesos_i(14493) := b"0000000000000000_0000000000000000_0000010010010101_0010101101001010"; -- 0.017901139761624354
	pesos_i(14494) := b"0000000000000000_0000000000000000_0000110100101011_0100110111010011"; -- 0.051442016640329824
	pesos_i(14495) := b"1111111111111111_1111111111111111_1110011101111100_1000011110000010"; -- -0.09575608315993249
	pesos_i(14496) := b"1111111111111111_1111111111111111_1110001001100011_1011010100000101"; -- -0.11566609035849784
	pesos_i(14497) := b"1111111111111111_1111111111111111_1110100011101110_1100110111000011"; -- -0.09010614395307326
	pesos_i(14498) := b"0000000000000000_0000000000000000_0001000000010011_0011111101011001"; -- 0.0627936927111173
	pesos_i(14499) := b"1111111111111111_1111111111111111_1110101010010010_1110011100000111"; -- -0.0836959465949571
	pesos_i(14500) := b"1111111111111111_1111111111111111_1101111100101100_1101010111101011"; -- -0.12822211283626428
	pesos_i(14501) := b"1111111111111111_1111111111111111_1111010110000000_0011000110001000"; -- -0.041012672739450126
	pesos_i(14502) := b"0000000000000000_0000000000000000_0000111101010101_0100000111111111"; -- 0.05989468079803638
	pesos_i(14503) := b"1111111111111111_1111111111111111_1110000111111101_1111100110100110"; -- -0.11721839621556186
	pesos_i(14504) := b"1111111111111111_1111111111111111_1110001111101010_1101110011001100"; -- -0.10969753278989212
	pesos_i(14505) := b"1111111111111111_1111111111111111_1110001100000110_0110011100100110"; -- -0.11318354921409675
	pesos_i(14506) := b"0000000000000000_0000000000000000_0000001100001010_1011111010011011"; -- 0.01188269890204015
	pesos_i(14507) := b"0000000000000000_0000000000000000_0000000101101010_0011100010110110"; -- 0.005527061890729264
	pesos_i(14508) := b"1111111111111111_1111111111111111_1111010111110111_0001101000110100"; -- -0.039198267265241324
	pesos_i(14509) := b"1111111111111111_1111111111111111_1111001111111000_0001111100001100"; -- -0.0469952198557922
	pesos_i(14510) := b"0000000000000000_0000000000000000_0000111001010011_1000100110100110"; -- 0.05596218393641623
	pesos_i(14511) := b"0000000000000000_0000000000000000_0001001110011111_1101101100101001"; -- 0.07665796049267953
	pesos_i(14512) := b"0000000000000000_0000000000000000_0001110100001110_1100101010011110"; -- 0.11350695001424743
	pesos_i(14513) := b"1111111111111111_1111111111111111_1101100111100001_0011000111101101"; -- -0.1489075467011873
	pesos_i(14514) := b"0000000000000000_0000000000000000_0001000100000000_1100111110110101"; -- 0.06641863029473828
	pesos_i(14515) := b"0000000000000000_0000000000000000_0010000000011111_1010000110010111"; -- 0.1254826540795719
	pesos_i(14516) := b"1111111111111111_1111111111111111_1110000101110011_0010100010110001"; -- -0.11933656388972226
	pesos_i(14517) := b"1111111111111111_1111111111111111_1111101001110001_1110010011011100"; -- -0.021699615840171486
	pesos_i(14518) := b"1111111111111111_1111111111111111_1111101100000100_1010011111000010"; -- -0.019460215746256095
	pesos_i(14519) := b"1111111111111111_1111111111111111_1111010101111001_0000101111011100"; -- -0.04112172973811903
	pesos_i(14520) := b"0000000000000000_0000000000000000_0010001001111010_1100110000001010"; -- 0.1346862338362922
	pesos_i(14521) := b"0000000000000000_0000000000000000_0000110111110001_1100100000001101"; -- 0.054470542010678705
	pesos_i(14522) := b"1111111111111111_1111111111111111_1110011001100000_0000101010101100"; -- -0.10009702026397559
	pesos_i(14523) := b"0000000000000000_0000000000000000_0000011001000111_1010111010101101"; -- 0.02453128540215583
	pesos_i(14524) := b"1111111111111111_1111111111111111_1101110110100011_0000001010010010"; -- -0.13423141412136644
	pesos_i(14525) := b"0000000000000000_0000000000000000_0001111001011101_1000101000101110"; -- 0.11861480358844718
	pesos_i(14526) := b"0000000000000000_0000000000000000_0000000010010000_0001100011110101"; -- 0.0021987531163761187
	pesos_i(14527) := b"0000000000000000_0000000000000000_0000011000000001_1000101001100000"; -- 0.023461006645553673
	pesos_i(14528) := b"0000000000000000_0000000000000000_0001010100010110_0011100110111000"; -- 0.08237038357125098
	pesos_i(14529) := b"0000000000000000_0000000000000000_0001001100111110_0111110101000001"; -- 0.07517226053144165
	pesos_i(14530) := b"1111111111111111_1111111111111111_1101110001110101_1011001111011111"; -- -0.13882900047181534
	pesos_i(14531) := b"0000000000000000_0000000000000000_0000011111011010_1000011110011011"; -- 0.030678248633372603
	pesos_i(14532) := b"0000000000000000_0000000000000000_0000101100011001_0011001100010011"; -- 0.04335326389366918
	pesos_i(14533) := b"0000000000000000_0000000000000000_0000101100011101_1010110101110101"; -- 0.04342159374624115
	pesos_i(14534) := b"1111111111111111_1111111111111111_1110001101110001_0101101100011001"; -- -0.11155157703512925
	pesos_i(14535) := b"1111111111111111_1111111111111111_1110001100111010_1100001110011010"; -- -0.11238458142232681
	pesos_i(14536) := b"1111111111111111_1111111111111111_1110011001101010_0010100110011000"; -- -0.09994258910833112
	pesos_i(14537) := b"1111111111111111_1111111111111111_1110010000000001_0010110110111101"; -- -0.10935701489425943
	pesos_i(14538) := b"1111111111111111_1111111111111111_1111010011101110_0001110000000010"; -- -0.04324173881006454
	pesos_i(14539) := b"0000000000000000_0000000000000000_0000111011100001_0111100100000100"; -- 0.05812794067529205
	pesos_i(14540) := b"0000000000000000_0000000000000000_0001000010010000_0000110010001110"; -- 0.06469801386835504
	pesos_i(14541) := b"1111111111111111_1111111111111111_1101111000110111_1001011000101100"; -- -0.13196431571058442
	pesos_i(14542) := b"1111111111111111_1111111111111111_1110111110110101_1100110100110000"; -- -0.06363217904131194
	pesos_i(14543) := b"1111111111111111_1111111111111111_1111011101010110_1100111101100100"; -- -0.033831632676624944
	pesos_i(14544) := b"1111111111111111_1111111111111111_1110111110011010_0000011101101100"; -- -0.06405595401983084
	pesos_i(14545) := b"1111111111111111_1111111111111111_1110011111010100_1010110110010011"; -- -0.09441104087461497
	pesos_i(14546) := b"1111111111111111_1111111111111111_1111101101100100_1100001001010011"; -- -0.017993788489018902
	pesos_i(14547) := b"1111111111111111_1111111111111111_1101110011111000_0000110111101011"; -- -0.13683999072783917
	pesos_i(14548) := b"0000000000000000_0000000000000000_0010000001100001_0000011101111111"; -- 0.12648054940701414
	pesos_i(14549) := b"1111111111111111_1111111111111111_1101110111000000_0100111001101000"; -- -0.133784389162771
	pesos_i(14550) := b"1111111111111111_1111111111111111_1110110011100011_0110010000010000"; -- -0.07465529074560144
	pesos_i(14551) := b"1111111111111111_1111111111111111_1110001101001000_1100000111000011"; -- -0.1121710680085728
	pesos_i(14552) := b"1111111111111111_1111111111111111_1101100010101100_1001001100111110"; -- -0.153616711886447
	pesos_i(14553) := b"0000000000000000_0000000000000000_0001010100001010_0111100110001000"; -- 0.08219108171679512
	pesos_i(14554) := b"0000000000000000_0000000000000000_0000010101111011_0010000011010110"; -- 0.021410038123995036
	pesos_i(14555) := b"0000000000000000_0000000000000000_0000110011111110_0010110101001111"; -- 0.05075343307203431
	pesos_i(14556) := b"1111111111111111_1111111111111111_1101110100000101_0110001111110011"; -- -0.1366364987260986
	pesos_i(14557) := b"1111111111111111_1111111111111111_1110011010100001_1110001001011010"; -- -0.09909234336431097
	pesos_i(14558) := b"1111111111111111_1111111111111111_1101011011101110_0101010111010001"; -- -0.16042579314017033
	pesos_i(14559) := b"0000000000000000_0000000000000000_0000110001111011_0111010100111111"; -- 0.04875881954136963
	pesos_i(14560) := b"0000000000000000_0000000000000000_0000110011010000_0101000001111011"; -- 0.050053625113229853
	pesos_i(14561) := b"0000000000000000_0000000000000000_0000110110010001_0000010011001111"; -- 0.05299406103371408
	pesos_i(14562) := b"0000000000000000_0000000000000000_0001101010110101_0011011010101101"; -- 0.10432759978171183
	pesos_i(14563) := b"1111111111111111_1111111111111111_1110111101000111_1010011110000100"; -- -0.0653128911599004
	pesos_i(14564) := b"1111111111111111_1111111111111111_1111101110110011_1010111100100100"; -- -0.01678948764048004
	pesos_i(14565) := b"1111111111111111_1111111111111111_1101011101011010_1101001111000101"; -- -0.1587703366367863
	pesos_i(14566) := b"1111111111111111_1111111111111111_1110011010011110_0000000100101010"; -- -0.09915154198279469
	pesos_i(14567) := b"0000000000000000_0000000000000000_0001100011111110_1110000001001100"; -- 0.09763910156274686
	pesos_i(14568) := b"0000000000000000_0000000000000000_0010000000000010_1011111000011101"; -- 0.12504184922672004
	pesos_i(14569) := b"0000000000000000_0000000000000000_0000100110011011_0101110010000110"; -- 0.03752687702909971
	pesos_i(14570) := b"0000000000000000_0000000000000000_0001010111110011_1010010111111100"; -- 0.08574902928915305
	pesos_i(14571) := b"0000000000000000_0000000000000000_0000000110101001_1100100010010001"; -- 0.006496940011448581
	pesos_i(14572) := b"0000000000000000_0000000000000000_0010010001101001_1010110110001010"; -- 0.14223751650246702
	pesos_i(14573) := b"1111111111111111_1111111111111111_1110000010100010_0101101111101101"; -- -0.12252259687794606
	pesos_i(14574) := b"1111111111111111_1111111111111111_1111101110100101_0111100110111010"; -- -0.017006294320775665
	pesos_i(14575) := b"0000000000000000_0000000000000000_0001100111101110_1000011011011011"; -- 0.10129587977058983
	pesos_i(14576) := b"1111111111111111_1111111111111111_1110000010111010_1011101101111111"; -- -0.12215068953769037
	pesos_i(14577) := b"1111111111111111_1111111111111111_1101101011101011_0100000111010000"; -- -0.1448477618032725
	pesos_i(14578) := b"0000000000000000_0000000000000000_0000110100100001_1011001001010101"; -- 0.051295419389856836
	pesos_i(14579) := b"0000000000000000_0000000000000000_0000101001100110_1101010110011100"; -- 0.04063162856693927
	pesos_i(14580) := b"0000000000000000_0000000000000000_0000101011101000_0100101100001100"; -- 0.04260701227229929
	pesos_i(14581) := b"1111111111111111_1111111111111111_1111111101100011_1001110111011100"; -- -0.0023862208459303033
	pesos_i(14582) := b"0000000000000000_0000000000000000_0001001100100000_0100101101001011"; -- 0.0747115191173145
	pesos_i(14583) := b"1111111111111111_1111111111111111_1111101011100001_0110011100001100"; -- -0.019998130279026752
	pesos_i(14584) := b"1111111111111111_1111111111111111_1110001110100100_1011100011101110"; -- -0.11076778586062391
	pesos_i(14585) := b"1111111111111111_1111111111111111_1111011000000011_0101000110001001"; -- -0.03901186378929832
	pesos_i(14586) := b"0000000000000000_0000000000000000_0001000011010100_1110100110100100"; -- 0.0657487893942231
	pesos_i(14587) := b"0000000000000000_0000000000000000_0000001110010001_0000010011111100"; -- 0.013931571456610597
	pesos_i(14588) := b"1111111111111111_1111111111111111_1110111100111111_1000110110010010"; -- -0.06543650800041122
	pesos_i(14589) := b"0000000000000000_0000000000000000_0000010001111010_0001100011010001"; -- 0.017488051400232456
	pesos_i(14590) := b"0000000000000000_0000000000000000_0000111111001011_0010111010111011"; -- 0.061694069429199236
	pesos_i(14591) := b"1111111111111111_1111111111111111_1111000111111110_1110011101011011"; -- -0.054704227642994124
	pesos_i(14592) := b"1111111111111111_1111111111111111_1110101101101110_0100010111000111"; -- -0.08034862405865918
	pesos_i(14593) := b"0000000000000000_0000000000000000_0000000101111000_1111101011011100"; -- 0.005752257137094415
	pesos_i(14594) := b"0000000000000000_0000000000000000_0010000101011001_1010011001101001"; -- 0.13027420095114234
	pesos_i(14595) := b"0000000000000000_0000000000000000_0001001011111011_1000010110000101"; -- 0.07415041446033022
	pesos_i(14596) := b"1111111111111111_1111111111111111_1110010000110111_1111000011111010"; -- -0.10852140336533414
	pesos_i(14597) := b"0000000000000000_0000000000000000_0001111011110101_0111011111011110"; -- 0.12093304804276572
	pesos_i(14598) := b"1111111111111111_1111111111111111_1111111101000001_0111011001001110"; -- -0.002907377216387258
	pesos_i(14599) := b"0000000000000000_0000000000000000_0001010110000101_0011000011001001"; -- 0.08406357677546106
	pesos_i(14600) := b"0000000000000000_0000000000000000_0001100100101011_1110100110101110"; -- 0.09832630639565001
	pesos_i(14601) := b"1111111111111111_1111111111111111_1111001011011100_0111110101011101"; -- -0.05132309411165387
	pesos_i(14602) := b"1111111111111111_1111111111111111_1110000010000001_0011000101110111"; -- -0.12302866794290283
	pesos_i(14603) := b"1111111111111111_1111111111111111_1110110111101100_0010101101011001"; -- -0.07061509211425313
	pesos_i(14604) := b"1111111111111111_1111111111111111_1111101010001110_0111101001101110"; -- -0.021263454594073895
	pesos_i(14605) := b"0000000000000000_0000000000000000_0001100101010011_1110110000111011"; -- 0.09893681001612654
	pesos_i(14606) := b"0000000000000000_0000000000000000_0010000111100011_0010111000111001"; -- 0.1323727501357347
	pesos_i(14607) := b"1111111111111111_1111111111111111_1110010111001011_0001010000011011"; -- -0.10237001734646314
	pesos_i(14608) := b"0000000000000000_0000000000000000_0000010100010001_0001000100111001"; -- 0.019791675893789926
	pesos_i(14609) := b"0000000000000000_0000000000000000_0001110010100000_1000100011010011"; -- 0.11182456172269634
	pesos_i(14610) := b"1111111111111111_1111111111111111_1111101100101001_1001011011110111"; -- -0.0188966414506763
	pesos_i(14611) := b"1111111111111111_1111111111111111_1110001111111101_0101000000101001"; -- -0.1094159983435806
	pesos_i(14612) := b"1111111111111111_1111111111111111_1111011111000011_0110110100000111"; -- -0.03217428754783904
	pesos_i(14613) := b"1111111111111111_1111111111111111_1111111000110000_0110100011111011"; -- -0.007073820752981273
	pesos_i(14614) := b"0000000000000000_0000000000000000_0001111010001110_1110110011100111"; -- 0.11936836843263744
	pesos_i(14615) := b"0000000000000000_0000000000000000_0001110011101111_0101010100100001"; -- 0.1130269246395397
	pesos_i(14616) := b"0000000000000000_0000000000000000_0001010100111010_0111100111111100"; -- 0.08292353062081786
	pesos_i(14617) := b"0000000000000000_0000000000000000_0000001010011101_0101010111001010"; -- 0.010213243205425054
	pesos_i(14618) := b"0000000000000000_0000000000000000_0000010111010101_1001010010001000"; -- 0.022790225225382352
	pesos_i(14619) := b"0000000000000000_0000000000000000_0000001000001001_1101110100010011"; -- 0.007963006245892615
	pesos_i(14620) := b"1111111111111111_1111111111111111_1111010000010101_0101001001001100"; -- -0.046549660175718786
	pesos_i(14621) := b"1111111111111111_1111111111111111_1101001101101011_1010001111111110"; -- -0.17413878490941753
	pesos_i(14622) := b"1111111111111111_1111111111111111_1101111100001100_0011111011110101"; -- -0.1287193919365192
	pesos_i(14623) := b"0000000000000000_0000000000000000_0010001101111100_0110010110101010"; -- 0.13861689950260458
	pesos_i(14624) := b"1111111111111111_1111111111111111_1111011000110100_1011110100000111"; -- -0.03825777602264203
	pesos_i(14625) := b"1111111111111111_1111111111111111_1110110010100110_1011000010011000"; -- -0.07558151510708547
	pesos_i(14626) := b"1111111111111111_1111111111111111_1110111010100101_0100001011101101"; -- -0.0677908106504976
	pesos_i(14627) := b"1111111111111111_1111111111111111_1111110011001111_1101011000000101"; -- -0.01245367404972822
	pesos_i(14628) := b"0000000000000000_0000000000000000_0010001010110101_0000000101000000"; -- 0.1355744153214428
	pesos_i(14629) := b"0000000000000000_0000000000000000_0000110011100111_0111010101010110"; -- 0.05040677404151986
	pesos_i(14630) := b"1111111111111111_1111111111111111_1111000010110000_1100011011111000"; -- -0.059802593586472906
	pesos_i(14631) := b"1111111111111111_1111111111111111_1111100110011110_1111100111110100"; -- -0.02491796285000079
	pesos_i(14632) := b"0000000000000000_0000000000000000_0000011111111010_0010101000111011"; -- 0.0311609645073305
	pesos_i(14633) := b"0000000000000000_0000000000000000_0001011011010100_1011111101110000"; -- 0.08918377392673406
	pesos_i(14634) := b"0000000000000000_0000000000000000_0001010000000011_0101000100010000"; -- 0.07817560801963505
	pesos_i(14635) := b"1111111111111111_1111111111111111_1110100010001111_0011000010101111"; -- -0.09156509133436319
	pesos_i(14636) := b"1111111111111111_1111111111111111_1111101011100101_0001010010110001"; -- -0.019942004063877056
	pesos_i(14637) := b"1111111111111111_1111111111111111_1111011011001110_1111010101110011"; -- -0.035904559602597856
	pesos_i(14638) := b"0000000000000000_0000000000000000_0001110011111000_1110100011100000"; -- 0.11317306001964944
	pesos_i(14639) := b"1111111111111111_1111111111111111_1111000101000100_0110011000101010"; -- -0.05755006289922892
	pesos_i(14640) := b"0000000000000000_0000000000000000_0001100101000111_1101101111001000"; -- 0.09875272399445766
	pesos_i(14641) := b"1111111111111111_1111111111111111_1110101110110011_1101000111100111"; -- -0.0792874155459764
	pesos_i(14642) := b"0000000000000000_0000000000000000_0001000111000000_0101101100110001"; -- 0.06934137285343717
	pesos_i(14643) := b"1111111111111111_1111111111111111_1111011011110011_1011000011000101"; -- -0.03534407806561163
	pesos_i(14644) := b"1111111111111111_1111111111111111_1110001110010101_1010001110000100"; -- -0.11099794402447288
	pesos_i(14645) := b"1111111111111111_1111111111111111_1101101011101111_0000010101011111"; -- -0.14479032936179778
	pesos_i(14646) := b"1111111111111111_1111111111111111_1101100000100010_0111001001011100"; -- -0.15572438472748518
	pesos_i(14647) := b"1111111111111111_1111111111111111_1110010000000011_1111110111010000"; -- -0.10931409529402439
	pesos_i(14648) := b"0000000000000000_0000000000000000_0001110000010000_1000100110111111"; -- 0.10962735100330914
	pesos_i(14649) := b"1111111111111111_1111111111111111_1101110011011010_1010101001000101"; -- -0.13728843522160308
	pesos_i(14650) := b"1111111111111111_1111111111111111_1110100000010111_1110010010100101"; -- -0.09338541950220167
	pesos_i(14651) := b"0000000000000000_0000000000000000_0000011110110011_0001010000110000"; -- 0.03007627652104376
	pesos_i(14652) := b"0000000000000000_0000000000000000_0001100010010101_1110000000101100"; -- 0.09603692129796175
	pesos_i(14653) := b"1111111111111111_1111111111111111_1111010111010010_1010100100101111"; -- -0.0397543200739857
	pesos_i(14654) := b"0000000000000000_0000000000000000_0010011010100011_0000001100011011"; -- 0.15092486764633217
	pesos_i(14655) := b"0000000000000000_0000000000000000_0000011100011111_1011011010111110"; -- 0.027827664741663618
	pesos_i(14656) := b"1111111111111111_1111111111111111_1110000100101010_1111111011000111"; -- -0.12043769494824326
	pesos_i(14657) := b"1111111111111111_1111111111111111_1101111000111100_1110000001110000"; -- -0.1318835951293636
	pesos_i(14658) := b"1111111111111111_1111111111111111_1110000000110100_1101010010111101"; -- -0.12419386286530623
	pesos_i(14659) := b"1111111111111111_1111111111111111_1111010011001111_1100000110111111"; -- -0.04370488258409595
	pesos_i(14660) := b"0000000000000000_0000000000000000_0001110100011011_1111100011100100"; -- 0.11370807226908064
	pesos_i(14661) := b"1111111111111111_1111111111111111_1111000010011101_1010100010100011"; -- -0.06009431849352433
	pesos_i(14662) := b"0000000000000000_0000000000000000_0010100011101111_0011001111010110"; -- 0.15989994019293755
	pesos_i(14663) := b"0000000000000000_0000000000000000_0001101010011101_0101100010000010"; -- 0.10396340536079132
	pesos_i(14664) := b"0000000000000000_0000000000000000_0000111111011011_1011101010101000"; -- 0.06194655027695227
	pesos_i(14665) := b"1111111111111111_1111111111111111_1110011000001111_1101111001100101"; -- -0.1013203625155161
	pesos_i(14666) := b"0000000000000000_0000000000000000_0001110100001011_1111011010011000"; -- 0.11346379471853482
	pesos_i(14667) := b"1111111111111111_1111111111111111_1101101010001001_0110001000100000"; -- -0.14634119727359027
	pesos_i(14668) := b"0000000000000000_0000000000000000_0001010001011110_0011001111101000"; -- 0.07956241996611271
	pesos_i(14669) := b"1111111111111111_1111111111111111_1110010010111101_1000011001110010"; -- -0.10648307531094274
	pesos_i(14670) := b"1111111111111111_1111111111111111_1110110100010101_1111000100000111"; -- -0.07388394908425604
	pesos_i(14671) := b"0000000000000000_0000000000000000_0010011000110101_1001110101110000"; -- 0.14925559976287678
	pesos_i(14672) := b"1111111111111111_1111111111111111_1111001000000111_1111010011010001"; -- -0.05456609627206003
	pesos_i(14673) := b"1111111111111111_1111111111111111_1111101010110000_1011110011101101"; -- -0.02074069231715258
	pesos_i(14674) := b"1111111111111111_1111111111111111_1110110001100101_0101100110111110"; -- -0.07657851324055549
	pesos_i(14675) := b"1111111111111111_1111111111111111_1111010101000111_1101101000001001"; -- -0.04187238008932231
	pesos_i(14676) := b"0000000000000000_0000000000000000_0000001100101000_0100110100011001"; -- 0.012333696872370663
	pesos_i(14677) := b"0000000000000000_0000000000000000_0000000101101101_0010010101010001"; -- 0.005571682341537056
	pesos_i(14678) := b"0000000000000000_0000000000000000_0010000101001000_0001101100011010"; -- 0.13000649828846428
	pesos_i(14679) := b"1111111111111111_1111111111111111_1111110100011101_0001100011100001"; -- -0.011274762293966088
	pesos_i(14680) := b"0000000000000000_0000000000000000_0010001011001110_1111111111001011"; -- 0.1359710570266713
	pesos_i(14681) := b"1111111111111111_1111111111111111_1111011100000001_1001011010001110"; -- -0.03513201746772055
	pesos_i(14682) := b"0000000000000000_0000000000000000_0010010100101111_1000111010011101"; -- 0.14525691352763942
	pesos_i(14683) := b"1111111111111111_1111111111111111_1110100010110111_1100110000101010"; -- -0.0909454724829211
	pesos_i(14684) := b"1111111111111111_1111111111111111_1111111000010011_0111011100100110"; -- -0.007515481154188176
	pesos_i(14685) := b"0000000000000000_0000000000000000_0000010100110001_0100010001011111"; -- 0.020283006003429197
	pesos_i(14686) := b"1111111111111111_1111111111111111_1101111101111011_0101110111111100"; -- -0.12702381711119493
	pesos_i(14687) := b"0000000000000000_0000000000000000_0000100100011100_0101100111000011"; -- 0.035588846380605034
	pesos_i(14688) := b"0000000000000000_0000000000000000_0001101101001101_1100101010000011"; -- 0.10665574739922946
	pesos_i(14689) := b"1111111111111111_1111111111111111_1110001010100101_1010110101110101"; -- -0.11465946100881784
	pesos_i(14690) := b"0000000000000000_0000000000000000_0000110010101111_0111011011010110"; -- 0.04955237128919452
	pesos_i(14691) := b"1111111111111111_1111111111111111_1111010001100110_0011101001110010"; -- -0.045315119864616164
	pesos_i(14692) := b"0000000000000000_0000000000000000_0010001011100000_0010000101100001"; -- 0.13623245826197197
	pesos_i(14693) := b"0000000000000000_0000000000000000_0001100011000110_0000101111101101"; -- 0.0967719510111749
	pesos_i(14694) := b"1111111111111111_1111111111111111_1111101110110110_1001110010000001"; -- -0.01674482208984693
	pesos_i(14695) := b"0000000000000000_0000000000000000_0001000100000101_1001100110100000"; -- 0.06649170062145354
	pesos_i(14696) := b"0000000000000000_0000000000000000_0000100111011011_1011111001011100"; -- 0.03850927108729279
	pesos_i(14697) := b"0000000000000000_0000000000000000_0000110011011001_0000110101000010"; -- 0.05018694742187849
	pesos_i(14698) := b"1111111111111111_1111111111111111_1110111111110000_1100010001110000"; -- -0.06273243209183758
	pesos_i(14699) := b"0000000000000000_0000000000000000_0000100110001111_0010001110111001"; -- 0.03734038603446434
	pesos_i(14700) := b"0000000000000000_0000000000000000_0001000101110001_0111101101111011"; -- 0.06813785317422763
	pesos_i(14701) := b"1111111111111111_1111111111111111_1110101000110110_1000111000110000"; -- -0.08510505039388422
	pesos_i(14702) := b"0000000000000000_0000000000000000_0000000001010111_0100001110100000"; -- 0.0013315454986810946
	pesos_i(14703) := b"1111111111111111_1111111111111111_1111001001011000_0001010001010110"; -- -0.05334351440085276
	pesos_i(14704) := b"0000000000000000_0000000000000000_0010010110110100_1010101000100010"; -- 0.14728797280549955
	pesos_i(14705) := b"0000000000000000_0000000000000000_0000111000010110_0001110110110010"; -- 0.05502496333841773
	pesos_i(14706) := b"1111111111111111_1111111111111111_1111101110010100_1000100011100111"; -- -0.017264789288298034
	pesos_i(14707) := b"1111111111111111_1111111111111111_1111001110111111_1111100010001010"; -- -0.047852007228505106
	pesos_i(14708) := b"1111111111111111_1111111111111111_1111101111110101_1111010100011000"; -- -0.015778237845738605
	pesos_i(14709) := b"0000000000000000_0000000000000000_0010001110000110_1111110101110110"; -- 0.13877853513061816
	pesos_i(14710) := b"0000000000000000_0000000000000000_0001100111101111_0000101110101110"; -- 0.10130379667644344
	pesos_i(14711) := b"0000000000000000_0000000000000000_0001000001101011_0001111110010001"; -- 0.06413457187125365
	pesos_i(14712) := b"1111111111111111_1111111111111111_1111111000011001_0010011011110010"; -- -0.007428708980645728
	pesos_i(14713) := b"1111111111111111_1111111111111111_1110000010100011_1011011011010101"; -- -0.12250191967249802
	pesos_i(14714) := b"0000000000000000_0000000000000000_0000000101001100_0000100100100000"; -- 0.0050664619401936525
	pesos_i(14715) := b"0000000000000000_0000000000000000_0000101000111010_0110011100010100"; -- 0.039953653678542554
	pesos_i(14716) := b"1111111111111111_1111111111111111_1111100000100101_0100011100000100"; -- -0.030681191950943553
	pesos_i(14717) := b"0000000000000000_0000000000000000_0001010001101110_0010100100010001"; -- 0.07980591445063853
	pesos_i(14718) := b"0000000000000000_0000000000000000_0000110000001010_0001001100110011"; -- 0.0470287322831645
	pesos_i(14719) := b"1111111111111111_1111111111111111_1101111101100010_0100111110001001"; -- -0.12740614809224352
	pesos_i(14720) := b"1111111111111111_1111111111111111_1111100001100000_1001000000100100"; -- -0.029776564832011423
	pesos_i(14721) := b"1111111111111111_1111111111111111_1111000110011110_0011110100000101"; -- -0.0561792242405117
	pesos_i(14722) := b"1111111111111111_1111111111111111_1110000100000010_1111100100100000"; -- -0.12104838352871271
	pesos_i(14723) := b"1111111111111111_1111111111111111_1111101011101010_1001010100111010"; -- -0.019858048878424555
	pesos_i(14724) := b"0000000000000000_0000000000000000_0001010100011001_0110010001111001"; -- 0.08241870825051127
	pesos_i(14725) := b"1111111111111111_1111111111111111_1110101111011111_0000111111101101"; -- -0.07862759073065122
	pesos_i(14726) := b"1111111111111111_1111111111111111_1111000010001010_0001001001110001"; -- -0.060393187813610624
	pesos_i(14727) := b"0000000000000000_0000000000000000_0001110110001111_1101000011000111"; -- 0.1154757009774149
	pesos_i(14728) := b"0000000000000000_0000000000000000_0001010011100111_1001010001100010"; -- 0.08165862465916608
	pesos_i(14729) := b"1111111111111111_1111111111111111_1110010000010111_1001000110000101"; -- -0.10901537412733507
	pesos_i(14730) := b"1111111111111111_1111111111111111_1101011101111000_0110100110011101"; -- -0.15831890018842704
	pesos_i(14731) := b"0000000000000000_0000000000000000_0000000001001100_0001100011001011"; -- 0.0011611457545128271
	pesos_i(14732) := b"0000000000000000_0000000000000000_0001001101111100_1010100010011101"; -- 0.07612088993063465
	pesos_i(14733) := b"0000000000000000_0000000000000000_0000010001000100_0000100010001101"; -- 0.01666310723787583
	pesos_i(14734) := b"0000000000000000_0000000000000000_0000101100111110_1010010111101111"; -- 0.04392468533867235
	pesos_i(14735) := b"0000000000000000_0000000000000000_0000101110101110_0101110001010110"; -- 0.04562928301123146
	pesos_i(14736) := b"0000000000000000_0000000000000000_0000011001001100_0010001010000000"; -- 0.02459922436211324
	pesos_i(14737) := b"1111111111111111_1111111111111111_1111000000010100_0000111110011101"; -- -0.06219389359996707
	pesos_i(14738) := b"1111111111111111_1111111111111111_1101101010101110_1010011100100011"; -- -0.14577250853935808
	pesos_i(14739) := b"1111111111111111_1111111111111111_1110110000100110_1011101011000000"; -- -0.07753403482360326
	pesos_i(14740) := b"0000000000000000_0000000000000000_0000010011001100_0010001011011100"; -- 0.018739870824183085
	pesos_i(14741) := b"1111111111111111_1111111111111111_1101111011000100_1011110101011101"; -- -0.1298104903424819
	pesos_i(14742) := b"1111111111111111_1111111111111111_1110010110001110_0011000111011101"; -- -0.10329902976265128
	pesos_i(14743) := b"0000000000000000_0000000000000000_0001100100000011_0001001111111100"; -- 0.0977032175761114
	pesos_i(14744) := b"0000000000000000_0000000000000000_0010001100010110_1010011010111000"; -- 0.13706438062225265
	pesos_i(14745) := b"0000000000000000_0000000000000000_0000110011101000_1110100001111000"; -- 0.0504288952412719
	pesos_i(14746) := b"0000000000000000_0000000000000000_0001000010011110_1101011001001011"; -- 0.0649236614815467
	pesos_i(14747) := b"0000000000000000_0000000000000000_0000110110000011_1101011100100110"; -- 0.05279297530539395
	pesos_i(14748) := b"1111111111111111_1111111111111111_1111111001101001_1111001010110110"; -- -0.006195860562696662
	pesos_i(14749) := b"0000000000000000_0000000000000000_0010001010011101_1101000110110001"; -- 0.1352206285366296
	pesos_i(14750) := b"1111111111111111_1111111111111111_1111101110001011_0000010101000001"; -- -0.0174099652773019
	pesos_i(14751) := b"0000000000000000_0000000000000000_0001101100011000_0010111100100110"; -- 0.10583777114617002
	pesos_i(14752) := b"1111111111111111_1111111111111111_1111101000100001_0100010001010111"; -- -0.022929886488418174
	pesos_i(14753) := b"1111111111111111_1111111111111111_1110100100010101_0110110101100100"; -- -0.0895167952103466
	pesos_i(14754) := b"0000000000000000_0000000000000000_0001001101010101_1110111111010001"; -- 0.07553004116843125
	pesos_i(14755) := b"1111111111111111_1111111111111111_1101110010000001_0100101010111100"; -- -0.1386521616231669
	pesos_i(14756) := b"0000000000000000_0000000000000000_0000111001011100_1001101001001001"; -- 0.05610050468494577
	pesos_i(14757) := b"1111111111111111_1111111111111111_1110010001000010_0001101110000001"; -- -0.10836628064639907
	pesos_i(14758) := b"0000000000000000_0000000000000000_0001101111011010_1110100011101011"; -- 0.1088090489207355
	pesos_i(14759) := b"0000000000000000_0000000000000000_0001100010100011_0000110010000010"; -- 0.09623792803614285
	pesos_i(14760) := b"1111111111111111_1111111111111111_1111010000011000_0100100010110111"; -- -0.046504454935602596
	pesos_i(14761) := b"0000000000000000_0000000000000000_0010001111000101_1001001010110001"; -- 0.1397334749962222
	pesos_i(14762) := b"1111111111111111_1111111111111111_1111001010000000_0100111110001011"; -- -0.052729633817263116
	pesos_i(14763) := b"0000000000000000_0000000000000000_0000111001111010_1110100100010010"; -- 0.05656296426834519
	pesos_i(14764) := b"0000000000000000_0000000000000000_0001001100011111_0100000010011000"; -- 0.07469562259070296
	pesos_i(14765) := b"1111111111111111_1111111111111111_1111011000011001_1110000110111111"; -- -0.03866757483492167
	pesos_i(14766) := b"1111111111111111_1111111111111111_1101111110010110_0001101011111001"; -- -0.12661582390909257
	pesos_i(14767) := b"1111111111111111_1111111111111111_1111001010110100_1011001001011111"; -- -0.051930286200753864
	pesos_i(14768) := b"1111111111111111_1111111111111111_1110100101010001_1011100001000011"; -- -0.08859680520179342
	pesos_i(14769) := b"0000000000000000_0000000000000000_0001010010100110_0100110011110010"; -- 0.08066254522933353
	pesos_i(14770) := b"1111111111111111_1111111111111111_1110100101100100_1001001010001000"; -- -0.08830913704269512
	pesos_i(14771) := b"1111111111111111_1111111111111111_1101101110010011_0010000111101110"; -- -0.14228618568958845
	pesos_i(14772) := b"1111111111111111_1111111111111111_1111111110010110_0111011011111011"; -- -0.0016103397404795266
	pesos_i(14773) := b"0000000000000000_0000000000000000_0001001110101010_1010001000011101"; -- 0.07682240681189481
	pesos_i(14774) := b"0000000000000000_0000000000000000_0000100101100010_0101101111010111"; -- 0.0366570854164382
	pesos_i(14775) := b"0000000000000000_0000000000000000_0001000011000110_0110010010110001"; -- 0.06552724183709564
	pesos_i(14776) := b"0000000000000000_0000000000000000_0001110101100101_1110100011111010"; -- 0.11483627409601437
	pesos_i(14777) := b"1111111111111111_1111111111111111_1110010001101100_0011001111001100"; -- -0.10772396335335621
	pesos_i(14778) := b"0000000000000000_0000000000000000_0001001101111110_1010101111101001"; -- 0.07615160398282764
	pesos_i(14779) := b"0000000000000000_0000000000000000_0001001110110111_1011010110010110"; -- 0.07702193171734005
	pesos_i(14780) := b"1111111111111111_1111111111111111_1111010011010001_0011110100000010"; -- -0.043682276742680486
	pesos_i(14781) := b"0000000000000000_0000000000000000_0000011100101101_1100110101010001"; -- 0.02804263334255601
	pesos_i(14782) := b"0000000000000000_0000000000000000_0000110101111010_0011011010100100"; -- 0.05264607909835352
	pesos_i(14783) := b"0000000000000000_0000000000000000_0000101101110111_0110000101010011"; -- 0.04479034696698352
	pesos_i(14784) := b"1111111111111111_1111111111111111_1110100010000100_0101100001011001"; -- -0.09173057395783087
	pesos_i(14785) := b"1111111111111111_1111111111111111_1111011000110001_1010101011100110"; -- -0.03830463301492663
	pesos_i(14786) := b"1111111111111111_1111111111111111_1110011111111010_0111011100010011"; -- -0.09383445542688555
	pesos_i(14787) := b"1111111111111111_1111111111111111_1110111000001000_0010010011111010"; -- -0.07018822570444161
	pesos_i(14788) := b"1111111111111111_1111111111111111_1111010101110100_1011010001011100"; -- -0.04118798017661733
	pesos_i(14789) := b"0000000000000000_0000000000000000_0010001000010101_0100010101100110"; -- 0.13313707111391518
	pesos_i(14790) := b"0000000000000000_0000000000000000_0000001100110011_1111000110000111"; -- 0.012511344478762166
	pesos_i(14791) := b"1111111111111111_1111111111111111_1110100001110101_0110011000101110"; -- -0.09195863120111408
	pesos_i(14792) := b"1111111111111111_1111111111111111_1110111011101010_0111111011011110"; -- -0.06673438151658564
	pesos_i(14793) := b"0000000000000000_0000000000000000_0000110000001110_1111011010010001"; -- 0.04710331953930816
	pesos_i(14794) := b"1111111111111111_1111111111111111_1110111011111110_0101111110110001"; -- -0.06643106395979656
	pesos_i(14795) := b"0000000000000000_0000000000000000_0001000000110010_1001110000100010"; -- 0.06327224558792877
	pesos_i(14796) := b"0000000000000000_0000000000000000_0010001011010110_1000010000111110"; -- 0.13608576316013857
	pesos_i(14797) := b"1111111111111111_1111111111111111_1101101010010011_1000101000110010"; -- -0.1461862209703997
	pesos_i(14798) := b"1111111111111111_1111111111111111_1101100101001111_0001101100100000"; -- -0.15113668894833923
	pesos_i(14799) := b"1111111111111111_1111111111111111_1101110110110010_1111100110001010"; -- -0.13398781176651256
	pesos_i(14800) := b"0000000000000000_0000000000000000_0000011100000110_0001101000100000"; -- 0.02743685994548539
	pesos_i(14801) := b"1111111111111111_1111111111111111_1111100111011010_0101010001100011"; -- -0.024012304064566104
	pesos_i(14802) := b"0000000000000000_0000000000000000_0000000011010001_0101101001010110"; -- 0.003194471349533364
	pesos_i(14803) := b"1111111111111111_1111111111111111_1111010111011101_0111011001001000"; -- -0.03958950753239567
	pesos_i(14804) := b"1111111111111111_1111111111111111_1110001001100111_1001001000000101"; -- -0.11560714123553154
	pesos_i(14805) := b"0000000000000000_0000000000000000_0001111000010011_0010100110111111"; -- 0.1174799052251677
	pesos_i(14806) := b"0000000000000000_0000000000000000_0001010000100000_1000101000010111"; -- 0.07862151204450259
	pesos_i(14807) := b"1111111111111111_1111111111111111_1110111011010111_0001010111110010"; -- -0.06703055226810674
	pesos_i(14808) := b"1111111111111111_1111111111111111_1110101000110001_0100100001101010"; -- -0.08518550301830397
	pesos_i(14809) := b"1111111111111111_1111111111111111_1111101010001010_1110001011011000"; -- -0.021318266216059468
	pesos_i(14810) := b"0000000000000000_0000000000000000_0000111011110010_0101010111100101"; -- 0.058385246667516925
	pesos_i(14811) := b"1111111111111111_1111111111111111_1101110010011000_0110011101100110"; -- -0.13829950104646418
	pesos_i(14812) := b"1111111111111111_1111111111111111_1110010110100110_1001111011000001"; -- -0.10292632848021087
	pesos_i(14813) := b"0000000000000000_0000000000000000_0001110000111011_0101101100101010"; -- 0.11028070241302992
	pesos_i(14814) := b"1111111111111111_1111111111111111_1101011101100101_0101001110011111"; -- -0.15861012806177974
	pesos_i(14815) := b"1111111111111111_1111111111111111_1110111100001001_1100100001001001"; -- -0.06625698292602486
	pesos_i(14816) := b"1111111111111111_1111111111111111_1111010111100100_1010010000110111"; -- -0.03947995823254318
	pesos_i(14817) := b"1111111111111111_1111111111111111_1111100110000100_1101100001011100"; -- -0.025316693722607104
	pesos_i(14818) := b"1111111111111111_1111111111111111_1101110011010000_1101000011100011"; -- -0.13743872120383624
	pesos_i(14819) := b"0000000000000000_0000000000000000_0000110101101110_0011010000100010"; -- 0.05246282423188259
	pesos_i(14820) := b"0000000000000000_0000000000000000_0010000101101001_0101111100100011"; -- 0.130514093373984
	pesos_i(14821) := b"0000000000000000_0000000000000000_0010100000010000_0100110001111110"; -- 0.15649869984773848
	pesos_i(14822) := b"0000000000000000_0000000000000000_0000011101000000_0000111111001011"; -- 0.028321253784300095
	pesos_i(14823) := b"1111111111111111_1111111111111111_1101101101000100_1110001011001010"; -- -0.14348013466948456
	pesos_i(14824) := b"0000000000000000_0000000000000000_0001001000101011_0010101101011001"; -- 0.07097121174336984
	pesos_i(14825) := b"1111111111111111_1111111111111111_1110011101011101_1101010000100110"; -- -0.09622453753970563
	pesos_i(14826) := b"0000000000000000_0000000000000000_0000000111110010_1101100010111111"; -- 0.007611796079586448
	pesos_i(14827) := b"0000000000000000_0000000000000000_0001010010100010_1110001001101100"; -- 0.08061041959760429
	pesos_i(14828) := b"0000000000000000_0000000000000000_0000010000100100_0001011100011000"; -- 0.016175692808545715
	pesos_i(14829) := b"0000000000000000_0000000000000000_0000011010100110_0100001000010110"; -- 0.025974398030522733
	pesos_i(14830) := b"1111111111111111_1111111111111111_1110000000010001_1111100001001111"; -- -0.12472580016531488
	pesos_i(14831) := b"1111111111111111_1111111111111111_1110100111011000_0011001110100000"; -- -0.08654477457865485
	pesos_i(14832) := b"1111111111111111_1111111111111111_1110001000001100_1010001011000001"; -- -0.11699469356142324
	pesos_i(14833) := b"0000000000000000_0000000000000000_0010001111101001_1100010110001110"; -- 0.14028582310547238
	pesos_i(14834) := b"1111111111111111_1111111111111111_1110110000010011_1111010001111100"; -- -0.07782051068080255
	pesos_i(14835) := b"1111111111111111_1111111111111111_1111000110100100_1011000010001101"; -- -0.056080785388965784
	pesos_i(14836) := b"0000000000000000_0000000000000000_0001011110100011_1111001000001001"; -- 0.09234535898087236
	pesos_i(14837) := b"1111111111111111_1111111111111111_1111111001100100_1000110110011110"; -- -0.006278180038319767
	pesos_i(14838) := b"1111111111111111_1111111111111111_1111110110100010_1010000000001111"; -- -0.009237286002708796
	pesos_i(14839) := b"1111111111111111_1111111111111111_1111010010010110_0111010010001010"; -- -0.044579235393156356
	pesos_i(14840) := b"1111111111111111_1111111111111111_1111010011110110_0111010000010001"; -- -0.043114419720575343
	pesos_i(14841) := b"0000000000000000_0000000000000000_0010010011000011_0010101010101011"; -- 0.14360300709481336
	pesos_i(14842) := b"0000000000000000_0000000000000000_0010001001101110_0110001111011111"; -- 0.13449691963980906
	pesos_i(14843) := b"1111111111111111_1111111111111111_1110010101110011_0011100100011001"; -- -0.103710585942551
	pesos_i(14844) := b"1111111111111111_1111111111111111_1110001110110100_0001000000011101"; -- -0.11053370753878772
	pesos_i(14845) := b"1111111111111111_1111111111111111_1111000111100000_0011011100010011"; -- -0.055172498625933944
	pesos_i(14846) := b"1111111111111111_1111111111111111_1101111111110100_0111111100111011"; -- -0.1251755220343689
	pesos_i(14847) := b"1111111111111111_1111111111111111_1110010010000000_1110110110100010"; -- -0.10740771098922902
	pesos_i(14848) := b"1111111111111111_1111111111111111_1111001111000101_1010000010110011"; -- -0.04776569023075203
	pesos_i(14849) := b"1111111111111111_1111111111111111_1111101100011010_0101000000011101"; -- -0.019129746268110457
	pesos_i(14850) := b"1111111111111111_1111111111111111_1111111110101100_1000100101011101"; -- -0.0012735508952002735
	pesos_i(14851) := b"0000000000000000_0000000000000000_0001110000110111_1111010101011000"; -- 0.11022885711555258
	pesos_i(14852) := b"1111111111111111_1111111111111111_1110001001111010_0001100111101011"; -- -0.11532438285545543
	pesos_i(14853) := b"0000000000000000_0000000000000000_0001100011111001_1011000000101100"; -- 0.09755993902618533
	pesos_i(14854) := b"0000000000000000_0000000000000000_0000100100110001_1101110111011100"; -- 0.035917154467709766
	pesos_i(14855) := b"1111111111111111_1111111111111111_1111000110110101_0100010111111010"; -- -0.05582773825807941
	pesos_i(14856) := b"0000000000000000_0000000000000000_0001011110101100_0011110101001010"; -- 0.09247191474647314
	pesos_i(14857) := b"0000000000000000_0000000000000000_0001001101100000_1100011000001100"; -- 0.0756953983744821
	pesos_i(14858) := b"1111111111111111_1111111111111111_1110000110110011_1110101110001100"; -- -0.11834838710353962
	pesos_i(14859) := b"0000000000000000_0000000000000000_0001000010000110_1100010100010011"; -- 0.06455642416178052
	pesos_i(14860) := b"0000000000000000_0000000000000000_0001000010110001_1010010000010100"; -- 0.06521058543148604
	pesos_i(14861) := b"1111111111111111_1111111111111111_1110011011111111_0011011010111111"; -- -0.09766824568710082
	pesos_i(14862) := b"1111111111111111_1111111111111111_1111010010010100_1010010010001100"; -- -0.0446068915477749
	pesos_i(14863) := b"0000000000000000_0000000000000000_0000100001110001_0000100111100111"; -- 0.03297483336157174
	pesos_i(14864) := b"1111111111111111_1111111111111111_1111101110010111_0111011100100001"; -- -0.017220072254297523
	pesos_i(14865) := b"1111111111111111_1111111111111111_1111011001010001_1101111101000110"; -- -0.03781322998780189
	pesos_i(14866) := b"1111111111111111_1111111111111111_1110001110010000_1110101110011011"; -- -0.11106994109043133
	pesos_i(14867) := b"0000000000000000_0000000000000000_0000100010111010_0100010011100111"; -- 0.03409224159539192
	pesos_i(14868) := b"0000000000000000_0000000000000000_0001011111000110_1011101001101011"; -- 0.0928761016767581
	pesos_i(14869) := b"1111111111111111_1111111111111111_1111001111101010_1010110001000000"; -- -0.04720042637736298
	pesos_i(14870) := b"1111111111111111_1111111111111111_1111001101110011_1010100101001101"; -- -0.04901639820011789
	pesos_i(14871) := b"0000000000000000_0000000000000000_0001001010101000_0001011001011110"; -- 0.07287730985508865
	pesos_i(14872) := b"1111111111111111_1111111111111111_1110101011110110_1111100100110000"; -- -0.08216898510384582
	pesos_i(14873) := b"1111111111111111_1111111111111111_1110111101100100_0110001111100111"; -- -0.06487441645085891
	pesos_i(14874) := b"0000000000000000_0000000000000000_0000110111000110_0101010011011001"; -- 0.05380754758608703
	pesos_i(14875) := b"0000000000000000_0000000000000000_0001100010110001_0001110101001101"; -- 0.09645255203891263
	pesos_i(14876) := b"1111111111111111_1111111111111111_1101011000101110_0000111010110010"; -- -0.16335971968301072
	pesos_i(14877) := b"1111111111111111_1111111111111111_1110101010001100_0101110101110101"; -- -0.08379569912769197
	pesos_i(14878) := b"0000000000000000_0000000000000000_0001011110011010_0010001100000100"; -- 0.092195690566124
	pesos_i(14879) := b"0000000000000000_0000000000000000_0001111010000111_1100011101110011"; -- 0.11925932460718261
	pesos_i(14880) := b"1111111111111111_1111111111111111_1110110110011011_1010100100011000"; -- -0.07184355884678778
	pesos_i(14881) := b"1111111111111111_1111111111111111_1110000101110000_0101111101000110"; -- -0.1193790868349204
	pesos_i(14882) := b"0000000000000000_0000000000000000_0001111101011000_1110000000010110"; -- 0.12244988004500199
	pesos_i(14883) := b"1111111111111111_1111111111111111_1110111011010110_0101000011001111"; -- -0.06704230267662716
	pesos_i(14884) := b"1111111111111111_1111111111111111_1111010110001110_0100011101000011"; -- -0.04079775442671467
	pesos_i(14885) := b"1111111111111111_1111111111111111_1111101010010000_0001101110110001"; -- -0.021238583763509022
	pesos_i(14886) := b"1111111111111111_1111111111111111_1111000001010010_1100010001000111"; -- -0.06123708015925426
	pesos_i(14887) := b"0000000000000000_0000000000000000_0001110010011001_0111010110100111"; -- 0.11171660723946591
	pesos_i(14888) := b"1111111111111111_1111111111111111_1111000111110001_0110110001001100"; -- -0.05490992695013552
	pesos_i(14889) := b"1111111111111111_1111111111111111_1110010001100001_0110111001010001"; -- -0.10788832212333772
	pesos_i(14890) := b"0000000000000000_0000000000000000_0000110110110010_0110010101110000"; -- 0.053503360493869404
	pesos_i(14891) := b"0000000000000000_0000000000000000_0001100110110101_0110101010111000"; -- 0.10042445186178553
	pesos_i(14892) := b"1111111111111111_1111111111111111_1111111000110001_1111111100000111"; -- -0.007049618555251885
	pesos_i(14893) := b"0000000000000000_0000000000000000_0001101101110011_1010010110001000"; -- 0.10723337715587322
	pesos_i(14894) := b"1111111111111111_1111111111111111_1110001111011110_0101001001100011"; -- -0.10988888813636288
	pesos_i(14895) := b"0000000000000000_0000000000000000_0001111011000011_1111111101001101"; -- 0.12017818091785352
	pesos_i(14896) := b"1111111111111111_1111111111111111_1110100010111000_0000110011011110"; -- -0.09094161579005729
	pesos_i(14897) := b"0000000000000000_0000000000000000_0000010000111010_1100100000101101"; -- 0.01652194124116497
	pesos_i(14898) := b"0000000000000000_0000000000000000_0010001101101000_1001111010111110"; -- 0.13831512593951645
	pesos_i(14899) := b"0000000000000000_0000000000000000_0010001100010110_1101001100011101"; -- 0.1370670267376732
	pesos_i(14900) := b"0000000000000000_0000000000000000_0001001001110010_1101100100110001"; -- 0.07206494760149872
	pesos_i(14901) := b"0000000000000000_0000000000000000_0001001011111011_1101110010100110"; -- 0.07415560761977039
	pesos_i(14902) := b"1111111111111111_1111111111111111_1110010100010011_0100000011001100"; -- -0.10517497071674861
	pesos_i(14903) := b"1111111111111111_1111111111111111_1111111011111010_0000100000000111"; -- -0.003997324245234295
	pesos_i(14904) := b"1111111111111111_1111111111111111_1101111111000010_0011101010010011"; -- -0.1259425537058004
	pesos_i(14905) := b"0000000000000000_0000000000000000_0000001100111100_1010100011100011"; -- 0.012644343878212339
	pesos_i(14906) := b"0000000000000000_0000000000000000_0001000001100111_1000110001001110"; -- 0.06408001811838494
	pesos_i(14907) := b"1111111111111111_1111111111111111_1111101111000001_1011110100000010"; -- -0.01657503797587356
	pesos_i(14908) := b"1111111111111111_1111111111111111_1101110100100000_1001111111111100"; -- -0.13622093303977936
	pesos_i(14909) := b"0000000000000000_0000000000000000_0001011111000100_1111100111011010"; -- 0.09284936487455758
	pesos_i(14910) := b"0000000000000000_0000000000000000_0000111101011011_1100000110101111"; -- 0.059993844344664635
	pesos_i(14911) := b"1111111111111111_1111111111111111_1110101110010011_1111100111011110"; -- -0.07977331471824062
	pesos_i(14912) := b"0000000000000000_0000000000000000_0000001101001001_0110100001111011"; -- 0.012838869058503035
	pesos_i(14913) := b"1111111111111111_1111111111111111_1111010011110000_0101010010011101"; -- -0.04320784720764908
	pesos_i(14914) := b"1111111111111111_1111111111111111_1101110010011000_1100000110111110"; -- -0.13829411609744136
	pesos_i(14915) := b"0000000000000000_0000000000000000_0001100111111000_1011101011011000"; -- 0.1014515664035038
	pesos_i(14916) := b"0000000000000000_0000000000000000_0001000000111101_0100010110101011"; -- 0.06343493877066544
	pesos_i(14917) := b"0000000000000000_0000000000000000_0010001111010111_1011101000011000"; -- 0.14001048174066874
	pesos_i(14918) := b"0000000000000000_0000000000000000_0000110010111001_1111111101001010"; -- 0.049713092422032354
	pesos_i(14919) := b"0000000000000000_0000000000000000_0001001110111100_1101000001000000"; -- 0.07709981509102339
	pesos_i(14920) := b"0000000000000000_0000000000000000_0010010101000110_1000010101011011"; -- 0.14560731373442826
	pesos_i(14921) := b"1111111111111111_1111111111111111_1110101101001000_0100001111111000"; -- -0.08092856600583943
	pesos_i(14922) := b"0000000000000000_0000000000000000_0001001011001010_0101000111110001"; -- 0.07339965951224182
	pesos_i(14923) := b"1111111111111111_1111111111111111_1111010011010110_1100011010100111"; -- -0.043597778556615334
	pesos_i(14924) := b"0000000000000000_0000000000000000_0000101100011111_0101001101001010"; -- 0.04344673686140296
	pesos_i(14925) := b"1111111111111111_1111111111111111_1110001101010100_0001101111011000"; -- -0.11199785210713883
	pesos_i(14926) := b"1111111111111111_1111111111111111_1111001001010101_1011110100110001"; -- -0.053379226169674124
	pesos_i(14927) := b"1111111111111111_1111111111111111_1111011001011011_1111000110111110"; -- -0.03765954112508133
	pesos_i(14928) := b"1111111111111111_1111111111111111_1101111011001000_0011011011000110"; -- -0.1297574774103737
	pesos_i(14929) := b"1111111111111111_1111111111111111_1101111011001011_0001111101010101"; -- -0.129713098281852
	pesos_i(14930) := b"1111111111111111_1111111111111111_1111000111011011_1111101111010001"; -- -0.05523706585675522
	pesos_i(14931) := b"1111111111111111_1111111111111111_1111111110010101_1111101010101101"; -- -0.0016177490244349934
	pesos_i(14932) := b"0000000000000000_0000000000000000_0000100000011001_1001101111011100"; -- 0.031640759671605276
	pesos_i(14933) := b"0000000000000000_0000000000000000_0001110100110100_0001011001100001"; -- 0.11407604100179192
	pesos_i(14934) := b"1111111111111111_1111111111111111_1110011101011000_1000111010010100"; -- -0.09630497829071791
	pesos_i(14935) := b"0000000000000000_0000000000000000_0001100100000001_0010001110011010"; -- 0.09767363079162635
	pesos_i(14936) := b"1111111111111111_1111111111111111_1111100111000110_0110101010110000"; -- -0.024316150712473786
	pesos_i(14937) := b"0000000000000000_0000000000000000_0000011000101100_0111100010111011"; -- 0.024116082720957346
	pesos_i(14938) := b"0000000000000000_0000000000000000_0000000000100110_1100001100000001"; -- 0.0005914571645369686
	pesos_i(14939) := b"0000000000000000_0000000000000000_0010000101111110_0011100111101110"; -- 0.13083231028097583
	pesos_i(14940) := b"1111111111111111_1111111111111111_1110001001110011_0000110010001010"; -- -0.11543199197312905
	pesos_i(14941) := b"1111111111111111_1111111111111111_1111011011110010_0001000111000100"; -- -0.03536881422714226
	pesos_i(14942) := b"1111111111111111_1111111111111111_1110100001011010_1011010011000110"; -- -0.09236593415769992
	pesos_i(14943) := b"1111111111111111_1111111111111111_1110111000000100_0010001000110000"; -- -0.07024942711893403
	pesos_i(14944) := b"1111111111111111_1111111111111111_1111110100011101_0100011011011101"; -- -0.011272021246555464
	pesos_i(14945) := b"0000000000000000_0000000000000000_0001100100101101_0000010110011111"; -- 0.09834323052960148
	pesos_i(14946) := b"1111111111111111_1111111111111111_1101111000101100_1100101101101001"; -- -0.13212898919476193
	pesos_i(14947) := b"0000000000000000_0000000000000000_0001101111100101_1100011101011110"; -- 0.10897489580653323
	pesos_i(14948) := b"1111111111111111_1111111111111111_1111110010111000_0011100111001111"; -- -0.012813937200518918
	pesos_i(14949) := b"0000000000000000_0000000000000000_0000010110010010_1110100111000101"; -- 0.021772967045137523
	pesos_i(14950) := b"1111111111111111_1111111111111111_1110011010001001_0000011100000011"; -- -0.09947162799994948
	pesos_i(14951) := b"0000000000000000_0000000000000000_0000001000011100_0101010001101001"; -- 0.008244777258188703
	pesos_i(14952) := b"0000000000000000_0000000000000000_0001111110111000_1001000011100101"; -- 0.12391000365607122
	pesos_i(14953) := b"0000000000000000_0000000000000000_0000010011110010_1000001000110110"; -- 0.01932538804475522
	pesos_i(14954) := b"1111111111111111_1111111111111111_1110100111101101_1110100101010000"; -- -0.08621351051015229
	pesos_i(14955) := b"0000000000000000_0000000000000000_0001100111001111_1011101111011100"; -- 0.1008260165383107
	pesos_i(14956) := b"1111111111111111_1111111111111111_1111100011101010_1011010010100000"; -- -0.02766867725773046
	pesos_i(14957) := b"0000000000000000_0000000000000000_0001010110110001_0001110011011011"; -- 0.08473377554675461
	pesos_i(14958) := b"1111111111111111_1111111111111111_1111110110100111_0110010001001110"; -- -0.009164553572635365
	pesos_i(14959) := b"1111111111111111_1111111111111111_1101110100011011_0011010100111101"; -- -0.1363035895090753
	pesos_i(14960) := b"0000000000000000_0000000000000000_0001101010010010_0111100000101011"; -- 0.10379744579266213
	pesos_i(14961) := b"1111111111111111_1111111111111111_1111100110100010_0101011001101100"; -- -0.024866675104530927
	pesos_i(14962) := b"1111111111111111_1111111111111111_1111000010111000_0101000001110000"; -- -0.05968758831192646
	pesos_i(14963) := b"1111111111111111_1111111111111111_1111010010000010_0000110011110010"; -- -0.04489058587434039
	pesos_i(14964) := b"0000000000000000_0000000000000000_0000010100011010_0110000011000001"; -- 0.01993374545752883
	pesos_i(14965) := b"0000000000000000_0000000000000000_0000100100110000_0100011001001000"; -- 0.03589286088900842
	pesos_i(14966) := b"1111111111111111_1111111111111111_1111001101100110_1001100110111100"; -- -0.049215690292271054
	pesos_i(14967) := b"0000000000000000_0000000000000000_0010000101110111_1101010101011011"; -- 0.13073476287955804
	pesos_i(14968) := b"1111111111111111_1111111111111111_1111110000111010_1011010011101110"; -- -0.014729205919686746
	pesos_i(14969) := b"0000000000000000_0000000000000000_0000100000001100_0100101100110000"; -- 0.03143758701484326
	pesos_i(14970) := b"1111111111111111_1111111111111111_1110011111000001_0010101111010110"; -- -0.09470869093059694
	pesos_i(14971) := b"0000000000000000_0000000000000000_0001000010000010_0010110011011001"; -- 0.06448631571859396
	pesos_i(14972) := b"0000000000000000_0000000000000000_0010001000000001_0101011000000100"; -- 0.1328328856198849
	pesos_i(14973) := b"0000000000000000_0000000000000000_0001110000101110_1101111111110110"; -- 0.11009025350544535
	pesos_i(14974) := b"0000000000000000_0000000000000000_0010000101001110_1101111011101001"; -- 0.13010972195202566
	pesos_i(14975) := b"1111111111111111_1111111111111111_1110011101001110_1110100001111100"; -- -0.09645220720175944
	pesos_i(14976) := b"0000000000000000_0000000000000000_0001100111011011_1110001100110110"; -- 0.10101146772877319
	pesos_i(14977) := b"0000000000000000_0000000000000000_0001001100010100_0000010100000011"; -- 0.07452422455336184
	pesos_i(14978) := b"1111111111111111_1111111111111111_1111110110011011_1010110111011110"; -- -0.009343274483713795
	pesos_i(14979) := b"1111111111111111_1111111111111111_1111110011010011_0100100101110110"; -- -0.012401016892556967
	pesos_i(14980) := b"1111111111111111_1111111111111111_1110111000110110_1000111101000101"; -- -0.06947998593449584
	pesos_i(14981) := b"1111111111111111_1111111111111111_1110011110010111_0111100100101111"; -- -0.09534494976146034
	pesos_i(14982) := b"0000000000000000_0000000000000000_0010100101000101_1011101100110001"; -- 0.1612202638241388
	pesos_i(14983) := b"0000000000000000_0000000000000000_0000010010000110_0010101110100111"; -- 0.017672279514410447
	pesos_i(14984) := b"1111111111111111_1111111111111111_1111000100010100_1101110111001111"; -- -0.05827535347875812
	pesos_i(14985) := b"0000000000000000_0000000000000000_0000001100111110_0011101000001110"; -- 0.012668255291982499
	pesos_i(14986) := b"1111111111111111_1111111111111111_1110000101101101_0000001100100001"; -- -0.11943035539247389
	pesos_i(14987) := b"1111111111111111_1111111111111111_1110010110100001_1111101101111110"; -- -0.1029970949553788
	pesos_i(14988) := b"0000000000000000_0000000000000000_0000111010010111_0111010110101011"; -- 0.05699859080123176
	pesos_i(14989) := b"1111111111111111_1111111111111111_1101011101110000_1000110001001000"; -- -0.15843890422296567
	pesos_i(14990) := b"0000000000000000_0000000000000000_0001110001100011_0000000000111000"; -- 0.11088563316887737
	pesos_i(14991) := b"0000000000000000_0000000000000000_0000111010110010_1011111100001111"; -- 0.05741495251599762
	pesos_i(14992) := b"0000000000000000_0000000000000000_0001000101011001_0011100110001111"; -- 0.06776771302252399
	pesos_i(14993) := b"0000000000000000_0000000000000000_0001101110100110_1000111010010011"; -- 0.1080102070978051
	pesos_i(14994) := b"1111111111111111_1111111111111111_1111101110000010_0111110010000111"; -- -0.017540185081419937
	pesos_i(14995) := b"1111111111111111_1111111111111111_1101101110110001_0100110110011001"; -- -0.14182581921939974
	pesos_i(14996) := b"0000000000000000_0000000000000000_0010011101010000_0011001011000101"; -- 0.15356747932482992
	pesos_i(14997) := b"1111111111111111_1111111111111111_1111100001001010_1101001110001010"; -- -0.03010824081603409
	pesos_i(14998) := b"1111111111111111_1111111111111111_1110000101110101_1110110111110101"; -- -0.11929428838310568
	pesos_i(14999) := b"1111111111111111_1111111111111111_1101111010010100_0000001000110000"; -- -0.13055406889795498
	pesos_i(15000) := b"0000000000000000_0000000000000000_0001010011001100_1011010011000100"; -- 0.08124856748981395
	pesos_i(15001) := b"1111111111111111_1111111111111111_1101101100010000_1011001101110010"; -- -0.14427641350379541
	pesos_i(15002) := b"0000000000000000_0000000000000000_0000010101010011_1010110000110101"; -- 0.02080799389296916
	pesos_i(15003) := b"0000000000000000_0000000000000000_0000011100011111_1111000001111001"; -- 0.027831105854971623
	pesos_i(15004) := b"0000000000000000_0000000000000000_0000000000001000_1110101001011110"; -- 0.00013603978675578353
	pesos_i(15005) := b"1111111111111111_1111111111111111_1110000001011110_1011000111110110"; -- -0.12355506654142397
	pesos_i(15006) := b"1111111111111111_1111111111111111_1111100011010010_1111101100011010"; -- -0.028030687530051814
	pesos_i(15007) := b"1111111111111111_1111111111111111_1110100111101100_1100010100001001"; -- -0.08623093154958389
	pesos_i(15008) := b"1111111111111111_1111111111111111_1111011100000110_1110011110011001"; -- -0.0350508928543002
	pesos_i(15009) := b"0000000000000000_0000000000000000_0000110101100101_0001000111101010"; -- 0.05232345557215084
	pesos_i(15010) := b"1111111111111111_1111111111111111_1101110111100110_1000001110100000"; -- -0.13320138307962162
	pesos_i(15011) := b"1111111111111111_1111111111111111_1110001001001101_1000101001011000"; -- -0.11600432727369349
	pesos_i(15012) := b"0000000000000000_0000000000000000_0000001101001010_0001101000100110"; -- 0.012849459065539987
	pesos_i(15013) := b"0000000000000000_0000000000000000_0010100100101100_0011011001000011"; -- 0.16083087105504323
	pesos_i(15014) := b"1111111111111111_1111111111111111_1110011001001110_1100001010110000"; -- -0.10036071009751366
	pesos_i(15015) := b"1111111111111111_1111111111111111_1111000010010111_1110111110010111"; -- -0.06018164228529884
	pesos_i(15016) := b"0000000000000000_0000000000000000_0001101110000100_0010110100111010"; -- 0.10748560584996358
	pesos_i(15017) := b"1111111111111111_1111111111111111_1111000010101110_1001111010111010"; -- -0.0598355099199709
	pesos_i(15018) := b"1111111111111111_1111111111111111_1101111000000100_1011101000000110"; -- -0.13274037689920715
	pesos_i(15019) := b"0000000000000000_0000000000000000_0010000010111110_1010100001110001"; -- 0.12790920971733588
	pesos_i(15020) := b"1111111111111111_1111111111111111_1101011011000110_1001110000100111"; -- -0.1610319524487131
	pesos_i(15021) := b"0000000000000000_0000000000000000_0010001010001111_0101100101110001"; -- 0.134999837953936
	pesos_i(15022) := b"0000000000000000_0000000000000000_0001111100011111_0001000110110110"; -- 0.1215678281179077
	pesos_i(15023) := b"1111111111111111_1111111111111111_1111110010100000_0111010011111011"; -- -0.013176621097261127
	pesos_i(15024) := b"0000000000000000_0000000000000000_0000010001100100_1000101011011011"; -- 0.017159155431678095
	pesos_i(15025) := b"0000000000000000_0000000000000000_0001011100111100_0110000100000110"; -- 0.09076506041052998
	pesos_i(15026) := b"0000000000000000_0000000000000000_0001110010001110_0000000101001001"; -- 0.11154182454568942
	pesos_i(15027) := b"1111111111111111_1111111111111111_1111100101011110_0111110111111010"; -- -0.02590191514010734
	pesos_i(15028) := b"0000000000000000_0000000000000000_0001111110010011_1111100010110011"; -- 0.12335161554211242
	pesos_i(15029) := b"1111111111111111_1111111111111111_1111101011110100_1100100010001111"; -- -0.019702401300969535
	pesos_i(15030) := b"0000000000000000_0000000000000000_0000010111010011_1110101101011010"; -- 0.022764882476247077
	pesos_i(15031) := b"0000000000000000_0000000000000000_0000010011101111_0011110001110000"; -- 0.019275452842692373
	pesos_i(15032) := b"1111111111111111_1111111111111111_1110111111101001_0001000000110010"; -- -0.06284998683625413
	pesos_i(15033) := b"1111111111111111_1111111111111111_1110101000111100_1110101100101110"; -- -0.08500795491404753
	pesos_i(15034) := b"1111111111111111_1111111111111111_1110000001110101_0001111101010000"; -- -0.12321285522283883
	pesos_i(15035) := b"0000000000000000_0000000000000000_0000111101111101_1001011001001110"; -- 0.06051005741065921
	pesos_i(15036) := b"1111111111111111_1111111111111111_1111010101100100_1010101010110110"; -- -0.04143269590046024
	pesos_i(15037) := b"0000000000000000_0000000000000000_0001000010111101_0000110011111011"; -- 0.06538468482776592
	pesos_i(15038) := b"1111111111111111_1111111111111111_1111001011011011_0111011101011011"; -- -0.05133871095450697
	pesos_i(15039) := b"1111111111111111_1111111111111111_1111111100101100_0110110101000110"; -- -0.0032283499968632605
	pesos_i(15040) := b"1111111111111111_1111111111111111_1110011011111001_0010100000010000"; -- -0.09776067366327733
	pesos_i(15041) := b"1111111111111111_1111111111111111_1110101010110011_0010100110101100"; -- -0.08320369300583004
	pesos_i(15042) := b"1111111111111111_1111111111111111_1110100110001010_0010100000111001"; -- -0.08773563974635949
	pesos_i(15043) := b"0000000000000000_0000000000000000_0001100001111111_1101101110111111"; -- 0.09570096403533392
	pesos_i(15044) := b"1111111111111111_1111111111111111_1111010011001001_1001000010010110"; -- -0.0437993654661946
	pesos_i(15045) := b"0000000000000000_0000000000000000_0000100001001110_1010011010111110"; -- 0.03245012416925054
	pesos_i(15046) := b"1111111111111111_1111111111111111_1111100111001110_1010110110110010"; -- -0.024190086436523518
	pesos_i(15047) := b"0000000000000000_0000000000000000_0000110100110011_0110110110100110"; -- 0.05156598375279759
	pesos_i(15048) := b"0000000000000000_0000000000000000_0001000000000100_1111110101010110"; -- 0.06257613526116045
	pesos_i(15049) := b"0000000000000000_0000000000000000_0010000101000100_1111101010100111"; -- 0.1299587876059392
	pesos_i(15050) := b"0000000000000000_0000000000000000_0000111011000000_0001000111111010"; -- 0.057618259066976665
	pesos_i(15051) := b"0000000000000000_0000000000000000_0000110011111011_0101111111110101"; -- 0.05071067546279155
	pesos_i(15052) := b"1111111111111111_1111111111111111_1110111111111100_0000011110000111"; -- -0.06256058653526946
	pesos_i(15053) := b"1111111111111111_1111111111111111_1111011011111000_0110011111010001"; -- -0.03527213232751417
	pesos_i(15054) := b"1111111111111111_1111111111111111_1110010000000110_1101001110010011"; -- -0.10927083655190148
	pesos_i(15055) := b"1111111111111111_1111111111111111_1101011100010010_1010101000111111"; -- -0.15987144427366543
	pesos_i(15056) := b"1111111111111111_1111111111111111_1110111111001110_0101100011010110"; -- -0.06325764444150489
	pesos_i(15057) := b"0000000000000000_0000000000000000_0000101101111000_0100101000101110"; -- 0.04480422611995992
	pesos_i(15058) := b"0000000000000000_0000000000000000_0001000000100101_0100111001010011"; -- 0.06306924358508251
	pesos_i(15059) := b"1111111111111111_1111111111111111_1101100000001010_1001010101111101"; -- -0.1560885019086486
	pesos_i(15060) := b"0000000000000000_0000000000000000_0010001111110010_0111010011111010"; -- 0.1404183492117584
	pesos_i(15061) := b"0000000000000000_0000000000000000_0001001111011010_0010111010111010"; -- 0.07754795121603861
	pesos_i(15062) := b"0000000000000000_0000000000000000_0000101110000001_1011001101010110"; -- 0.044947823044844626
	pesos_i(15063) := b"0000000000000000_0000000000000000_0000010100101011_1110100000010111"; -- 0.020201211534875366
	pesos_i(15064) := b"1111111111111111_1111111111111111_1101110111110001_1111111010001011"; -- -0.13302620990429967
	pesos_i(15065) := b"0000000000000000_0000000000000000_0010000110101011_1100110001001110"; -- 0.13152768050908734
	pesos_i(15066) := b"1111111111111111_1111111111111111_1110000001000010_1110101000111010"; -- -0.12397895894844882
	pesos_i(15067) := b"1111111111111111_1111111111111111_1110011110011001_1010111101011111"; -- -0.095311202230857
	pesos_i(15068) := b"1111111111111111_1111111111111111_1111110100011011_1001010000100011"; -- -0.011297932959729143
	pesos_i(15069) := b"1111111111111111_1111111111111111_1111000101011111_0111111101100100"; -- -0.05713657189893108
	pesos_i(15070) := b"1111111111111111_1111111111111111_1111011001101001_1110101111100110"; -- -0.03744626640844234
	pesos_i(15071) := b"0000000000000000_0000000000000000_0000101111100110_0101000100010000"; -- 0.04648310325379121
	pesos_i(15072) := b"0000000000000000_0000000000000000_0001001001001110_0001010011111111"; -- 0.07150393709236137
	pesos_i(15073) := b"1111111111111111_1111111111111111_1110100100011010_1000101100000000"; -- -0.08943873653759647
	pesos_i(15074) := b"0000000000000000_0000000000000000_0000001001000000_1011100110111010"; -- 0.008800132767980046
	pesos_i(15075) := b"0000000000000000_0000000000000000_0000101100001001_1100110011100001"; -- 0.04311829079165264
	pesos_i(15076) := b"1111111111111111_1111111111111111_1111011001100000_1100010011010111"; -- -0.03758592362128145
	pesos_i(15077) := b"1111111111111111_1111111111111111_1111011110111101_0010110110010011"; -- -0.03226962237257056
	pesos_i(15078) := b"1111111111111111_1111111111111111_1101111001100001_1001000100100101"; -- -0.13132374625534735
	pesos_i(15079) := b"1111111111111111_1111111111111111_1111011011111010_0001001100100101"; -- -0.035246661587651315
	pesos_i(15080) := b"1111111111111111_1111111111111111_1110000001100111_1111010110010111"; -- -0.12341370642842608
	pesos_i(15081) := b"1111111111111111_1111111111111111_1110011111110001_0011101100010010"; -- -0.0939753609892308
	pesos_i(15082) := b"1111111111111111_1111111111111111_1111110001100100_1110010101010110"; -- -0.014085451565773519
	pesos_i(15083) := b"0000000000000000_0000000000000000_0010010001100100_0111001000111111"; -- 0.14215768839292342
	pesos_i(15084) := b"1111111111111111_1111111111111111_1111001101011001_0000101111110001"; -- -0.049422506046344655
	pesos_i(15085) := b"1111111111111111_1111111111111111_1111011111011000_0000110011011110"; -- -0.03185958464538683
	pesos_i(15086) := b"1111111111111111_1111111111111111_1110011000010101_0000101001010000"; -- -0.10124145078478591
	pesos_i(15087) := b"0000000000000000_0000000000000000_0000111010010011_0110111101110101"; -- 0.056937185233958736
	pesos_i(15088) := b"0000000000000000_0000000000000000_0000011001110000_0101110000100101"; -- 0.02515197669050326
	pesos_i(15089) := b"1111111111111111_1111111111111111_1111001110010100_1110111101111111"; -- -0.04850867403309175
	pesos_i(15090) := b"0000000000000000_0000000000000000_0010010111110000_1001111011000010"; -- 0.14820282196487394
	pesos_i(15091) := b"1111111111111111_1111111111111111_1111000000101000_0110000001011000"; -- -0.061883905924781005
	pesos_i(15092) := b"1111111111111111_1111111111111111_1110100100110110_0001111101111110"; -- -0.08901789835209106
	pesos_i(15093) := b"1111111111111111_1111111111111111_1110011011101000_0110100011011101"; -- -0.09801621058026598
	pesos_i(15094) := b"0000000000000000_0000000000000000_0000110101000000_0111001000111110"; -- 0.05176462189656354
	pesos_i(15095) := b"1111111111111111_1111111111111111_1111011100001110_1011100110011011"; -- -0.03493156407859757
	pesos_i(15096) := b"1111111111111111_1111111111111111_1111010110001011_0010101010101110"; -- -0.04084523433656918
	pesos_i(15097) := b"0000000000000000_0000000000000000_0000101000010001_0010101001100000"; -- 0.03932442514359801
	pesos_i(15098) := b"1111111111111111_1111111111111111_1101110001101110_0010100010010000"; -- -0.1389441155943388
	pesos_i(15099) := b"1111111111111111_1111111111111111_1111100111111100_0101101000010010"; -- -0.023493166483722266
	pesos_i(15100) := b"0000000000000000_0000000000000000_0010000110101110_1011001001111001"; -- 0.1315719169816006
	pesos_i(15101) := b"1111111111111111_1111111111111111_1111100110110101_1011000110000100"; -- -0.024571328444703708
	pesos_i(15102) := b"0000000000000000_0000000000000000_0000010010110011_1101100111101100"; -- 0.01836931228295751
	pesos_i(15103) := b"0000000000000000_0000000000000000_0000101010101001_0110101000011111"; -- 0.04164756058878344
	pesos_i(15104) := b"1111111111111111_1111111111111111_1110100011000011_0010001011011011"; -- -0.09077245863160963
	pesos_i(15105) := b"1111111111111111_1111111111111111_1110001111110101_1011100111011110"; -- -0.10953176823934672
	pesos_i(15106) := b"0000000000000000_0000000000000000_0001010110100101_1001011001010011"; -- 0.08455791032486153
	pesos_i(15107) := b"1111111111111111_1111111111111111_1110011001111000_1101101111111001"; -- -0.09971833393209877
	pesos_i(15108) := b"1111111111111111_1111111111111111_1101110100101111_0111100100000110"; -- -0.13599437330413475
	pesos_i(15109) := b"1111111111111111_1111111111111111_1110011010100001_0110011001011101"; -- -0.09909973369000726
	pesos_i(15110) := b"1111111111111111_1111111111111111_1110000111111101_1111101101110110"; -- -0.11721828816352484
	pesos_i(15111) := b"1111111111111111_1111111111111111_1111001011001010_0010011011011100"; -- -0.05160290835780976
	pesos_i(15112) := b"0000000000000000_0000000000000000_0010001100010000_0001100010011001"; -- 0.13696435676334592
	pesos_i(15113) := b"1111111111111111_1111111111111111_1110011110010000_0001110011111110"; -- -0.09545725641490496
	pesos_i(15114) := b"0000000000000000_0000000000000000_0010000001011000_0011011101010010"; -- 0.12634607083402946
	pesos_i(15115) := b"1111111111111111_1111111111111111_1110111000011100_0101110010010010"; -- -0.0698797363473254
	pesos_i(15116) := b"1111111111111111_1111111111111111_1110110110100011_1111101110010100"; -- -0.07171657221616837
	pesos_i(15117) := b"1111111111111111_1111111111111111_1101101011100000_1100001001011100"; -- -0.1450079464991756
	pesos_i(15118) := b"1111111111111111_1111111111111111_1111001000001100_0001000100001100"; -- -0.05450337843241499
	pesos_i(15119) := b"1111111111111111_1111111111111111_1111110110011000_1110110011010101"; -- -0.009385297877983815
	pesos_i(15120) := b"1111111111111111_1111111111111111_1111101101000000_1110100110011111"; -- -0.018540762526331384
	pesos_i(15121) := b"0000000000000000_0000000000000000_0001111010001010_1000001100110100"; -- 0.1193010332384225
	pesos_i(15122) := b"1111111111111111_1111111111111111_1110011101110101_0000011110001000"; -- -0.09587052277664522
	pesos_i(15123) := b"1111111111111111_1111111111111111_1101101101101011_0101100111111000"; -- -0.14289319694865651
	pesos_i(15124) := b"0000000000000000_0000000000000000_0000000011111001_0001011000100100"; -- 0.0038007580741093545
	pesos_i(15125) := b"1111111111111111_1111111111111111_1111110010111100_0010001011000001"; -- -0.01275427618674326
	pesos_i(15126) := b"0000000000000000_0000000000000000_0001110110101001_1100011010000011"; -- 0.11587181746485188
	pesos_i(15127) := b"1111111111111111_1111111111111111_1111100111010001_1111111110000111"; -- -0.02413943248857157
	pesos_i(15128) := b"0000000000000000_0000000000000000_0000000101010100_1101000000001011"; -- 0.005200388714410023
	pesos_i(15129) := b"1111111111111111_1111111111111111_1110011100101111_0011011111001111"; -- -0.0969357605721562
	pesos_i(15130) := b"0000000000000000_0000000000000000_0001101001100110_0101111111010110"; -- 0.10312460881671917
	pesos_i(15131) := b"1111111111111111_1111111111111111_1101100011100110_0011000100111000"; -- -0.15273754492476146
	pesos_i(15132) := b"1111111111111111_1111111111111111_1111101001011000_0000110101000111"; -- -0.022093935172606247
	pesos_i(15133) := b"1111111111111111_1111111111111111_1110000011111110_0100011001000000"; -- -0.1211200802721777
	pesos_i(15134) := b"0000000000000000_0000000000000000_0000001000011011_1100010000011111"; -- 0.008236176923931162
	pesos_i(15135) := b"0000000000000000_0000000000000000_0010011101001001_0110000010011011"; -- 0.15346339984839766
	pesos_i(15136) := b"0000000000000000_0000000000000000_0000111110011000_1111010111101000"; -- 0.06092774305675384
	pesos_i(15137) := b"1111111111111111_1111111111111111_1110011011111101_1100010001101100"; -- -0.09769031881538681
	pesos_i(15138) := b"1111111111111111_1111111111111111_1111110110101100_1100110000100111"; -- -0.009082069889613159
	pesos_i(15139) := b"1111111111111111_1111111111111111_1101100110110000_1100101001010000"; -- -0.14964614433359408
	pesos_i(15140) := b"1111111111111111_1111111111111111_1101110001011100_1101100001111011"; -- -0.13920828807703797
	pesos_i(15141) := b"0000000000000000_0000000000000000_0000100101111101_0111000001011110"; -- 0.0370702961242343
	pesos_i(15142) := b"0000000000000000_0000000000000000_0010010001100110_0101110111110000"; -- 0.14218699555104836
	pesos_i(15143) := b"0000000000000000_0000000000000000_0001111001011010_0110011111000010"; -- 0.1185669754722105
	pesos_i(15144) := b"0000000000000000_0000000000000000_0000001100100100_0100000101011100"; -- 0.012271962171361037
	pesos_i(15145) := b"0000000000000000_0000000000000000_0001000111001101_1101111101101011"; -- 0.06954761840020114
	pesos_i(15146) := b"0000000000000000_0000000000000000_0001101011001100_0000000010000001"; -- 0.10467532290308044
	pesos_i(15147) := b"1111111111111111_1111111111111111_1110000010100000_0011101011101101"; -- -0.12255508146671915
	pesos_i(15148) := b"1111111111111111_1111111111111111_1111000011101001_1110101000110001"; -- -0.058930743294162834
	pesos_i(15149) := b"0000000000000000_0000000000000000_0010001110111111_0100010111000000"; -- 0.1396373360221222
	pesos_i(15150) := b"1111111111111111_1111111111111111_1110100010100111_0100111110100101"; -- -0.09119703507353906
	pesos_i(15151) := b"1111111111111111_1111111111111111_1110000010110010_1101110110001111"; -- -0.1222707295659443
	pesos_i(15152) := b"0000000000000000_0000000000000000_0001101011110001_1100011011101111"; -- 0.10525172560117371
	pesos_i(15153) := b"0000000000000000_0000000000000000_0000010000100000_0101101101110110"; -- 0.01611873266382557
	pesos_i(15154) := b"1111111111111111_1111111111111111_1110111110100000_0000000001000001"; -- -0.06396482857731188
	pesos_i(15155) := b"0000000000000000_0000000000000000_0000001000011010_0110001011000000"; -- 0.008215114472301116
	pesos_i(15156) := b"1111111111111111_1111111111111111_1101100001111010_1110010000111101"; -- -0.15437482360764165
	pesos_i(15157) := b"1111111111111111_1111111111111111_1101101011000001_0000111001000000"; -- -0.1454917042583777
	pesos_i(15158) := b"1111111111111111_1111111111111111_1110001010011010_0111111101110111"; -- -0.11483004909333318
	pesos_i(15159) := b"1111111111111111_1111111111111111_1101110100000001_1111001110011011"; -- -0.1366889710837288
	pesos_i(15160) := b"1111111111111111_1111111111111111_1110100000110110_1100101001111001"; -- -0.09291395700240815
	pesos_i(15161) := b"1111111111111111_1111111111111111_1111001100001110_0110110101100001"; -- -0.050561107509314106
	pesos_i(15162) := b"1111111111111111_1111111111111111_1110100100000101_0001110101000110"; -- -0.08976571118121016
	pesos_i(15163) := b"0000000000000000_0000000000000000_0000000000000000_0011000110000000"; -- 2.9504245683426027e-06
	pesos_i(15164) := b"0000000000000000_0000000000000000_0001010110010100_1111001001010001"; -- 0.08430399391870264
	pesos_i(15165) := b"0000000000000000_0000000000000000_0000000011000100_0001010111100011"; -- 0.002992027249615366
	pesos_i(15166) := b"0000000000000000_0000000000000000_0001111001010000_1101111010001100"; -- 0.11842146785766089
	pesos_i(15167) := b"0000000000000000_0000000000000000_0010001101100100_0110100110000000"; -- 0.13825091713261412
	pesos_i(15168) := b"1111111111111111_1111111111111111_1101110101001100_1100100011000110"; -- -0.13554711503954978
	pesos_i(15169) := b"1111111111111111_1111111111111111_1110001001010000_1110010010010110"; -- -0.11595317206119679
	pesos_i(15170) := b"0000000000000000_0000000000000000_0000011110100110_1110101100101110"; -- 0.029890726751485845
	pesos_i(15171) := b"1111111111111111_1111111111111111_1110101011100101_0001111001110101"; -- -0.08244142184232946
	pesos_i(15172) := b"0000000000000000_0000000000000000_0000100110110001_0101000011000101"; -- 0.03786186985166941
	pesos_i(15173) := b"0000000000000000_0000000000000000_0010000100111100_0011001110010110"; -- 0.12982485211185701
	pesos_i(15174) := b"1111111111111111_1111111111111111_1110010011001111_0001000110111011"; -- -0.10621537373827367
	pesos_i(15175) := b"0000000000000000_0000000000000000_0010001111111111_0110010000000000"; -- 0.14061570173255125
	pesos_i(15176) := b"0000000000000000_0000000000000000_0001010111000011_1000001011010001"; -- 0.08501451121517457
	pesos_i(15177) := b"0000000000000000_0000000000000000_0010000110011100_1111000111111111"; -- 0.13130104507568163
	pesos_i(15178) := b"1111111111111111_1111111111111111_1111101111110100_1011011011110100"; -- -0.015797200726428817
	pesos_i(15179) := b"1111111111111111_1111111111111111_1110111100001100_1100100100011000"; -- -0.06621115844921832
	pesos_i(15180) := b"1111111111111111_1111111111111111_1101111101011001_0111101110010010"; -- -0.12754085248049032
	pesos_i(15181) := b"0000000000000000_0000000000000000_0001010111111111_1100110110110111"; -- 0.08593450271585037
	pesos_i(15182) := b"1111111111111111_1111111111111111_1110000100011111_1001110111000010"; -- -0.12061132452778618
	pesos_i(15183) := b"0000000000000000_0000000000000000_0001111100100000_1111101000010100"; -- 0.12159693707394152
	pesos_i(15184) := b"0000000000000000_0000000000000000_0001001100001011_0011111101000001"; -- 0.07439036701144121
	pesos_i(15185) := b"0000000000000000_0000000000000000_0000011011100011_0001110100101110"; -- 0.02690298446288662
	pesos_i(15186) := b"1111111111111111_1111111111111111_1110110101101001_0100100011110000"; -- -0.07261222978601657
	pesos_i(15187) := b"0000000000000000_0000000000000000_0001001110100111_1001101100100001"; -- 0.07677621424423689
	pesos_i(15188) := b"0000000000000000_0000000000000000_0001111111010110_1100000010011011"; -- 0.12437061103172006
	pesos_i(15189) := b"0000000000000000_0000000000000000_0000010100000001_1110010101110111"; -- 0.019560185937416704
	pesos_i(15190) := b"1111111111111111_1111111111111111_1111100110100000_0011110011011001"; -- -0.024898716995673743
	pesos_i(15191) := b"0000000000000000_0000000000000000_0000101100011111_1111101011010000"; -- 0.04345672205682857
	pesos_i(15192) := b"0000000000000000_0000000000000000_0001100101100110_1010110100000100"; -- 0.09922295907911609
	pesos_i(15193) := b"0000000000000000_0000000000000000_0001001001000111_0101011111011110"; -- 0.07140111133471727
	pesos_i(15194) := b"1111111111111111_1111111111111111_1110010110001110_0110111010001001"; -- -0.10329541359976402
	pesos_i(15195) := b"0000000000000000_0000000000000000_0010010111110010_0110111111011001"; -- 0.1482305435200401
	pesos_i(15196) := b"0000000000000000_0000000000000000_0010010010011011_0101110001100101"; -- 0.14299561953378406
	pesos_i(15197) := b"0000000000000000_0000000000000000_0001111100111000_0001011001000000"; -- 0.12194956844850226
	pesos_i(15198) := b"0000000000000000_0000000000000000_0001001101100110_1000111110011001"; -- 0.07578370567997988
	pesos_i(15199) := b"1111111111111111_1111111111111111_1101101001001010_1111101011101011"; -- -0.14729339370326677
	pesos_i(15200) := b"0000000000000000_0000000000000000_0000010100011100_0010111101010011"; -- 0.019961316894349174
	pesos_i(15201) := b"0000000000000000_0000000000000000_0000111010111101_1110110000001000"; -- 0.05758547968947894
	pesos_i(15202) := b"0000000000000000_0000000000000000_0000011100000010_1011100111111010"; -- 0.027385352723827774
	pesos_i(15203) := b"1111111111111111_1111111111111111_1101111101010110_0111100011111110"; -- -0.12758678241482807
	pesos_i(15204) := b"0000000000000000_0000000000000000_0000111100100100_1010010010111100"; -- 0.059152885381033825
	pesos_i(15205) := b"0000000000000000_0000000000000000_0001101001101011_0001010000010000"; -- 0.10319638614685221
	pesos_i(15206) := b"1111111111111111_1111111111111111_1110011011101011_1110111000000001"; -- -0.09796249847244713
	pesos_i(15207) := b"0000000000000000_0000000000000000_0001110111001111_1101111001011111"; -- 0.11645307364343813
	pesos_i(15208) := b"1111111111111111_1111111111111111_1110100101100010_1110000101001101"; -- -0.08833495979797307
	pesos_i(15209) := b"0000000000000000_0000000000000000_0000110000101011_1110111001001111"; -- 0.047545332323256674
	pesos_i(15210) := b"1111111111111111_1111111111111111_1111111011111010_0011101110110111"; -- -0.003994243401514209
	pesos_i(15211) := b"0000000000000000_0000000000000000_0010000001010110_1110001111110110"; -- 0.1263258433341319
	pesos_i(15212) := b"0000000000000000_0000000000000000_0001111000100001_0100000001111010"; -- 0.117694883254297
	pesos_i(15213) := b"0000000000000000_0000000000000000_0000010000111000_0010111010101111"; -- 0.016482274795475902
	pesos_i(15214) := b"0000000000000000_0000000000000000_0001100110000011_0100011010001100"; -- 0.09965935639778296
	pesos_i(15215) := b"0000000000000000_0000000000000000_0000010110111110_1101011000100101"; -- 0.022443183961549942
	pesos_i(15216) := b"0000000000000000_0000000000000000_0000001011010110_1001110100101111"; -- 0.011087249737073257
	pesos_i(15217) := b"1111111111111111_1111111111111111_1111111100111101_0101111100000010"; -- -0.002969800952992859
	pesos_i(15218) := b"1111111111111111_1111111111111111_1111110101101100_0111011010010101"; -- -0.010063732755579284
	pesos_i(15219) := b"1111111111111111_1111111111111111_1110001111110011_1010011100101011"; -- -0.10956340036149456
	pesos_i(15220) := b"1111111111111111_1111111111111111_1111100111101111_0101011111001000"; -- -0.02369166718443208
	pesos_i(15221) := b"0000000000000000_0000000000000000_0010010100010111_1010011110110011"; -- 0.1448921977483987
	pesos_i(15222) := b"1111111111111111_1111111111111111_1110111010001111_0000011110001000"; -- -0.06813004420679133
	pesos_i(15223) := b"0000000000000000_0000000000000000_0010011111101110_1001010110110001"; -- 0.15598426413580005
	pesos_i(15224) := b"0000000000000000_0000000000000000_0000100101110111_0111000000110111"; -- 0.03697873451932398
	pesos_i(15225) := b"1111111111111111_1111111111111111_1101111011010110_1101111000001111"; -- -0.1295338833976236
	pesos_i(15226) := b"0000000000000000_0000000000000000_0010000110100001_1000001111111010"; -- 0.13137078145921
	pesos_i(15227) := b"1111111111111111_1111111111111111_1101100101001011_0110001000000110"; -- -0.15119349819477276
	pesos_i(15228) := b"1111111111111111_1111111111111111_1111010010101010_1111110001101100"; -- -0.04426596039638661
	pesos_i(15229) := b"0000000000000000_0000000000000000_0001100011101011_1111011000000100"; -- 0.09735047920537673
	pesos_i(15230) := b"1111111111111111_1111111111111111_1111100100111111_0110110010111110"; -- -0.026375964701530485
	pesos_i(15231) := b"0000000000000000_0000000000000000_0000001011100000_1111000001111001"; -- 0.01124480204236313
	pesos_i(15232) := b"0000000000000000_0000000000000000_0010000000100101_1010010100011111"; -- 0.1255744171706717
	pesos_i(15233) := b"0000000000000000_0000000000000000_0000100101011010_0101100001100001"; -- 0.03653480885574359
	pesos_i(15234) := b"0000000000000000_0000000000000000_0010010100100110_0001010100000011"; -- 0.14511233643485785
	pesos_i(15235) := b"1111111111111111_1111111111111111_1111111000010000_0000000101010001"; -- -0.007568280881671062
	pesos_i(15236) := b"1111111111111111_1111111111111111_1110111001100100_1111110111011011"; -- -0.06877149007166215
	pesos_i(15237) := b"0000000000000000_0000000000000000_0001001010110010_0010010010101011"; -- 0.0730307501327683
	pesos_i(15238) := b"0000000000000000_0000000000000000_0000110010001010_0000101010110111"; -- 0.048981351531327245
	pesos_i(15239) := b"0000000000000000_0000000000000000_0000000100000111_0000110001001011"; -- 0.004013794237106524
	pesos_i(15240) := b"1111111111111111_1111111111111111_1110110011100011_0111010100100000"; -- -0.0746542735751049
	pesos_i(15241) := b"1111111111111111_1111111111111111_1111111001011001_1111111110100010"; -- -0.00643923081560555
	pesos_i(15242) := b"1111111111111111_1111111111111111_1110001000100000_1000000110101000"; -- -0.11669149073879845
	pesos_i(15243) := b"1111111111111111_1111111111111111_1110001011010110_1100100101100110"; -- -0.11391011491393478
	pesos_i(15244) := b"1111111111111111_1111111111111111_1110110100001100_1110011110000111"; -- -0.07402184451007425
	pesos_i(15245) := b"1111111111111111_1111111111111111_1111010100111100_1011010101110111"; -- -0.042042406603946585
	pesos_i(15246) := b"0000000000000000_0000000000000000_0000101000011111_0010110001011000"; -- 0.039538165623405695
	pesos_i(15247) := b"0000000000000000_0000000000000000_0001000000110000_0110110111011000"; -- 0.06323896903162135
	pesos_i(15248) := b"0000000000000000_0000000000000000_0001010001000110_1010000110111000"; -- 0.07920275447676085
	pesos_i(15249) := b"1111111111111111_1111111111111111_1110000100010111_1100000000111010"; -- -0.12073134018920918
	pesos_i(15250) := b"1111111111111111_1111111111111111_1110110110010011_0110110101011001"; -- -0.07196919048059335
	pesos_i(15251) := b"0000000000000000_0000000000000000_0000100100011110_0010001000000001"; -- 0.03561604039560172
	pesos_i(15252) := b"1111111111111111_1111111111111111_1110000111011010_0001001100001010"; -- -0.11776619913475263
	pesos_i(15253) := b"0000000000000000_0000000000000000_0010000010100001_0110111111000110"; -- 0.1274633271457356
	pesos_i(15254) := b"0000000000000000_0000000000000000_0010000000111000_0010100010010001"; -- 0.12585691010976308
	pesos_i(15255) := b"1111111111111111_1111111111111111_1110000000110011_1100011111101011"; -- -0.12420988565261734
	pesos_i(15256) := b"0000000000000000_0000000000000000_0010010010110111_0100010100100010"; -- 0.14342147898999977
	pesos_i(15257) := b"0000000000000000_0000000000000000_0000111011011001_0001000101110101"; -- 0.057999697778514304
	pesos_i(15258) := b"1111111111111111_1111111111111111_1111011011110010_0010110010101001"; -- -0.035367210984233524
	pesos_i(15259) := b"1111111111111111_1111111111111111_1110101101011100_0010010011111111"; -- -0.0806252361642757
	pesos_i(15260) := b"0000000000000000_0000000000000000_0010000110001000_1101110010111000"; -- 0.1309946011474064
	pesos_i(15261) := b"0000000000000000_0000000000000000_0000101101000001_0010011101000100"; -- 0.04396291162254709
	pesos_i(15262) := b"0000000000000000_0000000000000000_0000111011110111_0110111010010001"; -- 0.058463011133357876
	pesos_i(15263) := b"0000000000000000_0000000000000000_0000111101001100_0001010000001011"; -- 0.05975461260218813
	pesos_i(15264) := b"1111111111111111_1111111111111111_1110111001011011_1111101011100100"; -- -0.06890899588959518
	pesos_i(15265) := b"0000000000000000_0000000000000000_0001010111111010_1111100101111000"; -- 0.08586081671294285
	pesos_i(15266) := b"0000000000000000_0000000000000000_0001010100010111_0001100001001100"; -- 0.08238365024894057
	pesos_i(15267) := b"1111111111111111_1111111111111111_1111100010110001_0001100101001001"; -- -0.028547687210405754
	pesos_i(15268) := b"1111111111111111_1111111111111111_1110110001011110_0001011101110110"; -- -0.0766892754297723
	pesos_i(15269) := b"1111111111111111_1111111111111111_1111110000001111_1110010000100001"; -- -0.015382520532519059
	pesos_i(15270) := b"0000000000000000_0000000000000000_0000010110101001_1111100101110111"; -- 0.022124854646073847
	pesos_i(15271) := b"1111111111111111_1111111111111111_1111001100100110_0011100111111010"; -- -0.05019796035614114
	pesos_i(15272) := b"1111111111111111_1111111111111111_1101011001111111_1010011010100000"; -- -0.16211470214180504
	pesos_i(15273) := b"0000000000000000_0000000000000000_0001110001111010_1100010111111101"; -- 0.11124837336248118
	pesos_i(15274) := b"1111111111111111_1111111111111111_1111010101011011_0001011101101000"; -- -0.041578805109102196
	pesos_i(15275) := b"1111111111111111_1111111111111111_1111011000111010_0100001011011010"; -- -0.038173505602860376
	pesos_i(15276) := b"0000000000000000_0000000000000000_0001011101000011_0001001011011001"; -- 0.0908672122668248
	pesos_i(15277) := b"0000000000000000_0000000000000000_0001101101000001_0001010111001100"; -- 0.10646187047944414
	pesos_i(15278) := b"1111111111111111_1111111111111111_1110000101011001_0101100101010100"; -- -0.119730393395365
	pesos_i(15279) := b"1111111111111111_1111111111111111_1110111000000111_0000101001011011"; -- -0.07020507127720543
	pesos_i(15280) := b"0000000000000000_0000000000000000_0001100101101000_0111011101110000"; -- 0.09925028317187451
	pesos_i(15281) := b"0000000000000000_0000000000000000_0010001010001101_1111110001011110"; -- 0.13497903154033417
	pesos_i(15282) := b"1111111111111111_1111111111111111_1110101001000110_0100101001000110"; -- -0.08486495768461289
	pesos_i(15283) := b"1111111111111111_1111111111111111_1111011101100110_0001111001011010"; -- -0.033598044521467675
	pesos_i(15284) := b"0000000000000000_0000000000000000_0001010011100110_1001110000011000"; -- 0.08164382546204363
	pesos_i(15285) := b"0000000000000000_0000000000000000_0010000011001010_0101110010011001"; -- 0.12808779463852613
	pesos_i(15286) := b"1111111111111111_1111111111111111_1101110011111000_1011010111000110"; -- -0.13682998584640005
	pesos_i(15287) := b"0000000000000000_0000000000000000_0001000100110111_1000101110101100"; -- 0.0672538085843555
	pesos_i(15288) := b"1111111111111111_1111111111111111_1101011111011000_0001001111101110"; -- -0.15685916369570432
	pesos_i(15289) := b"0000000000000000_0000000000000000_0001101010011001_0100110111101001"; -- 0.10390173864163826
	pesos_i(15290) := b"1111111111111111_1111111111111111_1110010000111100_0000111100000000"; -- -0.10845857848724064
	pesos_i(15291) := b"0000000000000000_0000000000000000_0001011000111111_1010001101101100"; -- 0.08690854438598936
	pesos_i(15292) := b"0000000000000000_0000000000000000_0000000001010110_0111110111001111"; -- 0.0013197545749027814
	pesos_i(15293) := b"0000000000000000_0000000000000000_0000111110101000_1100110010000101"; -- 0.06116941693044329
	pesos_i(15294) := b"0000000000000000_0000000000000000_0001101010111011_0110110000111000"; -- 0.1044223438091618
	pesos_i(15295) := b"1111111111111111_1111111111111111_1110100101101111_1010010101101010"; -- -0.08814016490802228
	pesos_i(15296) := b"1111111111111111_1111111111111111_1110011011011011_1100101110110011"; -- -0.0982086837585865
	pesos_i(15297) := b"1111111111111111_1111111111111111_1111110111110001_0110000000000110"; -- -0.008035658427381022
	pesos_i(15298) := b"0000000000000000_0000000000000000_0010010110001110_1011101011000101"; -- 0.14670913037658226
	pesos_i(15299) := b"0000000000000000_0000000000000000_0001110111110101_1101010001111111"; -- 0.11703231912694204
	pesos_i(15300) := b"0000000000000000_0000000000000000_0001011011100001_0111100011001000"; -- 0.08937792673682333
	pesos_i(15301) := b"1111111111111111_1111111111111111_1111000011110101_1000101010111111"; -- -0.058753326755322875
	pesos_i(15302) := b"0000000000000000_0000000000000000_0001101101011111_1011111110101111"; -- 0.10692976026165427
	pesos_i(15303) := b"0000000000000000_0000000000000000_0000001010110011_1000001110001011"; -- 0.010551663926496138
	pesos_i(15304) := b"1111111111111111_1111111111111111_1111000010100000_0011100010011001"; -- -0.060055220268604145
	pesos_i(15305) := b"0000000000000000_0000000000000000_0000010011000100_0110001110111001"; -- 0.018621666516551245
	pesos_i(15306) := b"0000000000000000_0000000000000000_0010001111010001_1110101001110011"; -- 0.13992181128081146
	pesos_i(15307) := b"0000000000000000_0000000000000000_0010010111100010_1000101001011000"; -- 0.14798798237335045
	pesos_i(15308) := b"0000000000000000_0000000000000000_0000000101011001_0111000001011000"; -- 0.0052709784474247335
	pesos_i(15309) := b"0000000000000000_0000000000000000_0001100011101010_1010111110111000"; -- 0.09733103039418972
	pesos_i(15310) := b"0000000000000000_0000000000000000_0010001001001101_0000111011101000"; -- 0.13398831522154817
	pesos_i(15311) := b"1111111111111111_1111111111111111_1110010110001110_0000001101100001"; -- -0.1033018006098553
	pesos_i(15312) := b"1111111111111111_1111111111111111_1101011011011011_1111000001001000"; -- -0.16070650331151748
	pesos_i(15313) := b"1111111111111111_1111111111111111_1110111001100001_1011000101000001"; -- -0.06882183221790752
	pesos_i(15314) := b"0000000000000000_0000000000000000_0000110000010001_1001000001001001"; -- 0.04714299945136337
	pesos_i(15315) := b"0000000000000000_0000000000000000_0000001011110100_0010110011000100"; -- 0.011538312712336327
	pesos_i(15316) := b"0000000000000000_0000000000000000_0000101010111101_0111001001011010"; -- 0.0419532270984947
	pesos_i(15317) := b"1111111111111111_1111111111111111_1111001001001100_1000101111010111"; -- -0.05351949681281109
	pesos_i(15318) := b"0000000000000000_0000000000000000_0000001010110010_1001110010110001"; -- 0.010537904063347979
	pesos_i(15319) := b"1111111111111111_1111111111111111_1110101010100011_0011110111101110"; -- -0.08344662600032135
	pesos_i(15320) := b"1111111111111111_1111111111111111_1101100100111011_1001101101010110"; -- -0.15143422271749976
	pesos_i(15321) := b"0000000000000000_0000000000000000_0010001100101100_1101010101100000"; -- 0.1374028549316481
	pesos_i(15322) := b"1111111111111111_1111111111111111_1111000100011001_1100000000110101"; -- -0.05820082377689291
	pesos_i(15323) := b"1111111111111111_1111111111111111_1111000000010101_0101001010011111"; -- -0.06217464081342346
	pesos_i(15324) := b"0000000000000000_0000000000000000_0000100001100100_1011000101101101"; -- 0.03278645431655611
	pesos_i(15325) := b"0000000000000000_0000000000000000_0001100001000011_0111110011010000"; -- 0.09477977835906426
	pesos_i(15326) := b"0000000000000000_0000000000000000_0001101110100011_1001111100011101"; -- 0.10796541659500544
	pesos_i(15327) := b"1111111111111111_1111111111111111_1111110101000111_1110101100001000"; -- -0.010621366950217963
	pesos_i(15328) := b"0000000000000000_0000000000000000_0000111100110110_0101011111001110"; -- 0.05942295820518562
	pesos_i(15329) := b"0000000000000000_0000000000000000_0001011011011000_1001011000110010"; -- 0.0892423507962128
	pesos_i(15330) := b"0000000000000000_0000000000000000_0010010110101100_1011111011110110"; -- 0.1471671439560508
	pesos_i(15331) := b"0000000000000000_0000000000000000_0001110111011111_1111001111010111"; -- 0.11669849395226067
	pesos_i(15332) := b"0000000000000000_0000000000000000_0000101011000110_0100010110111000"; -- 0.042087895761627345
	pesos_i(15333) := b"0000000000000000_0000000000000000_0001000001111010_1010110111001101"; -- 0.06437193157804705
	pesos_i(15334) := b"1111111111111111_1111111111111111_1110001011011010_1110100011011111"; -- -0.11384720368909969
	pesos_i(15335) := b"1111111111111111_1111111111111111_1110100101100111_1011011100111100"; -- -0.08826117315283091
	pesos_i(15336) := b"0000000000000000_0000000000000000_0010001100001000_1110100100010011"; -- 0.13685471260963555
	pesos_i(15337) := b"0000000000000000_0000000000000000_0010011011100010_1111100110101110"; -- 0.15190086839336028
	pesos_i(15338) := b"1111111111111111_1111111111111111_1101111001111001_0000011110010001"; -- -0.13096573549333496
	pesos_i(15339) := b"0000000000000000_0000000000000000_0010010100100101_0101010101100011"; -- 0.1451009146660318
	pesos_i(15340) := b"1111111111111111_1111111111111111_1110101111101101_0100100000100111"; -- -0.07841061643946806
	pesos_i(15341) := b"1111111111111111_1111111111111111_1111100011011101_1101110010001001"; -- -0.027864662729803428
	pesos_i(15342) := b"1111111111111111_1111111111111111_1111110100010011_1110101010000001"; -- -0.011414855416809361
	pesos_i(15343) := b"0000000000000000_0000000000000000_0001101011001101_1011001000111010"; -- 0.10470117484590205
	pesos_i(15344) := b"0000000000000000_0000000000000000_0001001011000100_1101100101111111"; -- 0.073316186352272
	pesos_i(15345) := b"1111111111111111_1111111111111111_1110000110111001_1010000001100100"; -- -0.11826131405445107
	pesos_i(15346) := b"1111111111111111_1111111111111111_1101110110100100_1111010110000001"; -- -0.13420167540372285
	pesos_i(15347) := b"1111111111111111_1111111111111111_1110100101100000_1000000101111000"; -- -0.08837118922857114
	pesos_i(15348) := b"1111111111111111_1111111111111111_1111001001111101_0011010010011101"; -- -0.05277701528396675
	pesos_i(15349) := b"0000000000000000_0000000000000000_0001001100010100_1001111111111110"; -- 0.07453346210331371
	pesos_i(15350) := b"0000000000000000_0000000000000000_0010000000110111_0111011001111110"; -- 0.12584629606453104
	pesos_i(15351) := b"0000000000000000_0000000000000000_0001000100100000_1010101111010111"; -- 0.06690477378797549
	pesos_i(15352) := b"1111111111111111_1111111111111111_1111011100111011_1010110110001111"; -- -0.03424563646563903
	pesos_i(15353) := b"1111111111111111_1111111111111111_1111101010110011_1100101101110110"; -- -0.020694049577273162
	pesos_i(15354) := b"0000000000000000_0000000000000000_0010001010110101_1100010000010110"; -- 0.1355860284295206
	pesos_i(15355) := b"0000000000000000_0000000000000000_0000000110010110_1001100101111001"; -- 0.006204215978763734
	pesos_i(15356) := b"0000000000000000_0000000000000000_0000010000011011_0000110111000011"; -- 0.016037807669327594
	pesos_i(15357) := b"1111111111111111_1111111111111111_1110000010111100_1101010111001001"; -- -0.12211860516059952
	pesos_i(15358) := b"0000000000000000_0000000000000000_0000111011101000_1011010011101101"; -- 0.058238323096033794
	pesos_i(15359) := b"0000000000000000_0000000000000000_0000000111101010_1000101000010100"; -- 0.0074850368433270744
	pesos_i(15360) := b"0000000000000000_0000000000000000_0001000100011110_0110110011111001"; -- 0.06687050888133964
	pesos_i(15361) := b"1111111111111111_1111111111111111_1110110101010100_1110011011010110"; -- -0.0729232528553983
	pesos_i(15362) := b"1111111111111111_1111111111111111_1111110000000111_1110010001110011"; -- -0.015504571748568318
	pesos_i(15363) := b"0000000000000000_0000000000000000_0001100101101100_1100001110111110"; -- 0.09931586627150467
	pesos_i(15364) := b"1111111111111111_1111111111111111_1101100001101110_1110010000001011"; -- -0.1545579408473243
	pesos_i(15365) := b"0000000000000000_0000000000000000_0001110101110010_0101100011110010"; -- 0.11502605342784643
	pesos_i(15366) := b"1111111111111111_1111111111111111_1111011000000000_0001011100011001"; -- -0.0390611232912701
	pesos_i(15367) := b"1111111111111111_1111111111111111_1101110010010001_0000000001111101"; -- -0.13841244647021372
	pesos_i(15368) := b"1111111111111111_1111111111111111_1110001111010011_0010101110001011"; -- -0.11005905012798645
	pesos_i(15369) := b"1111111111111111_1111111111111111_1110100010100011_1000010111101101"; -- -0.09125483478212862
	pesos_i(15370) := b"0000000000000000_0000000000000000_0000000001010110_0101101000010101"; -- 0.0013176250507528642
	pesos_i(15371) := b"1111111111111111_1111111111111111_1110011011010000_0000100101000000"; -- -0.09838812043887142
	pesos_i(15372) := b"0000000000000000_0000000000000000_0001011100111100_0101000011010110"; -- 0.09076409559196832
	pesos_i(15373) := b"0000000000000000_0000000000000000_0001111010111010_1000001011111111"; -- 0.12003344263734436
	pesos_i(15374) := b"1111111111111111_1111111111111111_1110110101000110_1001001001111100"; -- -0.07314190364326832
	pesos_i(15375) := b"1111111111111111_1111111111111111_1111011100111101_0101101101111000"; -- -0.03422001199897155
	pesos_i(15376) := b"1111111111111111_1111111111111111_1111111000110010_1001010011111100"; -- -0.007040680478491622
	pesos_i(15377) := b"0000000000000000_0000000000000000_0001110001011010_0001111111011010"; -- 0.11075018940211391
	pesos_i(15378) := b"1111111111111111_1111111111111111_1111011100011011_0001110000100011"; -- -0.03474258568137401
	pesos_i(15379) := b"1111111111111111_1111111111111111_1110001001110111_0011010111000110"; -- -0.1153684989680222
	pesos_i(15380) := b"0000000000000000_0000000000000000_0000001110000011_0001111100001001"; -- 0.013719501191250491
	pesos_i(15381) := b"1111111111111111_1111111111111111_1101110001101000_0010001010010110"; -- -0.13903602443229038
	pesos_i(15382) := b"0000000000000000_0000000000000000_0000110011011100_1001000010100101"; -- 0.050240555177018684
	pesos_i(15383) := b"1111111111111111_1111111111111111_1111110111011111_0000011101110001"; -- -0.008315596499720388
	pesos_i(15384) := b"1111111111111111_1111111111111111_1111110001100001_0110001110010110"; -- -0.01413896175487011
	pesos_i(15385) := b"0000000000000000_0000000000000000_0000101111011010_1110001011101001"; -- 0.04630869102415155
	pesos_i(15386) := b"1111111111111111_1111111111111111_1110100101011101_1001111100001111"; -- -0.08841520194348293
	pesos_i(15387) := b"1111111111111111_1111111111111111_1111101100111111_0000110010010000"; -- -0.018569197439789593
	pesos_i(15388) := b"0000000000000000_0000000000000000_0000011101110100_0000101001011011"; -- 0.02911438677897622
	pesos_i(15389) := b"0000000000000000_0000000000000000_0001010100100110_0000001110100011"; -- 0.08261130076077079
	pesos_i(15390) := b"0000000000000000_0000000000000000_0000110010010110_1111000101000001"; -- 0.0491781983017314
	pesos_i(15391) := b"1111111111111111_1111111111111111_1101110011001000_0011001111101111"; -- -0.13757014662256298
	pesos_i(15392) := b"0000000000000000_0000000000000000_0001111110111111_0100010100100001"; -- 0.12401229908161646
	pesos_i(15393) := b"0000000000000000_0000000000000000_0001100101011110_1110100100011110"; -- 0.09910447095541776
	pesos_i(15394) := b"0000000000000000_0000000000000000_0001001110110011_1000000001110110"; -- 0.07695773019079598
	pesos_i(15395) := b"0000000000000000_0000000000000000_0001001101010110_1101010101110111"; -- 0.07554372928236991
	pesos_i(15396) := b"0000000000000000_0000000000000000_0010010111111101_1110010110100101"; -- 0.14840541154670153
	pesos_i(15397) := b"0000000000000000_0000000000000000_0000010011000001_0001000100000100"; -- 0.018570960424453185
	pesos_i(15398) := b"0000000000000000_0000000000000000_0001101111111001_0000110111000010"; -- 0.10926900846570804
	pesos_i(15399) := b"1111111111111111_1111111111111111_1111101110011100_0000100011100010"; -- -0.01715034955494039
	pesos_i(15400) := b"0000000000000000_0000000000000000_0000110101101011_0011101000010010"; -- 0.05241740179344854
	pesos_i(15401) := b"1111111111111111_1111111111111111_1110010101110011_1000100100001000"; -- -0.10370582145715831
	pesos_i(15402) := b"0000000000000000_0000000000000000_0010010011100111_0100010110100101"; -- 0.14415393135726326
	pesos_i(15403) := b"0000000000000000_0000000000000000_0001010010110011_1000010110001110"; -- 0.08086428364237175
	pesos_i(15404) := b"0000000000000000_0000000000000000_0000100011011001_1010110010011001"; -- 0.0345714448495512
	pesos_i(15405) := b"0000000000000000_0000000000000000_0000101010111011_0111111000111000"; -- 0.04192341687038482
	pesos_i(15406) := b"0000000000000000_0000000000000000_0010010001101101_0101001111100100"; -- 0.14229320828179823
	pesos_i(15407) := b"0000000000000000_0000000000000000_0000010101101111_1011000010011101"; -- 0.021235502542677816
	pesos_i(15408) := b"0000000000000000_0000000000000000_0000111000001010_0110010000011110"; -- 0.05484605541609326
	pesos_i(15409) := b"1111111111111111_1111111111111111_1111100101100001_0101101010010001"; -- -0.025858249281621407
	pesos_i(15410) := b"1111111111111111_1111111111111111_1111000100011011_1010010011110111"; -- -0.05817193009792994
	pesos_i(15411) := b"1111111111111111_1111111111111111_1111110010000001_1110111010100001"; -- -0.013642392714009069
	pesos_i(15412) := b"1111111111111111_1111111111111111_1101101010000111_0110101100010110"; -- -0.14637118077284716
	pesos_i(15413) := b"0000000000000000_0000000000000000_0010010010100110_1101000000111011"; -- 0.14317037058109283
	pesos_i(15414) := b"0000000000000000_0000000000000000_0000011100000001_1100011110011001"; -- 0.02737090567315777
	pesos_i(15415) := b"1111111111111111_1111111111111111_1110110011010000_1000100000001111"; -- -0.07494306222579934
	pesos_i(15416) := b"1111111111111111_1111111111111111_1110011110001110_0000011001001001"; -- -0.09548912739843733
	pesos_i(15417) := b"1111111111111111_1111111111111111_1111010100011001_1111001011110110"; -- -0.04257279867608931
	pesos_i(15418) := b"0000000000000000_0000000000000000_0001011110110010_1100101100110111"; -- 0.09257192694795993
	pesos_i(15419) := b"0000000000000000_0000000000000000_0000000011100111_0101010001011011"; -- 0.003529808258083461
	pesos_i(15420) := b"1111111111111111_1111111111111111_1111100000000110_1101111010111100"; -- -0.031145171198140913
	pesos_i(15421) := b"0000000000000000_0000000000000000_0001101000100011_0100100011101001"; -- 0.10210090337739965
	pesos_i(15422) := b"0000000000000000_0000000000000000_0000001010101101_0100111001000110"; -- 0.010456935878489075
	pesos_i(15423) := b"1111111111111111_1111111111111111_1111001010010110_1110001101101100"; -- -0.05238512634515635
	pesos_i(15424) := b"0000000000000000_0000000000000000_0001001010101010_0100000001100001"; -- 0.07291033130807333
	pesos_i(15425) := b"0000000000000000_0000000000000000_0001000010001001_1101111010101111"; -- 0.0646037271210522
	pesos_i(15426) := b"1111111111111111_1111111111111111_1111100010000000_1010100011100010"; -- -0.02928680887997899
	pesos_i(15427) := b"1111111111111111_1111111111111111_1110101001000011_1111000101000000"; -- -0.0849007815624668
	pesos_i(15428) := b"0000000000000000_0000000000000000_0001100111111111_1011001101110010"; -- 0.10155793693722323
	pesos_i(15429) := b"1111111111111111_1111111111111111_1110111110101010_0111000000101111"; -- -0.06380556929096452
	pesos_i(15430) := b"0000000000000000_0000000000000000_0010100011111100_1111010011000000"; -- 0.1601098030598047
	pesos_i(15431) := b"1111111111111111_1111111111111111_1101101010010001_0011101110011110"; -- -0.1462214221525318
	pesos_i(15432) := b"0000000000000000_0000000000000000_0001010011010100_1001001000101100"; -- 0.08136857576338374
	pesos_i(15433) := b"1111111111111111_1111111111111111_1111101011001111_1110001011011100"; -- -0.020265408767499403
	pesos_i(15434) := b"0000000000000000_0000000000000000_0000100101110000_1101111011100101"; -- 0.03687851987181526
	pesos_i(15435) := b"0000000000000000_0000000000000000_0010010001101011_0101011101001101"; -- 0.14226289402311326
	pesos_i(15436) := b"1111111111111111_1111111111111111_1101110100011110_0011010110000010"; -- -0.13625779707804894
	pesos_i(15437) := b"1111111111111111_1111111111111111_1101010000010000_0110000001111110"; -- -0.17162510797360842
	pesos_i(15438) := b"0000000000000000_0000000000000000_0010001110001010_0010011100011001"; -- 0.13882679318475974
	pesos_i(15439) := b"0000000000000000_0000000000000000_0001101001101001_0010011001110101"; -- 0.10316696509693277
	pesos_i(15440) := b"1111111111111111_1111111111111111_1110101101011110_0010010010110011"; -- -0.08059473634267315
	pesos_i(15441) := b"1111111111111111_1111111111111111_1111011111111110_0000110100010010"; -- -0.03127973851453704
	pesos_i(15442) := b"1111111111111111_1111111111111111_1111110011001101_0000110000110110"; -- -0.012496220376584374
	pesos_i(15443) := b"1111111111111111_1111111111111111_1101111010100101_1101011001110111"; -- -0.1302820166279927
	pesos_i(15444) := b"1111111111111111_1111111111111111_1110100001110001_1101001010011110"; -- -0.09201320310518733
	pesos_i(15445) := b"0000000000000000_0000000000000000_0010100100010101_0010101001110111"; -- 0.16047921560527534
	pesos_i(15446) := b"1111111111111111_1111111111111111_1111111001111111_1111001100001110"; -- -0.005860146594133379
	pesos_i(15447) := b"1111111111111111_1111111111111111_1110101111000110_1000010010110100"; -- -0.07900209999544083
	pesos_i(15448) := b"1111111111111111_1111111111111111_1110011011111101_0011101011101001"; -- -0.09769851509498616
	pesos_i(15449) := b"0000000000000000_0000000000000000_0001001011000100_1001100101001111"; -- 0.07331236053005023
	pesos_i(15450) := b"1111111111111111_1111111111111111_1110101001011111_0100011001000001"; -- -0.08448372753637579
	pesos_i(15451) := b"0000000000000000_0000000000000000_0000000110111100_0011101111000110"; -- 0.006778465013942695
	pesos_i(15452) := b"0000000000000000_0000000000000000_0000100000001110_1110010101001111"; -- 0.03147729098950412
	pesos_i(15453) := b"0000000000000000_0000000000000000_0001001000101001_1100011100101100"; -- 0.07094998191406911
	pesos_i(15454) := b"0000000000000000_0000000000000000_0000001000101100_0100010010001001"; -- 0.008487971830759175
	pesos_i(15455) := b"1111111111111111_1111111111111111_1111111001000101_1111011000011101"; -- -0.006744974092161243
	pesos_i(15456) := b"1111111111111111_1111111111111111_1110111000000011_1100110000110101"; -- -0.07025455199506728
	pesos_i(15457) := b"0000000000000000_0000000000000000_0010001111000101_1001111011000000"; -- 0.13973419358518377
	pesos_i(15458) := b"0000000000000000_0000000000000000_0001100010010000_1000100001001011"; -- 0.09595538928456022
	pesos_i(15459) := b"1111111111111111_1111111111111111_1110010001100011_1011000010100110"; -- -0.10785385071199548
	pesos_i(15460) := b"1111111111111111_1111111111111111_1110001111101111_1111110110001110"; -- -0.10961928638562775
	pesos_i(15461) := b"0000000000000000_0000000000000000_0001101011001001_0011000110001101"; -- 0.10463247013553237
	pesos_i(15462) := b"0000000000000000_0000000000000000_0011001101011101_0010100111111011"; -- 0.20064031960737136
	pesos_i(15463) := b"1111111111111111_1111111111111111_1111110001000100_1111010110011101"; -- -0.014572762593346791
	pesos_i(15464) := b"0000000000000000_0000000000000000_0001000001011111_0001100101111111"; -- 0.06395110458086949
	pesos_i(15465) := b"0000000000000000_0000000000000000_0000001100011010_0100011001100010"; -- 0.01211967359810202
	pesos_i(15466) := b"1111111111111111_1111111111111111_1111100011000111_1100001101110101"; -- -0.028201850915507594
	pesos_i(15467) := b"0000000000000000_0000000000000000_0000100101101110_0100011101000010"; -- 0.03683896407805856
	pesos_i(15468) := b"1111111111111111_1111111111111111_1110000110100011_1010001111000111"; -- -0.11859680541020394
	pesos_i(15469) := b"1111111111111111_1111111111111111_1110100110111111_1001111111100100"; -- -0.0869197910688791
	pesos_i(15470) := b"0000000000000000_0000000000000000_0000110000000010_0010010001101000"; -- 0.046907687557631916
	pesos_i(15471) := b"1111111111111111_1111111111111111_1110110000011111_0000111001111011"; -- -0.07765111438715071
	pesos_i(15472) := b"1111111111111111_1111111111111111_1110101111110100_1101110101111000"; -- -0.07829490484979643
	pesos_i(15473) := b"0000000000000000_0000000000000000_0001011110000110_1111010011010001"; -- 0.09190301983608624
	pesos_i(15474) := b"1111111111111111_1111111111111111_1111001011001010_1110000001000010"; -- -0.05159185790313579
	pesos_i(15475) := b"0000000000000000_0000000000000000_0001110111111000_1110000000001100"; -- 0.11707878384883011
	pesos_i(15476) := b"1111111111111111_1111111111111111_1111110010001100_0110111011111101"; -- -0.01348215406684044
	pesos_i(15477) := b"1111111111111111_1111111111111111_1111001000010101_0000101011100011"; -- -0.05436641655949959
	pesos_i(15478) := b"0000000000000000_0000000000000000_0000010101100110_0010100100111100"; -- 0.021090104277060047
	pesos_i(15479) := b"0000000000000000_0000000000000000_0010000010100110_0100001000100010"; -- 0.12753690083743136
	pesos_i(15480) := b"0000000000000000_0000000000000000_0010000011000011_0110001101110001"; -- 0.12798139104735523
	pesos_i(15481) := b"0000000000000000_0000000000000000_0010011000011011_1010011101000011"; -- 0.14885945685222912
	pesos_i(15482) := b"1111111111111111_1111111111111111_1111000110100101_0110000100110010"; -- -0.05607025662369449
	pesos_i(15483) := b"1111111111111111_1111111111111111_1101010101100111_1101011111100101"; -- -0.1663842263910117
	pesos_i(15484) := b"0000000000000000_0000000000000000_0000011000110101_0100000101010110"; -- 0.024250110098840042
	pesos_i(15485) := b"1111111111111111_1111111111111111_1110001011111010_0110100111111001"; -- -0.11336648627434683
	pesos_i(15486) := b"0000000000000000_0000000000000000_0001111101010001_1100000001101010"; -- 0.12234118077790299
	pesos_i(15487) := b"0000000000000000_0000000000000000_0001101011100110_0000011110110010"; -- 0.10507248019412367
	pesos_i(15488) := b"0000000000000000_0000000000000000_0001001011100101_0110110110000000"; -- 0.07381328937915985
	pesos_i(15489) := b"0000000000000000_0000000000000000_0000010110000101_0101110110010001"; -- 0.02156624592140035
	pesos_i(15490) := b"1111111111111111_1111111111111111_1111110111001110_0011110101001001"; -- -0.008571786613524717
	pesos_i(15491) := b"0000000000000000_0000000000000000_0000001110111010_0011011001100100"; -- 0.014560126813329254
	pesos_i(15492) := b"1111111111111111_1111111111111111_1110101010100100_1100110110001011"; -- -0.08342280724990268
	pesos_i(15493) := b"1111111111111111_1111111111111111_1111000100101011_1101110010110100"; -- -0.057924467046064715
	pesos_i(15494) := b"1111111111111111_1111111111111111_1101110010011110_0000000000110111"; -- -0.13821409850755584
	pesos_i(15495) := b"1111111111111111_1111111111111111_1111001001101111_0111000100110011"; -- -0.05298702709952446
	pesos_i(15496) := b"0000000000000000_0000000000000000_0001001001100010_1111111110100110"; -- 0.07182309915713256
	pesos_i(15497) := b"0000000000000000_0000000000000000_0001000001101010_1101000010111111"; -- 0.06412987387297797
	pesos_i(15498) := b"1111111111111111_1111111111111111_1110101001010001_1001011111000000"; -- -0.08469249299131358
	pesos_i(15499) := b"1111111111111111_1111111111111111_1111001101000011_1100111101100000"; -- -0.049746550600865906
	pesos_i(15500) := b"1111111111111111_1111111111111111_1111000010000001_1111010001101001"; -- -0.06051704812944044
	pesos_i(15501) := b"1111111111111111_1111111111111111_1110101010100000_0000100101110110"; -- -0.08349552972339927
	pesos_i(15502) := b"1111111111111111_1111111111111111_1111011001101110_0110011100010001"; -- -0.037377889928301565
	pesos_i(15503) := b"1111111111111111_1111111111111111_1110110101001101_0000001101110001"; -- -0.07304361806961558
	pesos_i(15504) := b"0000000000000000_0000000000000000_0000011011011001_0100000001011110"; -- 0.026752493868638087
	pesos_i(15505) := b"0000000000000000_0000000000000000_0010000000101111_0011110010011100"; -- 0.12572077564297507
	pesos_i(15506) := b"1111111111111111_1111111111111111_1101100001010010_1000110001011101"; -- -0.15499041308205846
	pesos_i(15507) := b"0000000000000000_0000000000000000_0000111000110100_0000001011100011"; -- 0.05548112904287321
	pesos_i(15508) := b"1111111111111111_1111111111111111_1110011001101011_0100100101101100"; -- -0.09992543326946798
	pesos_i(15509) := b"1111111111111111_1111111111111111_1110001001110010_0001010101111000"; -- -0.1154467184667696
	pesos_i(15510) := b"1111111111111111_1111111111111111_1111101101001110_1110100111111001"; -- -0.018327118599621522
	pesos_i(15511) := b"0000000000000000_0000000000000000_0000100011110000_1101110111101111"; -- 0.034925337688563124
	pesos_i(15512) := b"0000000000000000_0000000000000000_0000110110111111_0001011101100111"; -- 0.0536970735044433
	pesos_i(15513) := b"0000000000000000_0000000000000000_0010011001110000_0111111000100010"; -- 0.15015400255250358
	pesos_i(15514) := b"1111111111111111_1111111111111111_1111110100100010_1011001101011000"; -- -0.01118926136694152
	pesos_i(15515) := b"1111111111111111_1111111111111111_1111000111011000_0110111111101000"; -- -0.055291181433362424
	pesos_i(15516) := b"0000000000000000_0000000000000000_0001111011000111_1001101010011101"; -- 0.12023321480376703
	pesos_i(15517) := b"0000000000000000_0000000000000000_0001101111110110_1010011011111110"; -- 0.10923236554769694
	pesos_i(15518) := b"1111111111111111_1111111111111111_1101110000011011_1101011100011111"; -- -0.1402001905748892
	pesos_i(15519) := b"1111111111111111_1111111111111111_1111101111001001_0011101100001001"; -- -0.016460714521564217
	pesos_i(15520) := b"0000000000000000_0000000000000000_0001010100011000_0111001101000101"; -- 0.08240433157824388
	pesos_i(15521) := b"0000000000000000_0000000000000000_0000010110011000_1011011011011010"; -- 0.021861484652740997
	pesos_i(15522) := b"1111111111111111_1111111111111111_1110001000010010_1010011101011010"; -- -0.11690286691822656
	pesos_i(15523) := b"1111111111111111_1111111111111111_1101100110101110_1110010111011010"; -- -0.14967502055278356
	pesos_i(15524) := b"1111111111111111_1111111111111111_1111001110100011_1000011011100101"; -- -0.048286027148416275
	pesos_i(15525) := b"1111111111111111_1111111111111111_1101111101100001_0100101001011101"; -- -0.12742171498953242
	pesos_i(15526) := b"1111111111111111_1111111111111111_1111110011001011_1111101100010001"; -- -0.012512501168113161
	pesos_i(15527) := b"1111111111111111_1111111111111111_1111001101101010_1000100011100110"; -- -0.0491556585016076
	pesos_i(15528) := b"0000000000000000_0000000000000000_0010000001001000_1110011001000010"; -- 0.12611235718206396
	pesos_i(15529) := b"1111111111111111_1111111111111111_1111011111010011_0000100010011001"; -- -0.03193613301157626
	pesos_i(15530) := b"0000000000000000_0000000000000000_0001110011010101_0101101100001000"; -- 0.11263054790206524
	pesos_i(15531) := b"1111111111111111_1111111111111111_1111100111010010_1111010010000100"; -- -0.024124829917541685
	pesos_i(15532) := b"1111111111111111_1111111111111111_1110111011110100_0110010110000000"; -- -0.06658330560482142
	pesos_i(15533) := b"0000000000000000_0000000000000000_0000100111100111_1101101010001100"; -- 0.038694056665823984
	pesos_i(15534) := b"0000000000000000_0000000000000000_0001101101100110_0001100001011110"; -- 0.10702659877201165
	pesos_i(15535) := b"0000000000000000_0000000000000000_0001110101010011_1100001000111101"; -- 0.11455930693727596
	pesos_i(15536) := b"1111111111111111_1111111111111111_1110100100101011_0101001011100101"; -- -0.08918268126021202
	pesos_i(15537) := b"1111111111111111_1111111111111111_1111100110010110_1010011100100101"; -- -0.025044968966711316
	pesos_i(15538) := b"0000000000000000_0000000000000000_0001111011010110_1111101000101111"; -- 0.12046779305052062
	pesos_i(15539) := b"0000000000000000_0000000000000000_0010000001010000_1100100000100101"; -- 0.12623263256466546
	pesos_i(15540) := b"1111111111111111_1111111111111111_1101101111011010_1000110100110101"; -- -0.14119641733186727
	pesos_i(15541) := b"0000000000000000_0000000000000000_0010100011111011_1001100110100100"; -- 0.16008911368853385
	pesos_i(15542) := b"1111111111111111_1111111111111111_1101101101001111_0110110010111000"; -- -0.14331932543399975
	pesos_i(15543) := b"1111111111111111_1111111111111111_1110010000110001_0010000101111110"; -- -0.10862532312558344
	pesos_i(15544) := b"0000000000000000_0000000000000000_0000011101100111_0101010100111011"; -- 0.028920485367588254
	pesos_i(15545) := b"0000000000000000_0000000000000000_0001011010110111_1010100100010101"; -- 0.08873993653747038
	pesos_i(15546) := b"1111111111111111_1111111111111111_1110011111001000_1101111011111010"; -- -0.0945912017917333
	pesos_i(15547) := b"1111111111111111_1111111111111111_1110101110110000_1000001000000101"; -- -0.07933795344235914
	pesos_i(15548) := b"0000000000000000_0000000000000000_0000100011010110_1001111010010010"; -- 0.0345248323988163
	pesos_i(15549) := b"1111111111111111_1111111111111111_1111100000010101_0100100101111111"; -- -0.0309251847486521
	pesos_i(15550) := b"1111111111111111_1111111111111111_1111101110110110_0010110011010100"; -- -0.016751478524861804
	pesos_i(15551) := b"0000000000000000_0000000000000000_0001000011101010_0000111011100111"; -- 0.06607144479205165
	pesos_i(15552) := b"1111111111111111_1111111111111111_1111100110011011_1011100101001111"; -- -0.024967592444635135
	pesos_i(15553) := b"1111111111111111_1111111111111111_1110011001100001_1101110110011100"; -- -0.10006918847139906
	pesos_i(15554) := b"1111111111111111_1111111111111111_1101110010000000_0100100000000110"; -- -0.13866758215336325
	pesos_i(15555) := b"0000000000000000_0000000000000000_0001101000110001_1000111101001111"; -- 0.10231872256823381
	pesos_i(15556) := b"0000000000000000_0000000000000000_0001000110001101_1000100001000110"; -- 0.06856586180320162
	pesos_i(15557) := b"1111111111111111_1111111111111111_1101101111101101_0001010000010110"; -- -0.1409137196836307
	pesos_i(15558) := b"1111111111111111_1111111111111111_1111111110001011_0000011110101001"; -- -0.001784821685038268
	pesos_i(15559) := b"1111111111111111_1111111111111111_1110101010100101_0100001001101101"; -- -0.08341584045552472
	pesos_i(15560) := b"0000000000000000_0000000000000000_0001011001110101_0001011101011001"; -- 0.08772417002981427
	pesos_i(15561) := b"0000000000000000_0000000000000000_0010001011001111_1101101011111011"; -- 0.1359841215724197
	pesos_i(15562) := b"0000000000000000_0000000000000000_0001010000001110_0000011111000101"; -- 0.07833908626297235
	pesos_i(15563) := b"0000000000000000_0000000000000000_0000011011000111_0110111010011001"; -- 0.026480591195082864
	pesos_i(15564) := b"0000000000000000_0000000000000000_0001110011101110_1110001100011100"; -- 0.11302012852227512
	pesos_i(15565) := b"0000000000000000_0000000000000000_0010000000100111_0001011001110001"; -- 0.12559643039497703
	pesos_i(15566) := b"1111111111111111_1111111111111111_1110010011111011_1000100000001100"; -- -0.10553693499894581
	pesos_i(15567) := b"0000000000000000_0000000000000000_0000011110000111_1001110011111010"; -- 0.02941304314147352
	pesos_i(15568) := b"0000000000000000_0000000000000000_0001100101010111_0110010110111001"; -- 0.0989898277454933
	pesos_i(15569) := b"1111111111111111_1111111111111111_1101111101111001_0110110000100110"; -- -0.1270534904384392
	pesos_i(15570) := b"1111111111111111_1111111111111111_1110010100101101_0000010000100100"; -- -0.10478185769641749
	pesos_i(15571) := b"0000000000000000_0000000000000000_0001011100110001_1001001011001010"; -- 0.09060018006604323
	pesos_i(15572) := b"1111111111111111_1111111111111111_1101110101011100_0101110010111001"; -- -0.13530941467460347
	pesos_i(15573) := b"0000000000000000_0000000000000000_0001111001100111_0111011010011010"; -- 0.11876622445534515
	pesos_i(15574) := b"0000000000000000_0000000000000000_0000111000001001_1110011010111011"; -- 0.05483858162782882
	pesos_i(15575) := b"1111111111111111_1111111111111111_1111011100000001_1101110100001110"; -- -0.035127815346740233
	pesos_i(15576) := b"1111111111111111_1111111111111111_1111111010011010_1100011010111101"; -- -0.005450800808568608
	pesos_i(15577) := b"0000000000000000_0000000000000000_0001010111110000_0011111101000101"; -- 0.08569713044695458
	pesos_i(15578) := b"0000000000000000_0000000000000000_0000101101110110_0000101001010011"; -- 0.04476990240561585
	pesos_i(15579) := b"1111111111111111_1111111111111111_1111110100101010_1010101010100111"; -- -0.011067709262319527
	pesos_i(15580) := b"0000000000000000_0000000000000000_0000000001001101_0111101111110001"; -- 0.0011823141251827106
	pesos_i(15581) := b"1111111111111111_1111111111111111_1110101110000001_1100100000110000"; -- -0.08005093410944032
	pesos_i(15582) := b"1111111111111111_1111111111111111_1110101000101101_0100011110101010"; -- -0.08524658293624587
	pesos_i(15583) := b"1111111111111111_1111111111111111_1111111011011001_0100011000110011"; -- -0.004497158583214698
	pesos_i(15584) := b"1111111111111111_1111111111111111_1101101010111011_1000010111001110"; -- -0.14557613115856377
	pesos_i(15585) := b"0000000000000000_0000000000000000_0000000001101011_1100100000000100"; -- 0.0016446122036502559
	pesos_i(15586) := b"1111111111111111_1111111111111111_1111010110111010_1111001101001101"; -- -0.04011611335996295
	pesos_i(15587) := b"1111111111111111_1111111111111111_1111000001110100_1010000111110001"; -- -0.06072032799347883
	pesos_i(15588) := b"0000000000000000_0000000000000000_0001111001001011_1000100100010011"; -- 0.11834007953198485
	pesos_i(15589) := b"1111111111111111_1111111111111111_1110100001001010_0100110110100101"; -- -0.09261622169951546
	pesos_i(15590) := b"1111111111111111_1111111111111111_1110100110110110_0000000110110000"; -- -0.08706654989885919
	pesos_i(15591) := b"1111111111111111_1111111111111111_1111100000101001_0111001000000111"; -- -0.030617592987088778
	pesos_i(15592) := b"0000000000000000_0000000000000000_0001000001011101_1001100111100111"; -- 0.06392824056133821
	pesos_i(15593) := b"1111111111111111_1111111111111111_1101111010110111_0101001100011011"; -- -0.1300151882125175
	pesos_i(15594) := b"1111111111111111_1111111111111111_1111011100101111_1111110101010100"; -- -0.03442398732387136
	pesos_i(15595) := b"1111111111111111_1111111111111111_1111001100001000_1001001010011111"; -- -0.05065044042192909
	pesos_i(15596) := b"0000000000000000_0000000000000000_0000111111010110_0000011010100001"; -- 0.06185952586518159
	pesos_i(15597) := b"1111111111111111_1111111111111111_1110100010010010_0110101000111001"; -- -0.09151588533966734
	pesos_i(15598) := b"0000000000000000_0000000000000000_0000101111001010_0110011100000010"; -- 0.04605716516335882
	pesos_i(15599) := b"0000000000000000_0000000000000000_0001011011010011_1000001111001110"; -- 0.08916496070918181
	pesos_i(15600) := b"1111111111111111_1111111111111111_1110110110000000_0000101001111100"; -- -0.07226500016841045
	pesos_i(15601) := b"1111111111111111_1111111111111111_1111111111110011_1101000100110110"; -- -0.0001858942350979701
	pesos_i(15602) := b"0000000000000000_0000000000000000_0000100100110111_1111100000100100"; -- 0.03601027372899973
	pesos_i(15603) := b"0000000000000000_0000000000000000_0010010011101010_0101010101111001"; -- 0.14420065125887402
	pesos_i(15604) := b"0000000000000000_0000000000000000_0001001101100111_1000000010110011"; -- 0.0757980764509908
	pesos_i(15605) := b"1111111111111111_1111111111111111_1111010000111010_1001010111110011"; -- -0.045981052600011105
	pesos_i(15606) := b"0000000000000000_0000000000000000_0001110000110101_1011100011101011"; -- 0.11019473790053673
	pesos_i(15607) := b"1111111111111111_1111111111111111_1111010011000011_1011101110010100"; -- -0.04388835553398914
	pesos_i(15608) := b"1111111111111111_1111111111111111_1110000010110100_0011111010000000"; -- -0.12224969278086964
	pesos_i(15609) := b"0000000000000000_0000000000000000_0000001101111000_1010000110101001"; -- 0.01355944035353268
	pesos_i(15610) := b"0000000000000000_0000000000000000_0001111001111001_0001100101010011"; -- 0.1190353229746203
	pesos_i(15611) := b"1111111111111111_1111111111111111_1111101101010101_1101010001011001"; -- -0.01822159609321731
	pesos_i(15612) := b"1111111111111111_1111111111111111_1111000000000000_1011111000010000"; -- -0.06248867139776552
	pesos_i(15613) := b"1111111111111111_1111111111111111_1101110001011110_1110110000010001"; -- -0.13917660306041948
	pesos_i(15614) := b"1111111111111111_1111111111111111_1111000100010100_1110010101100101"; -- -0.058274901277019585
	pesos_i(15615) := b"1111111111111111_1111111111111111_1110101111001011_1011000111110111"; -- -0.07892310828423442
	pesos_i(15616) := b"0000000000000000_0000000000000000_0000110100010010_0011011010000011"; -- 0.051059157445195714
	pesos_i(15617) := b"0000000000000000_0000000000000000_0000101110010111_0010100110110110"; -- 0.04527531332025092
	pesos_i(15618) := b"1111111111111111_1111111111111111_1111001100000010_0001001011001110"; -- -0.050749611504672394
	pesos_i(15619) := b"1111111111111111_1111111111111111_1110011010000101_0111011010010101"; -- -0.09952601300831035
	pesos_i(15620) := b"0000000000000000_0000000000000000_0010000100100000_1101100101111100"; -- 0.12940749435161977
	pesos_i(15621) := b"1111111111111111_1111111111111111_1111001100001110_0101110111000110"; -- -0.050562037562933364
	pesos_i(15622) := b"1111111111111111_1111111111111111_1110111100111110_0001010111101110"; -- -0.0654588979668331
	pesos_i(15623) := b"0000000000000000_0000000000000000_0001110101000010_1011110111010011"; -- 0.11429964440622835
	pesos_i(15624) := b"0000000000000000_0000000000000000_0000110100111010_0000001101011110"; -- 0.05166646056336929
	pesos_i(15625) := b"1111111111111111_1111111111111111_1110000000110101_0101101100110101"; -- -0.12418584779764763
	pesos_i(15626) := b"1111111111111111_1111111111111111_1111110011111101_1001111101011011"; -- -0.01175502812477664
	pesos_i(15627) := b"0000000000000000_0000000000000000_0001100111110111_0111100010101110"; -- 0.10143236404213987
	pesos_i(15628) := b"0000000000000000_0000000000000000_0010000000101101_1101011000100101"; -- 0.12569940942641292
	pesos_i(15629) := b"1111111111111111_1111111111111111_1111111011000111_1000101110010111"; -- -0.004767680750420157
	pesos_i(15630) := b"1111111111111111_1111111111111111_1111011110000000_1101011111101011"; -- -0.03319025534330437
	pesos_i(15631) := b"1111111111111111_1111111111111111_1110101100011000_1001111010010000"; -- -0.08165558802382321
	pesos_i(15632) := b"1111111111111111_1111111111111111_1111010000001001_0000101100001000"; -- -0.046737013378207785
	pesos_i(15633) := b"1111111111111111_1111111111111111_1101011111010011_1110100001101111"; -- -0.1569227913906045
	pesos_i(15634) := b"1111111111111111_1111111111111111_1111000011101000_0011101010111011"; -- -0.05895646022408815
	pesos_i(15635) := b"1111111111111111_1111111111111111_1111000000110101_0010010011111000"; -- -0.0616890807470648
	pesos_i(15636) := b"1111111111111111_1111111111111111_1110111001001010_0100110011111001"; -- -0.06917876164989911
	pesos_i(15637) := b"1111111111111111_1111111111111111_1110001010101010_0000110001111110"; -- -0.11459276134139972
	pesos_i(15638) := b"1111111111111111_1111111111111111_1111000111110111_0110101100001001"; -- -0.05481844926505485
	pesos_i(15639) := b"0000000000000000_0000000000000000_0000001010100000_1100001110001001"; -- 0.01026556110350269
	pesos_i(15640) := b"1111111111111111_1111111111111111_1110001011010001_1010010000100101"; -- -0.11398862935861541
	pesos_i(15641) := b"1111111111111111_1111111111111111_1111000010010000_1001100110111001"; -- -0.060293571749948406
	pesos_i(15642) := b"0000000000000000_0000000000000000_0001000101111111_0101000100110000"; -- 0.06834895531628492
	pesos_i(15643) := b"0000000000000000_0000000000000000_0010001000001011_0011000001011100"; -- 0.13298322905779866
	pesos_i(15644) := b"0000000000000000_0000000000000000_0000011000011000_1010010000011101"; -- 0.02381349296435319
	pesos_i(15645) := b"0000000000000000_0000000000000000_0001101001000101_1100100011001111"; -- 0.10262732552287196
	pesos_i(15646) := b"1111111111111111_1111111111111111_1101110101101111_0100110000000110"; -- -0.13502049298046442
	pesos_i(15647) := b"0000000000000000_0000000000000000_0010011001010010_1000110011110001"; -- 0.14969712136821758
	pesos_i(15648) := b"0000000000000000_0000000000000000_0001010111110101_1100011001011111"; -- 0.08578147720411768
	pesos_i(15649) := b"1111111111111111_1111111111111111_1111110000001100_1011111010110110"; -- -0.015430527334304852
	pesos_i(15650) := b"0000000000000000_0000000000000000_0010010000011011_1111110000011000"; -- 0.1410520132302416
	pesos_i(15651) := b"0000000000000000_0000000000000000_0000001111111100_0110100001011100"; -- 0.01557018503413514
	pesos_i(15652) := b"0000000000000000_0000000000000000_0000111100010000_0001111010111011"; -- 0.05883972230513611
	pesos_i(15653) := b"1111111111111111_1111111111111111_1111011101001011_1100000111011010"; -- -0.03400028641123489
	pesos_i(15654) := b"0000000000000000_0000000000000000_0001010110111110_0101110111100111"; -- 0.08493601696470066
	pesos_i(15655) := b"1111111111111111_1111111111111111_1110110011100001_1100011101000001"; -- -0.07467989609954202
	pesos_i(15656) := b"1111111111111111_1111111111111111_1101100110000001_0101011101010111"; -- -0.1503701602650682
	pesos_i(15657) := b"0000000000000000_0000000000000000_0000001111011101_0011001111111001"; -- 0.01509404024538272
	pesos_i(15658) := b"1111111111111111_1111111111111111_1111010000111100_0101111111111101"; -- -0.04595375128057509
	pesos_i(15659) := b"0000000000000000_0000000000000000_0000000111100110_1101111010011010"; -- 0.007429039625966309
	pesos_i(15660) := b"1111111111111111_1111111111111111_1110110110010100_1111001110011100"; -- -0.07194592889543627
	pesos_i(15661) := b"1111111111111111_1111111111111111_1110101011100101_1010101111010011"; -- -0.08243299589949007
	pesos_i(15662) := b"1111111111111111_1111111111111111_1101111111101001_1111111100000010"; -- -0.12533575260930396
	pesos_i(15663) := b"1111111111111111_1111111111111111_1101101010011011_0100101110100001"; -- -0.14606787977032487
	pesos_i(15664) := b"0000000000000000_0000000000000000_0001000011011010_0110001010010011"; -- 0.0658322915059379
	pesos_i(15665) := b"0000000000000000_0000000000000000_0001010011000101_0100010100011011"; -- 0.08113510046905101
	pesos_i(15666) := b"1111111111111111_1111111111111111_1110100110010001_0110111000001100"; -- -0.08762466619740404
	pesos_i(15667) := b"0000000000000000_0000000000000000_0000111101001111_0000001011010000"; -- 0.05979936194670791
	pesos_i(15668) := b"0000000000000000_0000000000000000_0001100101010101_0000110001100001"; -- 0.0989539849870394
	pesos_i(15669) := b"1111111111111111_1111111111111111_1110101100110001_1100011111101111"; -- -0.08127165231927885
	pesos_i(15670) := b"1111111111111111_1111111111111111_1111101101110111_0111000001111101"; -- -0.017708749234492813
	pesos_i(15671) := b"1111111111111111_1111111111111111_1111110000100101_1111110100101011"; -- -0.015045334842264857
	pesos_i(15672) := b"0000000000000000_0000000000000000_0001100111111000_0111001000101110"; -- 0.10144723530745313
	pesos_i(15673) := b"0000000000000000_0000000000000000_0001000010011110_0000100111110010"; -- 0.06491148140921008
	pesos_i(15674) := b"1111111111111111_1111111111111111_1111110111011101_1000000111101000"; -- -0.008338814583062976
	pesos_i(15675) := b"1111111111111111_1111111111111111_1110100011110110_0101011001010111"; -- -0.08999119155837143
	pesos_i(15676) := b"1111111111111111_1111111111111111_1101100100011111_1110100100100001"; -- -0.15185683199371194
	pesos_i(15677) := b"0000000000000000_0000000000000000_0010000010110101_1001101100101000"; -- 0.12777108894144312
	pesos_i(15678) := b"0000000000000000_0000000000000000_0000001001010101_0101000000001111"; -- 0.00911426884646197
	pesos_i(15679) := b"0000000000000000_0000000000000000_0001001011101101_1100001010001101"; -- 0.07394042924575209
	pesos_i(15680) := b"0000000000000000_0000000000000000_0001101100010101_1100100011001110"; -- 0.10580115342063909
	pesos_i(15681) := b"0000000000000000_0000000000000000_0000010110011001_0000011100000101"; -- 0.021866263166433357
	pesos_i(15682) := b"0000000000000000_0000000000000000_0001011000110101_0010100110011011"; -- 0.0867486956459658
	pesos_i(15683) := b"0000000000000000_0000000000000000_0010001110010001_0110100011111110"; -- 0.13893753238077727
	pesos_i(15684) := b"0000000000000000_0000000000000000_0000111011111010_1001000010100001"; -- 0.05851081778450897
	pesos_i(15685) := b"0000000000000000_0000000000000000_0001011011010110_0111001101010000"; -- 0.08920975412741311
	pesos_i(15686) := b"1111111111111111_1111111111111111_1110110100000101_1011000010110001"; -- -0.0741319244660353
	pesos_i(15687) := b"1111111111111111_1111111111111111_1101110110100110_0111100000110011"; -- -0.13417862653103843
	pesos_i(15688) := b"1111111111111111_1111111111111111_1110000010100111_1101110001100100"; -- -0.12243864586980076
	pesos_i(15689) := b"0000000000000000_0000000000000000_0001100010110101_1001110011010011"; -- 0.09652118837465759
	pesos_i(15690) := b"1111111111111111_1111111111111111_1110111010001101_1010100011011001"; -- -0.06815094667579771
	pesos_i(15691) := b"0000000000000000_0000000000000000_0001001000010011_0101000010100000"; -- 0.07060722262649771
	pesos_i(15692) := b"0000000000000000_0000000000000000_0001101000101001_1100111000010001"; -- 0.10220039275628684
	pesos_i(15693) := b"1111111111111111_1111111111111111_1110011001010110_1001000011110110"; -- -0.10024160381970171
	pesos_i(15694) := b"0000000000000000_0000000000000000_0000001010101001_0100000100101110"; -- 0.010395120344168713
	pesos_i(15695) := b"0000000000000000_0000000000000000_0010001101110000_0010110111010111"; -- 0.13843046670564077
	pesos_i(15696) := b"0000000000000000_0000000000000000_0001010001001101_1010110111101001"; -- 0.07931029252081784
	pesos_i(15697) := b"0000000000000000_0000000000000000_0000000010110010_0101000101001111"; -- 0.0027209107469001194
	pesos_i(15698) := b"1111111111111111_1111111111111111_1110010010111100_0000000000001100"; -- -0.10650634475725339
	pesos_i(15699) := b"0000000000000000_0000000000000000_0000111001000111_1001101101001101"; -- 0.05578013059504499
	pesos_i(15700) := b"0000000000000000_0000000000000000_0001110100110110_1011111100011011"; -- 0.11411661526940944
	pesos_i(15701) := b"0000000000000000_0000000000000000_0000010100000100_0010100110000100"; -- 0.019594759599868665
	pesos_i(15702) := b"1111111111111111_1111111111111111_1101110011100101_1111011100011001"; -- -0.13711600907905516
	pesos_i(15703) := b"1111111111111111_1111111111111111_1111101100101101_0110110110100010"; -- -0.01883806978262989
	pesos_i(15704) := b"1111111111111111_1111111111111111_1110010111111100_1001110001001100"; -- -0.10161421914548767
	pesos_i(15705) := b"1111111111111111_1111111111111111_1110110101100011_0111110011001010"; -- -0.07270069176832378
	pesos_i(15706) := b"0000000000000000_0000000000000000_0001000111101110_1001010110011011"; -- 0.07004675898899665
	pesos_i(15707) := b"0000000000000000_0000000000000000_0001101010011101_1011001100011011"; -- 0.1039688054263811
	pesos_i(15708) := b"0000000000000000_0000000000000000_0010010010101011_0000111001010111"; -- 0.14323510773055737
	pesos_i(15709) := b"1111111111111111_1111111111111111_1101110101000110_1101011001100000"; -- -0.13563785701224088
	pesos_i(15710) := b"0000000000000000_0000000000000000_0000010101111010_0101100001100100"; -- 0.02139809064826673
	pesos_i(15711) := b"1111111111111111_1111111111111111_1110101111110100_0110100110011001"; -- -0.07830181134432994
	pesos_i(15712) := b"0000000000000000_0000000000000000_0000100011111001_1001101111000011"; -- 0.035058722667360424
	pesos_i(15713) := b"0000000000000000_0000000000000000_0001011111010011_0110110011111011"; -- 0.09306985025459336
	pesos_i(15714) := b"1111111111111111_1111111111111111_1110001001010000_1010010000001000"; -- -0.11595701975169011
	pesos_i(15715) := b"0000000000000000_0000000000000000_0001011001010010_1000010111100110"; -- 0.08719670164345251
	pesos_i(15716) := b"1111111111111111_1111111111111111_1110100110100001_0011110100101001"; -- -0.08738343948447654
	pesos_i(15717) := b"1111111111111111_1111111111111111_1111010110000100_0000101010001010"; -- -0.04095396158700838
	pesos_i(15718) := b"1111111111111111_1111111111111111_1110110101000101_1110010011000000"; -- -0.07315225891191485
	pesos_i(15719) := b"1111111111111111_1111111111111111_1110101100011110_1011100100000001"; -- -0.08156245923742753
	pesos_i(15720) := b"0000000000000000_0000000000000000_0001010101000111_0011010001101101"; -- 0.08311774892767429
	pesos_i(15721) := b"0000000000000000_0000000000000000_0000101001001011_0001101110001101"; -- 0.040208551337365096
	pesos_i(15722) := b"1111111111111111_1111111111111111_1111110111010110_1111011001101000"; -- -0.00843868212580374
	pesos_i(15723) := b"1111111111111111_1111111111111111_1110100100101111_0011101001100101"; -- -0.08912310630306033
	pesos_i(15724) := b"0000000000000000_0000000000000000_0000101010100001_1010111111000110"; -- 0.041529642015080345
	pesos_i(15725) := b"1111111111111111_1111111111111111_1111010011110000_0010110101011011"; -- -0.04321018727022053
	pesos_i(15726) := b"0000000000000000_0000000000000000_0000111100000110_1000101101100111"; -- 0.05869361167139842
	pesos_i(15727) := b"1111111111111111_1111111111111111_1111010010100011_1100111101100010"; -- -0.044375456511579585
	pesos_i(15728) := b"0000000000000000_0000000000000000_0001111000100001_1110001111011000"; -- 0.1177046206284123
	pesos_i(15729) := b"1111111111111111_1111111111111111_1101111110000110_0010001000110111"; -- -0.12685953284028342
	pesos_i(15730) := b"0000000000000000_0000000000000000_0000111101001110_1010010001110011"; -- 0.059793737486276956
	pesos_i(15731) := b"0000000000000000_0000000000000000_0000101100000110_0110001010101010"; -- 0.04306618350595566
	pesos_i(15732) := b"1111111111111111_1111111111111111_1111110001000000_1110101001010011"; -- -0.014634470652505224
	pesos_i(15733) := b"1111111111111111_1111111111111111_1101011101011110_1011101000110000"; -- -0.1587108261301081
	pesos_i(15734) := b"0000000000000000_0000000000000000_0001101011110000_0110100011111011"; -- 0.10523086678529202
	pesos_i(15735) := b"1111111111111111_1111111111111111_1110100110001110_0101001100101001"; -- -0.08767204511483515
	pesos_i(15736) := b"1111111111111111_1111111111111111_1110101010111010_1010101000000000"; -- -0.08308923250350932
	pesos_i(15737) := b"1111111111111111_1111111111111111_1111100001110111_1111111111011110"; -- -0.0294189532833627
	pesos_i(15738) := b"1111111111111111_1111111111111111_1101101100100000_1100101101010110"; -- -0.14403084894205728
	pesos_i(15739) := b"0000000000000000_0000000000000000_0001010110101110_1001000110010001"; -- 0.08469495584166264
	pesos_i(15740) := b"0000000000000000_0000000000000000_0001010001110000_0000110011100111"; -- 0.07983475340406737
	pesos_i(15741) := b"0000000000000000_0000000000000000_0000001110010110_1000001011001100"; -- 0.014015364457596708
	pesos_i(15742) := b"0000000000000000_0000000000000000_0010011001111010_1101100010100001"; -- 0.1503119842778029
	pesos_i(15743) := b"1111111111111111_1111111111111111_1110011110101111_1100011011101001"; -- -0.09497410592402936
	pesos_i(15744) := b"1111111111111111_1111111111111111_1110101110001000_1111001100100110"; -- -0.07994156179944328
	pesos_i(15745) := b"0000000000000000_0000000000000000_0001111001110011_1011010000011110"; -- 0.11895299654061314
	pesos_i(15746) := b"0000000000000000_0000000000000000_0000111111110110_1111001111001011"; -- 0.06236194330666338
	pesos_i(15747) := b"0000000000000000_0000000000000000_0000011100010101_0000001101100000"; -- 0.027664385702911333
	pesos_i(15748) := b"0000000000000000_0000000000000000_0000110110110011_0100110001000110"; -- 0.05351711957017938
	pesos_i(15749) := b"1111111111111111_1111111111111111_1111110000000110_1001010010010011"; -- -0.015524591478153093
	pesos_i(15750) := b"0000000000000000_0000000000000000_0001110010011100_0111101011000100"; -- 0.11176268855245207
	pesos_i(15751) := b"1111111111111111_1111111111111111_1111001101001100_0100001000010110"; -- -0.04961764294182034
	pesos_i(15752) := b"1111111111111111_1111111111111111_1110100001010011_1000000000111001"; -- -0.09247587773717715
	pesos_i(15753) := b"1111111111111111_1111111111111111_1101100110010110_1000111010011011"; -- -0.15004643167215453
	pesos_i(15754) := b"0000000000000000_0000000000000000_0010000111010010_0010010011110010"; -- 0.13211279773453652
	pesos_i(15755) := b"1111111111111111_1111111111111111_1110001100011010_0010011110101100"; -- -0.112882156893593
	pesos_i(15756) := b"1111111111111111_1111111111111111_1110101110101000_0101110101011101"; -- -0.0794622086399381
	pesos_i(15757) := b"1111111111111111_1111111111111111_1111011111000010_1101011011110011"; -- -0.032183232926017824
	pesos_i(15758) := b"0000000000000000_0000000000000000_0001110000001101_1010100000010010"; -- 0.10958338211093976
	pesos_i(15759) := b"0000000000000000_0000000000000000_0000100001011000_1001101001110010"; -- 0.032601979076207044
	pesos_i(15760) := b"0000000000000000_0000000000000000_0000000111110001_0111111100011000"; -- 0.007591193646550365
	pesos_i(15761) := b"0000000000000000_0000000000000000_0000110111001101_0000101000110110"; -- 0.05390991027600597
	pesos_i(15762) := b"0000000000000000_0000000000000000_0001000111001000_1100110100001011"; -- 0.0694702292114
	pesos_i(15763) := b"0000000000000000_0000000000000000_0000011010101101_1101011001011010"; -- 0.0260900467898956
	pesos_i(15764) := b"1111111111111111_1111111111111111_1101100100110000_1101110111010100"; -- -0.15159810611565744
	pesos_i(15765) := b"0000000000000000_0000000000000000_0000111110001111_1111111110010010"; -- 0.060790990114249266
	pesos_i(15766) := b"1111111111111111_1111111111111111_1110110000101101_1100000101000101"; -- -0.07742683480489135
	pesos_i(15767) := b"1111111111111111_1111111111111111_1110010100100000_1010010011001000"; -- -0.10497064710207539
	pesos_i(15768) := b"0000000000000000_0000000000000000_0001001010101001_1100010110011110"; -- 0.0729030143673837
	pesos_i(15769) := b"1111111111111111_1111111111111111_1110100100101000_1001110110110001"; -- -0.08922399934368859
	pesos_i(15770) := b"1111111111111111_1111111111111111_1110110000111110_0110000010000001"; -- -0.07717320289421914
	pesos_i(15771) := b"0000000000000000_0000000000000000_0001000101111110_1101100110110100"; -- 0.06834183352842514
	pesos_i(15772) := b"0000000000000000_0000000000000000_0010000110010100_1111010100011111"; -- 0.13117916117806847
	pesos_i(15773) := b"0000000000000000_0000000000000000_0001001000000001_1011100000111110"; -- 0.07033874038512555
	pesos_i(15774) := b"1111111111111111_1111111111111111_1110101101100110_1101001111101001"; -- -0.0804622227675707
	pesos_i(15775) := b"1111111111111111_1111111111111111_1110101011100111_0111101001000000"; -- -0.08240543310759012
	pesos_i(15776) := b"0000000000000000_0000000000000000_0010010001010011_0101101110100001"; -- 0.14189694093725358
	pesos_i(15777) := b"0000000000000000_0000000000000000_0001001100101001_0110010000110000"; -- 0.07485033191627503
	pesos_i(15778) := b"1111111111111111_1111111111111111_1111010111010000_1101111100000011"; -- -0.03978162930908356
	pesos_i(15779) := b"1111111111111111_1111111111111111_1111010101010100_0011000001010010"; -- -0.041684131580190076
	pesos_i(15780) := b"0000000000000000_0000000000000000_0001111000101010_0101111001110001"; -- 0.1178339983792856
	pesos_i(15781) := b"0000000000000000_0000000000000000_0010000000101100_0110101000011011"; -- 0.12567771109845058
	pesos_i(15782) := b"1111111111111111_1111111111111111_1110001001001010_0011110100001111"; -- -0.11605471021789275
	pesos_i(15783) := b"0000000000000000_0000000000000000_0000110010011000_0100001110101100"; -- 0.04919836955438773
	pesos_i(15784) := b"1111111111111111_1111111111111111_1101111100001000_1011011111010101"; -- -0.12877322241709546
	pesos_i(15785) := b"0000000000000000_0000000000000000_0001110110010000_0111101000011110"; -- 0.11548579440374894
	pesos_i(15786) := b"0000000000000000_0000000000000000_0001110010110111_0110011101101011"; -- 0.11217352247840166
	pesos_i(15787) := b"0000000000000000_0000000000000000_0000001000001101_1001001110010100"; -- 0.008019660701257633
	pesos_i(15788) := b"0000000000000000_0000000000000000_0010011010000011_0101010011100010"; -- 0.15044146073220555
	pesos_i(15789) := b"0000000000000000_0000000000000000_0001011110011110_1101010111000100"; -- 0.09226738002311875
	pesos_i(15790) := b"0000000000000000_0000000000000000_0001100001000010_1001010011001100"; -- 0.09476594906322967
	pesos_i(15791) := b"1111111111111111_1111111111111111_1110101010000100_0000111011110100"; -- -0.083922448493496
	pesos_i(15792) := b"1111111111111111_1111111111111111_1111001111110011_0001111101001001"; -- -0.04707149949891621
	pesos_i(15793) := b"0000000000000000_0000000000000000_0001111010110110_1001010101100011"; -- 0.11997350371471337
	pesos_i(15794) := b"1111111111111111_1111111111111111_1111001110110101_1010001011110000"; -- -0.0480096972765649
	pesos_i(15795) := b"1111111111111111_1111111111111111_1101110000100010_0110000110011100"; -- -0.14010038313540052
	pesos_i(15796) := b"0000000000000000_0000000000000000_0001010011110101_1001010111110111"; -- 0.08187234185466367
	pesos_i(15797) := b"0000000000000000_0000000000000000_0000000100010011_1101001100001010"; -- 0.004208745975791252
	pesos_i(15798) := b"1111111111111111_1111111111111111_1101111001000101_0000011111011100"; -- -0.1317591751167544
	pesos_i(15799) := b"1111111111111111_1111111111111111_1110010001011010_1101110111101101"; -- -0.10798848117083851
	pesos_i(15800) := b"0000000000000000_0000000000000000_0001011111011100_1111111100100000"; -- 0.09321589013022794
	pesos_i(15801) := b"0000000000000000_0000000000000000_0010001011101011_0100001101111111"; -- 0.13640233846616207
	pesos_i(15802) := b"0000000000000000_0000000000000000_0000001100110111_1001100100010010"; -- 0.012567107097617833
	pesos_i(15803) := b"1111111111111111_1111111111111111_1110000000011101_1001011001001000"; -- -0.12454853757514954
	pesos_i(15804) := b"0000000000000000_0000000000000000_0000011000101100_1110111110000100"; -- 0.024123163056561835
	pesos_i(15805) := b"0000000000000000_0000000000000000_0000001001101010_1111010001011101"; -- 0.009444496777728625
	pesos_i(15806) := b"1111111111111111_1111111111111111_1110111000100111_1110101100001100"; -- -0.06970339727711035
	pesos_i(15807) := b"1111111111111111_1111111111111111_1110011010010001_1101110110111010"; -- -0.09933675972399272
	pesos_i(15808) := b"0000000000000000_0000000000000000_0001001010011100_1101011100101001"; -- 0.07270569572926495
	pesos_i(15809) := b"0000000000000000_0000000000000000_0010001011110110_1000101111110010"; -- 0.13657450339002317
	pesos_i(15810) := b"0000000000000000_0000000000000000_0001110110101000_1010110010001100"; -- 0.11585501109247398
	pesos_i(15811) := b"1111111111111111_1111111111111111_1110100011100010_0010010000001110"; -- -0.09029936469768844
	pesos_i(15812) := b"1111111111111111_1111111111111111_1110000100010011_0101101011100000"; -- -0.12079841633345312
	pesos_i(15813) := b"1111111111111111_1111111111111111_1110100111111100_1101111010011001"; -- -0.08598526720163151
	pesos_i(15814) := b"1111111111111111_1111111111111111_1110110101101000_0000101111000001"; -- -0.07263113534665203
	pesos_i(15815) := b"1111111111111111_1111111111111111_1110111110010010_0001011011011000"; -- -0.064177105264052
	pesos_i(15816) := b"1111111111111111_1111111111111111_1110011111110101_0111001011101110"; -- -0.0939109964280735
	pesos_i(15817) := b"1111111111111111_1111111111111111_1110011000001100_1111100001101111"; -- -0.1013645866790313
	pesos_i(15818) := b"1111111111111111_1111111111111111_1110101011011011_0110011100010111"; -- -0.08258968064504957
	pesos_i(15819) := b"0000000000000000_0000000000000000_0001001111001111_1100010100100101"; -- 0.0773890701021509
	pesos_i(15820) := b"1111111111111111_1111111111111111_1101101100111010_1010010110111100"; -- -0.14363636168379745
	pesos_i(15821) := b"1111111111111111_1111111111111111_1110100010000011_0101100001001111"; -- -0.0917458349264082
	pesos_i(15822) := b"0000000000000000_0000000000000000_0000111011101110_1110110110101101"; -- 0.058333258330700764
	pesos_i(15823) := b"1111111111111111_1111111111111111_1110111001001100_0001101111110101"; -- -0.0691511657637018
	pesos_i(15824) := b"0000000000000000_0000000000000000_0000000000011101_0000001101100000"; -- 0.0004427060028765929
	pesos_i(15825) := b"0000000000000000_0000000000000000_0000011010100000_1101111101010001"; -- 0.025892216926747466
	pesos_i(15826) := b"0000000000000000_0000000000000000_0001000110111010_0111111111111001"; -- 0.06925201250940359
	pesos_i(15827) := b"1111111111111111_1111111111111111_1111001001110000_1000110110111110"; -- -0.05297006710831322
	pesos_i(15828) := b"1111111111111111_1111111111111111_1110100010000100_0101110111000101"; -- -0.09173025080433148
	pesos_i(15829) := b"1111111111111111_1111111111111111_1110100110010011_1101100000110001"; -- -0.08758782201209693
	pesos_i(15830) := b"0000000000000000_0000000000000000_0001110111001011_1001001111100101"; -- 0.11638759926793313
	pesos_i(15831) := b"1111111111111111_1111111111111111_1110101001011011_0010100110100011"; -- -0.08454646841166766
	pesos_i(15832) := b"0000000000000000_0000000000000000_0000111000111000_0010011111110100"; -- 0.055544373514179145
	pesos_i(15833) := b"1111111111111111_1111111111111111_1101110111111100_1000110001101111"; -- -0.13286516470599402
	pesos_i(15834) := b"0000000000000000_0000000000000000_0001111100001100_1111111001110100"; -- 0.1212920220622233
	pesos_i(15835) := b"0000000000000000_0000000000000000_0001110000100100_1100101001000101"; -- 0.10993637270206198
	pesos_i(15836) := b"0000000000000000_0000000000000000_0000110001011001_0100110000000011"; -- 0.04823756298436288
	pesos_i(15837) := b"0000000000000000_0000000000000000_0000110101101011_1111100011110111"; -- 0.05242878000647839
	pesos_i(15838) := b"0000000000000000_0000000000000000_0010000111011110_0000000010101111"; -- 0.132293741976149
	pesos_i(15839) := b"1111111111111111_1111111111111111_1101011010001111_0111111111111110"; -- -0.16187286422447436
	pesos_i(15840) := b"1111111111111111_1111111111111111_1110111011010000_0110001110100101"; -- -0.06713273271212722
	pesos_i(15841) := b"1111111111111111_1111111111111111_1111110000001111_1100011001111011"; -- -0.0153842877100147
	pesos_i(15842) := b"0000000000000000_0000000000000000_0001000001100011_1010111100100101"; -- 0.06402105957695396
	pesos_i(15843) := b"1111111111111111_1111111111111111_1111111110101110_1000000100000010"; -- -0.0012435311343774963
	pesos_i(15844) := b"0000000000000000_0000000000000000_0000101000000000_1101010001000010"; -- 0.039075151622373454
	pesos_i(15845) := b"0000000000000000_0000000000000000_0010010110110001_1011011001110100"; -- 0.14724293073940944
	pesos_i(15846) := b"0000000000000000_0000000000000000_0010101000101010_1001001110101010"; -- 0.16471217071130212
	pesos_i(15847) := b"1111111111111111_1111111111111111_1101011100101010_1100001001011101"; -- -0.15950379580349042
	pesos_i(15848) := b"0000000000000000_0000000000000000_0001000110011100_1011010010010011"; -- 0.06879738414669566
	pesos_i(15849) := b"1111111111111111_1111111111111111_1110101101000110_1101110001100100"; -- -0.08094999844315373
	pesos_i(15850) := b"0000000000000000_0000000000000000_0010000101111111_0111001000011011"; -- 0.13085091732196055
	pesos_i(15851) := b"0000000000000000_0000000000000000_0001101010000010_0010101010010111"; -- 0.10354868113141368
	pesos_i(15852) := b"0000000000000000_0000000000000000_0000011101101001_1001001001110100"; -- 0.028954652229312164
	pesos_i(15853) := b"0000000000000000_0000000000000000_0000011010101101_1010011110101111"; -- 0.026087265246552808
	pesos_i(15854) := b"1111111111111111_1111111111111111_1101111110110010_0111111101100001"; -- -0.12618259305718754
	pesos_i(15855) := b"0000000000000000_0000000000000000_0001110100101101_0001100010000100"; -- 0.11396935669713586
	pesos_i(15856) := b"1111111111111111_1111111111111111_1111110101000110_0010110011011101"; -- -0.010647960707782478
	pesos_i(15857) := b"1111111111111111_1111111111111111_1110110100101110_1110110000101001"; -- -0.07350276951845582
	pesos_i(15858) := b"0000000000000000_0000000000000000_0001011011000001_1110111011111001"; -- 0.08889669023604804
	pesos_i(15859) := b"1111111111111111_1111111111111111_1111000111101000_1001000011001010"; -- -0.05504508089032463
	pesos_i(15860) := b"1111111111111111_1111111111111111_1111110001101000_0100111010110110"; -- -0.014033394436524028
	pesos_i(15861) := b"1111111111111111_1111111111111111_1111110011101100_0110001111100111"; -- -0.012017971242800319
	pesos_i(15862) := b"1111111111111111_1111111111111111_1110001011000000_0111101000100101"; -- -0.1142505321230199
	pesos_i(15863) := b"1111111111111111_1111111111111111_1111110101011101_1101111101111100"; -- -0.010286361980708182
	pesos_i(15864) := b"0000000000000000_0000000000000000_0001000111000010_1111000010001101"; -- 0.0693807930128672
	pesos_i(15865) := b"0000000000000000_0000000000000000_0000111100100100_1100111010111111"; -- 0.05915538940246003
	pesos_i(15866) := b"0000000000000000_0000000000000000_0001111011100110_1110011010111010"; -- 0.12071077386289539
	pesos_i(15867) := b"1111111111111111_1111111111111111_1110111111001101_1100010110000001"; -- -0.06326642597832173
	pesos_i(15868) := b"1111111111111111_1111111111111111_1111011000011100_1111010001110011"; -- -0.03862068368207226
	pesos_i(15869) := b"1111111111111111_1111111111111111_1110011011100100_1000010001100011"; -- -0.09807560521773019
	pesos_i(15870) := b"1111111111111111_1111111111111111_1111100110110100_0110111111000110"; -- -0.02459050573947326
	pesos_i(15871) := b"0000000000000000_0000000000000000_0001000110100001_1010001110110010"; -- 0.06887267197342375
	pesos_i(15872) := b"1111111111111111_1111111111111111_1101110101011100_0100000101100110"; -- -0.1353110434097423
	pesos_i(15873) := b"0000000000000000_0000000000000000_0000111111000110_0100011100110100"; -- 0.06161923416095
	pesos_i(15874) := b"0000000000000000_0000000000000000_0000111011111110_1110010000001101"; -- 0.05857682540303246
	pesos_i(15875) := b"0000000000000000_0000000000000000_0001111000000001_0110111101101110"; -- 0.11720940050282933
	pesos_i(15876) := b"0000000000000000_0000000000000000_0010011011001000_1001000010100001"; -- 0.15149787841987736
	pesos_i(15877) := b"0000000000000000_0000000000000000_0001011101101011_0010011010010110"; -- 0.09147874039343205
	pesos_i(15878) := b"0000000000000000_0000000000000000_0000110110001110_1111000101011111"; -- 0.052962384933843254
	pesos_i(15879) := b"1111111111111111_1111111111111111_1111110111111100_0000110101011000"; -- -0.007872739799122732
	pesos_i(15880) := b"1111111111111111_1111111111111111_1101111101011101_1100101001011111"; -- -0.1274751202819827
	pesos_i(15881) := b"1111111111111111_1111111111111111_1101101000100010_0001101110001100"; -- -0.14791705916597686
	pesos_i(15882) := b"0000000000000000_0000000000000000_0000001100000000_1101110010010010"; -- 0.011731897085265817
	pesos_i(15883) := b"1111111111111111_1111111111111111_1110001101010000_0100011011000001"; -- -0.11205632952137852
	pesos_i(15884) := b"0000000000000000_0000000000000000_0000011010100111_0011111101110000"; -- 0.02598949897535796
	pesos_i(15885) := b"1111111111111111_1111111111111111_1101111110001101_0011101101101001"; -- -0.1267512195306099
	pesos_i(15886) := b"1111111111111111_1111111111111111_1110001000011111_0111110010110101"; -- -0.11670704441025713
	pesos_i(15887) := b"0000000000000000_0000000000000000_0000100110010101_1101110110001001"; -- 0.03744301414476058
	pesos_i(15888) := b"0000000000000000_0000000000000000_0000101111000100_0000111101011100"; -- 0.04596038816318909
	pesos_i(15889) := b"1111111111111111_1111111111111111_1111000101001000_1000100011110001"; -- -0.05748695483963528
	pesos_i(15890) := b"1111111111111111_1111111111111111_1101101111011111_0110101101100001"; -- -0.1411221398400923
	pesos_i(15891) := b"1111111111111111_1111111111111111_1111110101110010_0100011010110101"; -- -0.009975033511606148
	pesos_i(15892) := b"0000000000000000_0000000000000000_0001100010101011_1111111000100001"; -- 0.09637440023582823
	pesos_i(15893) := b"1111111111111111_1111111111111111_1110000011111100_1000001000000001"; -- -0.12114703631635187
	pesos_i(15894) := b"1111111111111111_1111111111111111_1111001010111110_0101111000111011"; -- -0.05178271341827129
	pesos_i(15895) := b"1111111111111111_1111111111111111_1111010011010011_0010100101011001"; -- -0.043652931000742225
	pesos_i(15896) := b"0000000000000000_0000000000000000_0000111000101101_0100000001101010"; -- 0.0553779847964151
	pesos_i(15897) := b"0000000000000000_0000000000000000_0001000011010110_1101011001101101"; -- 0.06577816152014641
	pesos_i(15898) := b"1111111111111111_1111111111111111_1101111100101000_1101111110111000"; -- -0.1282825638020775
	pesos_i(15899) := b"1111111111111111_1111111111111111_1110001011000011_0000101101111000"; -- -0.11421135264707673
	pesos_i(15900) := b"1111111111111111_1111111111111111_1111010111111010_1011111001011100"; -- -0.03914270638894924
	pesos_i(15901) := b"0000000000000000_0000000000000000_0001111111010101_0111110100000011"; -- 0.1243513233541209
	pesos_i(15902) := b"0000000000000000_0000000000000000_0001111001111110_1010011111000001"; -- 0.11912010630596598
	pesos_i(15903) := b"0000000000000000_0000000000000000_0010011111010001_0100010111111001"; -- 0.15553700751749971
	pesos_i(15904) := b"1111111111111111_1111111111111111_1101100110001111_1001100001100110"; -- -0.15015265949037665
	pesos_i(15905) := b"1111111111111111_1111111111111111_1110100110000010_1001110000011100"; -- -0.08785080257023473
	pesos_i(15906) := b"0000000000000000_0000000000000000_0000100011011011_1011110111111011"; -- 0.03460299856193635
	pesos_i(15907) := b"0000000000000000_0000000000000000_0000100110001111_0011101010110100"; -- 0.03734175586835735
	pesos_i(15908) := b"1111111111111111_1111111111111111_1111000111001010_1010011101011000"; -- -0.055501500097151414
	pesos_i(15909) := b"1111111111111111_1111111111111111_1101110010101111_1001100100110110"; -- -0.13794557971900162
	pesos_i(15910) := b"1111111111111111_1111111111111111_1111010011001011_0000111001011101"; -- -0.043776609700295926
	pesos_i(15911) := b"1111111111111111_1111111111111111_1110010001110110_1110000001010010"; -- -0.10756109227774752
	pesos_i(15912) := b"1111111111111111_1111111111111111_1110001101100011_1010011101100010"; -- -0.11176065298593364
	pesos_i(15913) := b"1111111111111111_1111111111111111_1111011010010001_0000101101010011"; -- -0.03684930070724672
	pesos_i(15914) := b"0000000000000000_0000000000000000_0001010111010000_1100001010111101"; -- 0.08521668550875103
	pesos_i(15915) := b"0000000000000000_0000000000000000_0010001011110110_0100011110011101"; -- 0.13657043053104362
	pesos_i(15916) := b"0000000000000000_0000000000000000_0001111010011110_0010011100001001"; -- 0.11960071526692648
	pesos_i(15917) := b"1111111111111111_1111111111111111_1111000000100100_1110001000011010"; -- -0.06193720686944071
	pesos_i(15918) := b"0000000000000000_0000000000000000_0010010100100101_1101100111110111"; -- 0.1451088169958191
	pesos_i(15919) := b"1111111111111111_1111111111111111_1110111101010010_1110111010000100"; -- -0.06514081256204013
	pesos_i(15920) := b"1111111111111111_1111111111111111_1110000101010011_0111001111000010"; -- -0.11982037088646126
	pesos_i(15921) := b"0000000000000000_0000000000000000_0001110000001101_1101100000010110"; -- 0.1095862439301492
	pesos_i(15922) := b"1111111111111111_1111111111111111_1111110001110001_1001010010010010"; -- -0.01389190125959203
	pesos_i(15923) := b"0000000000000000_0000000000000000_0010001101111110_1011101001011100"; -- 0.138652465390284
	pesos_i(15924) := b"1111111111111111_1111111111111111_1110110101100001_0010010101010101"; -- -0.0727364223305945
	pesos_i(15925) := b"0000000000000000_0000000000000000_0000110010001110_0111110110111011"; -- 0.049049242196556125
	pesos_i(15926) := b"1111111111111111_1111111111111111_1110010000111110_1001111110111110"; -- -0.10841943381724567
	pesos_i(15927) := b"1111111111111111_1111111111111111_1110000011110001_1010101110000001"; -- -0.12131240946433505
	pesos_i(15928) := b"1111111111111111_1111111111111111_1111101100101110_0010111110010010"; -- -0.018826510363941198
	pesos_i(15929) := b"0000000000000000_0000000000000000_0000111010010101_0000101110101110"; -- 0.05696175572680586
	pesos_i(15930) := b"1111111111111111_1111111111111111_1111000101000010_1100010001111100"; -- -0.05757495855712455
	pesos_i(15931) := b"1111111111111111_1111111111111111_1101111010100100_1011100010010001"; -- -0.1302990575225926
	pesos_i(15932) := b"1111111111111111_1111111111111111_1111001101100101_1111101011010011"; -- -0.049225161936870834
	pesos_i(15933) := b"0000000000000000_0000000000000000_0000111011011001_1001000111010010"; -- 0.058007348696098686
	pesos_i(15934) := b"1111111111111111_1111111111111111_1111010001001110_0010111011100011"; -- -0.0456820197031719
	pesos_i(15935) := b"1111111111111111_1111111111111111_1111000110100110_0101100001110111"; -- -0.056055518137393685
	pesos_i(15936) := b"0000000000000000_0000000000000000_0001101101101101_0111101001101000"; -- 0.10713925401228522
	pesos_i(15937) := b"1111111111111111_1111111111111111_1111001010000011_0011010100001001"; -- -0.052685437465315274
	pesos_i(15938) := b"0000000000000000_0000000000000000_0000111010001100_0101110110000111"; -- 0.056829305137030425
	pesos_i(15939) := b"0000000000000000_0000000000000000_0000101001100001_0001000010001000"; -- 0.04054358795584703
	pesos_i(15940) := b"1111111111111111_1111111111111111_1110111111010010_1010000110110101"; -- -0.06319226588310618
	pesos_i(15941) := b"1111111111111111_1111111111111111_1101101111010000_1111100100001100"; -- -0.1413425774895411
	pesos_i(15942) := b"0000000000000000_0000000000000000_0000101101001001_1000000110010000"; -- 0.04409036413999396
	pesos_i(15943) := b"1111111111111111_1111111111111111_1111101000101111_0101001011101110"; -- -0.02271539384663192
	pesos_i(15944) := b"1111111111111111_1111111111111111_1110100101100000_0001110001010011"; -- -0.08837721804310847
	pesos_i(15945) := b"1111111111111111_1111111111111111_1110100110110001_1000011101001100"; -- -0.08713487992032173
	pesos_i(15946) := b"1111111111111111_1111111111111111_1110000010101100_0100010001100010"; -- -0.12237141224101007
	pesos_i(15947) := b"1111111111111111_1111111111111111_1110010000111100_1111101001111100"; -- -0.10844454255636146
	pesos_i(15948) := b"0000000000000000_0000000000000000_0010001001110011_1010101110101010"; -- 0.1345774928024886
	pesos_i(15949) := b"1111111111111111_1111111111111111_1111111101110111_1000001011000111"; -- -0.0020826592482719487
	pesos_i(15950) := b"1111111111111111_1111111111111111_1110101110001110_0110100100010111"; -- -0.0798582381137631
	pesos_i(15951) := b"0000000000000000_0000000000000000_0000010101000101_0100000010010110"; -- 0.0205879559608054
	pesos_i(15952) := b"0000000000000000_0000000000000000_0001100100101111_0110101110000110"; -- 0.0983798220236217
	pesos_i(15953) := b"1111111111111111_1111111111111111_1110101101110110_0111110011110011"; -- -0.0802232653084179
	pesos_i(15954) := b"0000000000000000_0000000000000000_0001110101001110_1000001110100010"; -- 0.11447928142195007
	pesos_i(15955) := b"0000000000000000_0000000000000000_0000110011101100_0110011111101011"; -- 0.05048226823868917
	pesos_i(15956) := b"0000000000000000_0000000000000000_0000000111010010_0100010100101010"; -- 0.0071147182388358425
	pesos_i(15957) := b"0000000000000000_0000000000000000_0000001110011111_1010101111011001"; -- 0.014155140325450098
	pesos_i(15958) := b"1111111111111111_1111111111111111_1101111011101000_1111001011001000"; -- -0.12925799012205264
	pesos_i(15959) := b"0000000000000000_0000000000000000_0000001100100110_0100111110001010"; -- 0.012303324838249342
	pesos_i(15960) := b"1111111111111111_1111111111111111_1111000010010010_1111110100110111"; -- -0.06025712390514212
	pesos_i(15961) := b"1111111111111111_1111111111111111_1111111011100110_1001000111011111"; -- -0.004294283849156374
	pesos_i(15962) := b"1111111111111111_1111111111111111_1101101010010100_0011000010001011"; -- -0.14617630582046517
	pesos_i(15963) := b"0000000000000000_0000000000000000_0000110000011001_0001001000110010"; -- 0.04725755430077865
	pesos_i(15964) := b"0000000000000000_0000000000000000_0001101001110100_0110100110000101"; -- 0.10333880906291612
	pesos_i(15965) := b"1111111111111111_1111111111111111_1110000100100000_0000110110010101"; -- -0.12060465930910089
	pesos_i(15966) := b"0000000000000000_0000000000000000_0010010000100101_0010000110110110"; -- 0.14119158441062196
	pesos_i(15967) := b"0000000000000000_0000000000000000_0001011010110101_1001011101100111"; -- 0.08870836517657585
	pesos_i(15968) := b"0000000000000000_0000000000000000_0000110100010011_1110011111100010"; -- 0.051084988366221835
	pesos_i(15969) := b"1111111111111111_1111111111111111_1111010110100010_0101010001110000"; -- -0.040491793403273454
	pesos_i(15970) := b"0000000000000000_0000000000000000_0000111101001001_1111001111100111"; -- 0.059722179358939885
	pesos_i(15971) := b"0000000000000000_0000000000000000_0000110100111000_0010111011101000"; -- 0.051638537924001686
	pesos_i(15972) := b"0000000000000000_0000000000000000_0001110110101100_1010000101000010"; -- 0.11591537352963631
	pesos_i(15973) := b"0000000000000000_0000000000000000_0000010110110011_0111110011111001"; -- 0.02227002220573458
	pesos_i(15974) := b"0000000000000000_0000000000000000_0000010111101011_0000100110000110"; -- 0.0231176331560737
	pesos_i(15975) := b"0000000000000000_0000000000000000_0001111101100000_0010111100011010"; -- 0.12256140121638967
	pesos_i(15976) := b"0000000000000000_0000000000000000_0010010010001111_0011111100101101"; -- 0.14281077241419896
	pesos_i(15977) := b"1111111111111111_1111111111111111_1101110010100111_0011100100111100"; -- -0.13807337079284965
	pesos_i(15978) := b"0000000000000000_0000000000000000_0000001101000100_1100011001001100"; -- 0.012768167112266799
	pesos_i(15979) := b"0000000000000000_0000000000000000_0000100110100011_0110010100100100"; -- 0.037649460977789886
	pesos_i(15980) := b"1111111111111111_1111111111111111_1110101111001011_0100000110101010"; -- -0.07892980184367612
	pesos_i(15981) := b"0000000000000000_0000000000000000_0010011000011100_0111100100010010"; -- 0.1488719623990634
	pesos_i(15982) := b"0000000000000000_0000000000000000_0000001111101110_1110010001010010"; -- 0.015363950707555118
	pesos_i(15983) := b"1111111111111111_1111111111111111_1110010010011101_1111101000111111"; -- -0.1069644542119621
	pesos_i(15984) := b"1111111111111111_1111111111111111_1111001010110100_0000100011111011"; -- -0.05194038279933887
	pesos_i(15985) := b"1111111111111111_1111111111111111_1110111001000101_1100111110101011"; -- -0.0692472656828624
	pesos_i(15986) := b"0000000000000000_0000000000000000_0000100100100101_1111001011011001"; -- 0.035735300055672006
	pesos_i(15987) := b"0000000000000000_0000000000000000_0000110100101010_0101010111110111"; -- 0.051427243140267094
	pesos_i(15988) := b"0000000000000000_0000000000000000_0000110010010111_1010001100010110"; -- 0.049188797783735874
	pesos_i(15989) := b"0000000000000000_0000000000000000_0001100100001110_0000100101110100"; -- 0.09787043646040172
	pesos_i(15990) := b"0000000000000000_0000000000000000_0000100011110000_0001001011110101"; -- 0.03491323922817009
	pesos_i(15991) := b"1111111111111111_1111111111111111_1110001011010010_1010010011011000"; -- -0.11397332886137479
	pesos_i(15992) := b"0000000000000000_0000000000000000_0000000000000001_0010011100001111"; -- 1.758683374121679e-05
	pesos_i(15993) := b"1111111111111111_1111111111111111_1111011011001100_0111000011010111"; -- -0.03594298129351095
	pesos_i(15994) := b"0000000000000000_0000000000000000_0001100011110010_1100010110000100"; -- 0.09745439991006205
	pesos_i(15995) := b"0000000000000000_0000000000000000_0001111011100001_1100100001110000"; -- 0.12063267443464043
	pesos_i(15996) := b"0000000000000000_0000000000000000_0001001011001010_1001101101111111"; -- 0.07340404363927568
	pesos_i(15997) := b"1111111111111111_1111111111111111_1111000101111101_0111010101110001"; -- -0.056679401385993124
	pesos_i(15998) := b"1111111111111111_1111111111111111_1111011000000111_0010010011111111"; -- -0.03895348345210675
	pesos_i(15999) := b"0000000000000000_0000000000000000_0001111011100010_1011101010111111"; -- 0.12064711717535341
	pesos_i(16000) := b"1111111111111111_1111111111111111_1111011100001100_0001010000001010"; -- -0.034971950157224554
	pesos_i(16001) := b"1111111111111111_1111111111111111_1111111011011011_1001001011000001"; -- -0.0044620780578894246
	pesos_i(16002) := b"1111111111111111_1111111111111111_1110010101111101_0000000101100101"; -- -0.10356131822553152
	pesos_i(16003) := b"0000000000000000_0000000000000000_0001011011110011_0110100110000001"; -- 0.08965167437923648
	pesos_i(16004) := b"0000000000000000_0000000000000000_0000000111001010_0101110110011010"; -- 0.0069941045393488825
	pesos_i(16005) := b"0000000000000000_0000000000000000_0001010001110011_0100010100100111"; -- 0.07988388259224607
	pesos_i(16006) := b"1111111111111111_1111111111111111_1111110111011110_1000111000011111"; -- -0.008322827809738333
	pesos_i(16007) := b"1111111111111111_1111111111111111_1111010011000000_0011101110101010"; -- -0.043941756194729814
	pesos_i(16008) := b"1111111111111111_1111111111111111_1111001110011100_1011010001111111"; -- -0.048390120449281385
	pesos_i(16009) := b"1111111111111111_1111111111111111_1111010011010110_0110101011101001"; -- -0.043603246815122725
	pesos_i(16010) := b"1111111111111111_1111111111111111_1111111011100100_1011011000011110"; -- -0.004322641110585699
	pesos_i(16011) := b"0000000000000000_0000000000000000_0000010111100001_1111001100011100"; -- 0.02297896788353164
	pesos_i(16012) := b"0000000000000000_0000000000000000_0000101100110010_1101100010001011"; -- 0.04374459634677932
	pesos_i(16013) := b"1111111111111111_1111111111111111_1111010101000001_1100100000000000"; -- -0.041965007876049766
	pesos_i(16014) := b"1111111111111111_1111111111111111_1111000011100100_1101001110000111"; -- -0.059008387994765356
	pesos_i(16015) := b"1111111111111111_1111111111111111_1111100100101000_0011111100100011"; -- -0.026729635094229674
	pesos_i(16016) := b"0000000000000000_0000000000000000_0000001101100001_1110000110110101"; -- 0.013212305696203793
	pesos_i(16017) := b"0000000000000000_0000000000000000_0001010111101110_0100110100010100"; -- 0.08566743605631551
	pesos_i(16018) := b"1111111111111111_1111111111111111_1110101110001111_0001110101011100"; -- -0.0798474932296856
	pesos_i(16019) := b"1111111111111111_1111111111111111_1110101000000010_1011011111001010"; -- -0.08589602771004137
	pesos_i(16020) := b"1111111111111111_1111111111111111_1110000001110110_0010001010111010"; -- -0.12319739309934659
	pesos_i(16021) := b"1111111111111111_1111111111111111_1110110100100101_1101001000000010"; -- -0.073641657341007
	pesos_i(16022) := b"1111111111111111_1111111111111111_1111001001110000_0111100101100000"; -- -0.052971281125246746
	pesos_i(16023) := b"1111111111111111_1111111111111111_1111010111101011_1000111001011011"; -- -0.03937444945950671
	pesos_i(16024) := b"0000000000000000_0000000000000000_0001111010011101_1001011011101001"; -- 0.11959212478439535
	pesos_i(16025) := b"0000000000000000_0000000000000000_0000001001101011_1110001110010110"; -- 0.009458755682131947
	pesos_i(16026) := b"1111111111111111_1111111111111111_1110101100010000_1010010011101111"; -- -0.08177727857624137
	pesos_i(16027) := b"0000000000000000_0000000000000000_0010011000010001_0011000001000011"; -- 0.148699776103197
	pesos_i(16028) := b"1111111111111111_1111111111111111_1101110001011100_0001110010110101"; -- -0.1392194804429103
	pesos_i(16029) := b"1111111111111111_1111111111111111_1111111111001101_1100011011101001"; -- -0.0007663421893426647
	pesos_i(16030) := b"1111111111111111_1111111111111111_1111111000100100_1001111011001000"; -- -0.007253719526737344
	pesos_i(16031) := b"1111111111111111_1111111111111111_1101100100111101_1100100010110010"; -- -0.15140100159847503
	pesos_i(16032) := b"1111111111111111_1111111111111111_1111101001100100_1100111101101011"; -- -0.021899258060001963
	pesos_i(16033) := b"0000000000000000_0000000000000000_0000110110000000_1111001011000101"; -- 0.05274884523950841
	pesos_i(16034) := b"1111111111111111_1111111111111111_1111011111010010_1101100000011011"; -- -0.031939023371940996
	pesos_i(16035) := b"0000000000000000_0000000000000000_0000111100001100_0011110001000100"; -- 0.05878044768599975
	pesos_i(16036) := b"0000000000000000_0000000000000000_0000101110111101_1110111000011111"; -- 0.045866854257858046
	pesos_i(16037) := b"1111111111111111_1111111111111111_1110000001010011_1111101001001100"; -- -0.1237186017327975
	pesos_i(16038) := b"0000000000000000_0000000000000000_0010011011111001_0100100111010110"; -- 0.1522413394920494
	pesos_i(16039) := b"0000000000000000_0000000000000000_0000001000100001_0110010110110001"; -- 0.008322101425803164
	pesos_i(16040) := b"1111111111111111_1111111111111111_1111111101000110_1000100001011111"; -- -0.002830006522366791
	pesos_i(16041) := b"0000000000000000_0000000000000000_0000110110100101_0000110101001011"; -- 0.053299742420865284
	pesos_i(16042) := b"0000000000000000_0000000000000000_0001100001100101_1110101100100000"; -- 0.09530515217980055
	pesos_i(16043) := b"1111111111111111_1111111111111111_1110111100001000_0110110010111000"; -- -0.06627769950678769
	pesos_i(16044) := b"1111111111111111_1111111111111111_1110001011111011_1100110000100100"; -- -0.11334537616430829
	pesos_i(16045) := b"0000000000000000_0000000000000000_0010010000110111_0111111100111010"; -- 0.14147181676889775
	pesos_i(16046) := b"1111111111111111_1111111111111111_1110001010010011_1011111000110011"; -- -0.11493312125618618
	pesos_i(16047) := b"0000000000000000_0000000000000000_0000000101100011_0110101010010110"; -- 0.00542322313209973
	pesos_i(16048) := b"1111111111111111_1111111111111111_1111100111010101_1101010101101011"; -- -0.02408090719138733
	pesos_i(16049) := b"0000000000000000_0000000000000000_0000111011011000_1100101001111111"; -- 0.057995468259417954
	pesos_i(16050) := b"0000000000000000_0000000000000000_0000001110011101_1111100111001100"; -- 0.014129268912872207
	pesos_i(16051) := b"0000000000000000_0000000000000000_0000101111101100_0110100010110010"; -- 0.04657606448367548
	pesos_i(16052) := b"0000000000000000_0000000000000000_0000111001010010_1000001010001001"; -- 0.055946501301248557
	pesos_i(16053) := b"1111111111111111_1111111111111111_1110010011010011_0000101100100011"; -- -0.10615473180444437
	pesos_i(16054) := b"0000000000000000_0000000000000000_0001101110001111_1111101001010101"; -- 0.10766567788257711
	pesos_i(16055) := b"1111111111111111_1111111111111111_1101110111011101_1000000000010010"; -- -0.1333389239446319
	pesos_i(16056) := b"0000000000000000_0000000000000000_0001010111100110_0011000011100111"; -- 0.08554368632282049
	pesos_i(16057) := b"0000000000000000_0000000000000000_0001101001110111_0111011101011111"; -- 0.10338541101190775
	pesos_i(16058) := b"0000000000000000_0000000000000000_0010001001001011_0111010011010101"; -- 0.1339638728211115
	pesos_i(16059) := b"1111111111111111_1111111111111111_1111001000110101_1100011010100101"; -- -0.05386694396689524
	pesos_i(16060) := b"0000000000000000_0000000000000000_0000101010001101_1111001111001110"; -- 0.04122852107172996
	pesos_i(16061) := b"0000000000000000_0000000000000000_0001101011111010_1001110011011011"; -- 0.1053865466644247
	pesos_i(16062) := b"1111111111111111_1111111111111111_1111111100010000_0100100101111011"; -- -0.003657729566882354
	pesos_i(16063) := b"1111111111111111_1111111111111111_1111100000111101_1010100101010110"; -- -0.030309120560500356
	pesos_i(16064) := b"0000000000000000_0000000000000000_0000110111011101_1101100000110011"; -- 0.05416632889841135
	pesos_i(16065) := b"1111111111111111_1111111111111111_1111000110111011_1000111101101001"; -- -0.055731808482259046
	pesos_i(16066) := b"0000000000000000_0000000000000000_0000111111010001_1101111101101111"; -- 0.0617961545879442
	pesos_i(16067) := b"0000000000000000_0000000000000000_0001100110111100_1010111010101000"; -- 0.10053531258527912
	pesos_i(16068) := b"1111111111111111_1111111111111111_1101111010001110_0111011011110111"; -- -0.13063866104055177
	pesos_i(16069) := b"0000000000000000_0000000000000000_0010000000011111_1111110110110001"; -- 0.12548814366875244
	pesos_i(16070) := b"0000000000000000_0000000000000000_0000111010111101_0010011110010001"; -- 0.057573769545349776
	pesos_i(16071) := b"0000000000000000_0000000000000000_0001101010001110_1101000010111010"; -- 0.10374168905619517
	pesos_i(16072) := b"0000000000000000_0000000000000000_0000000111010110_1000010010100100"; -- 0.007179536784259317
	pesos_i(16073) := b"0000000000000000_0000000000000000_0000011100100110_1010100010110101"; -- 0.027933639822874935
	pesos_i(16074) := b"1111111111111111_1111111111111111_1111101001011010_1001010001100101"; -- -0.022055364045577584
	pesos_i(16075) := b"0000000000000000_0000000000000000_0001110010000010_1100100110010100"; -- 0.1113706576431942
	pesos_i(16076) := b"0000000000000000_0000000000000000_0001010000111111_1101100111000010"; -- 0.07909928319508651
	pesos_i(16077) := b"0000000000000000_0000000000000000_0000000111100110_0001101000100111"; -- 0.007417330226440697
	pesos_i(16078) := b"0000000000000000_0000000000000000_0000010111001111_0111000001100001"; -- 0.022696517634324464
	pesos_i(16079) := b"1111111111111111_1111111111111111_1101101010100110_1001101100000000"; -- -0.1458953023630952
	pesos_i(16080) := b"0000000000000000_0000000000000000_0010010101010000_1110111000001000"; -- 0.14576614092333012
	pesos_i(16081) := b"1111111111111111_1111111111111111_1110000000110101_0110100010110001"; -- -0.12418504406895163
	pesos_i(16082) := b"0000000000000000_0000000000000000_0000011000100010_0100001011100100"; -- 0.02396028592555993
	pesos_i(16083) := b"0000000000000000_0000000000000000_0000000010111011_0010010000111101"; -- 0.0028555536316208054
	pesos_i(16084) := b"1111111111111111_1111111111111111_1101110101101000_1100011110100010"; -- -0.13511993684528822
	pesos_i(16085) := b"0000000000000000_0000000000000000_0000000010110100_1000100101010110"; -- 0.0027547679130324526
	pesos_i(16086) := b"0000000000000000_0000000000000000_0000100000110110_0100001011010000"; -- 0.032077957040571176
	pesos_i(16087) := b"0000000000000000_0000000000000000_0000101101000100_0001001001000000"; -- 0.044007435527455736
	pesos_i(16088) := b"0000000000000000_0000000000000000_0000000010111111_1110010011001100"; -- 0.0029280661766610625
	pesos_i(16089) := b"0000000000000000_0000000000000000_0001010001101100_1011011011000111"; -- 0.07978384359688477
	pesos_i(16090) := b"1111111111111111_1111111111111111_1110000110111000_1000110010001110"; -- -0.11827775511495504
	pesos_i(16091) := b"0000000000000000_0000000000000000_0000011110100010_0101000101001000"; -- 0.029820518586738225
	pesos_i(16092) := b"1111111111111111_1111111111111111_1110111010110111_0111100111110111"; -- -0.06751287182072593
	pesos_i(16093) := b"0000000000000000_0000000000000000_0001100100101010_1110010000100011"; -- 0.09831071717346809
	pesos_i(16094) := b"1111111111111111_1111111111111111_1110011011101100_1101011010110011"; -- -0.09794862870759771
	pesos_i(16095) := b"0000000000000000_0000000000000000_0010010000100000_1000101010101010"; -- 0.14112154634172067
	pesos_i(16096) := b"0000000000000000_0000000000000000_0001110000010000_1111110001110001"; -- 0.1096341874161713
	pesos_i(16097) := b"0000000000000000_0000000000000000_0000010111010011_0010010000010101"; -- 0.0227530052427726
	pesos_i(16098) := b"1111111111111111_1111111111111111_1110100101110011_1001100011010011"; -- -0.0880798802202228
	pesos_i(16099) := b"0000000000000000_0000000000000000_0000100010100010_1001111100110000"; -- 0.03373141212326491
	pesos_i(16100) := b"0000000000000000_0000000000000000_0000101111111011_1100011101111110"; -- 0.046810596751320085
	pesos_i(16101) := b"1111111111111111_1111111111111111_1101110000111100_0110110001100111"; -- -0.13970301129457474
	pesos_i(16102) := b"0000000000000000_0000000000000000_0010111011111100_0010001110111010"; -- 0.18353484437288373
	pesos_i(16103) := b"1111111111111111_1111111111111111_1111101010000101_0001110001100100"; -- -0.02140638891828951
	pesos_i(16104) := b"1111111111111111_1111111111111111_1101101100101110_0100000010110110"; -- -0.14382548852700727
	pesos_i(16105) := b"1111111111111111_1111111111111111_1110000000111001_1001100000100010"; -- -0.12412118130278992
	pesos_i(16106) := b"1111111111111111_1111111111111111_1110011100110010_1100100110000110"; -- -0.09688129877523842
	pesos_i(16107) := b"1111111111111111_1111111111111111_1110110000000110_0010101000111111"; -- -0.07803092913738285
	pesos_i(16108) := b"0000000000000000_0000000000000000_0010011110111111_0000110111101111"; -- 0.1552590092947661
	pesos_i(16109) := b"0000000000000000_0000000000000000_0001001001110111_0101110110011100"; -- 0.07213387539715962
	pesos_i(16110) := b"0000000000000000_0000000000000000_0010000000111110_1110010011101101"; -- 0.12595968988634396
	pesos_i(16111) := b"0000000000000000_0000000000000000_0010000010000010_1010010100001101"; -- 0.12699348043160227
	pesos_i(16112) := b"1111111111111111_1111111111111111_1111010011110101_0010001010010011"; -- -0.04313453577979498
	pesos_i(16113) := b"1111111111111111_1111111111111111_1101100110100111_0101101100010111"; -- -0.14979010279175237
	pesos_i(16114) := b"0000000000000000_0000000000000000_0001000000011101_1010110110011101"; -- 0.06295285293771638
	pesos_i(16115) := b"0000000000000000_0000000000000000_0010010000010110_0000101100011111"; -- 0.14096135619162803
	pesos_i(16116) := b"0000000000000000_0000000000000000_0001100011010011_0100000110100001"; -- 0.09697351629474002
	pesos_i(16117) := b"1111111111111111_1111111111111111_1110111001010010_1010000010011001"; -- -0.0690517068361011
	pesos_i(16118) := b"1111111111111111_1111111111111111_1111101011011111_1101111101010100"; -- -0.020021478594362326
	pesos_i(16119) := b"0000000000000000_0000000000000000_0010000100111101_1100011000111000"; -- 0.1298488508714702
	pesos_i(16120) := b"1111111111111111_1111111111111111_1110100110000111_1000101111101100"; -- -0.08777547338523506
	pesos_i(16121) := b"1111111111111111_1111111111111111_1111001101000001_0010010000000111"; -- -0.04978728129305405
	pesos_i(16122) := b"1111111111111111_1111111111111111_1101011111110000_1111010011100010"; -- -0.15647954440116021
	pesos_i(16123) := b"0000000000000000_0000000000000000_0001110111000100_0110111100000100"; -- 0.11627858963746178
	pesos_i(16124) := b"0000000000000000_0000000000000000_0001011101011100_1101010110011101"; -- 0.09126029096344782
	pesos_i(16125) := b"1111111111111111_1111111111111111_1111010100101110_0011000001010010"; -- -0.04226396567560677
	pesos_i(16126) := b"0000000000000000_0000000000000000_0010000001111000_1111111000111111"; -- 0.12684620894230633
	pesos_i(16127) := b"0000000000000000_0000000000000000_0001101011000100_0100000111101101"; -- 0.10455715217129116
	pesos_i(16128) := b"1111111111111111_1111111111111111_1101111001001010_1110001110011111"; -- -0.13166978223182788
	pesos_i(16129) := b"0000000000000000_0000000000000000_0000010100101101_0111000000001110"; -- 0.02022457450747942
	pesos_i(16130) := b"0000000000000000_0000000000000000_0010010101001111_0100001100011010"; -- 0.14574069391870834
	pesos_i(16131) := b"0000000000000000_0000000000000000_0001100011111111_0011100010100001"; -- 0.09764436663877936
	pesos_i(16132) := b"0000000000000000_0000000000000000_0001001101100010_0101111000001010"; -- 0.07571971657943115
	pesos_i(16133) := b"1111111111111111_1111111111111111_1110101100100111_1011011011100011"; -- -0.08142525644192732
	pesos_i(16134) := b"0000000000000000_0000000000000000_0000010011010110_0110111001000000"; -- 0.01889695218519261
	pesos_i(16135) := b"1111111111111111_1111111111111111_1111010100001010_0001000010010101"; -- -0.04281517371626373
	pesos_i(16136) := b"1111111111111111_1111111111111111_1101111111111000_0011111101000110"; -- -0.125118298904054
	pesos_i(16137) := b"0000000000000000_0000000000000000_0001011001011100_0000111011011001"; -- 0.08734219351080715
	pesos_i(16138) := b"0000000000000000_0000000000000000_0001110101001101_1101001110111011"; -- 0.11446879685859895
	pesos_i(16139) := b"1111111111111111_1111111111111111_1110010110011100_1000101001111100"; -- -0.10308012448485307
	pesos_i(16140) := b"0000000000000000_0000000000000000_0010000001001100_0101001101011100"; -- 0.12616463648178494
	pesos_i(16141) := b"1111111111111111_1111111111111111_1110101001100001_0011100110001100"; -- -0.08445396728592587
	pesos_i(16142) := b"0000000000000000_0000000000000000_0000010010110010_1011001001001111"; -- 0.018351692537247857
	pesos_i(16143) := b"1111111111111111_1111111111111111_1111100000100001_1110101100100000"; -- -0.03073244531032781
	pesos_i(16144) := b"0000000000000000_0000000000000000_0000001111101100_1011111111010111"; -- 0.015331258839615437
	pesos_i(16145) := b"1111111111111111_1111111111111111_1111011000100011_0000111100010000"; -- -0.038527544699938604
	pesos_i(16146) := b"0000000000000000_0000000000000000_0001101010110000_1001010000110111"; -- 0.10425688107262802
	pesos_i(16147) := b"1111111111111111_1111111111111111_1110110110000110_0111011000100001"; -- -0.07216703125437036
	pesos_i(16148) := b"0000000000000000_0000000000000000_0000010111011101_0000001000011100"; -- 0.022903568000318945
	pesos_i(16149) := b"0000000000000000_0000000000000000_0001100010010100_0110110110011010"; -- 0.09601483351273914
	pesos_i(16150) := b"1111111111111111_1111111111111111_1111001000010111_0011011001001010"; -- -0.05433331204708496
	pesos_i(16151) := b"1111111111111111_1111111111111111_1110000011000001_1110011000001101"; -- -0.12204134154850696
	pesos_i(16152) := b"1111111111111111_1111111111111111_1111010101011001_1010110000011011"; -- -0.04160045958584517
	pesos_i(16153) := b"1111111111111111_1111111111111111_1111101101011111_1101110111011001"; -- -0.01806844180970038
	pesos_i(16154) := b"0000000000000000_0000000000000000_0000101100000100_0110010001111010"; -- 0.04303577414028241
	pesos_i(16155) := b"1111111111111111_1111111111111111_1101110000010001_1101101111010101"; -- -0.1403524976660692
	pesos_i(16156) := b"1111111111111111_1111111111111111_1111100011011101_1101001001011111"; -- -0.027865268508539067
	pesos_i(16157) := b"0000000000000000_0000000000000000_0010001011101101_0000100110111000"; -- 0.13642941230088435
	pesos_i(16158) := b"0000000000000000_0000000000000000_0001110100000000_1110001100000011"; -- 0.11329478099029011
	pesos_i(16159) := b"1111111111111111_1111111111111111_1111111010000001_1111010011111001"; -- -0.005829514783127288
	pesos_i(16160) := b"0000000000000000_0000000000000000_0001100111010010_0100000010101101"; -- 0.10086445068584253
	pesos_i(16161) := b"1111111111111111_1111111111111111_1110001001011000_1001000111100101"; -- -0.11583603061684436
	pesos_i(16162) := b"1111111111111111_1111111111111111_1111010100110001_0011100111100000"; -- -0.04221761977685327
	pesos_i(16163) := b"0000000000000000_0000000000000000_0000111101011101_0010001010100101"; -- 0.060014882358368764
	pesos_i(16164) := b"1111111111111111_1111111111111111_1110001101011100_0101111100000000"; -- -0.11187177888541978
	pesos_i(16165) := b"0000000000000000_0000000000000000_0010001100101010_0011111110110110"; -- 0.13736341657559997
	pesos_i(16166) := b"1111111111111111_1111111111111111_1110111100110110_1000101010001111"; -- -0.06557401657296254
	pesos_i(16167) := b"0000000000000000_0000000000000000_0000101000111010_1011100011101000"; -- 0.03995853114143062
	pesos_i(16168) := b"1111111111111111_1111111111111111_1110010010000101_0000011000101011"; -- -0.10734521334552789
	pesos_i(16169) := b"0000000000000000_0000000000000000_0010001100110111_1000110001011100"; -- 0.13756634955683386
	pesos_i(16170) := b"1111111111111111_1111111111111111_1110100011010111_0100101011011111"; -- -0.09046489762428749
	pesos_i(16171) := b"0000000000000000_0000000000000000_0000101110011111_0011111011100111"; -- 0.04539864666863553
	pesos_i(16172) := b"0000000000000000_0000000000000000_0001001110110111_1110101100110001"; -- 0.07702512681362224
	pesos_i(16173) := b"1111111111111111_1111111111111111_1111111011010000_1100000011000100"; -- -0.004627182138529182
	pesos_i(16174) := b"0000000000000000_0000000000000000_0000110010001000_0100000110110111"; -- 0.04895411211265877
	pesos_i(16175) := b"0000000000000000_0000000000000000_0001111111011000_1000110011011110"; -- 0.12439804486630981
	pesos_i(16176) := b"1111111111111111_1111111111111111_1110101110011100_1101001100000010"; -- -0.07963830197581905
	pesos_i(16177) := b"1111111111111111_1111111111111111_1110110110001111_0001100011010101"; -- -0.07203526302163002
	pesos_i(16178) := b"1111111111111111_1111111111111111_1110000000010011_1100001001110100"; -- -0.12469849270883565
	pesos_i(16179) := b"1111111111111111_1111111111111111_1111110111100001_1100101110100000"; -- -0.008273385580508802
	pesos_i(16180) := b"0000000000000000_0000000000000000_0000000111111000_1001010100111110"; -- 0.007699325227958107
	pesos_i(16181) := b"0000000000000000_0000000000000000_0000100111101101_0101100101011000"; -- 0.03877790824120071
	pesos_i(16182) := b"0000000000000000_0000000000000000_0000011100111110_1010110011011110"; -- 0.028300098610973184
	pesos_i(16183) := b"0000000000000000_0000000000000000_0001100101111000_1100000100010010"; -- 0.09949881260046371
	pesos_i(16184) := b"1111111111111111_1111111111111111_1111000101101100_1011000001110011"; -- -0.056935283704612365
	pesos_i(16185) := b"1111111111111111_1111111111111111_1110010010110000_0101010010011100"; -- -0.10668441012547775
	pesos_i(16186) := b"0000000000000000_0000000000000000_0000110011111000_1000001101011100"; -- 0.05066700939937303
	pesos_i(16187) := b"0000000000000000_0000000000000000_0000111101101110_0101100101011111"; -- 0.06027754372064365
	pesos_i(16188) := b"1111111111111111_1111111111111111_1111101111010110_0010101100010011"; -- -0.016263301775895127
	pesos_i(16189) := b"1111111111111111_1111111111111111_1101110111101110_0001101111001101"; -- -0.13308550115279308
	pesos_i(16190) := b"0000000000000000_0000000000000000_0001011010010101_0010000011011011"; -- 0.08821301792027803
	pesos_i(16191) := b"0000000000000000_0000000000000000_0001101001001101_1000001001000000"; -- 0.10274519030052975
	pesos_i(16192) := b"1111111111111111_1111111111111111_1111100100111010_0110100101100101"; -- -0.026452458236075418
	pesos_i(16193) := b"1111111111111111_1111111111111111_1101111011101000_1110010010111110"; -- -0.1292588268749521
	pesos_i(16194) := b"0000000000000000_0000000000000000_0010011110001000_0110011000010100"; -- 0.15442502974769723
	pesos_i(16195) := b"1111111111111111_1111111111111111_1110100111010110_1000111011101110"; -- -0.08656984984617525
	pesos_i(16196) := b"0000000000000000_0000000000000000_0000011100010101_0001011011100001"; -- 0.02766554829198416
	pesos_i(16197) := b"1111111111111111_1111111111111111_1110110101001110_1001101100010011"; -- -0.07301932128663782
	pesos_i(16198) := b"0000000000000000_0000000000000000_0000111000001110_1100001010110110"; -- 0.05491272869790013
	pesos_i(16199) := b"0000000000000000_0000000000000000_0001111101111001_1011111001111101"; -- 0.12295141741428557
	pesos_i(16200) := b"1111111111111111_1111111111111111_1110000100111000_0111100100001011"; -- -0.12023204316471783
	pesos_i(16201) := b"0000000000000000_0000000000000000_0001001000111101_0110001011110001"; -- 0.07124918347609253
	pesos_i(16202) := b"0000000000000000_0000000000000000_0000011011111111_0100011000101000"; -- 0.027332672829428438
	pesos_i(16203) := b"1111111111111111_1111111111111111_1111110000001001_1010000010000011"; -- -0.01547810355948123
	pesos_i(16204) := b"0000000000000000_0000000000000000_0001011011011100_0000011010010110"; -- 0.08929482616664952
	pesos_i(16205) := b"1111111111111111_1111111111111111_1111100110011110_0110100111101010"; -- -0.02492654836864812
	pesos_i(16206) := b"1111111111111111_1111111111111111_1111110010100001_0101101101111001"; -- -0.013162882875101973
	pesos_i(16207) := b"0000000000000000_0000000000000000_0001001010100100_0011011111101010"; -- 0.0728182740771874
	pesos_i(16208) := b"0000000000000000_0000000000000000_0010001100001001_0011011101001010"; -- 0.13685937463329245
	pesos_i(16209) := b"0000000000000000_0000000000000000_0010010101000011_1011101010110110"; -- 0.14556471780734118
	pesos_i(16210) := b"0000000000000000_0000000000000000_0000100110101111_0000110111011011"; -- 0.037827363873722326
	pesos_i(16211) := b"0000000000000000_0000000000000000_0010010011110100_0111110100001001"; -- 0.14435559711199616
	pesos_i(16212) := b"1111111111111111_1111111111111111_1111101111011100_1010100100100000"; -- -0.01616423574973241
	pesos_i(16213) := b"1111111111111111_1111111111111111_1111000100011010_1100100110111101"; -- -0.05818499696795931
	pesos_i(16214) := b"1111111111111111_1111111111111111_1110011011010010_0011010010111000"; -- -0.09835501200525998
	pesos_i(16215) := b"1111111111111111_1111111111111111_1110010110001000_1110100010000100"; -- -0.10337969571226154
	pesos_i(16216) := b"1111111111111111_1111111111111111_1101101010110010_0111100100100011"; -- -0.1457142152634594
	pesos_i(16217) := b"1111111111111111_1111111111111111_1110100110111111_0011011101101111"; -- -0.0869260170763814
	pesos_i(16218) := b"0000000000000000_0000000000000000_0001110001010010_1010100001101111"; -- 0.11063626003587226
	pesos_i(16219) := b"0000000000000000_0000000000000000_0010000000110111_1110011111011010"; -- 0.1258530528255565
	pesos_i(16220) := b"0000000000000000_0000000000000000_0000100001111100_1111101010000101"; -- 0.03315702192756556
	pesos_i(16221) := b"1111111111111111_1111111111111111_1111011101111000_1101011011010000"; -- -0.033312391546999845
	pesos_i(16222) := b"0000000000000000_0000000000000000_0000010000010110_1011010010101000"; -- 0.01597146120852551
	pesos_i(16223) := b"1111111111111111_1111111111111111_1110100100110001_0111010111111100"; -- -0.08908903690285103
	pesos_i(16224) := b"1111111111111111_1111111111111111_1101110010010000_1111011010101110"; -- -0.1384130311847339
	pesos_i(16225) := b"1111111111111111_1111111111111111_1111110011101010_0010101011110000"; -- -0.01205188408659539
	pesos_i(16226) := b"1111111111111111_1111111111111111_1110110010101110_1000011101001101"; -- -0.07546190610352718
	pesos_i(16227) := b"1111111111111111_1111111111111111_1101111010100111_0110001101000001"; -- -0.1302583663056146
	pesos_i(16228) := b"0000000000000000_0000000000000000_0000110010110001_1010011011101000"; -- 0.04958575413639799
	pesos_i(16229) := b"1111111111111111_1111111111111111_1110001001011100_0101000110000110"; -- -0.11577883219526261
	pesos_i(16230) := b"1111111111111111_1111111111111111_1101011011100010_1010101111100011"; -- -0.16060376844068852
	pesos_i(16231) := b"1111111111111111_1111111111111111_1110100010001010_0011100101101100"; -- -0.09164086459203291
	pesos_i(16232) := b"0000000000000000_0000000000000000_0010010100011101_1000110001100110"; -- 0.14498212329942006
	pesos_i(16233) := b"1111111111111111_1111111111111111_1101110010010111_0100011111011111"; -- -0.13831663889113643
	pesos_i(16234) := b"0000000000000000_0000000000000000_0001011110101100_0110111000110000"; -- 0.0924748293574029
	pesos_i(16235) := b"1111111111111111_1111111111111111_1110001101001110_0011010111000001"; -- -0.11208786042496298
	pesos_i(16236) := b"0000000000000000_0000000000000000_0001001101000010_1010111011110100"; -- 0.07523625800229038
	pesos_i(16237) := b"0000000000000000_0000000000000000_0001001001101101_0110001010100011"; -- 0.07198158710587552
	pesos_i(16238) := b"0000000000000000_0000000000000000_0000100010001110_1111010111110010"; -- 0.03343140745957705
	pesos_i(16239) := b"1111111111111111_1111111111111111_1111101100001000_1101111000011011"; -- -0.019395941162713065
	pesos_i(16240) := b"0000000000000000_0000000000000000_0000110001011101_1111111100001001"; -- 0.048309268719569365
	pesos_i(16241) := b"1111111111111111_1111111111111111_1101101001110101_0000100101010100"; -- -0.1466516657722065
	pesos_i(16242) := b"1111111111111111_1111111111111111_1111111000100011_0110110010101101"; -- -0.007271964908700557
	pesos_i(16243) := b"1111111111111111_1111111111111111_1111111111110001_0100101000101100"; -- -0.0002244608062431868
	pesos_i(16244) := b"0000000000000000_0000000000000000_0001010100101001_0001110101111001"; -- 0.0826586170911282
	pesos_i(16245) := b"1111111111111111_1111111111111111_1110111011101011_1000010000111011"; -- -0.06671880306495094
	pesos_i(16246) := b"0000000000000000_0000000000000000_0001001000001101_1111010101111110"; -- 0.07052549677721927
	pesos_i(16247) := b"0000000000000000_0000000000000000_0000101001011101_0110000011000011"; -- 0.040487334932665243
	pesos_i(16248) := b"0000000000000000_0000000000000000_0001100010000000_0011011011001010"; -- 0.09570639058408477
	pesos_i(16249) := b"0000000000000000_0000000000000000_0001001111010111_1001110000101100"; -- 0.07750869813133002
	pesos_i(16250) := b"0000000000000000_0000000000000000_0000111010100101_1101010100010100"; -- 0.05721790068309217
	pesos_i(16251) := b"0000000000000000_0000000000000000_0001110001000000_0101001100001111"; -- 0.11035651321733407
	pesos_i(16252) := b"1111111111111111_1111111111111111_1111000000101011_1011100000111101"; -- -0.06183289065996474
	pesos_i(16253) := b"1111111111111111_1111111111111111_1101110000010100_0110000101001011"; -- -0.14031402504807444
	pesos_i(16254) := b"0000000000000000_0000000000000000_0000111010101001_1110010000110101"; -- 0.0572798374912951
	pesos_i(16255) := b"1111111111111111_1111111111111111_1110011101001001_1011110101011001"; -- -0.09653107241703696
	pesos_i(16256) := b"0000000000000000_0000000000000000_0001110000100011_0001100011111110"; -- 0.10991054715872749
	pesos_i(16257) := b"0000000000000000_0000000000000000_0010000010010111_1001001000010010"; -- 0.12731278366282
	pesos_i(16258) := b"1111111111111111_1111111111111111_1110001010011011_1101111111010001"; -- -0.11480904711911885
	pesos_i(16259) := b"0000000000000000_0000000000000000_0001000101010101_0110111000010111"; -- 0.0677098088723673
	pesos_i(16260) := b"1111111111111111_1111111111111111_1110000110010011_0101001011011001"; -- -0.11884576989703508
	pesos_i(16261) := b"0000000000000000_0000000000000000_0010110011111001_1011100100001100"; -- 0.17568546821737488
	pesos_i(16262) := b"1111111111111111_1111111111111111_1111100101101001_1100111010110000"; -- -0.025729257701042015
	pesos_i(16263) := b"0000000000000000_0000000000000000_0000000011011111_1110011100010000"; -- 0.0034164823088537397
	pesos_i(16264) := b"1111111111111111_1111111111111111_1110011100111011_1001101101111001"; -- -0.09674671445893879
	pesos_i(16265) := b"1111111111111111_1111111111111111_1111100001001100_1100111111100001"; -- -0.030077941423923265
	pesos_i(16266) := b"1111111111111111_1111111111111111_1110111101011001_1100100111000001"; -- -0.06503619234722204
	pesos_i(16267) := b"0000000000000000_0000000000000000_0000010110111000_0111101001010001"; -- 0.02234615781356801
	pesos_i(16268) := b"1111111111111111_1111111111111111_1110011011001000_0001010100100001"; -- -0.09850948288333909
	pesos_i(16269) := b"0000000000000000_0000000000000000_0001111011001110_1001001101000011"; -- 0.12033958804221144
	pesos_i(16270) := b"1111111111111111_1111111111111111_1111111001011010_1101010110001111"; -- -0.006426479995486372
	pesos_i(16271) := b"1111111111111111_1111111111111111_1110001010101101_1100011000000011"; -- -0.11453592706323858
	pesos_i(16272) := b"0000000000000000_0000000000000000_0000110100011111_1000111110101001"; -- 0.051262835372845796
	pesos_i(16273) := b"1111111111111111_1111111111111111_1110110110011001_1011101111000111"; -- -0.07187296287498275
	pesos_i(16274) := b"0000000000000000_0000000000000000_0010011011011000_1111100011011010"; -- 0.1517482310366335
	pesos_i(16275) := b"1111111111111111_1111111111111111_1111110000111001_0001100111101111"; -- -0.014753703348798695
	pesos_i(16276) := b"1111111111111111_1111111111111111_1110010110110001_0101011111101001"; -- -0.10276270455272053
	pesos_i(16277) := b"0000000000000000_0000000000000000_0001001000110010_1011001100000011"; -- 0.07108610941996865
	pesos_i(16278) := b"0000000000000000_0000000000000000_0000010001100110_1111000101001000"; -- 0.01719577785424629
	pesos_i(16279) := b"0000000000000000_0000000000000000_0001110100111000_0001100101010100"; -- 0.11413725178193405
	pesos_i(16280) := b"0000000000000000_0000000000000000_0010011000110001_0010101001111000"; -- 0.1491877118919734
	pesos_i(16281) := b"0000000000000000_0000000000000000_0000101010100011_0000011100100100"; -- 0.04155010829902778
	pesos_i(16282) := b"1111111111111111_1111111111111111_1111011100101101_1001100111101111"; -- -0.034460429393589946
	pesos_i(16283) := b"0000000000000000_0000000000000000_0001001110111100_0111010010101110"; -- 0.07709435697697897
	pesos_i(16284) := b"0000000000000000_0000000000000000_0010001100000001_0100001101011010"; -- 0.13673802333378376
	pesos_i(16285) := b"0000000000000000_0000000000000000_0000001111011011_0100111100101100"; -- 0.015065143799579475
	pesos_i(16286) := b"1111111111111111_1111111111111111_1111010000110111_0001011101000000"; -- -0.04603438071476045
	pesos_i(16287) := b"0000000000000000_0000000000000000_0001010010011011_0101100111011000"; -- 0.08049546749459852
	pesos_i(16288) := b"1111111111111111_1111111111111111_1110001111111111_1110001100101000"; -- -0.10937671912964199
	pesos_i(16289) := b"0000000000000000_0000000000000000_0000000100101111_0101011110111101"; -- 0.004628642697145623
	pesos_i(16290) := b"0000000000000000_0000000000000000_0001101111000100_0011001111111100"; -- 0.10846257122858788
	pesos_i(16291) := b"1111111111111111_1111111111111111_1111100100001100_1110010111001011"; -- -0.027146947696997405
	pesos_i(16292) := b"1111111111111111_1111111111111111_1110111100110011_0010100101111010"; -- -0.06562557965603168
	pesos_i(16293) := b"1111111111111111_1111111111111111_1110000110111101_0111111000101100"; -- -0.11820231842931811
	pesos_i(16294) := b"1111111111111111_1111111111111111_1111010000100011_1000010000001011"; -- -0.046333072100403806
	pesos_i(16295) := b"0000000000000000_0000000000000000_0001101011001111_1000011011111101"; -- 0.10472911535677809
	pesos_i(16296) := b"1111111111111111_1111111111111111_1110111111110001_1011100011111011"; -- -0.06271785624350236
	pesos_i(16297) := b"0000000000000000_0000000000000000_0010100000000101_0100000000011110"; -- 0.1563301157093586
	pesos_i(16298) := b"0000000000000000_0000000000000000_0001111010011000_1110101010000011"; -- 0.11952081382033206
	pesos_i(16299) := b"1111111111111111_1111111111111111_1111100100011011_0000001011101010"; -- -0.02693158910059445
	pesos_i(16300) := b"1111111111111111_1111111111111111_1110111001100000_1111110111000001"; -- -0.06883253144275797
	pesos_i(16301) := b"1111111111111111_1111111111111111_1111110011011011_1101010001110110"; -- -0.01227066161372656
	pesos_i(16302) := b"1111111111111111_1111111111111111_1110111110001111_0110000101011001"; -- -0.06421844086407007
	pesos_i(16303) := b"0000000000000000_0000000000000000_0000101111011101_0110100000111011"; -- 0.04634715507315354
	pesos_i(16304) := b"0000000000000000_0000000000000000_0010000010001001_0010010100000101"; -- 0.12709266060955016
	pesos_i(16305) := b"0000000000000000_0000000000000000_0001011011001001_0011011100011110"; -- 0.08900780174141729
	pesos_i(16306) := b"1111111111111111_1111111111111111_1111110010110111_0000111010101000"; -- -0.012831768080317494
	pesos_i(16307) := b"1111111111111111_1111111111111111_1101011011101010_1000001111111000"; -- -0.1604840774058801
	pesos_i(16308) := b"0000000000000000_0000000000000000_0010001100011001_0011001110000010"; -- 0.13710328976157857
	pesos_i(16309) := b"0000000000000000_0000000000000000_0001001101010001_0010110000000110"; -- 0.07545733586054001
	pesos_i(16310) := b"1111111111111111_1111111111111111_1110100101110101_0100010000110110"; -- -0.08805440602696625
	pesos_i(16311) := b"0000000000000000_0000000000000000_0000100010100011_1110100001101000"; -- 0.033751035095486576
	pesos_i(16312) := b"0000000000000000_0000000000000000_0000111000111100_0010100110011000"; -- 0.05560550662113152
	pesos_i(16313) := b"0000000000000000_0000000000000000_0000010010110100_0100111100100011"; -- 0.018376298874971136
	pesos_i(16314) := b"0000000000000000_0000000000000000_0010000110011110_1101011011001100"; -- 0.1313299414614337
	pesos_i(16315) := b"1111111111111111_1111111111111111_1111000010011110_0011011010110010"; -- -0.06008585125241617
	pesos_i(16316) := b"1111111111111111_1111111111111111_1110001011111101_0001000101010101"; -- -0.11332599323016429
	pesos_i(16317) := b"1111111111111111_1111111111111111_1101110010111001_1010100110100100"; -- -0.13779201262106355
	pesos_i(16318) := b"0000000000000000_0000000000000000_0010010001101010_0101000100110010"; -- 0.14224727131134782
	pesos_i(16319) := b"1111111111111111_1111111111111111_1101101110000000_1101110011011011"; -- -0.14256496097942306
	pesos_i(16320) := b"0000000000000000_0000000000000000_0001001101010101_0111001000001111"; -- 0.07552254555168006
	pesos_i(16321) := b"0000000000000000_0000000000000000_0001010111111000_0011100001101011"; -- 0.08581879255184462
	pesos_i(16322) := b"0000000000000000_0000000000000000_0000100001110111_0101001010011101"; -- 0.03307071991840155
	pesos_i(16323) := b"1111111111111111_1111111111111111_1111010001011111_1100101111110110"; -- -0.04541325797858829
	pesos_i(16324) := b"0000000000000000_0000000000000000_0001110011001010_0011111001010000"; -- 0.112460989456886
	pesos_i(16325) := b"1111111111111111_1111111111111111_1111000001101101_1010000010111011"; -- -0.06082721167450419
	pesos_i(16326) := b"1111111111111111_1111111111111111_1101101010101010_1100101110001001"; -- -0.14583137414154376
	pesos_i(16327) := b"0000000000000000_0000000000000000_0000111010101111_1100000110010100"; -- 0.057369326313938464
	pesos_i(16328) := b"0000000000000000_0000000000000000_0001010111001100_1000100100001011"; -- 0.08515221127785043
	pesos_i(16329) := b"1111111111111111_1111111111111111_1110001110010011_0110110110110001"; -- -0.11103166988653763
	pesos_i(16330) := b"1111111111111111_1111111111111111_1111011011000000_1001101111000011"; -- -0.03612352831568488
	pesos_i(16331) := b"0000000000000000_0000000000000000_0001111111101001_1001000100100011"; -- 0.1246576986184212
	pesos_i(16332) := b"0000000000000000_0000000000000000_0010000111111111_0001011101001101"; -- 0.13279862999984016
	pesos_i(16333) := b"0000000000000000_0000000000000000_0010010110010001_1011110000100110"; -- 0.14675498891038344
	pesos_i(16334) := b"1111111111111111_1111111111111111_1110101100101011_0111110111010001"; -- -0.08136762291295058
	pesos_i(16335) := b"1111111111111111_1111111111111111_1110001100101110_1110101111011010"; -- -0.112565287839402
	pesos_i(16336) := b"0000000000000000_0000000000000000_0001000101001110_0011100001001001"; -- 0.06759979039775094
	pesos_i(16337) := b"0000000000000000_0000000000000000_0001100000000010_1001000000101000"; -- 0.09378910997756842
	pesos_i(16338) := b"0000000000000000_0000000000000000_0000101001010000_0000110101101100"; -- 0.04028400306271786
	pesos_i(16339) := b"0000000000000000_0000000000000000_0001001001001011_1001010001111100"; -- 0.07146575945251997
	pesos_i(16340) := b"0000000000000000_0000000000000000_0000111010010111_0100100001100010"; -- 0.05699589146124064
	pesos_i(16341) := b"1111111111111111_1111111111111111_1110110000011011_0111010001100001"; -- -0.07770607602264847
	pesos_i(16342) := b"0000000000000000_0000000000000000_0001001010100111_1100000110110111"; -- 0.07287226399757261
	pesos_i(16343) := b"0000000000000000_0000000000000000_0000000110001010_0101001100110000"; -- 0.006016921189467852
	pesos_i(16344) := b"0000000000000000_0000000000000000_0010001010010010_1010011011111011"; -- 0.13505023591851928
	pesos_i(16345) := b"1111111111111111_1111111111111111_1111110110010100_1011000101111001"; -- -0.009449871126835601
	pesos_i(16346) := b"1111111111111111_1111111111111111_1111010110010000_1001000010010011"; -- -0.04076286714958246
	pesos_i(16347) := b"0000000000000000_0000000000000000_0000000000111000_0111001100110001"; -- 0.0008613581787155511
	pesos_i(16348) := b"0000000000000000_0000000000000000_0010010010101001_0000010000000110"; -- 0.14320397527774742
	pesos_i(16349) := b"0000000000000000_0000000000000000_0001000111011000_0010101010010110"; -- 0.06970468672295102
	pesos_i(16350) := b"0000000000000000_0000000000000000_0001111101011110_0011111000101100"; -- 0.1225317819679145
	pesos_i(16351) := b"0000000000000000_0000000000000000_0001110100011110_0000110100011100"; -- 0.11373979511991592
	pesos_i(16352) := b"1111111111111111_1111111111111111_1111110110001100_0011010000010110"; -- -0.00957941504089029
	pesos_i(16353) := b"1111111111111111_1111111111111111_1111101110000111_1110100000001000"; -- -0.017457483369297686
	pesos_i(16354) := b"0000000000000000_0000000000000000_0001111111001001_1101011010011000"; -- 0.1241735574073309
	pesos_i(16355) := b"1111111111111111_1111111111111111_1111111111000110_1101010110110000"; -- -0.0008722730521519918
	pesos_i(16356) := b"0000000000000000_0000000000000000_0001011010011011_1100000111101001"; -- 0.08831417029010212
	pesos_i(16357) := b"0000000000000000_0000000000000000_0010001010011111_1010011110110000"; -- 0.13524864240297135
	pesos_i(16358) := b"0000000000000000_0000000000000000_0001010110111101_1010100000001100"; -- 0.08492517739400351
	pesos_i(16359) := b"0000000000000000_0000000000000000_0010010110100111_0100111001110101"; -- 0.14708414411862744
	pesos_i(16360) := b"0000000000000000_0000000000000000_0001100100110001_1101011001001010"; -- 0.09841670327901175
	pesos_i(16361) := b"1111111111111111_1111111111111111_1111111011110100_0001001001011010"; -- -0.004088261699917109
	pesos_i(16362) := b"0000000000000000_0000000000000000_0010010001001011_0010100011011010"; -- 0.14177184409213048
	pesos_i(16363) := b"0000000000000000_0000000000000000_0000110100001101_1101101111001111"; -- 0.05099271578775702
	pesos_i(16364) := b"1111111111111111_1111111111111111_1101101110110110_0001100000111110"; -- -0.14175270550167124
	pesos_i(16365) := b"0000000000000000_0000000000000000_0000111101010110_1010111101110000"; -- 0.05991646266255306
	pesos_i(16366) := b"0000000000000000_0000000000000000_0001010001111101_1000110111111101"; -- 0.08004081179597973
	pesos_i(16367) := b"0000000000000000_0000000000000000_0000011010011100_1111101100001011"; -- 0.02583283446462427
	pesos_i(16368) := b"1111111111111111_1111111111111111_1111100101001001_1100011001101011"; -- -0.02621803169333297
	pesos_i(16369) := b"0000000000000000_0000000000000000_0010001111100010_0010011101011001"; -- 0.14016958166422847
	pesos_i(16370) := b"1111111111111111_1111111111111111_1110010011100111_0101011001000101"; -- -0.10584507765816718
	pesos_i(16371) := b"0000000000000000_0000000000000000_0001101011001010_0011110111001111"; -- 0.10464845944317637
	pesos_i(16372) := b"1111111111111111_1111111111111111_1111001001011110_0100001111011101"; -- -0.053249128917803014
	pesos_i(16373) := b"0000000000000000_0000000000000000_0000110100100001_0000100000100001"; -- 0.05128527455641377
	pesos_i(16374) := b"0000000000000000_0000000000000000_0000110101000000_0101111101001001"; -- 0.05176349187973626
	pesos_i(16375) := b"1111111111111111_1111111111111111_1111101000010001_0100110010001101"; -- -0.023173537898889283
	pesos_i(16376) := b"1111111111111111_1111111111111111_1110111100110101_0100011101010000"; -- -0.06559328360828666
	pesos_i(16377) := b"0000000000000000_0000000000000000_0001100000111101_0111011100011100"; -- 0.09468788561904914
	pesos_i(16378) := b"1111111111111111_1111111111111111_1111101000010011_1010000110000001"; -- -0.023137956734214055
	pesos_i(16379) := b"0000000000000000_0000000000000000_0001101101111110_0001111111101101"; -- 0.10739326024988453
	pesos_i(16380) := b"1111111111111111_1111111111111111_1111101000110110_1100100011010001"; -- -0.022601555862745645
	pesos_i(16381) := b"0000000000000000_0000000000000000_0001111110110111_1100011010110110"; -- 0.12389795241560386
	pesos_i(16382) := b"0000000000000000_0000000000000000_0001000100100011_0011110010111101"; -- 0.06694392783283477
	pesos_i(16383) := b"1111111111111111_1111111111111111_1111100001000100_1000000000010001"; -- -0.030204768964149073
	pesos_i(16384) := b"0000000000000000_0000000000000000_0010001011101000_1111101100001000"; -- 0.13636750164736944
	pesos_i(16385) := b"1111111111111111_1111111111111111_1111010011010100_0101011100101010"; -- -0.043634941320794006
	pesos_i(16386) := b"1111111111111111_1111111111111111_1110011111011011_1110000011100111"; -- -0.09430116995774926
	pesos_i(16387) := b"1111111111111111_1111111111111111_1110111000100010_1110100110000111"; -- -0.06977978196074691
	pesos_i(16388) := b"1111111111111111_1111111111111111_1101110000000100_1011011001001001"; -- -0.1405530997394161
	pesos_i(16389) := b"0000000000000000_0000000000000000_0000010100111110_1111010110000111"; -- 0.020491929559578455
	pesos_i(16390) := b"1111111111111111_1111111111111111_1110100111100110_0010111010010011"; -- -0.08633145255981318
	pesos_i(16391) := b"1111111111111111_1111111111111111_1101101111110101_0100101011000001"; -- -0.1407883910456841
	pesos_i(16392) := b"1111111111111111_1111111111111111_1110101010111100_1101101000001011"; -- -0.0830558512076606
	pesos_i(16393) := b"0000000000000000_0000000000000000_0000111011110111_0011111010001110"; -- 0.058460149363589224
	pesos_i(16394) := b"0000000000000000_0000000000000000_0000111111010000_1101000001101111"; -- 0.06178000163206689
	pesos_i(16395) := b"1111111111111111_1111111111111111_1110011010000001_1101000101111000"; -- -0.09958163086953159
	pesos_i(16396) := b"1111111111111111_1111111111111111_1110010101001010_1001011111101010"; -- -0.10433054477111867
	pesos_i(16397) := b"1111111111111111_1111111111111111_1111000011011110_0000101011110010"; -- -0.059111896451441444
	pesos_i(16398) := b"0000000000000000_0000000000000000_0001011110000101_0000011110110111"; -- 0.09187362881509643
	pesos_i(16399) := b"1111111111111111_1111111111111111_1111100110110111_1111110110101011"; -- -0.024536271739706295
	pesos_i(16400) := b"0000000000000000_0000000000000000_0001111000001100_0011110111101111"; -- 0.11737429703755449
	pesos_i(16401) := b"0000000000000000_0000000000000000_0001110100010010_0100010010001011"; -- 0.11355999371829319
	pesos_i(16402) := b"1111111111111111_1111111111111111_1101101101111011_1111110111100101"; -- -0.14263928561681305
	pesos_i(16403) := b"0000000000000000_0000000000000000_0001001001010010_0001111000100110"; -- 0.07156551779700353
	pesos_i(16404) := b"0000000000000000_0000000000000000_0001100000101101_1100011100000111"; -- 0.09444850853653142
	pesos_i(16405) := b"1111111111111111_1111111111111111_1110000110100001_1111011110011110"; -- -0.11862232579438466
	pesos_i(16406) := b"1111111111111111_1111111111111111_1111111110111001_1011111111010100"; -- -0.0010719400730325067
	pesos_i(16407) := b"0000000000000000_0000000000000000_0001011101000100_1100101100101111"; -- 0.09089345832911278
	pesos_i(16408) := b"0000000000000000_0000000000000000_0000100100011001_0100100011100011"; -- 0.035542064163044784
	pesos_i(16409) := b"1111111111111111_1111111111111111_1111000010110110_1000101011001010"; -- -0.05971462794924672
	pesos_i(16410) := b"0000000000000000_0000000000000000_0010000111111100_1110101000101110"; -- 0.13276542309547226
	pesos_i(16411) := b"0000000000000000_0000000000000000_0001100000011000_1000101011110010"; -- 0.09412449262729243
	pesos_i(16412) := b"0000000000000000_0000000000000000_0001100111100010_1101111101101111"; -- 0.10111805391176756
	pesos_i(16413) := b"1111111111111111_1111111111111111_1111111101000101_1110101010011101"; -- -0.002839409553004005
	pesos_i(16414) := b"0000000000000000_0000000000000000_0000011100101010_1011010001010001"; -- 0.027995366881101633
	pesos_i(16415) := b"0000000000000000_0000000000000000_0000011100111111_0111101100100001"; -- 0.028312392717063064
	pesos_i(16416) := b"0000000000000000_0000000000000000_0010000001110001_1011111000001000"; -- 0.12673556999178884
	pesos_i(16417) := b"0000000000000000_0000000000000000_0001000100010101_1110110111001110"; -- 0.06674085881789986
	pesos_i(16418) := b"0000000000000000_0000000000000000_0000110111101111_0111010001100000"; -- 0.054435036998217924
	pesos_i(16419) := b"0000000000000000_0000000000000000_0001110000110110_0110000100110101"; -- 0.11020476859784858
	pesos_i(16420) := b"0000000000000000_0000000000000000_0001010110101001_1010001101011011"; -- 0.0846197222080891
	pesos_i(16421) := b"0000000000000000_0000000000000000_0001001100011001_1101011010001001"; -- 0.07461300706045113
	pesos_i(16422) := b"1111111111111111_1111111111111111_1110000000000010_0111001110010110"; -- -0.12496259295745746
	pesos_i(16423) := b"0000000000000000_0000000000000000_0001101011011000_0101100110000001"; -- 0.10486373337744705
	pesos_i(16424) := b"1111111111111111_1111111111111111_1110100110111110_0011001010101001"; -- -0.08694156043569931
	pesos_i(16425) := b"1111111111111111_1111111111111111_1110010101101111_0110111111110011"; -- -0.10376835162722751
	pesos_i(16426) := b"0000000000000000_0000000000000000_0001110000010110_1110001001011111"; -- 0.10972418608871942
	pesos_i(16427) := b"0000000000000000_0000000000000000_0000101100011001_0001011100110110"; -- 0.04335160310371978
	pesos_i(16428) := b"0000000000000000_0000000000000000_0001101100001000_1001100110101100"; -- 0.10559997985638749
	pesos_i(16429) := b"1111111111111111_1111111111111111_1111110110001001_0000110101001001"; -- -0.009627504113474211
	pesos_i(16430) := b"1111111111111111_1111111111111111_1101101101011010_1100010100101001"; -- -0.14314620736580758
	pesos_i(16431) := b"0000000000000000_0000000000000000_0000001100001001_1011110011010111"; -- 0.011867334769373664
	pesos_i(16432) := b"0000000000000000_0000000000000000_0001011011001000_0100010011001110"; -- 0.08899335878557482
	pesos_i(16433) := b"1111111111111111_1111111111111111_1101111110000101_1011110001000001"; -- -0.12686561024356047
	pesos_i(16434) := b"0000000000000000_0000000000000000_0001010000011111_0010000011001110"; -- 0.07859997787076081
	pesos_i(16435) := b"0000000000000000_0000000000000000_0000010110101001_1011110110110000"; -- 0.02212129149358562
	pesos_i(16436) := b"0000000000000000_0000000000000000_0001100000010011_1101111100010001"; -- 0.09405321285813187
	pesos_i(16437) := b"1111111111111111_1111111111111111_1101111110101101_1100001111101000"; -- -0.12625480263437802
	pesos_i(16438) := b"0000000000000000_0000000000000000_0000010000011110_1000101100011001"; -- 0.01609105445497978
	pesos_i(16439) := b"1111111111111111_1111111111111111_1111001011111001_1111001100010101"; -- -0.05087357259524136
	pesos_i(16440) := b"1111111111111111_1111111111111111_1111111000111111_1101100110111011"; -- -0.0068382185313063315
	pesos_i(16441) := b"0000000000000000_0000000000000000_0001101110010100_0100001000100111"; -- 0.10773099379322891
	pesos_i(16442) := b"0000000000000000_0000000000000000_0010011001110111_1000110110010011"; -- 0.1502617344368243
	pesos_i(16443) := b"1111111111111111_1111111111111111_1110010000101111_0111010010110100"; -- -0.10865088077520291
	pesos_i(16444) := b"1111111111111111_1111111111111111_1110111010100100_0010000010011110"; -- -0.06780811441295913
	pesos_i(16445) := b"0000000000000000_0000000000000000_0000010010011110_0000110011111001"; -- 0.018036662007758088
	pesos_i(16446) := b"0000000000000000_0000000000000000_0001111001000010_0011001010011101"; -- 0.11819759698061201
	pesos_i(16447) := b"0000000000000000_0000000000000000_0000110101100011_0100001110001010"; -- 0.052295895828394445
	pesos_i(16448) := b"0000000000000000_0000000000000000_0000011111110101_1001101111011000"; -- 0.031091442272364295
	pesos_i(16449) := b"1111111111111111_1111111111111111_1111100010010000_0011001000100010"; -- -0.02904974633456201
	pesos_i(16450) := b"0000000000000000_0000000000000000_0000001001001101_0101100111100011"; -- 0.008992784534937775
	pesos_i(16451) := b"1111111111111111_1111111111111111_1110111101110001_0110000100111001"; -- -0.06467621202597
	pesos_i(16452) := b"0000000000000000_0000000000000000_0001001100101110_1011100011000101"; -- 0.07493166730941318
	pesos_i(16453) := b"0000000000000000_0000000000000000_0000001111000010_1001000111000011"; -- 0.014687643118119046
	pesos_i(16454) := b"0000000000000000_0000000000000000_0010000000010101_0100110000100111"; -- 0.12532497350304936
	pesos_i(16455) := b"0000000000000000_0000000000000000_0001111111110101_0110101011010001"; -- 0.12483852002158466
	pesos_i(16456) := b"1111111111111111_1111111111111111_1110101111100110_1101110111111111"; -- -0.0785084964354015
	pesos_i(16457) := b"0000000000000000_0000000000000000_0000011001000000_1101110101110011"; -- 0.02442726192603008
	pesos_i(16458) := b"0000000000000000_0000000000000000_0010010011111010_1111010001010100"; -- 0.14445426025585856
	pesos_i(16459) := b"1111111111111111_1111111111111111_1101101010000100_0101011100001101"; -- -0.1464181512260886
	pesos_i(16460) := b"1111111111111111_1111111111111111_1110000111111011_1101111110010001"; -- -0.11725046834775078
	pesos_i(16461) := b"1111111111111111_1111111111111111_1111110101011010_0011110111110011"; -- -0.010341766464846278
	pesos_i(16462) := b"1111111111111111_1111111111111111_1110010100010111_1100110111101010"; -- -0.1051055243777394
	pesos_i(16463) := b"1111111111111111_1111111111111111_1111001111011000_1000101110010101"; -- -0.04747703193273135
	pesos_i(16464) := b"1111111111111111_1111111111111111_1101111111001101_0011110011011001"; -- -0.1257745713266593
	pesos_i(16465) := b"0000000000000000_0000000000000000_0000000010011100_0010000010000010"; -- 0.0023823086162954284
	pesos_i(16466) := b"1111111111111111_1111111111111111_1110010110010011_0101111011010100"; -- -0.10322005578543426
	pesos_i(16467) := b"1111111111111111_1111111111111111_1111100110001100_0010010001101100"; -- -0.02520534866369858
	pesos_i(16468) := b"1111111111111111_1111111111111111_1111101110110110_1111000011100011"; -- -0.016739792421741315
	pesos_i(16469) := b"0000000000000000_0000000000000000_0001001011000001_0101110100000110"; -- 0.07326299094825857
	pesos_i(16470) := b"1111111111111111_1111111111111111_1101111010011010_1111011111101011"; -- -0.13044786935104571
	pesos_i(16471) := b"0000000000000000_0000000000000000_0001000111110010_1101110100111001"; -- 0.07011206281077631
	pesos_i(16472) := b"1111111111111111_1111111111111111_1101111110100001_1001011110111101"; -- -0.126440540638832
	pesos_i(16473) := b"1111111111111111_1111111111111111_1110101000010100_1010110001011101"; -- -0.08562205046621309
	pesos_i(16474) := b"0000000000000000_0000000000000000_0000100111001011_0011001011001011"; -- 0.038256811781899235
	pesos_i(16475) := b"1111111111111111_1111111111111111_1101110011010011_0101100101101011"; -- -0.137400065721921
	pesos_i(16476) := b"0000000000000000_0000000000000000_0000010100000010_0010010100101100"; -- 0.019563983250113406
	pesos_i(16477) := b"0000000000000000_0000000000000000_0000011110011001_1100100111110001"; -- 0.029690381401018318
	pesos_i(16478) := b"1111111111111111_1111111111111111_1111100100110000_1011001011000000"; -- -0.026600673769566555
	pesos_i(16479) := b"1111111111111111_1111111111111111_1111000101101110_1000100110110101"; -- -0.056907075323149384
	pesos_i(16480) := b"1111111111111111_1111111111111111_1111001011101001_0100110110110111"; -- -0.051127570043535076
	pesos_i(16481) := b"1111111111111111_1111111111111111_1111000011100001_0011000111111110"; -- -0.05906379264039063
	pesos_i(16482) := b"0000000000000000_0000000000000000_0000001010010001_0001011110110100"; -- 0.010026437123606957
	pesos_i(16483) := b"1111111111111111_1111111111111111_1110010001000011_1000101110111011"; -- -0.1083443324780933
	pesos_i(16484) := b"0000000000000000_0000000000000000_0001000001000101_1001001100101111"; -- 0.06356162935068943
	pesos_i(16485) := b"1111111111111111_1111111111111111_1111101110001110_0001010110101111"; -- -0.017363209434527384
	pesos_i(16486) := b"1111111111111111_1111111111111111_1101101110101100_0000001100110101"; -- -0.1419065470301567
	pesos_i(16487) := b"1111111111111111_1111111111111111_1111010101101110_1011110101111010"; -- -0.04127898963481354
	pesos_i(16488) := b"0000000000000000_0000000000000000_0000010000100001_0011001010110110"; -- 0.01613156273433986
	pesos_i(16489) := b"1111111111111111_1111111111111111_1111101101110000_1111000100010001"; -- -0.017807896955202473
	pesos_i(16490) := b"0000000000000000_0000000000000000_0010010011000000_0001000001101101"; -- 0.1435556666163143
	pesos_i(16491) := b"1111111111111111_1111111111111111_1111111111011011_0000000000010111"; -- -0.0005645697426964144
	pesos_i(16492) := b"0000000000000000_0000000000000000_0001111111001111_1110001110010011"; -- 0.12426588377538413
	pesos_i(16493) := b"1111111111111111_1111111111111111_1111001100101111_0110101111010111"; -- -0.05005765924162088
	pesos_i(16494) := b"1111111111111111_1111111111111111_1111010110011101_1011001100011111"; -- -0.04056244360448442
	pesos_i(16495) := b"0000000000000000_0000000000000000_0001000110101110_0010101100010111"; -- 0.06906384769326604
	pesos_i(16496) := b"0000000000000000_0000000000000000_0001101011001110_1111101111010001"; -- 0.10472081998014707
	pesos_i(16497) := b"1111111111111111_1111111111111111_1111000110110110_0010011011000111"; -- -0.05581433919688082
	pesos_i(16498) := b"0000000000000000_0000000000000000_0000000111100110_1001110100010111"; -- 0.007425134738996275
	pesos_i(16499) := b"0000000000000000_0000000000000000_0000010010111111_1101110011000011"; -- 0.0185525872415341
	pesos_i(16500) := b"1111111111111111_1111111111111111_1111011100111101_0011110100100000"; -- -0.03422182048684094
	pesos_i(16501) := b"1111111111111111_1111111111111111_1111010100011000_1101001111101111"; -- -0.04258990673160658
	pesos_i(16502) := b"0000000000000000_0000000000000000_0001100010001000_0001101100001011"; -- 0.0958268072438814
	pesos_i(16503) := b"0000000000000000_0000000000000000_0001010100010111_1001100101010110"; -- 0.08239134166334942
	pesos_i(16504) := b"0000000000000000_0000000000000000_0000100100010111_1110111010101100"; -- 0.03552142809059685
	pesos_i(16505) := b"0000000000000000_0000000000000000_0000011011010010_0010001100010101"; -- 0.026643936675980192
	pesos_i(16506) := b"0000000000000000_0000000000000000_0010000011100111_0111010001011011"; -- 0.12853171549313905
	pesos_i(16507) := b"1111111111111111_1111111111111111_1110111100111110_0101110100000010"; -- -0.0654546612897293
	pesos_i(16508) := b"0000000000000000_0000000000000000_0001011011100000_0111010011100101"; -- 0.08936243612047359
	pesos_i(16509) := b"1111111111111111_1111111111111111_1101111101010011_1010110010110110"; -- -0.1276294760602906
	pesos_i(16510) := b"1111111111111111_1111111111111111_1110010101100011_0111111110101000"; -- -0.10395052093435672
	pesos_i(16511) := b"0000000000000000_0000000000000000_0000010101011001_0000011101110100"; -- 0.020889726402932123
	pesos_i(16512) := b"0000000000000000_0000000000000000_0001100100110110_0111001010010010"; -- 0.09848705351962406
	pesos_i(16513) := b"1111111111111111_1111111111111111_1110011011111011_1101101010011011"; -- -0.09771951415227768
	pesos_i(16514) := b"0000000000000000_0000000000000000_0000000110011010_1000111111000100"; -- 0.00626467259693036
	pesos_i(16515) := b"0000000000000000_0000000000000000_0010010010111000_0100001111001101"; -- 0.1434366585310557
	pesos_i(16516) := b"0000000000000000_0000000000000000_0001110111011000_1110111000011011"; -- 0.11659134057969345
	pesos_i(16517) := b"1111111111111111_1111111111111111_1110100101101110_1100010000110010"; -- -0.08815358894939984
	pesos_i(16518) := b"1111111111111111_1111111111111111_1110010110101010_1010000110111000"; -- -0.10286511674749726
	pesos_i(16519) := b"0000000000000000_0000000000000000_0000011010010011_1000100001101000"; -- 0.025688672407776794
	pesos_i(16520) := b"1111111111111111_1111111111111111_1111001100000001_1100000100010100"; -- -0.05075448297223811
	pesos_i(16521) := b"0000000000000000_0000000000000000_0000000100011011_1000001010111011"; -- 0.0043260295065656665
	pesos_i(16522) := b"0000000000000000_0000000000000000_0001000111110011_0100001010111001"; -- 0.07011811265305981
	pesos_i(16523) := b"1111111111111111_1111111111111111_1110101110010001_0100111001101010"; -- -0.0798140517532643
	pesos_i(16524) := b"1111111111111111_1111111111111111_1110001100011011_1001110100100101"; -- -0.11285989612395973
	pesos_i(16525) := b"1111111111111111_1111111111111111_1110100001011101_1101001100110110"; -- -0.09231834341991661
	pesos_i(16526) := b"0000000000000000_0000000000000000_0000011110011010_0100000001111001"; -- 0.02969744634039083
	pesos_i(16527) := b"1111111111111111_1111111111111111_1111010010110110_0101010110111000"; -- -0.04409279120995935
	pesos_i(16528) := b"1111111111111111_1111111111111111_1110111000111110_0101001011100010"; -- -0.0693615148142287
	pesos_i(16529) := b"0000000000000000_0000000000000000_0001001111110001_1110111100011101"; -- 0.07791037050532088
	pesos_i(16530) := b"1111111111111111_1111111111111111_1111111010111101_0111001011010011"; -- -0.004921744870783264
	pesos_i(16531) := b"1111111111111111_1111111111111111_1110110110000100_1111110000001111"; -- -0.07218956587234727
	pesos_i(16532) := b"0000000000000000_0000000000000000_0000110001101100_0100000001101110"; -- 0.048526789617090026
	pesos_i(16533) := b"1111111111111111_1111111111111111_1111011011110111_0011010111100101"; -- -0.03529036682530472
	pesos_i(16534) := b"1111111111111111_1111111111111111_1101101000000101_1011111101011100"; -- -0.14834980023460695
	pesos_i(16535) := b"1111111111111111_1111111111111111_1110010001010111_0100000010001110"; -- -0.10804363757320672
	pesos_i(16536) := b"1111111111111111_1111111111111111_1110001101001010_1101110110010101"; -- -0.1121388922746201
	pesos_i(16537) := b"0000000000000000_0000000000000000_0010010101101101_1010010100010101"; -- 0.14620429772649954
	pesos_i(16538) := b"0000000000000000_0000000000000000_0001101111110110_1100001111010010"; -- 0.10923408390221734
	pesos_i(16539) := b"1111111111111111_1111111111111111_1101111110001010_1101001010100111"; -- -0.12678798135451563
	pesos_i(16540) := b"1111111111111111_1111111111111111_1110001110110100_0100010111100011"; -- -0.11053050238089848
	pesos_i(16541) := b"0000000000000000_0000000000000000_0000001101101100_1000000000100010"; -- 0.013374336542903015
	pesos_i(16542) := b"0000000000000000_0000000000000000_0001110010110111_0010000110101001"; -- 0.1121693646619483
	pesos_i(16543) := b"0000000000000000_0000000000000000_0000100001110110_0100000010010000"; -- 0.033054385249324025
	pesos_i(16544) := b"0000000000000000_0000000000000000_0010010000101000_0100100101100110"; -- 0.14123972638030638
	pesos_i(16545) := b"1111111111111111_1111111111111111_1111010011001111_0001010000000101"; -- -0.04371523730934627
	pesos_i(16546) := b"1111111111111111_1111111111111111_1101110000011111_1100101110000001"; -- -0.1401398478562532
	pesos_i(16547) := b"0000000000000000_0000000000000000_0000100001010101_0100010011001011"; -- 0.0325510975621643
	pesos_i(16548) := b"1111111111111111_1111111111111111_1110110100000110_1100010001101101"; -- -0.07411548941124234
	pesos_i(16549) := b"0000000000000000_0000000000000000_0001011010001100_0101101101101001"; -- 0.08807917899064593
	pesos_i(16550) := b"0000000000000000_0000000000000000_0001110111110111_0111000010010011"; -- 0.11705688089159218
	pesos_i(16551) := b"1111111111111111_1111111111111111_1110011111100100_1101010110110101"; -- -0.09416450822275647
	pesos_i(16552) := b"0000000000000000_0000000000000000_0001010111101001_1110000001111001"; -- 0.08559992753090045
	pesos_i(16553) := b"0000000000000000_0000000000000000_0001010101000010_0011100110011100"; -- 0.08304176386300557
	pesos_i(16554) := b"1111111111111111_1111111111111111_1111001101011110_1110011101101110"; -- -0.04933312962123694
	pesos_i(16555) := b"0000000000000000_0000000000000000_0000111001110000_1100011100111000"; -- 0.05640835884720226
	pesos_i(16556) := b"1111111111111111_1111111111111111_1111001011100011_1110111001100101"; -- -0.0512095453472169
	pesos_i(16557) := b"1111111111111111_1111111111111111_1111111101110010_1111010000111001"; -- -0.002152191251823215
	pesos_i(16558) := b"0000000000000000_0000000000000000_0001101010010100_0010010110101111"; -- 0.10382304699158805
	pesos_i(16559) := b"0000000000000000_0000000000000000_0001101101100010_0101100011011101"; -- 0.10696940807517474
	pesos_i(16560) := b"0000000000000000_0000000000000000_0001000000001011_0110011001010101"; -- 0.06267394609579967
	pesos_i(16561) := b"1111111111111111_1111111111111111_1111110110101110_0110011011010111"; -- -0.009057590972550506
	pesos_i(16562) := b"0000000000000000_0000000000000000_0001001010111000_0100010010101000"; -- 0.07312420938554745
	pesos_i(16563) := b"0000000000000000_0000000000000000_0000001111010010_1011111110001101"; -- 0.014934513107795335
	pesos_i(16564) := b"1111111111111111_1111111111111111_1110010110011001_0010101001111000"; -- -0.10313162393496078
	pesos_i(16565) := b"0000000000000000_0000000000000000_0000111011111000_0000010001100010"; -- 0.05847194100711605
	pesos_i(16566) := b"1111111111111111_1111111111111111_1110011011101100_1110100011111101"; -- -0.09794753850765556
	pesos_i(16567) := b"0000000000000000_0000000000000000_0000010101111100_0000101010100000"; -- 0.021423973081490525
	pesos_i(16568) := b"1111111111111111_1111111111111111_1110000100101010_0000110000111001"; -- -0.1204521522565311
	pesos_i(16569) := b"1111111111111111_1111111111111111_1110011110101000_0000100100110010"; -- -0.09509222526612886
	pesos_i(16570) := b"0000000000000000_0000000000000000_0001110010111110_1111010101111100"; -- 0.1122888018761993
	pesos_i(16571) := b"1111111111111111_1111111111111111_1111100000100100_1010101001100000"; -- -0.030690528381652916
	pesos_i(16572) := b"1111111111111111_1111111111111111_1111000110010001_1001000001111011"; -- -0.056372613897511234
	pesos_i(16573) := b"1111111111111111_1111111111111111_1110100101111111_1101101000010101"; -- -0.08789288511664534
	pesos_i(16574) := b"0000000000000000_0000000000000000_0001101100001000_1011101011000110"; -- 0.10560195283020433
	pesos_i(16575) := b"0000000000000000_0000000000000000_0001110110000111_1100000100101011"; -- 0.115352700143694
	pesos_i(16576) := b"0000000000000000_0000000000000000_0000010011111001_0001110000000110"; -- 0.01942610891343765
	pesos_i(16577) := b"0000000000000000_0000000000000000_0010010111001111_0010111001110101"; -- 0.1476925884508416
	pesos_i(16578) := b"0000000000000000_0000000000000000_0010010000101100_1011111001111111"; -- 0.14130774123326284
	pesos_i(16579) := b"1111111111111111_1111111111111111_1111001100101000_0010011100101101"; -- -0.050168563363351265
	pesos_i(16580) := b"0000000000000000_0000000000000000_0000111100000100_0111001011011111"; -- 0.05866163210360287
	pesos_i(16581) := b"0000000000000000_0000000000000000_0000101011111100_1000000011101010"; -- 0.04291539870232072
	pesos_i(16582) := b"0000000000000000_0000000000000000_0001110011111110_1110100000111110"; -- 0.11326457515105477
	pesos_i(16583) := b"1111111111111111_1111111111111111_1111100100100110_1010011011001000"; -- -0.026753975000777808
	pesos_i(16584) := b"0000000000000000_0000000000000000_0000000101010111_1110110110110110"; -- 0.00524793337821387
	pesos_i(16585) := b"1111111111111111_1111111111111111_1110000001001001_0000110110101011"; -- -0.12388529361571532
	pesos_i(16586) := b"0000000000000000_0000000000000000_0001011100101000_1110001011001010"; -- 0.09046761914093683
	pesos_i(16587) := b"1111111111111111_1111111111111111_1110110101110000_0010111110100011"; -- -0.07250692626279405
	pesos_i(16588) := b"1111111111111111_1111111111111111_1110000110100011_1100010000010110"; -- -0.11859487965380457
	pesos_i(16589) := b"1111111111111111_1111111111111111_1110111111101111_0110101001011100"; -- -0.06275305986190208
	pesos_i(16590) := b"0000000000000000_0000000000000000_0001001010000010_1011011010001011"; -- 0.07230702295539601
	pesos_i(16591) := b"0000000000000000_0000000000000000_0010101000000110_1001011000000100"; -- 0.16416299447540297
	pesos_i(16592) := b"1111111111111111_1111111111111111_1110001011100111_0101100000011101"; -- -0.11365746777615796
	pesos_i(16593) := b"1111111111111111_1111111111111111_1110110010011100_1011110011111100"; -- -0.07573336461014649
	pesos_i(16594) := b"1111111111111111_1111111111111111_1111010011001011_1100110111101110"; -- -0.04376519136024491
	pesos_i(16595) := b"0000000000000000_0000000000000000_0000000110000011_1011010000101011"; -- 0.0059158901645775044
	pesos_i(16596) := b"0000000000000000_0000000000000000_0000000100111111_1100110001000000"; -- 0.004879728056725786
	pesos_i(16597) := b"1111111111111111_1111111111111111_1111101001100001_0001101011001100"; -- -0.02195580027589065
	pesos_i(16598) := b"1111111111111111_1111111111111111_1101110011101000_1111110101101100"; -- -0.13706985579597664
	pesos_i(16599) := b"1111111111111111_1111111111111111_1111100000000010_1011001101101011"; -- -0.031208788184615456
	pesos_i(16600) := b"0000000000000000_0000000000000000_0000011000100010_0101110010000101"; -- 0.02396181335918595
	pesos_i(16601) := b"0000000000000000_0000000000000000_0000100100100100_1110000011111010"; -- 0.035718975987873845
	pesos_i(16602) := b"1111111111111111_1111111111111111_1111100110001001_0011101101000100"; -- -0.025249763493590684
	pesos_i(16603) := b"1111111111111111_1111111111111111_1111110110100100_0001110110000101"; -- -0.009214549133787215
	pesos_i(16604) := b"0000000000000000_0000000000000000_0000001100000110_0000110111110001"; -- 0.011811133769604566
	pesos_i(16605) := b"1111111111111111_1111111111111111_1110010100010100_0011100111100110"; -- -0.10516012310824975
	pesos_i(16606) := b"1111111111111111_1111111111111111_1110111010010111_0000000101101011"; -- -0.0680083383683145
	pesos_i(16607) := b"1111111111111111_1111111111111111_1110001000101010_0110111010100111"; -- -0.11654003556104164
	pesos_i(16608) := b"1111111111111111_1111111111111111_1110010001010111_0111110000000101"; -- -0.10804009322979792
	pesos_i(16609) := b"1111111111111111_1111111111111111_1110101100010111_1010111111110110"; -- -0.08166980966890988
	pesos_i(16610) := b"1111111111111111_1111111111111111_1110101001110010_0110100100100001"; -- -0.0841917319278368
	pesos_i(16611) := b"0000000000000000_0000000000000000_0000101011010110_0001001100110001"; -- 0.042329024814931275
	pesos_i(16612) := b"0000000000000000_0000000000000000_0001001111101100_1111101001101010"; -- 0.07783475003631406
	pesos_i(16613) := b"1111111111111111_1111111111111111_1110101010111110_0111011100000101"; -- -0.08303123604018751
	pesos_i(16614) := b"0000000000000000_0000000000000000_0000110000111010_1011001000110111"; -- 0.04777063208216941
	pesos_i(16615) := b"0000000000000000_0000000000000000_0010000110010100_0111011000101011"; -- 0.13117159417849464
	pesos_i(16616) := b"0000000000000000_0000000000000000_0000101001111110_0010100110010001"; -- 0.04098758501913188
	pesos_i(16617) := b"0000000000000000_0000000000000000_0000110000011111_0000010110010101"; -- 0.047348355285620196
	pesos_i(16618) := b"0000000000000000_0000000000000000_0000111011111011_1011011101000100"; -- 0.05852837965051234
	pesos_i(16619) := b"0000000000000000_0000000000000000_0000001111110010_1000100101110011"; -- 0.015419569626221517
	pesos_i(16620) := b"1111111111111111_1111111111111111_1111011011001011_0100111100101000"; -- -0.035960247760625105
	pesos_i(16621) := b"0000000000000000_0000000000000000_0000101001011101_1010101100001101"; -- 0.04049176278199332
	pesos_i(16622) := b"1111111111111111_1111111111111111_1110110011111001_0111101110111010"; -- -0.07431818685546358
	pesos_i(16623) := b"0000000000000000_0000000000000000_0000110111001010_0010011000000011"; -- 0.053865791002215405
	pesos_i(16624) := b"1111111111111111_1111111111111111_1111110000101100_1011100000101011"; -- -0.014942636001673969
	pesos_i(16625) := b"0000000000000000_0000000000000000_0001101011010000_1100010101001101"; -- 0.10474808812452062
	pesos_i(16626) := b"1111111111111111_1111111111111111_1110000101101111_0010101101111101"; -- -0.11939743227018133
	pesos_i(16627) := b"0000000000000000_0000000000000000_0001110010101010_1100100100100011"; -- 0.11198098290581278
	pesos_i(16628) := b"0000000000000000_0000000000000000_0001100111110010_0000010111101000"; -- 0.1013492290794871
	pesos_i(16629) := b"0000000000000000_0000000000000000_0001110010110111_1110110000011100"; -- 0.11218143155817986
	pesos_i(16630) := b"1111111111111111_1111111111111111_1111010110011100_1001111001011100"; -- -0.04057894000559582
	pesos_i(16631) := b"0000000000000000_0000000000000000_0000110111011010_1111111100111000"; -- 0.05412287815430367
	pesos_i(16632) := b"1111111111111111_1111111111111111_1111010000001010_1011110000010101"; -- -0.04671120144642026
	pesos_i(16633) := b"1111111111111111_1111111111111111_1110101110110010_1000011110110011"; -- -0.07930709729710828
	pesos_i(16634) := b"1111111111111111_1111111111111111_1111001011011011_0111001010011110"; -- -0.051338993409514866
	pesos_i(16635) := b"1111111111111111_1111111111111111_1101111110001110_0110101001111101"; -- -0.12673315472778923
	pesos_i(16636) := b"1111111111111111_1111111111111111_1110100001101101_0000110011100101"; -- -0.09208602333845181
	pesos_i(16637) := b"1111111111111111_1111111111111111_1110101100000010_0101000010110000"; -- -0.08199592302128056
	pesos_i(16638) := b"1111111111111111_1111111111111111_1110111110110001_0101100100111011"; -- -0.06370012578289311
	pesos_i(16639) := b"1111111111111111_1111111111111111_1111000110001101_1000111101010100"; -- -0.05643371773137998
	pesos_i(16640) := b"1111111111111111_1111111111111111_1110001101001100_0101000100001000"; -- -0.11211675208430967
	pesos_i(16641) := b"0000000000000000_0000000000000000_0000101011111011_0011001000111011"; -- 0.042895449924864985
	pesos_i(16642) := b"0000000000000000_0000000000000000_0000101011111101_1001101011001111"; -- 0.042932200837319114
	pesos_i(16643) := b"0000000000000000_0000000000000000_0000011001010010_0011100100001000"; -- 0.02469211994940085
	pesos_i(16644) := b"1111111111111111_1111111111111111_1111000110001111_0000001000111101"; -- -0.05641160985725038
	pesos_i(16645) := b"1111111111111111_1111111111111111_1111100111110111_1110000101000101"; -- -0.023561401940967078
	pesos_i(16646) := b"0000000000000000_0000000000000000_0010000111001010_0100110111111001"; -- 0.13199317303197644
	pesos_i(16647) := b"1111111111111111_1111111111111111_1111110100110110_0111101011111101"; -- -0.010887444646833857
	pesos_i(16648) := b"1111111111111111_1111111111111111_1110101101101111_0110001011100110"; -- -0.08033162950358584
	pesos_i(16649) := b"1111111111111111_1111111111111111_1110011000111110_1110011101011000"; -- -0.10060266580966452
	pesos_i(16650) := b"0000000000000000_0000000000000000_0010011100101000_0011011011011000"; -- 0.15295737054276215
	pesos_i(16651) := b"0000000000000000_0000000000000000_0000100000110111_0100001001010001"; -- 0.032093186191567785
	pesos_i(16652) := b"1111111111111111_1111111111111111_1111101100000001_0010100111110101"; -- -0.019513490460837887
	pesos_i(16653) := b"0000000000000000_0000000000000000_0010000110101001_0001001100010100"; -- 0.13148612242202154
	pesos_i(16654) := b"0000000000000000_0000000000000000_0001100110110101_0011010110110100"; -- 0.10042129180442637
	pesos_i(16655) := b"1111111111111111_1111111111111111_1111011000011101_0000001110001101"; -- -0.038619783584955644
	pesos_i(16656) := b"0000000000000000_0000000000000000_0000011000010010_0101011111111101"; -- 0.023717402718216783
	pesos_i(16657) := b"0000000000000000_0000000000000000_0000011100000011_0001100011011110"; -- 0.027391008605543672
	pesos_i(16658) := b"0000000000000000_0000000000000000_0000011110000100_0111100011000000"; -- 0.02936510732541518
	pesos_i(16659) := b"0000000000000000_0000000000000000_0000111111111100_1111110010000111"; -- 0.06245401672452252
	pesos_i(16660) := b"0000000000000000_0000000000000000_0001101011100011_0010101010111110"; -- 0.10502879271748666
	pesos_i(16661) := b"1111111111111111_1111111111111111_1101101100011001_0000111000110000"; -- -0.14414893455561678
	pesos_i(16662) := b"0000000000000000_0000000000000000_0010011001110010_0010010100110110"; -- 0.15017921993680233
	pesos_i(16663) := b"1111111111111111_1111111111111111_1111001001010011_1101100001010010"; -- -0.053408126810834775
	pesos_i(16664) := b"0000000000000000_0000000000000000_0001001001000101_0101010000110011"; -- 0.07137037507186746
	pesos_i(16665) := b"0000000000000000_0000000000000000_0001111110001111_0110100001011000"; -- 0.12328197616488071
	pesos_i(16666) := b"0000000000000000_0000000000000000_0010010001111100_0100111100110111"; -- 0.14252181142240605
	pesos_i(16667) := b"0000000000000000_0000000000000000_0001101011110101_1110001100001010"; -- 0.10531443585968539
	pesos_i(16668) := b"1111111111111111_1111111111111111_1111100010100010_1101010011110110"; -- -0.028765382708931975
	pesos_i(16669) := b"1111111111111111_1111111111111111_1111110010011010_1001110011001010"; -- -0.013265801100732697
	pesos_i(16670) := b"1111111111111111_1111111111111111_1111101011100010_1111000101000001"; -- -0.019974633702732825
	pesos_i(16671) := b"0000000000000000_0000000000000000_0001110010101001_0111001110100011"; -- 0.11196062787893922
	pesos_i(16672) := b"0000000000000000_0000000000000000_0001000110011000_0101000010010110"; -- 0.0687303891784171
	pesos_i(16673) := b"1111111111111111_1111111111111111_1111001100110010_0100111001111101"; -- -0.05001363221851123
	pesos_i(16674) := b"0000000000000000_0000000000000000_0001000010101111_1011000110110111"; -- 0.06518088069003104
	pesos_i(16675) := b"0000000000000000_0000000000000000_0001001110000011_0100110110000001"; -- 0.07622227096394776
	pesos_i(16676) := b"0000000000000000_0000000000000000_0000011100010100_0100011010011001"; -- 0.027653133768912343
	pesos_i(16677) := b"0000000000000000_0000000000000000_0000000000001110_1111111111001011"; -- 0.00022886950298743323
	pesos_i(16678) := b"0000000000000000_0000000000000000_0000101101001110_0011111000111101"; -- 0.044162645285490215
	pesos_i(16679) := b"0000000000000000_0000000000000000_0001000110000100_1111000100000010"; -- 0.0684347753767663
	pesos_i(16680) := b"0000000000000000_0000000000000000_0010000011010100_1110001011010110"; -- 0.1282483837072952
	pesos_i(16681) := b"0000000000000000_0000000000000000_0001100101101000_1001111011100011"; -- 0.09925263444677403
	pesos_i(16682) := b"1111111111111111_1111111111111111_1111010110101100_0000101101000110"; -- -0.04034356630795126
	pesos_i(16683) := b"1111111111111111_1111111111111111_1111000000001110_1110000100010110"; -- -0.06227296090149868
	pesos_i(16684) := b"1111111111111111_1111111111111111_1110110110001001_1010010110001010"; -- -0.07211842893150945
	pesos_i(16685) := b"1111111111111111_1111111111111111_1110010101110010_0001001101000100"; -- -0.1037280998011243
	pesos_i(16686) := b"1111111111111111_1111111111111111_1111101010000010_0100000101101000"; -- -0.021449958824990182
	pesos_i(16687) := b"0000000000000000_0000000000000000_0000000111010010_0110010011011111"; -- 0.0071166081114915165
	pesos_i(16688) := b"0000000000000000_0000000000000000_0000111010100000_0001010011101011"; -- 0.05713015306958364
	pesos_i(16689) := b"1111111111111111_1111111111111111_1110000111010001_0011101011001001"; -- -0.11790115920040818
	pesos_i(16690) := b"0000000000000000_0000000000000000_0000100110000010_1101110011101101"; -- 0.03715306074486974
	pesos_i(16691) := b"1111111111111111_1111111111111111_1111010010100011_0101011001100001"; -- -0.04438266869662436
	pesos_i(16692) := b"1111111111111111_1111111111111111_1101101111001001_1111011110010011"; -- -0.1414494769151344
	pesos_i(16693) := b"1111111111111111_1111111111111111_1111000101001100_0100100010010101"; -- -0.05742975581302636
	pesos_i(16694) := b"1111111111111111_1111111111111111_1110011101101111_1100110100010011"; -- -0.09595030103851401
	pesos_i(16695) := b"1111111111111111_1111111111111111_1110010011010100_0000100001001110"; -- -0.10613964162259824
	pesos_i(16696) := b"1111111111111111_1111111111111111_1110001000000111_0101100111010110"; -- -0.11707533379345474
	pesos_i(16697) := b"1111111111111111_1111111111111111_1111101110010000_1111101101110001"; -- -0.017318997261661882
	pesos_i(16698) := b"1111111111111111_1111111111111111_1110110101100000_0100001110010010"; -- -0.07274987877290608
	pesos_i(16699) := b"0000000000000000_0000000000000000_0000100011100000_0111101110000000"; -- 0.034675329848876765
	pesos_i(16700) := b"1111111111111111_1111111111111111_1111011001101111_1100000011101010"; -- -0.037357275734862375
	pesos_i(16701) := b"1111111111111111_1111111111111111_1110110011100011_0011110000100001"; -- -0.07465767098674791
	pesos_i(16702) := b"1111111111111111_1111111111111111_1110001110101110_0111100101011001"; -- -0.11061898781605313
	pesos_i(16703) := b"1111111111111111_1111111111111111_1110010000001000_1111000011101101"; -- -0.10923856950469038
	pesos_i(16704) := b"0000000000000000_0000000000000000_0010001001011001_0111110110111011"; -- 0.1341780262856337
	pesos_i(16705) := b"1111111111111111_1111111111111111_1110001110000101_1101010000001110"; -- -0.11123919152799903
	pesos_i(16706) := b"1111111111111111_1111111111111111_1110000100001011_1001110010101100"; -- -0.1209165648656923
	pesos_i(16707) := b"0000000000000000_0000000000000000_0001001001010011_0001110010001000"; -- 0.07158068002287926
	pesos_i(16708) := b"0000000000000000_0000000000000000_0000101011100011_0100001111011000"; -- 0.04253028900863526
	pesos_i(16709) := b"0000000000000000_0000000000000000_0001111111110111_0001000101110010"; -- 0.12486371080516907
	pesos_i(16710) := b"1111111111111111_1111111111111111_1111111100001101_0011110011111101"; -- -0.0037042504569934783
	pesos_i(16711) := b"0000000000000000_0000000000000000_0000100111001000_1010001110010010"; -- 0.03821775742241651
	pesos_i(16712) := b"0000000000000000_0000000000000000_0001101110011100_1011000010111010"; -- 0.10785965485682075
	pesos_i(16713) := b"1111111111111111_1111111111111111_1111100000100011_1111010011001100"; -- -0.030701351430662483
	pesos_i(16714) := b"1111111111111111_1111111111111111_1110101001100110_1010101011110110"; -- -0.08437091339062455
	pesos_i(16715) := b"0000000000000000_0000000000000000_0001101011001100_1100100001101111"; -- 0.10468723974011737
	pesos_i(16716) := b"1111111111111111_1111111111111111_1110110100100001_0101100101110011"; -- -0.07370987830889231
	pesos_i(16717) := b"0000000000000000_0000000000000000_0001010001101010_1010101001100001"; -- 0.07975258709024301
	pesos_i(16718) := b"0000000000000000_0000000000000000_0000111011011100_0110000111111000"; -- 0.058050272959980505
	pesos_i(16719) := b"1111111111111111_1111111111111111_1111000011111101_0110010010001110"; -- -0.05863353277086974
	pesos_i(16720) := b"0000000000000000_0000000000000000_0010000100111111_1111000010100100"; -- 0.1298818969487341
	pesos_i(16721) := b"1111111111111111_1111111111111111_1101101111100000_0000111101001100"; -- -0.14111236937268454
	pesos_i(16722) := b"0000000000000000_0000000000000000_0001110000110100_0100100111100000"; -- 0.11017286034646197
	pesos_i(16723) := b"0000000000000000_0000000000000000_0010000011111110_1001001110111001"; -- 0.12888453727682794
	pesos_i(16724) := b"1111111111111111_1111111111111111_1101100010111011_1101000100000111"; -- -0.1533841475109345
	pesos_i(16725) := b"1111111111111111_1111111111111111_1110110100011011_1101001110100100"; -- -0.07379414800175577
	pesos_i(16726) := b"1111111111111111_1111111111111111_1101111010001011_1000111101011001"; -- -0.13068298416722776
	pesos_i(16727) := b"1111111111111111_1111111111111111_1111010001111010_1110111101010000"; -- -0.04499916358510145
	pesos_i(16728) := b"1111111111111111_1111111111111111_1110011100000000_1110001110111010"; -- -0.09764267634520761
	pesos_i(16729) := b"0000000000000000_0000000000000000_0010001011011000_1000100110011000"; -- 0.1361165996721117
	pesos_i(16730) := b"0000000000000000_0000000000000000_0001011000100011_0110011110001100"; -- 0.08647772956091838
	pesos_i(16731) := b"0000000000000000_0000000000000000_0001101100111001_0110000100010100"; -- 0.10634428716930971
	pesos_i(16732) := b"1111111111111111_1111111111111111_1110010110011010_1001011111011101"; -- -0.10310984463682854
	pesos_i(16733) := b"1111111111111111_1111111111111111_1101111010000010_1100001011100000"; -- -0.13081724190114805
	pesos_i(16734) := b"1111111111111111_1111111111111111_1110001111000001_0111111100110101"; -- -0.11032872162706754
	pesos_i(16735) := b"1111111111111111_1111111111111111_1110100001000110_0011000100100110"; -- -0.09267895528315238
	pesos_i(16736) := b"1111111111111111_1111111111111111_1110000001001010_0100111011111000"; -- -0.12386614273174328
	pesos_i(16737) := b"1111111111111111_1111111111111111_1110110011011001_0101000101110111"; -- -0.0748089870805249
	pesos_i(16738) := b"1111111111111111_1111111111111111_1111011000001010_1101011000010111"; -- -0.03889715143765512
	pesos_i(16739) := b"1111111111111111_1111111111111111_1111111101110010_1101010101010110"; -- -0.00215403217402304
	pesos_i(16740) := b"1111111111111111_1111111111111111_1101110111000000_0111110110010001"; -- -0.13378157825007966
	pesos_i(16741) := b"1111111111111111_1111111111111111_1110101101011100_1011101111101010"; -- -0.08061624084058581
	pesos_i(16742) := b"1111111111111111_1111111111111111_1111011111100101_1111110010000000"; -- -0.031646937130918505
	pesos_i(16743) := b"1111111111111111_1111111111111111_1111010101100111_1100100011010000"; -- -0.041385125378343574
	pesos_i(16744) := b"1111111111111111_1111111111111111_1111110111000000_0111111011001101"; -- -0.008781504506620512
	pesos_i(16745) := b"1111111111111111_1111111111111111_1111000101011101_1110110111110111"; -- -0.05716049876638251
	pesos_i(16746) := b"1111111111111111_1111111111111111_1110010110101111_0100010111011100"; -- -0.10279429806921948
	pesos_i(16747) := b"0000000000000000_0000000000000000_0000001011010100_0011011100111111"; -- 0.011050656113531628
	pesos_i(16748) := b"0000000000000000_0000000000000000_0000000111011011_1111100001101110"; -- 0.0072627323074261445
	pesos_i(16749) := b"1111111111111111_1111111111111111_1110010110000110_0000111010110000"; -- -0.10342319677824047
	pesos_i(16750) := b"0000000000000000_0000000000000000_0000101100011100_0100110010001111"; -- 0.04340055942235824
	pesos_i(16751) := b"1111111111111111_1111111111111111_1110110010100001_1100010101010010"; -- -0.07565657384267645
	pesos_i(16752) := b"1111111111111111_1111111111111111_1110000101110111_0110010111101011"; -- -0.11927187943160679
	pesos_i(16753) := b"0000000000000000_0000000000000000_0001110101010110_1000000110001011"; -- 0.1146012271239355
	pesos_i(16754) := b"0000000000000000_0000000000000000_0001011000010111_0011101001011100"; -- 0.08629193054163134
	pesos_i(16755) := b"1111111111111111_1111111111111111_1101110010000101_1000110101011001"; -- -0.13858715600658048
	pesos_i(16756) := b"0000000000000000_0000000000000000_0000110111001110_1000100111010111"; -- 0.053932776349811584
	pesos_i(16757) := b"1111111111111111_1111111111111111_1110000101001110_0100000110100100"; -- -0.11989965190473205
	pesos_i(16758) := b"0000000000000000_0000000000000000_0010010100110110_1010100001001100"; -- 0.14536525587513183
	pesos_i(16759) := b"0000000000000000_0000000000000000_0000110100111110_0100001011111110"; -- 0.05173128807714602
	pesos_i(16760) := b"0000000000000000_0000000000000000_0000001110101010_0101000001010100"; -- 0.01431753201896585
	pesos_i(16761) := b"0000000000000000_0000000000000000_0010010101100110_1000001001100011"; -- 0.14609541820227176
	pesos_i(16762) := b"0000000000000000_0000000000000000_0001101011000101_0000010101111001"; -- 0.10456880753741554
	pesos_i(16763) := b"1111111111111111_1111111111111111_1110000011011001_0110111101100100"; -- -0.12168220343285828
	pesos_i(16764) := b"1111111111111111_1111111111111111_1111000100000011_0000011001001100"; -- -0.0585475983643927
	pesos_i(16765) := b"1111111111111111_1111111111111111_1111000011101110_1111100110001100"; -- -0.05885353395600872
	pesos_i(16766) := b"0000000000000000_0000000000000000_0000110010000111_1100010110010101"; -- 0.04894671340805481
	pesos_i(16767) := b"0000000000000000_0000000000000000_0001101000010110_0100111100001011"; -- 0.1019029047797198
	pesos_i(16768) := b"0000000000000000_0000000000000000_0001100010000110_0010011111001110"; -- 0.09579705030843011
	pesos_i(16769) := b"0000000000000000_0000000000000000_0001001110110001_0100010010101011"; -- 0.07692364857197474
	pesos_i(16770) := b"0000000000000000_0000000000000000_0010000101010100_1010001010100100"; -- 0.13019768241003785
	pesos_i(16771) := b"0000000000000000_0000000000000000_0001101101111010_1111111001111011"; -- 0.10734549053513776
	pesos_i(16772) := b"1111111111111111_1111111111111111_1101110110001100_0011000110100110"; -- -0.1345795601590617
	pesos_i(16773) := b"0000000000000000_0000000000000000_0001010000011101_0001100010111001"; -- 0.07856897835462472
	pesos_i(16774) := b"1111111111111111_1111111111111111_1110011100000101_1100011001000111"; -- -0.09756813771465082
	pesos_i(16775) := b"0000000000000000_0000000000000000_0000100001110110_1101111101111110"; -- 0.033063858197962426
	pesos_i(16776) := b"1111111111111111_1111111111111111_1110001010111100_0010101000100011"; -- -0.11431633615576411
	pesos_i(16777) := b"1111111111111111_1111111111111111_1110000110111111_0100111000100001"; -- -0.11817466450210173
	pesos_i(16778) := b"1111111111111111_1111111111111111_1111110101011010_1000001000001110"; -- -0.010337707115376887
	pesos_i(16779) := b"0000000000000000_0000000000000000_0000100110001100_0011000101100001"; -- 0.03729542373954148
	pesos_i(16780) := b"1111111111111111_1111111111111111_1110011110101100_1111010111100110"; -- -0.09501708154695111
	pesos_i(16781) := b"1111111111111111_1111111111111111_1110000010100100_1100101101101000"; -- -0.12248543467084984
	pesos_i(16782) := b"1111111111111111_1111111111111111_1110001000101010_0111110110000001"; -- -0.11653915023303313
	pesos_i(16783) := b"0000000000000000_0000000000000000_0010011110111010_0110011011001110"; -- 0.1551880123043378
	pesos_i(16784) := b"1111111111111111_1111111111111111_1111101100000111_1010101000011011"; -- -0.019414299336417508
	pesos_i(16785) := b"1111111111111111_1111111111111111_1111111111110111_0111010001101100"; -- -0.00013038979251497735
	pesos_i(16786) := b"1111111111111111_1111111111111111_1111011011001101_0011010111001110"; -- -0.03593124127601035
	pesos_i(16787) := b"1111111111111111_1111111111111111_1110001111100011_0111101111100010"; -- -0.10981012092028825
	pesos_i(16788) := b"1111111111111111_1111111111111111_1110000101000100_1010010100001001"; -- -0.12004631553517126
	pesos_i(16789) := b"1111111111111111_1111111111111111_1111111010011100_1001101010110001"; -- -0.005422908634374291
	pesos_i(16790) := b"0000000000000000_0000000000000000_0001011000000100_1101010010010110"; -- 0.0860112061845349
	pesos_i(16791) := b"0000000000000000_0000000000000000_0010011001100000_0100000000110010"; -- 0.1499061701331589
	pesos_i(16792) := b"1111111111111111_1111111111111111_1111011110100101_0101001110001000"; -- -0.032633570869699854
	pesos_i(16793) := b"0000000000000000_0000000000000000_0001111001100001_0100100110001110"; -- 0.11867198662553492
	pesos_i(16794) := b"0000000000000000_0000000000000000_0000000011100100_0010001100101110"; -- 0.003481100702583895
	pesos_i(16795) := b"0000000000000000_0000000000000000_0001011111111100_0011011101011110"; -- 0.09369226497582786
	pesos_i(16796) := b"1111111111111111_1111111111111111_1101110000010011_1010100101111001"; -- -0.14032498156070666
	pesos_i(16797) := b"1111111111111111_1111111111111111_1110100110011110_1010000010110011"; -- -0.08742328296963754
	pesos_i(16798) := b"1111111111111111_1111111111111111_1111111001010000_0110100000110110"; -- -0.006585585356123247
	pesos_i(16799) := b"0000000000000000_0000000000000000_0010010000010101_0010100100000101"; -- 0.14094787957044067
	pesos_i(16800) := b"1111111111111111_1111111111111111_1111000111111000_0110011010011110"; -- -0.054803453767459646
	pesos_i(16801) := b"0000000000000000_0000000000000000_0001100000111110_1110000111000111"; -- 0.09470950232344066
	pesos_i(16802) := b"1111111111111111_1111111111111111_1101110000011001_0001000111111110"; -- -0.1402424578237589
	pesos_i(16803) := b"1111111111111111_1111111111111111_1110110010011010_1100101000100111"; -- -0.07576309734115726
	pesos_i(16804) := b"1111111111111111_1111111111111111_1111111100001100_0011100100110001"; -- -0.003719735768541163
	pesos_i(16805) := b"1111111111111111_1111111111111111_1101110101101111_1100011101010111"; -- -0.13501314281944288
	pesos_i(16806) := b"0000000000000000_0000000000000000_0010100110111100_0101101110111110"; -- 0.16303037061473707
	pesos_i(16807) := b"0000000000000000_0000000000000000_0000100001010101_1001010011001111"; -- 0.03255586675748752
	pesos_i(16808) := b"0000000000000000_0000000000000000_0000100011010110_0010011110011100"; -- 0.03451774170575448
	pesos_i(16809) := b"1111111111111111_1111111111111111_1110001111100011_0100000011001101"; -- -0.10981364236741445
	pesos_i(16810) := b"0000000000000000_0000000000000000_0010001010011101_1101010001010011"; -- 0.13522078534530113
	pesos_i(16811) := b"0000000000000000_0000000000000000_0000000011010110_1111011010110100"; -- 0.003280085495045707
	pesos_i(16812) := b"1111111111111111_1111111111111111_1110001111110101_0111101000010011"; -- -0.10953557045309711
	pesos_i(16813) := b"0000000000000000_0000000000000000_0001000000100010_0000100111110101"; -- 0.06301939221634346
	pesos_i(16814) := b"1111111111111111_1111111111111111_1110100010100111_0110010110000000"; -- -0.09119573238940888
	pesos_i(16815) := b"0000000000000000_0000000000000000_0000101011101110_1111111011000001"; -- 0.042709276426572566
	pesos_i(16816) := b"1111111111111111_1111111111111111_1111010001001101_1010010001110011"; -- -0.045690271229836564
	pesos_i(16817) := b"1111111111111111_1111111111111111_1111101111010011_1000001011011000"; -- -0.016303846667546737
	pesos_i(16818) := b"0000000000000000_0000000000000000_0000001010110100_1111010111110110"; -- 0.0105737424507839
	pesos_i(16819) := b"0000000000000000_0000000000000000_0001110101011010_0101000101010100"; -- 0.11465938859379972
	pesos_i(16820) := b"0000000000000000_0000000000000000_0001111110110111_1111101111111111"; -- 0.12390112858485994
	pesos_i(16821) := b"1111111111111111_1111111111111111_1111011100000110_0111011011011111"; -- -0.035057612013611135
	pesos_i(16822) := b"1111111111111111_1111111111111111_1111111110001111_0101101100111111"; -- -0.0017188045585633954
	pesos_i(16823) := b"1111111111111111_1111111111111111_1111000111010100_1100011110011101"; -- -0.05534698880875822
	pesos_i(16824) := b"1111111111111111_1111111111111111_1110000010010100_1000101100101001"; -- -0.12273340469155748
	pesos_i(16825) := b"1111111111111111_1111111111111111_1110010000011000_1111000100100110"; -- -0.10899441539215111
	pesos_i(16826) := b"1111111111111111_1111111111111111_1111111001001010_1011111100111101"; -- -0.006671951035168545
	pesos_i(16827) := b"1111111111111111_1111111111111111_1111111000010011_1101110001011101"; -- -0.007509448432217776
	pesos_i(16828) := b"0000000000000000_0000000000000000_0000011101111001_1001111101110010"; -- 0.029199567256415333
	pesos_i(16829) := b"1111111111111111_1111111111111111_1110011110100001_1100100111000101"; -- -0.09518755855206165
	pesos_i(16830) := b"1111111111111111_1111111111111111_1101111111001100_0100110101110111"; -- -0.12578883976228478
	pesos_i(16831) := b"1111111111111111_1111111111111111_1111000010110100_0000000100010011"; -- -0.059753354030387305
	pesos_i(16832) := b"0000000000000000_0000000000000000_0001010011011110_1000110010111001"; -- 0.08152083877955385
	pesos_i(16833) := b"1111111111111111_1111111111111111_1110011011001101_0111101001010000"; -- -0.09842715788284208
	pesos_i(16834) := b"0000000000000000_0000000000000000_0000000010111100_0101011101111001"; -- 0.0028738661826251716
	pesos_i(16835) := b"1111111111111111_1111111111111111_1110000111101010_0011111001010000"; -- -0.1175194792688333
	pesos_i(16836) := b"0000000000000000_0000000000000000_0001001010001010_0010001011101110"; -- 0.07242029480307242
	pesos_i(16837) := b"1111111111111111_1111111111111111_1111110000000110_1011110001011101"; -- -0.015522220042035163
	pesos_i(16838) := b"0000000000000000_0000000000000000_0000010111111010_1100001110000001"; -- 0.023357600180597373
	pesos_i(16839) := b"1111111111111111_1111111111111111_1101101000100101_0101100001111000"; -- -0.1478676517088505
	pesos_i(16840) := b"1111111111111111_1111111111111111_1110001100101100_1000011101111010"; -- -0.11260178824051277
	pesos_i(16841) := b"1111111111111111_1111111111111111_1110110111011011_0100011101010001"; -- -0.07087282435508775
	pesos_i(16842) := b"1111111111111111_1111111111111111_1110100111011111_1100001000101101"; -- -0.08642946629484319
	pesos_i(16843) := b"1111111111111111_1111111111111111_1111000001010010_0100110001101001"; -- -0.061244224816400517
	pesos_i(16844) := b"1111111111111111_1111111111111111_1111011000111000_0010010010001101"; -- -0.038205829319740175
	pesos_i(16845) := b"0000000000000000_0000000000000000_0010011111100101_1001100001111001"; -- 0.15584710078220282
	pesos_i(16846) := b"1111111111111111_1111111111111111_1110100101100111_1100100010000010"; -- -0.08826014351620831
	pesos_i(16847) := b"1111111111111111_1111111111111111_1110100111001011_1000001100000001"; -- -0.0867384073206342
	pesos_i(16848) := b"1111111111111111_1111111111111111_1110001000011101_1010000101000101"; -- -0.11673538259117867
	pesos_i(16849) := b"0000000000000000_0000000000000000_0000110111010110_1010011101010100"; -- 0.05405660447248092
	pesos_i(16850) := b"1111111111111111_1111111111111111_1101110101010111_1001111110101110"; -- -0.13538171776273933
	pesos_i(16851) := b"0000000000000000_0000000000000000_0001101001101001_0011111101111000"; -- 0.10316845592015783
	pesos_i(16852) := b"1111111111111111_1111111111111111_1110001101001101_0000000001010110"; -- -0.1121063032477123
	pesos_i(16853) := b"1111111111111111_1111111111111111_1110001011000110_1001000001101001"; -- -0.11415765215058143
	pesos_i(16854) := b"1111111111111111_1111111111111111_1110010011000000_1011010011100010"; -- -0.10643453114752012
	pesos_i(16855) := b"1111111111111111_1111111111111111_1111010110110010_1101000011001100"; -- -0.040240240392839674
	pesos_i(16856) := b"0000000000000000_0000000000000000_0001010101111001_0010101100010001"; -- 0.08388013033075865
	pesos_i(16857) := b"1111111111111111_1111111111111111_1111010001001101_1000111000101111"; -- -0.04569159838273201
	pesos_i(16858) := b"0000000000000000_0000000000000000_0010001010100110_1001000000011110"; -- 0.13535404905605522
	pesos_i(16859) := b"0000000000000000_0000000000000000_0000101001001101_0100101110101010"; -- 0.04024193674868912
	pesos_i(16860) := b"0000000000000000_0000000000000000_0001100010111010_0011100110110101"; -- 0.09659157437507335
	pesos_i(16861) := b"0000000000000000_0000000000000000_0001000000100100_0110010001100001"; -- 0.06305529942330607
	pesos_i(16862) := b"1111111111111111_1111111111111111_1111011101101111_1100011100111101"; -- -0.03345064887321427
	pesos_i(16863) := b"1111111111111111_1111111111111111_1101111001110111_0011101000000110"; -- -0.13099324555248942
	pesos_i(16864) := b"1111111111111111_1111111111111111_1110110010010010_1110010111110110"; -- -0.07588351015091685
	pesos_i(16865) := b"1111111111111111_1111111111111111_1111100110100111_0000110111101001"; -- -0.02479470322304468
	pesos_i(16866) := b"1111111111111111_1111111111111111_1110110000010100_1111111001010101"; -- -0.07780466494347278
	pesos_i(16867) := b"0000000000000000_0000000000000000_0001111011101101_0011111111001000"; -- 0.12080763465288637
	pesos_i(16868) := b"1111111111111111_1111111111111111_1111010001100001_1000010111100010"; -- -0.045386917361078846
	pesos_i(16869) := b"1111111111111111_1111111111111111_1101110101011010_0010100010010110"; -- -0.13534303998201605
	pesos_i(16870) := b"1111111111111111_1111111111111111_1111101000000010_1011000101001100"; -- -0.02339641471872067
	pesos_i(16871) := b"0000000000000000_0000000000000000_0000111100011011_1100001100111001"; -- 0.05901737349824281
	pesos_i(16872) := b"0000000000000000_0000000000000000_0000110100011011_0110011110011011"; -- 0.05119941259603536
	pesos_i(16873) := b"0000000000000000_0000000000000000_0001011110000101_0001111000101000"; -- 0.09187496646224941
	pesos_i(16874) := b"1111111111111111_1111111111111111_1110000010001010_0100010010000110"; -- -0.12289020274096613
	pesos_i(16875) := b"0000000000000000_0000000000000000_0010101000011100_1010101010011011"; -- 0.16449991492362043
	pesos_i(16876) := b"0000000000000000_0000000000000000_0010001110101111_0110000011000000"; -- 0.13939480492718187
	pesos_i(16877) := b"0000000000000000_0000000000000000_0001111101010101_1011111101010101"; -- 0.12240215138151926
	pesos_i(16878) := b"1111111111111111_1111111111111111_1101011110011010_0000000100011100"; -- -0.15780633025886032
	pesos_i(16879) := b"1111111111111111_1111111111111111_1111100101011101_0100000000111010"; -- -0.025920854328594083
	pesos_i(16880) := b"1111111111111111_1111111111111111_1101111001101010_1001001110110101"; -- -0.13118626422229224
	pesos_i(16881) := b"0000000000000000_0000000000000000_0001110010001110_1000010100000000"; -- 0.11154967546639241
	pesos_i(16882) := b"1111111111111111_1111111111111111_1101101101001101_1101110100000110"; -- -0.1433431493118839
	pesos_i(16883) := b"1111111111111111_1111111111111111_1101110011000101_0100101101110111"; -- -0.1376145205194847
	pesos_i(16884) := b"1111111111111111_1111111111111111_1110011111001011_0010101111110000"; -- -0.09455609698156371
	pesos_i(16885) := b"1111111111111111_1111111111111111_1101101011001001_0011100001000011"; -- -0.14536712997546006
	pesos_i(16886) := b"1111111111111111_1111111111111111_1110000110000000_1001110010100101"; -- -0.11913128831633453
	pesos_i(16887) := b"0000000000000000_0000000000000000_0001011101011100_1000010101001111"; -- 0.09125550432267174
	pesos_i(16888) := b"0000000000000000_0000000000000000_0001101010000000_0010001000010110"; -- 0.10351765673887964
	pesos_i(16889) := b"0000000000000000_0000000000000000_0001001001011111_1010111001111011"; -- 0.07177248490151202
	pesos_i(16890) := b"0000000000000000_0000000000000000_0000111000100111_0100110100110001"; -- 0.05528719381338199
	pesos_i(16891) := b"0000000000000000_0000000000000000_0000001001100001_1011011000011001"; -- 0.009303456475934122
	pesos_i(16892) := b"0000000000000000_0000000000000000_0010000101001101_0100100010001010"; -- 0.1300855004173956
	pesos_i(16893) := b"1111111111111111_1111111111111111_1110100001111011_0100010111111001"; -- -0.09186899822070789
	pesos_i(16894) := b"1111111111111111_1111111111111111_1110010110000111_0001100110101000"; -- -0.1034072841849703
	pesos_i(16895) := b"1111111111111111_1111111111111111_1110111100100011_1110000100011110"; -- -0.06585877430884972
	pesos_i(16896) := b"0000000000000000_0000000000000000_0000000110011100_1000011101000001"; -- 0.0062946827842607
	pesos_i(16897) := b"1111111111111111_1111111111111111_1110110100000110_1001111011100110"; -- -0.07411772626768427
	pesos_i(16898) := b"0000000000000000_0000000000000000_0000010101100110_1000001111001010"; -- 0.021095501810644623
	pesos_i(16899) := b"0000000000000000_0000000000000000_0010000110001111_1111101100001110"; -- 0.13110322082232936
	pesos_i(16900) := b"1111111111111111_1111111111111111_1110000100111001_0110010000010101"; -- -0.1202180336346232
	pesos_i(16901) := b"0000000000000000_0000000000000000_0000010011100011_0001110110010010"; -- 0.019090507560449093
	pesos_i(16902) := b"0000000000000000_0000000000000000_0010000100011001_0110110011010100"; -- 0.12929420645070805
	pesos_i(16903) := b"0000000000000000_0000000000000000_0001011001100111_0011010101101110"; -- 0.0875123399836563
	pesos_i(16904) := b"0000000000000000_0000000000000000_0000100101100110_0100111111010111"; -- 0.03671740525430449
	pesos_i(16905) := b"1111111111111111_1111111111111111_1110010101110011_0000100000111110"; -- -0.1037134980189097
	pesos_i(16906) := b"0000000000000000_0000000000000000_0000100110101110_0110010110101010"; -- 0.03781733897628711
	pesos_i(16907) := b"0000000000000000_0000000000000000_0010010001001011_0100010101111100"; -- 0.14177355073148099
	pesos_i(16908) := b"1111111111111111_1111111111111111_1111000000000010_0111101010000111"; -- -0.062462179263515466
	pesos_i(16909) := b"1111111111111111_1111111111111111_1110101100000110_1000011111100011"; -- -0.08193159777797805
	pesos_i(16910) := b"1111111111111111_1111111111111111_1110111000111110_0110111001100111"; -- -0.06935987452533539
	pesos_i(16911) := b"0000000000000000_0000000000000000_0001001001001100_0101111010010011"; -- 0.07147780496272027
	pesos_i(16912) := b"1111111111111111_1111111111111111_1111001010001101_0111010010010011"; -- -0.052529062455362735
	pesos_i(16913) := b"0000000000000000_0000000000000000_0000001010110011_1001000001010101"; -- 0.010552426065291364
	pesos_i(16914) := b"0000000000000000_0000000000000000_0001000010000111_1000100111011010"; -- 0.06456815301156504
	pesos_i(16915) := b"1111111111111111_1111111111111111_1110100101100101_1111101001101101"; -- -0.08828768568161234
	pesos_i(16916) := b"1111111111111111_1111111111111111_1110111001111101_1010101001010001"; -- -0.06839499969818623
	pesos_i(16917) := b"1111111111111111_1111111111111111_1111101001111110_1100110000001100"; -- -0.02150273044373832
	pesos_i(16918) := b"0000000000000000_0000000000000000_0001100110001111_0111110010111110"; -- 0.09984569204658193
	pesos_i(16919) := b"0000000000000000_0000000000000000_0000010111100111_0101110010110001"; -- 0.023061555224469753
	pesos_i(16920) := b"1111111111111111_1111111111111111_1110100011111011_0101110100110000"; -- -0.08991448950559679
	pesos_i(16921) := b"1111111111111111_1111111111111111_1101101111110111_0011110110110000"; -- -0.14075865216005992
	pesos_i(16922) := b"0000000000000000_0000000000000000_0001010111010011_1110100111000110"; -- 0.08526478837320313
	pesos_i(16923) := b"1111111111111111_1111111111111111_1111100110111011_0100101010111010"; -- -0.024485902322424535
	pesos_i(16924) := b"1111111111111111_1111111111111111_1110010010100010_0100101101000001"; -- -0.10689859076761439
	pesos_i(16925) := b"1111111111111111_1111111111111111_1101110100011010_0101110110001111"; -- -0.13631644503037327
	pesos_i(16926) := b"0000000000000000_0000000000000000_0010010001110011_0000100001111000"; -- 0.1423802655029675
	pesos_i(16927) := b"0000000000000000_0000000000000000_0001000011011011_0111011010010100"; -- 0.06584874253198844
	pesos_i(16928) := b"0000000000000000_0000000000000000_0000100101110100_0001101010100110"; -- 0.03692785798097057
	pesos_i(16929) := b"1111111111111111_1111111111111111_1111001010011011_0011100111000011"; -- -0.052318944941903735
	pesos_i(16930) := b"1111111111111111_1111111111111111_1111001000101001_0010001110010010"; -- -0.05405976938574806
	pesos_i(16931) := b"0000000000000000_0000000000000000_0000111100111010_1101011000011111"; -- 0.05949152246556216
	pesos_i(16932) := b"1111111111111111_1111111111111111_1111110101010100_0101001110100101"; -- -0.010432026096867483
	pesos_i(16933) := b"0000000000000000_0000000000000000_0000111100100110_1110011101101101"; -- 0.05918737799987485
	pesos_i(16934) := b"0000000000000000_0000000000000000_0001000000100000_0010111100110101"; -- 0.06299109509220215
	pesos_i(16935) := b"0000000000000000_0000000000000000_0001010110000110_1001101011111001"; -- 0.08408516486036433
	pesos_i(16936) := b"0000000000000000_0000000000000000_0010001001101110_1011000111111101"; -- 0.13450157572224006
	pesos_i(16937) := b"0000000000000000_0000000000000000_0001110010001111_0100001001110001"; -- 0.11156096705262354
	pesos_i(16938) := b"0000000000000000_0000000000000000_0000000100100001_1111110101011110"; -- 0.004424891821536933
	pesos_i(16939) := b"0000000000000000_0000000000000000_0001100110101010_0011100010001100"; -- 0.10025361448467741
	pesos_i(16940) := b"0000000000000000_0000000000000000_0010010001000010_1110010000101000"; -- 0.1416456792541079
	pesos_i(16941) := b"1111111111111111_1111111111111111_1110101000100111_0001000010000110"; -- -0.08534142242572018
	pesos_i(16942) := b"1111111111111111_1111111111111111_1110000110100110_1010110001110100"; -- -0.11855051207406161
	pesos_i(16943) := b"1111111111111111_1111111111111111_1111111000011101_0000011101110011"; -- -0.007369551011884394
	pesos_i(16944) := b"0000000000000000_0000000000000000_0010001000101001_0001010101101100"; -- 0.13343938715492767
	pesos_i(16945) := b"1111111111111111_1111111111111111_1110011010001101_0101001111010101"; -- -0.09940601403936526
	pesos_i(16946) := b"1111111111111111_1111111111111111_1110011111011110_1111010100100100"; -- -0.09425418742046134
	pesos_i(16947) := b"1111111111111111_1111111111111111_1111011011000010_1000010010101101"; -- -0.0360943869024691
	pesos_i(16948) := b"1111111111111111_1111111111111111_1111100100110110_0110011100001000"; -- -0.02651363416055283
	pesos_i(16949) := b"1111111111111111_1111111111111111_1110110101000110_0111101101011010"; -- -0.07314328243374793
	pesos_i(16950) := b"0000000000000000_0000000000000000_0010000011101011_1111011011011011"; -- 0.12860052910569864
	pesos_i(16951) := b"0000000000000000_0000000000000000_0000100010110100_0011111110111100"; -- 0.03400038084074175
	pesos_i(16952) := b"0000000000000000_0000000000000000_0010011000110101_0011011100010111"; -- 0.1492494994384785
	pesos_i(16953) := b"0000000000000000_0000000000000000_0001001101101011_1111111110100101"; -- 0.07586667793532266
	pesos_i(16954) := b"0000000000000000_0000000000000000_0000000111100100_0110000011100100"; -- 0.00739102903239237
	pesos_i(16955) := b"1111111111111111_1111111111111111_1101100101111010_0111111100100010"; -- -0.1504746001301416
	pesos_i(16956) := b"1111111111111111_1111111111111111_1110110010010010_0111110010010110"; -- -0.07588979081719635
	pesos_i(16957) := b"1111111111111111_1111111111111111_1110000010000111_1111110110101011"; -- -0.12292494376969024
	pesos_i(16958) := b"0000000000000000_0000000000000000_0010000100100010_0000101110101101"; -- 0.1294257448384625
	pesos_i(16959) := b"0000000000000000_0000000000000000_0000001011000011_1111001111001111"; -- 0.010802495922426941
	pesos_i(16960) := b"1111111111111111_1111111111111111_1110111011100111_1100011011111011"; -- -0.06677585954141159
	pesos_i(16961) := b"1111111111111111_1111111111111111_1110001001101011_1001011100011000"; -- -0.11554580366749514
	pesos_i(16962) := b"1111111111111111_1111111111111111_1111101111001001_0100010000001000"; -- -0.01646017831942449
	pesos_i(16963) := b"1111111111111111_1111111111111111_1110000110000100_0111110110101110"; -- -0.11907209877320345
	pesos_i(16964) := b"1111111111111111_1111111111111111_1101101100111100_0010011011110111"; -- -0.1436134001944323
	pesos_i(16965) := b"1111111111111111_1111111111111111_1111101110111000_0000011101010110"; -- -0.016723195474382634
	pesos_i(16966) := b"0000000000000000_0000000000000000_0010010000010110_1000110100101111"; -- 0.14096910849028646
	pesos_i(16967) := b"1111111111111111_1111111111111111_1111010111011110_0110001110110001"; -- -0.03957535668878465
	pesos_i(16968) := b"1111111111111111_1111111111111111_1110101001100000_0101011101110111"; -- -0.08446744285578069
	pesos_i(16969) := b"1111111111111111_1111111111111111_1110110110110000_1101011000010111"; -- -0.0715204422605718
	pesos_i(16970) := b"1111111111111111_1111111111111111_1111010100000000_0001111111010100"; -- -0.042966852780487834
	pesos_i(16971) := b"1111111111111111_1111111111111111_1111111000111010_1100111010001001"; -- -0.006915179719636447
	pesos_i(16972) := b"0000000000000000_0000000000000000_0001001010010101_0110001111110111"; -- 0.07259201785748433
	pesos_i(16973) := b"0000000000000000_0000000000000000_0000101001000011_1001011100111110"; -- 0.040093853540373994
	pesos_i(16974) := b"1111111111111111_1111111111111111_1111011011110101_0101110011111011"; -- -0.03531855471449007
	pesos_i(16975) := b"1111111111111111_1111111111111111_1110111000100010_1001001001010011"; -- -0.06978497961941095
	pesos_i(16976) := b"0000000000000000_0000000000000000_0000010010110011_0010101001101100"; -- 0.018358851881854682
	pesos_i(16977) := b"1111111111111111_1111111111111111_1110100010111111_1001010010000011"; -- -0.09082671931219873
	pesos_i(16978) := b"0000000000000000_0000000000000000_0001101111000011_0111010010111001"; -- 0.10845117102465739
	pesos_i(16979) := b"1111111111111111_1111111111111111_1110111010011111_1100110101111101"; -- -0.06787410437077425
	pesos_i(16980) := b"1111111111111111_1111111111111111_1111011011001111_1000101001011101"; -- -0.035895683522613284
	pesos_i(16981) := b"0000000000000000_0000000000000000_0001010011000101_1001011100001101"; -- 0.08113998466662735
	pesos_i(16982) := b"1111111111111111_1111111111111111_1110011101101111_1001110011000110"; -- -0.09595318007152713
	pesos_i(16983) := b"0000000000000000_0000000000000000_0001111001001000_1000001101001101"; -- 0.1182939589009158
	pesos_i(16984) := b"1111111111111111_1111111111111111_1111010000001111_1111110011010100"; -- -0.04663104851835354
	pesos_i(16985) := b"1111111111111111_1111111111111111_1110110111001110_0000101110000111"; -- -0.07107475246702157
	pesos_i(16986) := b"1111111111111111_1111111111111111_1110110000111111_1010000100110010"; -- -0.07715408836030989
	pesos_i(16987) := b"1111111111111111_1111111111111111_1110100001011010_1111011111110011"; -- -0.09236193013473627
	pesos_i(16988) := b"0000000000000000_0000000000000000_0001000001000000_0001100000101111"; -- 0.06347800403620855
	pesos_i(16989) := b"0000000000000000_0000000000000000_0000001111111010_1011000110001011"; -- 0.01554402976739877
	pesos_i(16990) := b"1111111111111111_1111111111111111_1111101011011001_0011010100000101"; -- -0.02012318264801191
	pesos_i(16991) := b"0000000000000000_0000000000000000_0000111011001011_1000000100000101"; -- 0.057792724388886274
	pesos_i(16992) := b"1111111111111111_1111111111111111_1110010101100000_1110110011011010"; -- -0.10398978882797336
	pesos_i(16993) := b"0000000000000000_0000000000000000_0000101011000110_0000100100101011"; -- 0.04208428674235245
	pesos_i(16994) := b"1111111111111111_1111111111111111_1110100100011001_1110001001100010"; -- -0.08944878691388494
	pesos_i(16995) := b"0000000000000000_0000000000000000_0000111011001100_1000000010000100"; -- 0.05780795302429155
	pesos_i(16996) := b"0000000000000000_0000000000000000_0001001101100000_1100110011101110"; -- 0.07569580853615321
	pesos_i(16997) := b"1111111111111111_1111111111111111_1111011010110111_1111101010101100"; -- -0.036255200314093516
	pesos_i(16998) := b"1111111111111111_1111111111111111_1111110000010000_1001010000111110"; -- -0.015372023411420554
	pesos_i(16999) := b"0000000000000000_0000000000000000_0010011001100001_0000100011000010"; -- 0.14991812446479222
	pesos_i(17000) := b"0000000000000000_0000000000000000_0001101010111110_1001111000100011"; -- 0.10447109556811048
	pesos_i(17001) := b"1111111111111111_1111111111111111_1111110101101101_0110001000000000"; -- -0.010049700660332226
	pesos_i(17002) := b"0000000000000000_0000000000000000_0001010001001111_1100100101010011"; -- 0.07934244422134269
	pesos_i(17003) := b"0000000000000000_0000000000000000_0001111111011001_1101011001010011"; -- 0.12441768200609987
	pesos_i(17004) := b"1111111111111111_1111111111111111_1110011010000000_1110000000101111"; -- -0.09959601262183089
	pesos_i(17005) := b"0000000000000000_0000000000000000_0001000100011101_1000011000001010"; -- 0.06685674433388851
	pesos_i(17006) := b"1111111111111111_1111111111111111_1111011111011000_1010101010101011"; -- -0.03185017898750728
	pesos_i(17007) := b"0000000000000000_0000000000000000_0001100001100110_0101111000000101"; -- 0.09531200045828375
	pesos_i(17008) := b"1111111111111111_1111111111111111_1111011000011011_0110001111010101"; -- -0.03864456220492875
	pesos_i(17009) := b"0000000000000000_0000000000000000_0000100101000110_1111011110000100"; -- 0.03623911842782338
	pesos_i(17010) := b"0000000000000000_0000000000000000_0001000011011001_1100010000000110"; -- 0.06582284121485364
	pesos_i(17011) := b"1111111111111111_1111111111111111_1110011001101101_0101011011100100"; -- -0.0998941129306466
	pesos_i(17012) := b"0000000000000000_0000000000000000_0001100110100000_0111111000100001"; -- 0.10010517417954409
	pesos_i(17013) := b"0000000000000000_0000000000000000_0001000001100111_1000110101110111"; -- 0.06408008716159076
	pesos_i(17014) := b"0000000000000000_0000000000000000_0001010111010010_1110111000100010"; -- 0.08524978961516909
	pesos_i(17015) := b"1111111111111111_1111111111111111_1111110011000000_1011100100101011"; -- -0.012684275597082384
	pesos_i(17016) := b"1111111111111111_1111111111111111_1111010111001011_0001111111111000"; -- -0.039869310247980065
	pesos_i(17017) := b"1111111111111111_1111111111111111_1110101011001101_0111101000101010"; -- -0.08280216678294637
	pesos_i(17018) := b"0000000000000000_0000000000000000_0000011010110110_0001011110110000"; -- 0.02621601153314328
	pesos_i(17019) := b"1111111111111111_1111111111111111_1111101101110010_0111110101110111"; -- -0.01778426968881988
	pesos_i(17020) := b"1111111111111111_1111111111111111_1110000000110011_1111001100101000"; -- -0.12420730854695097
	pesos_i(17021) := b"0000000000000000_0000000000000000_0000100110010101_1101001100110111"; -- 0.037442399026316395
	pesos_i(17022) := b"1111111111111111_1111111111111111_1110011101110000_1100010010111111"; -- -0.09593553854922807
	pesos_i(17023) := b"1111111111111111_1111111111111111_1101100010011100_0111100101011110"; -- -0.1538623947502319
	pesos_i(17024) := b"0000000000000000_0000000000000000_0010001101100101_1001001101111000"; -- 0.13826867745184543
	pesos_i(17025) := b"1111111111111111_1111111111111111_1111100001000110_0100101101000001"; -- -0.030177399179761286
	pesos_i(17026) := b"1111111111111111_1111111111111111_1111111000111100_1101011001001100"; -- -0.006884199669928418
	pesos_i(17027) := b"0000000000000000_0000000000000000_0010001000100001_1010011100101000"; -- 0.13332600339972536
	pesos_i(17028) := b"1111111111111111_1111111111111111_1101110001111001_1010100101110011"; -- -0.13876858646408888
	pesos_i(17029) := b"1111111111111111_1111111111111111_1111000111011110_0010000011011111"; -- -0.05520433960355925
	pesos_i(17030) := b"0000000000000000_0000000000000000_0000101100110100_1110110100000001"; -- 0.04377633364754105
	pesos_i(17031) := b"0000000000000000_0000000000000000_0010100010010110_1111001001101001"; -- 0.15855326715642992
	pesos_i(17032) := b"0000000000000000_0000000000000000_0000011001100110_1011101010000011"; -- 0.025005013343747315
	pesos_i(17033) := b"0000000000000000_0000000000000000_0000000101000110_1100100101000100"; -- 0.004986361503792193
	pesos_i(17034) := b"0000000000000000_0000000000000000_0000100011110110_1111001001010001"; -- 0.0350181051940568
	pesos_i(17035) := b"1111111111111111_1111111111111111_1110001101010000_0101000010010101"; -- -0.11205574383652046
	pesos_i(17036) := b"0000000000000000_0000000000000000_0000110111110111_0011101001100011"; -- 0.05455365107916128
	pesos_i(17037) := b"0000000000000000_0000000000000000_0000110110001101_0101100110000010"; -- 0.0529380744546394
	pesos_i(17038) := b"1111111111111111_1111111111111111_1110100100110101_0110101000000110"; -- -0.08902871464539226
	pesos_i(17039) := b"0000000000000000_0000000000000000_0000010110010001_0100001000100100"; -- 0.02174771663190689
	pesos_i(17040) := b"0000000000000000_0000000000000000_0000011000100001_1111110110001111"; -- 0.023956153355504883
	pesos_i(17041) := b"0000000000000000_0000000000000000_0000100111001110_0000011011100100"; -- 0.03829997119152488
	pesos_i(17042) := b"0000000000000000_0000000000000000_0000000001001110_0011111000011010"; -- 0.0011938871088563725
	pesos_i(17043) := b"0000000000000000_0000000000000000_0000010111001000_0101110001111000"; -- 0.022588519420898685
	pesos_i(17044) := b"1111111111111111_1111111111111111_1110101011101101_1110001100100010"; -- -0.08230762871397583
	pesos_i(17045) := b"1111111111111111_1111111111111111_1111100011100001_1010010110100000"; -- -0.027806900372331588
	pesos_i(17046) := b"0000000000000000_0000000000000000_0000001010110111_0001111101101101"; -- 0.010606731478913275
	pesos_i(17047) := b"0000000000000000_0000000000000000_0000100111011001_1000101110000001"; -- 0.03847572224773509
	pesos_i(17048) := b"0000000000000000_0000000000000000_0000111111101111_1000001110001111"; -- 0.06224844210162471
	pesos_i(17049) := b"0000000000000000_0000000000000000_0001000010011011_0000010110010011"; -- 0.06486544458147504
	pesos_i(17050) := b"0000000000000000_0000000000000000_0001011011110110_0111110101101010"; -- 0.08969863737055753
	pesos_i(17051) := b"1111111111111111_1111111111111111_1111000011110011_0000011101110111"; -- -0.058791669305559235
	pesos_i(17052) := b"1111111111111111_1111111111111111_1101110101101000_1101101011101100"; -- -0.1351187871223364
	pesos_i(17053) := b"1111111111111111_1111111111111111_1110101001101001_1100100001100100"; -- -0.08432338302843045
	pesos_i(17054) := b"1111111111111111_1111111111111111_1111111111111010_0010000000011101"; -- -8.963867890573501e-05
	pesos_i(17055) := b"1111111111111111_1111111111111111_1111011010110111_1100000110101000"; -- -0.0362585987737636
	pesos_i(17056) := b"0000000000000000_0000000000000000_0001100010000000_0101010101111101"; -- 0.09570822052687188
	pesos_i(17057) := b"0000000000000000_0000000000000000_0010011111001111_1001101011101010"; -- 0.15551155291564794
	pesos_i(17058) := b"1111111111111111_1111111111111111_1110110010100001_1011000111001110"; -- -0.07565773694924238
	pesos_i(17059) := b"1111111111111111_1111111111111111_1110011100011101_0100000011001011"; -- -0.09720988316907915
	pesos_i(17060) := b"1111111111111111_1111111111111111_1110000111000000_0000011000110010"; -- -0.11816369330388543
	pesos_i(17061) := b"0000000000000000_0000000000000000_0001101101111000_1100101111011101"; -- 0.10731195594182207
	pesos_i(17062) := b"0000000000000000_0000000000000000_0010011110101010_1101111010100001"; -- 0.15495101383677076
	pesos_i(17063) := b"0000000000000000_0000000000000000_0010010111110100_1110011000001001"; -- 0.1482681057312134
	pesos_i(17064) := b"0000000000000000_0000000000000000_0000100110000010_1000010110111110"; -- 0.03714786419009964
	pesos_i(17065) := b"1111111111111111_1111111111111111_1101110111010101_1010010101000001"; -- -0.13345877798509906
	pesos_i(17066) := b"0000000000000000_0000000000000000_0010001100010011_0000111100101001"; -- 0.13700957057537555
	pesos_i(17067) := b"0000000000000000_0000000000000000_0001110101010110_0000001000111010"; -- 0.1145936386831057
	pesos_i(17068) := b"0000000000000000_0000000000000000_0001101000100101_0000010010011010"; -- 0.10212734958553743
	pesos_i(17069) := b"1111111111111111_1111111111111111_1110110100110100_1100001101011001"; -- -0.0734136492667704
	pesos_i(17070) := b"1111111111111111_1111111111111111_1111111000100110_0100100111110000"; -- -0.00722825889556551
	pesos_i(17071) := b"0000000000000000_0000000000000000_0001000000110001_1101000000100100"; -- 0.06326008670134697
	pesos_i(17072) := b"0000000000000000_0000000000000000_0001000000100111_1001100101001111"; -- 0.06310423059291691
	pesos_i(17073) := b"1111111111111111_1111111111111111_1110101111010000_0000111000100110"; -- -0.07885657853207421
	pesos_i(17074) := b"0000000000000000_0000000000000000_0001101100011010_0000001001010100"; -- 0.10586561730803028
	pesos_i(17075) := b"1111111111111111_1111111111111111_1110101011101110_1110000001011111"; -- -0.0822925345429267
	pesos_i(17076) := b"1111111111111111_1111111111111111_1110101000001100_1011000011101000"; -- -0.08574385015957948
	pesos_i(17077) := b"1111111111111111_1111111111111111_1110101111000000_1100001001111001"; -- -0.07908997099633366
	pesos_i(17078) := b"0000000000000000_0000000000000000_0000111111000101_0110010100010011"; -- 0.061605756004044075
	pesos_i(17079) := b"1111111111111111_1111111111111111_1111100000101000_1100001010101100"; -- -0.03062804514013026
	pesos_i(17080) := b"0000000000000000_0000000000000000_0010001001101001_0101010111100110"; -- 0.1344197928984017
	pesos_i(17081) := b"0000000000000000_0000000000000000_0010011011100101_1011010011110000"; -- 0.1519425474924545
	pesos_i(17082) := b"1111111111111111_1111111111111111_1111100011111100_1111111000111010"; -- -0.02738963202900002
	pesos_i(17083) := b"1111111111111111_1111111111111111_1111010000111000_0111000011001101"; -- -0.04601378427919271
	pesos_i(17084) := b"0000000000000000_0000000000000000_0001000011000110_1100000001011000"; -- 0.06553270472902373
	pesos_i(17085) := b"1111111111111111_1111111111111111_1110001011101111_0101110110011010"; -- -0.11353507040626826
	pesos_i(17086) := b"1111111111111111_1111111111111111_1110110011111111_1110000001010101"; -- -0.07422063751231331
	pesos_i(17087) := b"1111111111111111_1111111111111111_1110011111111011_0010110100111110"; -- -0.09382359739282956
	pesos_i(17088) := b"1111111111111111_1111111111111111_1110001101100100_0001011010100111"; -- -0.11175402100940665
	pesos_i(17089) := b"0000000000000000_0000000000000000_0000011111110101_1111100100100111"; -- 0.031097004073147947
	pesos_i(17090) := b"1111111111111111_1111111111111111_1110111001011111_0010101010011001"; -- -0.06886037599039961
	pesos_i(17091) := b"0000000000000000_0000000000000000_0010000101100100_1111111010110110"; -- 0.13044731086665246
	pesos_i(17092) := b"1111111111111111_1111111111111111_1111010001100011_0101000001000001"; -- -0.045359596423889405
	pesos_i(17093) := b"1111111111111111_1111111111111111_1111111010100001_1101000010011110"; -- -0.005343400418597215
	pesos_i(17094) := b"1111111111111111_1111111111111111_1111110001000001_0011001001100110"; -- -0.014630174839434783
	pesos_i(17095) := b"0000000000000000_0000000000000000_0001100110010101_1010000110101010"; -- 0.09993944541155428
	pesos_i(17096) := b"1111111111111111_1111111111111111_1111100001111111_1110010000100011"; -- -0.02929853576986548
	pesos_i(17097) := b"0000000000000000_0000000000000000_0001101101000100_0111101010001111"; -- 0.10651365274870792
	pesos_i(17098) := b"1111111111111111_1111111111111111_1111000010001100_1101111010010100"; -- -0.06035050277497344
	pesos_i(17099) := b"0000000000000000_0000000000000000_0000000000100100_1101111010111011"; -- 0.0005625922497827079
	pesos_i(17100) := b"1111111111111111_1111111111111111_1110111001111100_1101101011111110"; -- -0.0684073573153258
	pesos_i(17101) := b"0000000000000000_0000000000000000_0010001101100011_1100101010010110"; -- 0.1382414451323876
	pesos_i(17102) := b"1111111111111111_1111111111111111_1110011111110111_0100011110111000"; -- -0.09388305430414999
	pesos_i(17103) := b"1111111111111111_1111111111111111_1101111001000101_0111110100100110"; -- -0.13175218423154192
	pesos_i(17104) := b"1111111111111111_1111111111111111_1111111010010000_1000010010110101"; -- -0.0056073244087843895
	pesos_i(17105) := b"0000000000000000_0000000000000000_0010001101100100_0111100001111000"; -- 0.13825180946867102
	pesos_i(17106) := b"1111111111111111_1111111111111111_1111111110100000_1000010100010001"; -- -0.0014569124241963715
	pesos_i(17107) := b"0000000000000000_0000000000000000_0000000100101100_1111000011011010"; -- 0.00459199266463146
	pesos_i(17108) := b"1111111111111111_1111111111111111_1110101001110100_1111000110111001"; -- -0.08415307265767907
	pesos_i(17109) := b"0000000000000000_0000000000000000_0001111110110110_1110010000111100"; -- 0.12388445349772897
	pesos_i(17110) := b"0000000000000000_0000000000000000_0001100111111010_1110000001010100"; -- 0.10148431820530858
	pesos_i(17111) := b"0000000000000000_0000000000000000_0010011011010001_0111011100101010"; -- 0.1516336897122577
	pesos_i(17112) := b"1111111111111111_1111111111111111_1111010011011011_0110100010001111"; -- -0.0435270929699468
	pesos_i(17113) := b"1111111111111111_1111111111111111_1110000011000110_0010111010110000"; -- -0.12197597697098737
	pesos_i(17114) := b"0000000000000000_0000000000000000_0000010111011010_1000100011100011"; -- 0.02286582513177166
	pesos_i(17115) := b"1111111111111111_1111111111111111_1111110100101010_1010001001100011"; -- -0.011068201891804486
	pesos_i(17116) := b"1111111111111111_1111111111111111_1111011100000110_1110110010101010"; -- -0.035050591089802935
	pesos_i(17117) := b"1111111111111111_1111111111111111_1110110000010101_1101011101110001"; -- -0.07779172408352088
	pesos_i(17118) := b"1111111111111111_1111111111111111_1110000101001001_0111101010111010"; -- -0.11997254327535001
	pesos_i(17119) := b"1111111111111111_1111111111111111_1111100100011110_1111110110000011"; -- -0.026870875774199474
	pesos_i(17120) := b"1111111111111111_1111111111111111_1111100111100000_1100001010001100"; -- -0.02391418539543854
	pesos_i(17121) := b"1111111111111111_1111111111111111_1101110111101011_1000100110000100"; -- -0.1331247379401239
	pesos_i(17122) := b"1111111111111111_1111111111111111_1110010011110011_0101000010100000"; -- -0.1056623087052517
	pesos_i(17123) := b"0000000000000000_0000000000000000_0001000110011001_1011100010001111"; -- 0.06875184528078125
	pesos_i(17124) := b"1111111111111111_1111111111111111_1101100111000101_1000100101111001"; -- -0.14932957448331566
	pesos_i(17125) := b"1111111111111111_1111111111111111_1111010011001110_0111001111110100"; -- -0.04372477800787575
	pesos_i(17126) := b"1111111111111111_1111111111111111_1110110111000000_0011111001010001"; -- -0.07128534820551735
	pesos_i(17127) := b"0000000000000000_0000000000000000_0001100101111000_1100100101000001"; -- 0.09949930038057421
	pesos_i(17128) := b"1111111111111111_1111111111111111_1101111111100101_1001001010111110"; -- -0.12540324072978504
	pesos_i(17129) := b"0000000000000000_0000000000000000_0000010001010011_1011010101111101"; -- 0.01690229714537565
	pesos_i(17130) := b"1111111111111111_1111111111111111_1111110111010010_0000010000011010"; -- -0.00851415981046031
	pesos_i(17131) := b"1111111111111111_1111111111111111_1111000101001101_1100011100011000"; -- -0.05740695634081512
	pesos_i(17132) := b"1111111111111111_1111111111111111_1111001110011111_1100111101110001"; -- -0.048342738098092586
	pesos_i(17133) := b"1111111111111111_1111111111111111_1110001111101001_0110000010001111"; -- -0.10972019671055873
	pesos_i(17134) := b"1111111111111111_1111111111111111_1111110100100110_0111100110100000"; -- -0.011131666676564268
	pesos_i(17135) := b"1111111111111111_1111111111111111_1110101101110100_1011000011011100"; -- -0.08025068894258797
	pesos_i(17136) := b"0000000000000000_0000000000000000_0001100100111011_1001111000011110"; -- 0.0985659430332505
	pesos_i(17137) := b"1111111111111111_1111111111111111_1111001101001101_1110101011001110"; -- -0.04959232768112911
	pesos_i(17138) := b"0000000000000000_0000000000000000_0000110110101011_1001100111111101"; -- 0.053399681427699665
	pesos_i(17139) := b"0000000000000000_0000000000000000_0010010001011001_1010100000001101"; -- 0.14199304888009862
	pesos_i(17140) := b"0000000000000000_0000000000000000_0001001101011001_0010110110000100"; -- 0.07557949513558537
	pesos_i(17141) := b"0000000000000000_0000000000000000_0000000111111011_1100110010100011"; -- 0.007748403451755986
	pesos_i(17142) := b"1111111111111111_1111111111111111_1110011010010011_1011111100000110"; -- -0.09930807215201094
	pesos_i(17143) := b"0000000000000000_0000000000000000_0000011000100001_1101100100000000"; -- 0.023953974263234305
	pesos_i(17144) := b"0000000000000000_0000000000000000_0001111000001011_0011100100000000"; -- 0.11735874425814506
	pesos_i(17145) := b"1111111111111111_1111111111111111_1110110111110111_0101111111110111"; -- -0.0704441092584031
	pesos_i(17146) := b"0000000000000000_0000000000000000_0001100111110110_0011000111100110"; -- 0.10141288635708842
	pesos_i(17147) := b"1111111111111111_1111111111111111_1110001110101110_0000001001010010"; -- -0.11062608233286904
	pesos_i(17148) := b"0000000000000000_0000000000000000_0001010011010100_0011011000011101"; -- 0.08136308862101325
	pesos_i(17149) := b"0000000000000000_0000000000000000_0000000100001000_0100001001111101"; -- 0.004032283344722078
	pesos_i(17150) := b"0000000000000000_0000000000000000_0000111010010111_0001000010111111"; -- 0.05699257526726733
	pesos_i(17151) := b"1111111111111111_1111111111111111_1110010100111111_0101001111110010"; -- -0.10450244273420992
	pesos_i(17152) := b"0000000000000000_0000000000000000_0010000000101001_0000110110101110"; -- 0.12562642571411153
	pesos_i(17153) := b"1111111111111111_1111111111111111_1110100001100001_1010111010101100"; -- -0.09225948631107525
	pesos_i(17154) := b"1111111111111111_1111111111111111_1110111110001111_1111001000110000"; -- -0.06420980772399351
	pesos_i(17155) := b"1111111111111111_1111111111111111_1111100001010010_1010100111101110"; -- -0.029988650732448153
	pesos_i(17156) := b"1111111111111111_1111111111111111_1111111111110011_0110001110001101"; -- -0.00019243063252356548
	pesos_i(17157) := b"0000000000000000_0000000000000000_0000110101110000_1111010110000011"; -- 0.05250486805860182
	pesos_i(17158) := b"1111111111111111_1111111111111111_1110100110010000_0000100011000011"; -- -0.08764596220747947
	pesos_i(17159) := b"0000000000000000_0000000000000000_0001000000011001_1011111000000000"; -- 0.06289279452176677
	pesos_i(17160) := b"0000000000000000_0000000000000000_0001010011110110_0011011000100100"; -- 0.08188188906732362
	pesos_i(17161) := b"1111111111111111_1111111111111111_1111011101001000_1101100110010111"; -- -0.03404464771344827
	pesos_i(17162) := b"1111111111111111_1111111111111111_1111011010101011_1000011100110110"; -- -0.036445187862575536
	pesos_i(17163) := b"1111111111111111_1111111111111111_1101110011011110_0111000110011011"; -- -0.1372307774540459
	pesos_i(17164) := b"0000000000000000_0000000000000000_0000011010010101_1010010101011101"; -- 0.02572091588742699
	pesos_i(17165) := b"1111111111111111_1111111111111111_1101110011001101_0111010100000001"; -- -0.13748997432101512
	pesos_i(17166) := b"1111111111111111_1111111111111111_1111111111011001_1111110101001011"; -- -0.0005799952248578269
	pesos_i(17167) := b"0000000000000000_0000000000000000_0001011010011011_1010111111000110"; -- 0.08831308911953552
	pesos_i(17168) := b"1111111111111111_1111111111111111_1101101001010110_1110000110100101"; -- -0.14711179467996222
	pesos_i(17169) := b"1111111111111111_1111111111111111_1111010110011111_1111001001011110"; -- -0.04052815636044407
	pesos_i(17170) := b"1111111111111111_1111111111111111_1110000110111110_1011000101001101"; -- -0.11818401206867966
	pesos_i(17171) := b"0000000000000000_0000000000000000_0000010000110101_1101111000101011"; -- 0.01644695806775243
	pesos_i(17172) := b"1111111111111111_1111111111111111_1110100101010101_0011011000001110"; -- -0.08854353096418206
	pesos_i(17173) := b"1111111111111111_1111111111111111_1111111111001000_1010000010011010"; -- -0.0008449194947113544
	pesos_i(17174) := b"1111111111111111_1111111111111111_1111100010010001_1010111101001101"; -- -0.029027026848727776
	pesos_i(17175) := b"0000000000000000_0000000000000000_0001101011111000_0111000100100100"; -- 0.10535342339946117
	pesos_i(17176) := b"1111111111111111_1111111111111111_1111000100001010_1001001011101001"; -- -0.05843240546909718
	pesos_i(17177) := b"1111111111111111_1111111111111111_1110011011100010_0110111010100010"; -- -0.09810741948032052
	pesos_i(17178) := b"0000000000000000_0000000000000000_0001001111011101_0011000110011010"; -- 0.07759389889400971
	pesos_i(17179) := b"0000000000000000_0000000000000000_0001100100011111_1101101111111100"; -- 0.09814238462881486
	pesos_i(17180) := b"1111111111111111_1111111111111111_1101101101010010_1001100110110100"; -- -0.14327086788765778
	pesos_i(17181) := b"0000000000000000_0000000000000000_0000100101010001_0011010110101010"; -- 0.03639541057680653
	pesos_i(17182) := b"0000000000000000_0000000000000000_0000101001100110_0111100001000100"; -- 0.040626064862463215
	pesos_i(17183) := b"1111111111111111_1111111111111111_1101110011100011_0101001111111000"; -- -0.13715625004092158
	pesos_i(17184) := b"1111111111111111_1111111111111111_1111010111011000_0101000001100101"; -- -0.03966805956957664
	pesos_i(17185) := b"0000000000000000_0000000000000000_0001110101011001_0010101100010110"; -- 0.11464185034716654
	pesos_i(17186) := b"1111111111111111_1111111111111111_1110001110001001_0000010010110100"; -- -0.11119051554242611
	pesos_i(17187) := b"1111111111111111_1111111111111111_1111000101010101_0011001111101001"; -- -0.057293658798496835
	pesos_i(17188) := b"1111111111111111_1111111111111111_1111000100000010_0110010010000011"; -- -0.05855724144858544
	pesos_i(17189) := b"1111111111111111_1111111111111111_1111011110110101_0010010101111100"; -- -0.0323921749165357
	pesos_i(17190) := b"1111111111111111_1111111111111111_1110011010100111_0110100111100111"; -- -0.09900797004365969
	pesos_i(17191) := b"1111111111111111_1111111111111111_1101101100010111_1100011001011011"; -- -0.14416847487360346
	pesos_i(17192) := b"0000000000000000_0000000000000000_0001110001010001_0001100100111011"; -- 0.1106124656620524
	pesos_i(17193) := b"1111111111111111_1111111111111111_1110000110011111_0001110100011101"; -- -0.11866586729645051
	pesos_i(17194) := b"1111111111111111_1111111111111111_1110000011101010_1110001011001000"; -- -0.12141592612263316
	pesos_i(17195) := b"0000000000000000_0000000000000000_0000010101100101_0111010100010001"; -- 0.021079365466140497
	pesos_i(17196) := b"0000000000000000_0000000000000000_0001101110111011_0110000000010111"; -- 0.10832787097385503
	pesos_i(17197) := b"1111111111111111_1111111111111111_1110100100000101_1001101000111110"; -- -0.08975826248048549
	pesos_i(17198) := b"1111111111111111_1111111111111111_1111001000101100_0011010000001111"; -- -0.05401301041941515
	pesos_i(17199) := b"1111111111111111_1111111111111111_1101011111001101_1001001111010010"; -- -0.1570193875718594
	pesos_i(17200) := b"0000000000000000_0000000000000000_0010011101100110_0010111100001010"; -- 0.1539029502757182
	pesos_i(17201) := b"0000000000000000_0000000000000000_0010000111011100_0010010010101110"; -- 0.13226536997278646
	pesos_i(17202) := b"0000000000000000_0000000000000000_0001010110001100_1100100010001111"; -- 0.08417943465401369
	pesos_i(17203) := b"0000000000000000_0000000000000000_0010001101001011_1000100001101100"; -- 0.1378712906651632
	pesos_i(17204) := b"1111111111111111_1111111111111111_1111011110000101_0010001000001111"; -- -0.033124801054056914
	pesos_i(17205) := b"1111111111111111_1111111111111111_1111001010110011_0110101011000011"; -- -0.051949813297477006
	pesos_i(17206) := b"0000000000000000_0000000000000000_0001001111001110_1001110000011101"; -- 0.07737136573482734
	pesos_i(17207) := b"0000000000000000_0000000000000000_0001110011001001_1101111110101011"; -- 0.11245534817708203
	pesos_i(17208) := b"1111111111111111_1111111111111111_1101101110110011_1001110100001001"; -- -0.14179056668518347
	pesos_i(17209) := b"0000000000000000_0000000000000000_0010010100110111_1111010001111010"; -- 0.1453850554498789
	pesos_i(17210) := b"0000000000000000_0000000000000000_0001011011110100_1101000011001101"; -- 0.08967309011092155
	pesos_i(17211) := b"1111111111111111_1111111111111111_1110011000110111_1101100000010011"; -- -0.10071038747913667
	pesos_i(17212) := b"0000000000000000_0000000000000000_0001000010011110_1100111110100101"; -- 0.06492326524133755
	pesos_i(17213) := b"1111111111111111_1111111111111111_1110000011001000_0010100011100010"; -- -0.12194580528613261
	pesos_i(17214) := b"0000000000000000_0000000000000000_0000101101011110_0111000101111110"; -- 0.044409840834450834
	pesos_i(17215) := b"1111111111111111_1111111111111111_1111101010111001_1101000000011010"; -- -0.02060222031070527
	pesos_i(17216) := b"0000000000000000_0000000000000000_0001101000110001_1101001101000110"; -- 0.10232277351207586
	pesos_i(17217) := b"0000000000000000_0000000000000000_0010100010101110_1010111100100100"; -- 0.15891546860144673
	pesos_i(17218) := b"1111111111111111_1111111111111111_1110000001110111_1110100011011111"; -- -0.12317032380326177
	pesos_i(17219) := b"1111111111111111_1111111111111111_1110100100101110_0000110001101000"; -- -0.08914110618738955
	pesos_i(17220) := b"0000000000000000_0000000000000000_0010010000111001_1010000010001011"; -- 0.1415043201127424
	pesos_i(17221) := b"1111111111111111_1111111111111111_1110001100110001_1110110010000011"; -- -0.11251947217980382
	pesos_i(17222) := b"1111111111111111_1111111111111111_1111111010001101_0111001110011000"; -- -0.005654120767374183
	pesos_i(17223) := b"1111111111111111_1111111111111111_1111001111001011_0010011000001110"; -- -0.0476814474815851
	pesos_i(17224) := b"0000000000000000_0000000000000000_0001100101100011_0000010110001000"; -- 0.09916719981830985
	pesos_i(17225) := b"1111111111111111_1111111111111111_1111011010001000_1011100001000011"; -- -0.03697632188338688
	pesos_i(17226) := b"0000000000000000_0000000000000000_0001010001101000_1111100100001110"; -- 0.07972675889092452
	pesos_i(17227) := b"1111111111111111_1111111111111111_1110100100110001_0111000000100001"; -- -0.08908938593083299
	pesos_i(17228) := b"0000000000000000_0000000000000000_0001101111010011_1111100010100111"; -- 0.10870317543736939
	pesos_i(17229) := b"1111111111111111_1111111111111111_1101011111001111_0011111111101111"; -- -0.15699386982884694
	pesos_i(17230) := b"1111111111111111_1111111111111111_1111100111011101_0010100110100001"; -- -0.023969076228770085
	pesos_i(17231) := b"1111111111111111_1111111111111111_1110001101101110_1011111001101001"; -- -0.11159143389507431
	pesos_i(17232) := b"1111111111111111_1111111111111111_1110111011100101_1000000101110010"; -- -0.0668105217596903
	pesos_i(17233) := b"1111111111111111_1111111111111111_1101110010111000_1101100001110111"; -- -0.13780448041252702
	pesos_i(17234) := b"1111111111111111_1111111111111111_1110111010000101_1010101000000101"; -- -0.06827294708423698
	pesos_i(17235) := b"0000000000000000_0000000000000000_0000000110100100_1011110111100010"; -- 0.006420009274823302
	pesos_i(17236) := b"1111111111111111_1111111111111111_1101111001001011_0011110010100011"; -- -0.1316644765631977
	pesos_i(17237) := b"0000000000000000_0000000000000000_0001110001011011_0010100110010111"; -- 0.11076602872844976
	pesos_i(17238) := b"1111111111111111_1111111111111111_1111110010101100_0010001110100010"; -- -0.012998364284198082
	pesos_i(17239) := b"0000000000000000_0000000000000000_0001100000101001_0100111000110010"; -- 0.09438027125172685
	pesos_i(17240) := b"1111111111111111_1111111111111111_1110101100010101_1000110010001001"; -- -0.08170243882617967
	pesos_i(17241) := b"0000000000000000_0000000000000000_0001011000111011_0110010010100011"; -- 0.08684376687668612
	pesos_i(17242) := b"1111111111111111_1111111111111111_1111110011000110_0001111000000000"; -- -0.012601971683343954
	pesos_i(17243) := b"0000000000000000_0000000000000000_0001010010000001_1001111101010001"; -- 0.08010287985978568
	pesos_i(17244) := b"1111111111111111_1111111111111111_1110000100101011_1110101011011001"; -- -0.1204236239464552
	pesos_i(17245) := b"0000000000000000_0000000000000000_0001111110000111_0010100111110111"; -- 0.12315618786158532
	pesos_i(17246) := b"1111111111111111_1111111111111111_1110101111011110_0101101100100010"; -- -0.07863836683374104
	pesos_i(17247) := b"0000000000000000_0000000000000000_0010000000110000_0101011010000000"; -- 0.1257375777675927
	pesos_i(17248) := b"1111111111111111_1111111111111111_1110001110010100_1000010100001000"; -- -0.11101501998996714
	pesos_i(17249) := b"1111111111111111_1111111111111111_1111111010100010_1011110000101010"; -- -0.005329360808269405
	pesos_i(17250) := b"0000000000000000_0000000000000000_0000110100100010_1110011111111011"; -- 0.0513138760484187
	pesos_i(17251) := b"1111111111111111_1111111111111111_1110010100001001_0100100110001000"; -- -0.10532703813273983
	pesos_i(17252) := b"1111111111111111_1111111111111111_1110111100000011_0011100001100110"; -- -0.06635711196452232
	pesos_i(17253) := b"0000000000000000_0000000000000000_0001001011001101_1100110000001001"; -- 0.0734527131757977
	pesos_i(17254) := b"0000000000000000_0000000000000000_0001100101100100_1011001001110001"; -- 0.0991927647411793
	pesos_i(17255) := b"1111111111111111_1111111111111111_1110101110110000_0000001111101000"; -- -0.07934547021441798
	pesos_i(17256) := b"0000000000000000_0000000000000000_0000010001001001_1111001000010110"; -- 0.01675332114367601
	pesos_i(17257) := b"1111111111111111_1111111111111111_1110110001001010_1011011000101010"; -- -0.07698499186280139
	pesos_i(17258) := b"1111111111111111_1111111111111111_1111011110110001_1111010001111110"; -- -0.03244087139814126
	pesos_i(17259) := b"0000000000000000_0000000000000000_0001101111000011_1100010100011011"; -- 0.10845596216941393
	pesos_i(17260) := b"1111111111111111_1111111111111111_1110101011001010_0000010111001000"; -- -0.08285488006851188
	pesos_i(17261) := b"1111111111111111_1111111111111111_1111011011101001_0010011100011000"; -- -0.03550487200269228
	pesos_i(17262) := b"1111111111111111_1111111111111111_1110110101001010_0010111101101000"; -- -0.07308677387003279
	pesos_i(17263) := b"1111111111111111_1111111111111111_1111111000110100_0100010101110111"; -- -0.007014902608750302
	pesos_i(17264) := b"1111111111111111_1111111111111111_1111100110010001_1000110001000101"; -- -0.025122864896467555
	pesos_i(17265) := b"1111111111111111_1111111111111111_1110011110011111_0111001001000111"; -- -0.09522329106934925
	pesos_i(17266) := b"0000000000000000_0000000000000000_0010100111100010_1101101001001110"; -- 0.16361774824238884
	pesos_i(17267) := b"0000000000000000_0000000000000000_0000001101000101_0111011111010001"; -- 0.012778747992327035
	pesos_i(17268) := b"1111111111111111_1111111111111111_1110101110011100_1111010110001111"; -- -0.0796362424405988
	pesos_i(17269) := b"1111111111111111_1111111111111111_1101100100000011_0110110011001111"; -- -0.1522914881989989
	pesos_i(17270) := b"0000000000000000_0000000000000000_0001000001111111_1001000001010001"; -- 0.06444646803268245
	pesos_i(17271) := b"0000000000000000_0000000000000000_0001101001000001_1110010011111000"; -- 0.10256796881225255
	pesos_i(17272) := b"1111111111111111_1111111111111111_1111000111011110_0110000000010101"; -- -0.05520057183825652
	pesos_i(17273) := b"0000000000000000_0000000000000000_0000010001010110_1101101000000010"; -- 0.01695025020077992
	pesos_i(17274) := b"0000000000000000_0000000000000000_0000100100010100_1010010111010111"; -- 0.035471310539738836
	pesos_i(17275) := b"1111111111111111_1111111111111111_1111110001111111_1011110010000101"; -- -0.01367589718126466
	pesos_i(17276) := b"1111111111111111_1111111111111111_1111100000000100_1000111000110111"; -- -0.031180488076587017
	pesos_i(17277) := b"0000000000000000_0000000000000000_0000100001100001_0010011010011010"; -- 0.03273240336109972
	pesos_i(17278) := b"1111111111111111_1111111111111111_1110001111000100_0100010010110011"; -- -0.11028643266689772
	pesos_i(17279) := b"0000000000000000_0000000000000000_0001010000110100_1001101001100001"; -- 0.07892765883879009
	pesos_i(17280) := b"1111111111111111_1111111111111111_1111110000111111_1000100000110100"; -- -0.014655578004946827
	pesos_i(17281) := b"0000000000000000_0000000000000000_0001010111111011_1001000110000100"; -- 0.08586987944736915
	pesos_i(17282) := b"0000000000000000_0000000000000000_0001101111010110_0010110111011110"; -- 0.10873686466733755
	pesos_i(17283) := b"1111111111111111_1111111111111111_1110000010110011_1001011010100001"; -- -0.12225969865038187
	pesos_i(17284) := b"0000000000000000_0000000000000000_0010000110111111_0101100100000010"; -- 0.1318259840347013
	pesos_i(17285) := b"0000000000000000_0000000000000000_0010011001010101_0000110010110111"; -- 0.14973525498296195
	pesos_i(17286) := b"1111111111111111_1111111111111111_1110110111001101_0011001000110101"; -- -0.07108770563893613
	pesos_i(17287) := b"0000000000000000_0000000000000000_0001011011101110_0000000010010100"; -- 0.08956912637185271
	pesos_i(17288) := b"1111111111111111_1111111111111111_1110010000001101_0101010100111000"; -- -0.1091715562567146
	pesos_i(17289) := b"1111111111111111_1111111111111111_1111100111100010_1101011111000010"; -- -0.023882403453983878
	pesos_i(17290) := b"0000000000000000_0000000000000000_0000101011110001_0000010011110010"; -- 0.042740162832702155
	pesos_i(17291) := b"0000000000000000_0000000000000000_0000101010100100_0111110000000110"; -- 0.04157233371274573
	pesos_i(17292) := b"1111111111111111_1111111111111111_1111110001101000_1001110011100011"; -- -0.01402873469789723
	pesos_i(17293) := b"1111111111111111_1111111111111111_1111010000111111_1011010010100000"; -- -0.04590293031301243
	pesos_i(17294) := b"1111111111111111_1111111111111111_1101101111111011_0111001000100110"; -- -0.14069449006392362
	pesos_i(17295) := b"1111111111111111_1111111111111111_1101101100011110_1100100010101000"; -- -0.14406152638543265
	pesos_i(17296) := b"0000000000000000_0000000000000000_0000011110010111_1010110001001100"; -- 0.029658096881705846
	pesos_i(17297) := b"0000000000000000_0000000000000000_0000000000011001_0100100001000000"; -- 0.00038577617514881966
	pesos_i(17298) := b"1111111111111111_1111111111111111_1111111110010001_0110011001001100"; -- -0.0016876282329000645
	pesos_i(17299) := b"1111111111111111_1111111111111111_1101110100111110_1110110000011010"; -- -0.13575863238822966
	pesos_i(17300) := b"0000000000000000_0000000000000000_0001111100111111_0101010111001010"; -- 0.12206016704754487
	pesos_i(17301) := b"1111111111111111_1111111111111111_1111111010100001_0100110111010110"; -- -0.005351195665492708
	pesos_i(17302) := b"0000000000000000_0000000000000000_0000100100010010_1100010101101101"; -- 0.035442675674487216
	pesos_i(17303) := b"1111111111111111_1111111111111111_1110001011010100_0101000100110101"; -- -0.11394779629343574
	pesos_i(17304) := b"1111111111111111_1111111111111111_1111000000101001_0110001010001110"; -- -0.061868515335487276
	pesos_i(17305) := b"1111111111111111_1111111111111111_1111011110100101_0010101010010110"; -- -0.03263601149969583
	pesos_i(17306) := b"1111111111111111_1111111111111111_1110110110101110_0001011001011001"; -- -0.07156238873466572
	pesos_i(17307) := b"1111111111111111_1111111111111111_1110100100010101_1100111111101111"; -- -0.08951092173029207
	pesos_i(17308) := b"0000000000000000_0000000000000000_0000010110110010_0010111111100010"; -- 0.022250168451436403
	pesos_i(17309) := b"1111111111111111_1111111111111111_1101110011011000_1111110110010100"; -- -0.13731398703746256
	pesos_i(17310) := b"0000000000000000_0000000000000000_0000101010111001_0001000000000100"; -- 0.04188633066279632
	pesos_i(17311) := b"1111111111111111_1111111111111111_1110110001010100_0001011000011101"; -- -0.07684194359083053
	pesos_i(17312) := b"0000000000000000_0000000000000000_0010000000010110_0010001000011000"; -- 0.12533772544035407
	pesos_i(17313) := b"1111111111111111_1111111111111111_1101110001001000_0110110100000110"; -- -0.13951986889280582
	pesos_i(17314) := b"0000000000000000_0000000000000000_0001101010110101_0110100101011100"; -- 0.1043306207494045
	pesos_i(17315) := b"0000000000000000_0000000000000000_0001100111011100_1111110001101000"; -- 0.10102822810736456
	pesos_i(17316) := b"0000000000000000_0000000000000000_0000000110001001_1011011011111100"; -- 0.006007610721494705
	pesos_i(17317) := b"0000000000000000_0000000000000000_0000001000101100_1011011100000101"; -- 0.008494795562946234
	pesos_i(17318) := b"0000000000000000_0000000000000000_0001001011000101_0011110110000010"; -- 0.07332214770037158
	pesos_i(17319) := b"1111111111111111_1111111111111111_1111101000101001_1101100000011100"; -- -0.022799008485182688
	pesos_i(17320) := b"1111111111111111_1111111111111111_1101110011001000_0110011000001011"; -- -0.13756715988723942
	pesos_i(17321) := b"1111111111111111_1111111111111111_1110111110101101_1111000011100000"; -- -0.06375212227413739
	pesos_i(17322) := b"0000000000000000_0000000000000000_0001111000101010_0110100010110010"; -- 0.11783460939374865
	pesos_i(17323) := b"0000000000000000_0000000000000000_0001111011000110_1111101001010010"; -- 0.12022366056042033
	pesos_i(17324) := b"1111111111111111_1111111111111111_1110011000010101_0110001000111100"; -- -0.10123621027556666
	pesos_i(17325) := b"0000000000000000_0000000000000000_0000100111101000_0011100001110001"; -- 0.03869965318982092
	pesos_i(17326) := b"0000000000000000_0000000000000000_0001000001100100_1001011011010100"; -- 0.0640348689415244
	pesos_i(17327) := b"0000000000000000_0000000000000000_0000010010110111_1011010000001110"; -- 0.018428090576472007
	pesos_i(17328) := b"1111111111111111_1111111111111111_1110110101001101_1011110010111111"; -- -0.07303257305974874
	pesos_i(17329) := b"1111111111111111_1111111111111111_1110001001110100_1001001101010000"; -- -0.1154087000401046
	pesos_i(17330) := b"1111111111111111_1111111111111111_1110111100111001_0100000100100001"; -- -0.06553261694405292
	pesos_i(17331) := b"0000000000000000_0000000000000000_0001100100000110_1011100110100000"; -- 0.09775886695127443
	pesos_i(17332) := b"0000000000000000_0000000000000000_0000100101101000_0100111111110110"; -- 0.03674793000898747
	pesos_i(17333) := b"1111111111111111_1111111111111111_1111110111111000_1010111110111010"; -- -0.007924096096386887
	pesos_i(17334) := b"1111111111111111_1111111111111111_1110010111000000_1111100011110010"; -- -0.10252422412044393
	pesos_i(17335) := b"0000000000000000_0000000000000000_0001011011000110_1000001100101110"; -- 0.08896655906974596
	pesos_i(17336) := b"1111111111111111_1111111111111111_1111110000010000_1010011001000011"; -- -0.015370949380681282
	pesos_i(17337) := b"1111111111111111_1111111111111111_1111010110100000_0101111100011011"; -- -0.040521675109526735
	pesos_i(17338) := b"0000000000000000_0000000000000000_0001001011111101_0000010100010010"; -- 0.0741732757684535
	pesos_i(17339) := b"1111111111111111_1111111111111111_1110000110100001_1111110100110000"; -- -0.11862199373181015
	pesos_i(17340) := b"1111111111111111_1111111111111111_1110001011100101_1100101100101010"; -- -0.11368112769122285
	pesos_i(17341) := b"0000000000000000_0000000000000000_0010001001000110_1101100111011101"; -- 0.13389360094761213
	pesos_i(17342) := b"0000000000000000_0000000000000000_0000100001110110_0110110110010011"; -- 0.033057068319636604
	pesos_i(17343) := b"0000000000000000_0000000000000000_0010001010011110_0101111010011000"; -- 0.1352290268442793
	pesos_i(17344) := b"1111111111111111_1111111111111111_1110111011010000_0111100011001100"; -- -0.06713147190426402
	pesos_i(17345) := b"0000000000000000_0000000000000000_0001011011000101_1110010010111010"; -- 0.08895711460121886
	pesos_i(17346) := b"1111111111111111_1111111111111111_1111000100111111_1001000001111111"; -- -0.05762383361316648
	pesos_i(17347) := b"1111111111111111_1111111111111111_1111101101000000_0101011010000001"; -- -0.01854953135265454
	pesos_i(17348) := b"0000000000000000_0000000000000000_0001010000000100_0110110011001000"; -- 0.07819251907734631
	pesos_i(17349) := b"1111111111111111_1111111111111111_1111001110101101_1011011101101000"; -- -0.0481305475695877
	pesos_i(17350) := b"0000000000000000_0000000000000000_0001110110100000_1010101100111100"; -- 0.11573286265143662
	pesos_i(17351) := b"0000000000000000_0000000000000000_0000011001010100_0101010100110010"; -- 0.02472431636393287
	pesos_i(17352) := b"0000000000000000_0000000000000000_0001100111110001_1110100100010100"; -- 0.1013475107615115
	pesos_i(17353) := b"0000000000000000_0000000000000000_0000001001111111_1001101001111011"; -- 0.009759574016946876
	pesos_i(17354) := b"1111111111111111_1111111111111111_1110110100000101_1100110101100111"; -- -0.07413021305905441
	pesos_i(17355) := b"1111111111111111_1111111111111111_1110001101110111_0011000101111111"; -- -0.11146250400082483
	pesos_i(17356) := b"1111111111111111_1111111111111111_1110111001000111_1110000000110000"; -- -0.06921576345757671
	pesos_i(17357) := b"1111111111111111_1111111111111111_1110110000110011_1110101001000100"; -- -0.07733283853856812
	pesos_i(17358) := b"0000000000000000_0000000000000000_0000000111100100_1101001010001011"; -- 0.007397803315833109
	pesos_i(17359) := b"0000000000000000_0000000000000000_0001001001000100_0100110110110011"; -- 0.07135472881725886
	pesos_i(17360) := b"0000000000000000_0000000000000000_0001010100010100_0101001111011011"; -- 0.08234142397208727
	pesos_i(17361) := b"1111111111111111_1111111111111111_1110010001011000_1001001100100110"; -- -0.10802345576280363
	pesos_i(17362) := b"1111111111111111_1111111111111111_1110110011100100_1101010100100110"; -- -0.07463329156248695
	pesos_i(17363) := b"0000000000000000_0000000000000000_0000100100110001_0110000011101000"; -- 0.03590970663465731
	pesos_i(17364) := b"1111111111111111_1111111111111111_1110101011110010_1101101010111001"; -- -0.08223183623833381
	pesos_i(17365) := b"0000000000000000_0000000000000000_0001000001000000_1001100000000010"; -- 0.06348562296029861
	pesos_i(17366) := b"0000000000000000_0000000000000000_0000000110000010_1001001000110101"; -- 0.005898607287548953
	pesos_i(17367) := b"1111111111111111_1111111111111111_1111110010001011_1111100100100010"; -- -0.013489178944174968
	pesos_i(17368) := b"0000000000000000_0000000000000000_0001010001101110_0011100001010010"; -- 0.07980682364326165
	pesos_i(17369) := b"1111111111111111_1111111111111111_1111001010101011_0101110000010111"; -- -0.05207275798579031
	pesos_i(17370) := b"0000000000000000_0000000000000000_0000000110011011_1000001100010110"; -- 0.006279175721815099
	pesos_i(17371) := b"0000000000000000_0000000000000000_0010011111100110_0100110110011101"; -- 0.1558578976447155
	pesos_i(17372) := b"1111111111111111_1111111111111111_1101101111101011_1101010111010000"; -- -0.14093269033116457
	pesos_i(17373) := b"0000000000000000_0000000000000000_0000011100100100_0110100010110110"; -- 0.027899307593129263
	pesos_i(17374) := b"0000000000000000_0000000000000000_0001110010111101_1010010110100011"; -- 0.1122687838491241
	pesos_i(17375) := b"0000000000000000_0000000000000000_0000001100000100_0011100110000100"; -- 0.01178321327050383
	pesos_i(17376) := b"1111111111111111_1111111111111111_1110101100001011_1011001011111110"; -- -0.08185273464529141
	pesos_i(17377) := b"1111111111111111_1111111111111111_1111001101101111_0101001010110011"; -- -0.04908259526222863
	pesos_i(17378) := b"0000000000000000_0000000000000000_0000110110011010_0010001001101100"; -- 0.05313315511319301
	pesos_i(17379) := b"0000000000000000_0000000000000000_0010010100001101_1101010110010011"; -- 0.14474234430746177
	pesos_i(17380) := b"1111111111111111_1111111111111111_1111110011100011_0100011010001100"; -- -0.012157050022883384
	pesos_i(17381) := b"0000000000000000_0000000000000000_0001001101010010_1001110001110001"; -- 0.07547929534476823
	pesos_i(17382) := b"1111111111111111_1111111111111111_1110011001011001_0110001100110110"; -- -0.10019855430619422
	pesos_i(17383) := b"0000000000000000_0000000000000000_0001111100010000_1000011101111100"; -- 0.12134596606216916
	pesos_i(17384) := b"0000000000000000_0000000000000000_0000001001101101_0001100000110101"; -- 0.009477150901328498
	pesos_i(17385) := b"0000000000000000_0000000000000000_0000000100100010_0011110111110100"; -- 0.004428741448276514
	pesos_i(17386) := b"1111111111111111_1111111111111111_1110010000111101_0010111010100011"; -- -0.10844143400469816
	pesos_i(17387) := b"0000000000000000_0000000000000000_0000111111100100_0111111011011010"; -- 0.06208031483651432
	pesos_i(17388) := b"0000000000000000_0000000000000000_0010000100111001_0101010111011111"; -- 0.12978111928841915
	pesos_i(17389) := b"0000000000000000_0000000000000000_0001100101001001_1011001100011010"; -- 0.09878081693734599
	pesos_i(17390) := b"1111111111111111_1111111111111111_1110010100010100_1011100010010000"; -- -0.10515257345480439
	pesos_i(17391) := b"1111111111111111_1111111111111111_1110000010010111_0010010011100111"; -- -0.12269372336385609
	pesos_i(17392) := b"1111111111111111_1111111111111111_1111111110001011_0010010000110001"; -- -0.0017831212194327078
	pesos_i(17393) := b"1111111111111111_1111111111111111_1111000000011111_0110000010010101"; -- -0.062021220903400884
	pesos_i(17394) := b"0000000000000000_0000000000000000_0001100001001000_0000001000111000"; -- 0.09484876515733043
	pesos_i(17395) := b"0000000000000000_0000000000000000_0000001111101010_1000001000101101"; -- 0.0152970656123458
	pesos_i(17396) := b"0000000000000000_0000000000000000_0001100100110100_0100101110011100"; -- 0.0984542137743357
	pesos_i(17397) := b"1111111111111111_1111111111111111_1110110110011000_0101011110100001"; -- -0.07189419094724607
	pesos_i(17398) := b"1111111111111111_1111111111111111_1110111100100000_0110110110010111"; -- -0.06591143660431302
	pesos_i(17399) := b"1111111111111111_1111111111111111_1111111110000001_1100101000011100"; -- -0.0019258195701695434
	pesos_i(17400) := b"0000000000000000_0000000000000000_0000000100111110_0101000000001010"; -- 0.004857065577009012
	pesos_i(17401) := b"0000000000000000_0000000000000000_0000001111011101_1010111111001011"; -- 0.015101420422719872
	pesos_i(17402) := b"0000000000000000_0000000000000000_0001110000011111_1110101011111001"; -- 0.10986202802932798
	pesos_i(17403) := b"1111111111111111_1111111111111111_1110000111010110_1110001000111011"; -- -0.11781488465142774
	pesos_i(17404) := b"1111111111111111_1111111111111111_1101111100101100_1101001001000111"; -- -0.1282223296924688
	pesos_i(17405) := b"1111111111111111_1111111111111111_1111010110100100_0111110110110010"; -- -0.04045881646876348
	pesos_i(17406) := b"1111111111111111_1111111111111111_1110101000011000_0010111000001000"; -- -0.08556854539712566
	pesos_i(17407) := b"0000000000000000_0000000000000000_0000100010010010_0001110101101000"; -- 0.03347953590126209
	pesos_i(17408) := b"0000000000000000_0000000000000000_0000100000101001_1010011011111010"; -- 0.031885562892987454
	pesos_i(17409) := b"1111111111111111_1111111111111111_1101110011101000_1010001001100100"; -- -0.13707528160219046
	pesos_i(17410) := b"0000000000000000_0000000000000000_0001001000110011_1100111110111111"; -- 0.07110308086257532
	pesos_i(17411) := b"0000000000000000_0000000000000000_0001010110000100_1011101110011101"; -- 0.08405659273223216
	pesos_i(17412) := b"0000000000000000_0000000000000000_0000011010111111_0110011101000111"; -- 0.026358084420923876
	pesos_i(17413) := b"0000000000000000_0000000000000000_0000001101101111_0111101100011110"; -- 0.013419813945715049
	pesos_i(17414) := b"1111111111111111_1111111111111111_1111010110100111_1001100011000011"; -- -0.04041142686254065
	pesos_i(17415) := b"0000000000000000_0000000000000000_0000010110110100_1011010110011000"; -- 0.022288655917245163
	pesos_i(17416) := b"1111111111111111_1111111111111111_1101111011110110_1101001000100010"; -- -0.12904631309760892
	pesos_i(17417) := b"0000000000000000_0000000000000000_0001000001011100_0001111100100100"; -- 0.06390566477053429
	pesos_i(17418) := b"0000000000000000_0000000000000000_0001000101000001_1000010000101011"; -- 0.06740594907112404
	pesos_i(17419) := b"1111111111111111_1111111111111111_1110010000111001_0111001111110101"; -- -0.10849833741365
	pesos_i(17420) := b"1111111111111111_1111111111111111_1111001011010101_1000011101100100"; -- -0.051429307934761165
	pesos_i(17421) := b"1111111111111111_1111111111111111_1110001101010000_1011011011111111"; -- -0.11204963947493661
	pesos_i(17422) := b"1111111111111111_1111111111111111_1110011011101101_0101111001011110"; -- -0.0979405421755719
	pesos_i(17423) := b"0000000000000000_0000000000000000_0000100010101111_0011000101110000"; -- 0.0339232347919315
	pesos_i(17424) := b"0000000000000000_0000000000000000_0001011001000000_1110101010010110"; -- 0.08692804479883003
	pesos_i(17425) := b"0000000000000000_0000000000000000_0000101011100000_1111011110011101"; -- 0.04249522758484276
	pesos_i(17426) := b"1111111111111111_1111111111111111_1111101100111100_0101111000100010"; -- -0.01861011181394486
	pesos_i(17427) := b"0000000000000000_0000000000000000_0010000011001011_1000110110100010"; -- 0.12810597620419628
	pesos_i(17428) := b"0000000000000000_0000000000000000_0010010010000110_1101101110000001"; -- 0.1426827612661523
	pesos_i(17429) := b"0000000000000000_0000000000000000_0000110001010011_0010111100100110"; -- 0.04814428971014443
	pesos_i(17430) := b"0000000000000000_0000000000000000_0001001101000100_0111001111000100"; -- 0.0752632477593839
	pesos_i(17431) := b"0000000000000000_0000000000000000_0001110101100011_0110100110010100"; -- 0.11479816313788707
	pesos_i(17432) := b"0000000000000000_0000000000000000_0000111110101100_1000001111000110"; -- 0.06122611593155651
	pesos_i(17433) := b"1111111111111111_1111111111111111_1101100110010010_0110101100001000"; -- -0.150109587133991
	pesos_i(17434) := b"0000000000000000_0000000000000000_0010000011110100_0001110100111001"; -- 0.12872488635594512
	pesos_i(17435) := b"1111111111111111_1111111111111111_1111111000010111_0010110010110100"; -- -0.007458883236445156
	pesos_i(17436) := b"1111111111111111_1111111111111111_1111101101011111_1011000001101100"; -- -0.018071149552543197
	pesos_i(17437) := b"0000000000000000_0000000000000000_0000101001100101_1101110100000000"; -- 0.040616810217785834
	pesos_i(17438) := b"1111111111111111_1111111111111111_1110001111000100_0110001111111010"; -- -0.11028456819841527
	pesos_i(17439) := b"0000000000000000_0000000000000000_0010001000111000_1100010101101000"; -- 0.1336787585577173
	pesos_i(17440) := b"1111111111111111_1111111111111111_1111000011001110_1111101100100110"; -- -0.0593417199378
	pesos_i(17441) := b"0000000000000000_0000000000000000_0001110100000101_1101011010110000"; -- 0.11337034025816695
	pesos_i(17442) := b"1111111111111111_1111111111111111_1110010111001101_1010101001110010"; -- -0.10233053880839232
	pesos_i(17443) := b"0000000000000000_0000000000000000_0000111111001011_0101111100011111"; -- 0.061696953741067796
	pesos_i(17444) := b"0000000000000000_0000000000000000_0010001111000101_0101011000010110"; -- 0.13972986262059164
	pesos_i(17445) := b"1111111111111111_1111111111111111_1110101110001111_0101000000011000"; -- -0.07984446929926367
	pesos_i(17446) := b"0000000000000000_0000000000000000_0001110001010011_1101101110111011"; -- 0.11065457654009006
	pesos_i(17447) := b"1111111111111111_1111111111111111_1110101010010011_1011110100110110"; -- -0.08368318006188066
	pesos_i(17448) := b"1111111111111111_1111111111111111_1110000111010000_0110001100010001"; -- -0.11791401707443101
	pesos_i(17449) := b"0000000000000000_0000000000000000_0001101011111110_1101111101001001"; -- 0.10545154126794183
	pesos_i(17450) := b"0000000000000000_0000000000000000_0010000001100000_1011101011001110"; -- 0.1264759782868781
	pesos_i(17451) := b"1111111111111111_1111111111111111_1110001001001000_1110000010001101"; -- -0.11607548286615117
	pesos_i(17452) := b"0000000000000000_0000000000000000_0000101110111010_1001001111110111"; -- 0.04581570407177483
	pesos_i(17453) := b"0000000000000000_0000000000000000_0001111010101101_1011111111111110"; -- 0.11983871407519112
	pesos_i(17454) := b"0000000000000000_0000000000000000_0000011110101011_1011011011011110"; -- 0.029963902684893493
	pesos_i(17455) := b"0000000000000000_0000000000000000_0001010001100010_1010101011100001"; -- 0.07963054647440822
	pesos_i(17456) := b"1111111111111111_1111111111111111_1110001010011010_1011000111110001"; -- -0.114827040462422
	pesos_i(17457) := b"0000000000000000_0000000000000000_0010000111110001_1010101110101101"; -- 0.13259385080072283
	pesos_i(17458) := b"0000000000000000_0000000000000000_0010010000011000_0001011000001011"; -- 0.14099252478477706
	pesos_i(17459) := b"1111111111111111_1111111111111111_1111011111100011_0110010110111000"; -- -0.03168644196964467
	pesos_i(17460) := b"1111111111111111_1111111111111111_1111100100011011_1011111010011101"; -- -0.026920401164613982
	pesos_i(17461) := b"0000000000000000_0000000000000000_0000001010001010_1101010011000110"; -- 0.009930895256529184
	pesos_i(17462) := b"1111111111111111_1111111111111111_1111000101101111_1011100110100000"; -- -0.0568889602038185
	pesos_i(17463) := b"1111111111111111_1111111111111111_1110010000110110_1101011000001101"; -- -0.10853826694304229
	pesos_i(17464) := b"0000000000000000_0000000000000000_0001010111000001_1110111101111000"; -- 0.08499046963394244
	pesos_i(17465) := b"0000000000000000_0000000000000000_0001001010000000_1101001111101011"; -- 0.07227825622504296
	pesos_i(17466) := b"1111111111111111_1111111111111111_1111100110111011_0110000000100110"; -- -0.02448462547499737
	pesos_i(17467) := b"1111111111111111_1111111111111111_1110110110111110_0100011001001110"; -- -0.07131538956673251
	pesos_i(17468) := b"1111111111111111_1111111111111111_1101111110110110_1011100110100010"; -- -0.12611808578303055
	pesos_i(17469) := b"1111111111111111_1111111111111111_1110101110101100_1011101100110101"; -- -0.07939557992079657
	pesos_i(17470) := b"0000000000000000_0000000000000000_0000010010111100_0110011010010100"; -- 0.018499766586665765
	pesos_i(17471) := b"1111111111111111_1111111111111111_1110001001000101_0110111110010110"; -- -0.11612799261785607
	pesos_i(17472) := b"0000000000000000_0000000000000000_0010010110110010_0110100010101110"; -- 0.14725355392649828
	pesos_i(17473) := b"1111111111111111_1111111111111111_1110100101101100_0000101110101001"; -- -0.08819510589371975
	pesos_i(17474) := b"0000000000000000_0000000000000000_0001000001011001_1110010100111011"; -- 0.06387169548377993
	pesos_i(17475) := b"1111111111111111_1111111111111111_1110011000101001_0000011101111011"; -- -0.10093644387406693
	pesos_i(17476) := b"0000000000000000_0000000000000000_0000011110100100_1011000100101100"; -- 0.029856751579912726
	pesos_i(17477) := b"1111111111111111_1111111111111111_1110101011111110_0010101110001000"; -- -0.08205917283710584
	pesos_i(17478) := b"0000000000000000_0000000000000000_0010000010010001_0100100000101010"; -- 0.12721682575526935
	pesos_i(17479) := b"1111111111111111_1111111111111111_1111000111000001_1001110110100001"; -- -0.055639408185031596
	pesos_i(17480) := b"1111111111111111_1111111111111111_1111111101001001_1011111001000011"; -- -0.002781017929501164
	pesos_i(17481) := b"1111111111111111_1111111111111111_1110100001110110_1100001100011100"; -- -0.09193783346604695
	pesos_i(17482) := b"0000000000000000_0000000000000000_0001000101111101_0011100111000001"; -- 0.06831704091877495
	pesos_i(17483) := b"0000000000000000_0000000000000000_0001101100100001_0101001111101101"; -- 0.10597729233125247
	pesos_i(17484) := b"0000000000000000_0000000000000000_0000101111000000_1000110100101011"; -- 0.045906851878264064
	pesos_i(17485) := b"0000000000000000_0000000000000000_0001000111001000_1010001100001010"; -- 0.06946772581320687
	pesos_i(17486) := b"1111111111111111_1111111111111111_1110000101111111_1000100001110010"; -- -0.11914775098512768
	pesos_i(17487) := b"0000000000000000_0000000000000000_0001110100110011_1001101001011111"; -- 0.11406864943939658
	pesos_i(17488) := b"0000000000000000_0000000000000000_0000100010110101_0011010011010101"; -- 0.03401498977949074
	pesos_i(17489) := b"0000000000000000_0000000000000000_0001000111111100_1011111001011111"; -- 0.07026281173507443
	pesos_i(17490) := b"1111111111111111_1111111111111111_1111010001110010_1000100101010011"; -- -0.045127312792739946
	pesos_i(17491) := b"0000000000000000_0000000000000000_0001010011110001_0000111000101000"; -- 0.08180321194619768
	pesos_i(17492) := b"0000000000000000_0000000000000000_0010001010100011_0010010101111000"; -- 0.1353019160046425
	pesos_i(17493) := b"1111111111111111_1111111111111111_1111001010001011_1110100101101010"; -- -0.05255261568815086
	pesos_i(17494) := b"0000000000000000_0000000000000000_0000000011100111_0111110011110001"; -- 0.0035322274032635456
	pesos_i(17495) := b"0000000000000000_0000000000000000_0000011011100000_0001011010110100"; -- 0.02685682201644868
	pesos_i(17496) := b"0000000000000000_0000000000000000_0010000010001111_0000011111111010"; -- 0.12718248237075597
	pesos_i(17497) := b"0000000000000000_0000000000000000_0000111011011000_0111010101000011"; -- 0.05799038767077397
	pesos_i(17498) := b"0000000000000000_0000000000000000_0001101100100111_1000010001111001"; -- 0.10607173881405377
	pesos_i(17499) := b"0000000000000000_0000000000000000_0000001001010011_0100110001100110"; -- 0.009083533290644237
	pesos_i(17500) := b"1111111111111111_1111111111111111_1111001101111010_1010011111011101"; -- -0.04890967228281421
	pesos_i(17501) := b"1111111111111111_1111111111111111_1101111111010101_0111100001100001"; -- -0.12564895272601653
	pesos_i(17502) := b"1111111111111111_1111111111111111_1111001101000110_1001100011110001"; -- -0.049704018654970324
	pesos_i(17503) := b"0000000000000000_0000000000000000_0001101100011111_0011100110111100"; -- 0.10594521360056558
	pesos_i(17504) := b"1111111111111111_1111111111111111_1110001000011010_1100011100100010"; -- -0.11677890214466916
	pesos_i(17505) := b"1111111111111111_1111111111111111_1111011111101100_0011110111100011"; -- -0.03155148706802046
	pesos_i(17506) := b"0000000000000000_0000000000000000_0000111111010000_0110011000011000"; -- 0.061773663301185396
	pesos_i(17507) := b"0000000000000000_0000000000000000_0001010111000110_0110001101011111"; -- 0.08505841328833333
	pesos_i(17508) := b"0000000000000000_0000000000000000_0001110110011010_1100100000001011"; -- 0.11564302703668626
	pesos_i(17509) := b"1111111111111111_1111111111111111_1110000100111110_0110010111100000"; -- -0.12014163289485522
	pesos_i(17510) := b"1111111111111111_1111111111111111_1110000011000100_1100011001000111"; -- -0.12199745908342614
	pesos_i(17511) := b"0000000000000000_0000000000000000_0001010001100100_0011101000111100"; -- 0.07965435002674985
	pesos_i(17512) := b"0000000000000000_0000000000000000_0001100101000001_0011101000000011"; -- 0.0986515290478046
	pesos_i(17513) := b"0000000000000000_0000000000000000_0001011010111100_0101111100110011"; -- 0.08881182658375442
	pesos_i(17514) := b"0000000000000000_0000000000000000_0001001101110011_0111110101010110"; -- 0.0759809814013404
	pesos_i(17515) := b"0000000000000000_0000000000000000_0001000000111011_1010001011010100"; -- 0.06340997377951878
	pesos_i(17516) := b"1111111111111111_1111111111111111_1111110000001101_0011001010001111"; -- -0.015423622210415888
	pesos_i(17517) := b"0000000000000000_0000000000000000_0000001110000101_0110010110000110"; -- 0.013754220126217135
	pesos_i(17518) := b"0000000000000000_0000000000000000_0000111001100011_1100001001100010"; -- 0.05620970614687933
	pesos_i(17519) := b"0000000000000000_0000000000000000_0000111010111110_1011001001001000"; -- 0.057597296283436565
	pesos_i(17520) := b"0000000000000000_0000000000000000_0010000110111001_1111110000101001"; -- 0.13174415599461572
	pesos_i(17521) := b"1111111111111111_1111111111111111_1110010001110001_0101011100000101"; -- -0.10764557004193041
	pesos_i(17522) := b"0000000000000000_0000000000000000_0010010000100110_1100110011110010"; -- 0.14121704962406284
	pesos_i(17523) := b"0000000000000000_0000000000000000_0001000111101001_1010001011100111"; -- 0.06997125759984932
	pesos_i(17524) := b"0000000000000000_0000000000000000_0001100101000111_0111010100101001"; -- 0.09874660726619901
	pesos_i(17525) := b"0000000000000000_0000000000000000_0010000101000011_1000010100111001"; -- 0.12993652953415954
	pesos_i(17526) := b"0000000000000000_0000000000000000_0000101010111011_0010001101110001"; -- 0.04191800609809345
	pesos_i(17527) := b"1111111111111111_1111111111111111_1110010110100111_0011101100110011"; -- -0.10291700369740918
	pesos_i(17528) := b"1111111111111111_1111111111111111_1111111000110110_0100111001011011"; -- -0.006983855050407329
	pesos_i(17529) := b"0000000000000000_0000000000000000_0001001111011010_0011000100110011"; -- 0.07754809862182502
	pesos_i(17530) := b"1111111111111111_1111111111111111_1110010111111111_1111001000101101"; -- -0.10156332399564907
	pesos_i(17531) := b"1111111111111111_1111111111111111_1110100110001110_1111101110010110"; -- -0.08766200627813409
	pesos_i(17532) := b"1111111111111111_1111111111111111_1110011001100101_1011111001100001"; -- -0.10001001491416768
	pesos_i(17533) := b"0000000000000000_0000000000000000_0010000000001111_0101100101100010"; -- 0.1252342094739298
	pesos_i(17534) := b"0000000000000000_0000000000000000_0000001110101010_0001111111000001"; -- 0.014314636907116908
	pesos_i(17535) := b"1111111111111111_1111111111111111_1111000001100011_0000111001110010"; -- -0.060988518837224365
	pesos_i(17536) := b"1111111111111111_1111111111111111_1110111001111011_0101011100111000"; -- -0.06843047026726927
	pesos_i(17537) := b"1111111111111111_1111111111111111_1110100000101000_0110010010110000"; -- -0.09313364688812542
	pesos_i(17538) := b"0000000000000000_0000000000000000_0000110110000010_0111001010000000"; -- 0.05277171740113194
	pesos_i(17539) := b"0000000000000000_0000000000000000_0000110110010100_1000100000100101"; -- 0.053047665678987346
	pesos_i(17540) := b"1111111111111111_1111111111111111_1110010110111000_0101100101001011"; -- -0.10265581055765706
	pesos_i(17541) := b"1111111111111111_1111111111111111_1111100001101000_0101001010111011"; -- -0.0296581548896397
	pesos_i(17542) := b"1111111111111111_1111111111111111_1111110111000101_0010101111110101"; -- -0.00871014851950785
	pesos_i(17543) := b"0000000000000000_0000000000000000_0001110111010111_0001101000111101"; -- 0.11656345348334674
	pesos_i(17544) := b"0000000000000000_0000000000000000_0001110001011011_0111111110001010"; -- 0.11077115175775788
	pesos_i(17545) := b"1111111111111111_1111111111111111_1101100111010110_1000000101110100"; -- -0.1490706531076421
	pesos_i(17546) := b"1111111111111111_1111111111111111_1110111011111010_0011100010010010"; -- -0.06649443077456682
	pesos_i(17547) := b"1111111111111111_1111111111111111_1111101001001111_1101110001110000"; -- -0.022218916489020638
	pesos_i(17548) := b"1111111111111111_1111111111111111_1111010011110000_0011111111110011"; -- -0.043209078842758174
	pesos_i(17549) := b"0000000000000000_0000000000000000_0000011001111100_1000110011000011"; -- 0.02533797980367522
	pesos_i(17550) := b"1111111111111111_1111111111111111_1101111101100100_0001000000111101"; -- -0.1273794032867971
	pesos_i(17551) := b"0000000000000000_0000000000000000_0000010101111011_1100000101011110"; -- 0.021419606738668044
	pesos_i(17552) := b"1111111111111111_1111111111111111_1110001111010010_0011101010001011"; -- -0.11007341483442368
	pesos_i(17553) := b"1111111111111111_1111111111111111_1110011000101011_0101001000100010"; -- -0.100901476604094
	pesos_i(17554) := b"0000000000000000_0000000000000000_0010010011110101_1100100101111111"; -- 0.14437541350789163
	pesos_i(17555) := b"1111111111111111_1111111111111111_1111100100111100_0101101110110010"; -- -0.026422757291255317
	pesos_i(17556) := b"0000000000000000_0000000000000000_0010000011111111_1110010110001001"; -- 0.12890467260201233
	pesos_i(17557) := b"0000000000000000_0000000000000000_0001001111011110_0010001100010011"; -- 0.07760829177120557
	pesos_i(17558) := b"1111111111111111_1111111111111111_1101100010011011_0101110000011000"; -- -0.15387939852919505
	pesos_i(17559) := b"0000000000000000_0000000000000000_0010011001011011_1111101100110111"; -- 0.1498410234492596
	pesos_i(17560) := b"0000000000000000_0000000000000000_0001110100101011_0110101100001100"; -- 0.11394375840314788
	pesos_i(17561) := b"1111111111111111_1111111111111111_1110010000000101_0000010011100111"; -- -0.10929841376659101
	pesos_i(17562) := b"0000000000000000_0000000000000000_0010010000111101_1001010000000010"; -- 0.14156460818038186
	pesos_i(17563) := b"1111111111111111_1111111111111111_1101101110100011_1111000111001011"; -- -0.14202965535136977
	pesos_i(17564) := b"1111111111111111_1111111111111111_1110111101010000_0011111111000100"; -- -0.06518174604468252
	pesos_i(17565) := b"0000000000000000_0000000000000000_0001010001001101_1011010110010000"; -- 0.0793107487380995
	pesos_i(17566) := b"0000000000000000_0000000000000000_0000100100101000_1100101000001100"; -- 0.03577864443413691
	pesos_i(17567) := b"1111111111111111_1111111111111111_1111011011000100_0111000011010111"; -- -0.03606505163727594
	pesos_i(17568) := b"0000000000000000_0000000000000000_0001000111101110_1110011110111000"; -- 0.07005165327291969
	pesos_i(17569) := b"0000000000000000_0000000000000000_0001011111100100_0110000111111011"; -- 0.09332859390119591
	pesos_i(17570) := b"0000000000000000_0000000000000000_0010001001111010_0001011011011101"; -- 0.13467543511373023
	pesos_i(17571) := b"1111111111111111_1111111111111111_1111001101010010_0011101100010011"; -- -0.049526508140216675
	pesos_i(17572) := b"1111111111111111_1111111111111111_1110001010111001_1100000000111110"; -- -0.1143531655593858
	pesos_i(17573) := b"1111111111111111_1111111111111111_1111010100100000_1101111111001101"; -- -0.04246712927420275
	pesos_i(17574) := b"1111111111111111_1111111111111111_1110000000101000_1110000101100111"; -- -0.12437621351057244
	pesos_i(17575) := b"1111111111111111_1111111111111111_1111011100110011_0100001111110000"; -- -0.034374002373550455
	pesos_i(17576) := b"1111111111111111_1111111111111111_1110110101001101_1011101100011000"; -- -0.07303267155076218
	pesos_i(17577) := b"0000000000000000_0000000000000000_0000001101010100_0001011101011000"; -- 0.013001879637710486
	pesos_i(17578) := b"0000000000000000_0000000000000000_0000111011010000_0100110101010100"; -- 0.057865937215410466
	pesos_i(17579) := b"1111111111111111_1111111111111111_1110101110110010_1010110101000000"; -- -0.07930485903243649
	pesos_i(17580) := b"0000000000000000_0000000000000000_0001011100011111_1011010110101111"; -- 0.09032760153211317
	pesos_i(17581) := b"0000000000000000_0000000000000000_0001011110101000_0000101111010000"; -- 0.09240793068111039
	pesos_i(17582) := b"0000000000000000_0000000000000000_0000010110001011_0101000110111110"; -- 0.021657094006204563
	pesos_i(17583) := b"1111111111111111_1111111111111111_1111101111010001_1110101000010100"; -- -0.01632821091945036
	pesos_i(17584) := b"0000000000000000_0000000000000000_0000001101110000_1101110111110110"; -- 0.013440964368394953
	pesos_i(17585) := b"1111111111111111_1111111111111111_1110110011000010_0110000101100001"; -- -0.07515899059440585
	pesos_i(17586) := b"1111111111111111_1111111111111111_1110001000111010_1011010100001101"; -- -0.1162916987311751
	pesos_i(17587) := b"1111111111111111_1111111111111111_1101101000100010_1010101011111011"; -- -0.14790850989935078
	pesos_i(17588) := b"1111111111111111_1111111111111111_1110100001001000_1111100101010000"; -- -0.09263650694825526
	pesos_i(17589) := b"1111111111111111_1111111111111111_1110010011010010_1011010000001111"; -- -0.10615992199070669
	pesos_i(17590) := b"0000000000000000_0000000000000000_0000000111001000_0011100101011100"; -- 0.006961426586775765
	pesos_i(17591) := b"0000000000000000_0000000000000000_0010100001010001_1111110001011101"; -- 0.15750100394517458
	pesos_i(17592) := b"1111111111111111_1111111111111111_1110010011100010_0000100110001001"; -- -0.10592594534018344
	pesos_i(17593) := b"1111111111111111_1111111111111111_1101101011101001_0100010001011111"; -- -0.1448781269949601
	pesos_i(17594) := b"0000000000000000_0000000000000000_0010011101010110_0010001101010011"; -- 0.1536581113105054
	pesos_i(17595) := b"0000000000000000_0000000000000000_0001011110000000_1100000000001110"; -- 0.09180832232118455
	pesos_i(17596) := b"1111111111111111_1111111111111111_1101101000110100_1010100101111100"; -- -0.14763394089070486
	pesos_i(17597) := b"1111111111111111_1111111111111111_1110011010111011_1111110011100001"; -- -0.09869403365829334
	pesos_i(17598) := b"1111111111111111_1111111111111111_1111010010010001_1001001011100111"; -- -0.04465371956512144
	pesos_i(17599) := b"1111111111111111_1111111111111111_1111101001101100_0011100011011100"; -- -0.0217861617682058
	pesos_i(17600) := b"0000000000000000_0000000000000000_0001000110110110_1101011101011011"; -- 0.06919618571946264
	pesos_i(17601) := b"0000000000000000_0000000000000000_0000100001100110_0001010001010100"; -- 0.03280760811962268
	pesos_i(17602) := b"1111111111111111_1111111111111111_1111110110100011_0010110110111011"; -- -0.009228841687592892
	pesos_i(17603) := b"1111111111111111_1111111111111111_1110011001101011_0111110101000001"; -- -0.0999223437989798
	pesos_i(17604) := b"0000000000000000_0000000000000000_0001110011011110_0001010101101000"; -- 0.11276372705370866
	pesos_i(17605) := b"1111111111111111_1111111111111111_1111100010000100_1110011111011110"; -- -0.029222019455916636
	pesos_i(17606) := b"1111111111111111_1111111111111111_1111011101010010_0100010011101111"; -- -0.0339009204993333
	pesos_i(17607) := b"1111111111111111_1111111111111111_1110101000010100_0111000110100110"; -- -0.08562555035131655
	pesos_i(17608) := b"1111111111111111_1111111111111111_1101101001001000_0000101010001111"; -- -0.14733823774933014
	pesos_i(17609) := b"0000000000000000_0000000000000000_0000110111111000_1101000100111110"; -- 0.054577901598815176
	pesos_i(17610) := b"1111111111111111_1111111111111111_1111011011111010_1100110011111110"; -- -0.035235584337344784
	pesos_i(17611) := b"0000000000000000_0000000000000000_0001001011001101_0000010000010100"; -- 0.07344079477709099
	pesos_i(17612) := b"0000000000000000_0000000000000000_0000010110000000_1001101101110111"; -- 0.021493641415380068
	pesos_i(17613) := b"0000000000000000_0000000000000000_0000011111010000_0001010010011000"; -- 0.030518805623263923
	pesos_i(17614) := b"0000000000000000_0000000000000000_0010001010101100_1011110111011000"; -- 0.13544832725616462
	pesos_i(17615) := b"1111111111111111_1111111111111111_1111011100100000_1111001010100000"; -- -0.034653507269610265
	pesos_i(17616) := b"1111111111111111_1111111111111111_1110110100010100_1001110001001011"; -- -0.07390425852757616
	pesos_i(17617) := b"0000000000000000_0000000000000000_0000011010001001_0110010111111101"; -- 0.02553403308033263
	pesos_i(17618) := b"0000000000000000_0000000000000000_0001100001101000_0101000100101001"; -- 0.09534175153153504
	pesos_i(17619) := b"0000000000000000_0000000000000000_0000111100011110_1000101110101001"; -- 0.05905983805496516
	pesos_i(17620) := b"0000000000000000_0000000000000000_0000010011010000_1000001011000100"; -- 0.01880662236213048
	pesos_i(17621) := b"0000000000000000_0000000000000000_0000110001010010_0011110000010010"; -- 0.048129801141511615
	pesos_i(17622) := b"0000000000000000_0000000000000000_0000010010111111_0010010010001110"; -- 0.018541607496837892
	pesos_i(17623) := b"1111111111111111_1111111111111111_1110000110001001_0111000010010000"; -- -0.11899658658853651
	pesos_i(17624) := b"0000000000000000_0000000000000000_0000101011101110_0110100101111111"; -- 0.04270037996069416
	pesos_i(17625) := b"0000000000000000_0000000000000000_0001100000011101_0001110100110111"; -- 0.09419424611078335
	pesos_i(17626) := b"1111111111111111_1111111111111111_1111000111101110_1011101001100110"; -- -0.05495104805309808
	pesos_i(17627) := b"0000000000000000_0000000000000000_0001011000000100_1101100101111100"; -- 0.08601149824541603
	pesos_i(17628) := b"0000000000000000_0000000000000000_0000010110101000_0000101101111001"; -- 0.022095410429966728
	pesos_i(17629) := b"0000000000000000_0000000000000000_0001010111101100_0010011100000111"; -- 0.08563465053314953
	pesos_i(17630) := b"0000000000000000_0000000000000000_0001100101011001_0111101100010010"; -- 0.09902161773052474
	pesos_i(17631) := b"1111111111111111_1111111111111111_1111010001000100_1000101100111111"; -- -0.04582910268286892
	pesos_i(17632) := b"1111111111111111_1111111111111111_1101111101100111_1000101001001101"; -- -0.12732635144099014
	pesos_i(17633) := b"1111111111111111_1111111111111111_1110110010101100_1110011001101010"; -- -0.07548675451801433
	pesos_i(17634) := b"1111111111111111_1111111111111111_1110010110001100_0011101011111001"; -- -0.10332900451199292
	pesos_i(17635) := b"1111111111111111_1111111111111111_1110001110101000_1100010111010100"; -- -0.11070598203895289
	pesos_i(17636) := b"0000000000000000_0000000000000000_0001100000100000_0100111111010100"; -- 0.09424303938102989
	pesos_i(17637) := b"1111111111111111_1111111111111111_1111000101100010_0110010111100110"; -- -0.057092315109216626
	pesos_i(17638) := b"1111111111111111_1111111111111111_1111110101101000_0111010000000000"; -- -0.010124921771363206
	pesos_i(17639) := b"1111111111111111_1111111111111111_1110010110110010_1000111001011100"; -- -0.10274420016842371
	pesos_i(17640) := b"0000000000000000_0000000000000000_0000010011001011_1100101011001111"; -- 0.01873462246352045
	pesos_i(17641) := b"1111111111111111_1111111111111111_1111110101111001_1010100111001011"; -- -0.009862316087407983
	pesos_i(17642) := b"0000000000000000_0000000000000000_0000011101001110_0110010100010011"; -- 0.028539959984593504
	pesos_i(17643) := b"0000000000000000_0000000000000000_0001010100110101_1111110000010000"; -- 0.08285498991399833
	pesos_i(17644) := b"1111111111111111_1111111111111111_1110110000111011_1010001111100100"; -- -0.07721496283819622
	pesos_i(17645) := b"0000000000000000_0000000000000000_0010001101101000_1101111001110010"; -- 0.138318922856578
	pesos_i(17646) := b"1111111111111111_1111111111111111_1111101100111101_1010100001101010"; -- -0.018590425669463184
	pesos_i(17647) := b"1111111111111111_1111111111111111_1110011110001111_1001101101001011"; -- -0.09546498686749308
	pesos_i(17648) := b"0000000000000000_0000000000000000_0000010111100000_1010100000001100"; -- 0.022959235231776037
	pesos_i(17649) := b"1111111111111111_1111111111111111_1110110001000001_1001111111001110"; -- -0.07712365370374101
	pesos_i(17650) := b"0000000000000000_0000000000000000_0000010011001000_0000110110110110"; -- 0.018677575013089687
	pesos_i(17651) := b"0000000000000000_0000000000000000_0000000111111011_0111011111000100"; -- 0.007743344648935267
	pesos_i(17652) := b"0000000000000000_0000000000000000_0001100100000111_0011001110001100"; -- 0.09776613396213149
	pesos_i(17653) := b"1111111111111111_1111111111111111_1111011100011010_1000000001110010"; -- -0.034751865638246046
	pesos_i(17654) := b"1111111111111111_1111111111111111_1101100111000011_0000011101111010"; -- -0.14936784039080642
	pesos_i(17655) := b"0000000000000000_0000000000000000_0001001100001010_1011111011010100"; -- 0.07438271210848772
	pesos_i(17656) := b"1111111111111111_1111111111111111_1111110100001111_1111111001000100"; -- -0.011474712806871179
	pesos_i(17657) := b"1111111111111111_1111111111111111_1101101101011010_0101000111111001"; -- -0.14315307295136429
	pesos_i(17658) := b"0000000000000000_0000000000000000_0010000111010110_1101111111000101"; -- 0.13218496854578932
	pesos_i(17659) := b"1111111111111111_1111111111111111_1110001101100000_0101000101010110"; -- -0.11181155818106363
	pesos_i(17660) := b"0000000000000000_0000000000000000_0001010101100010_1000000100011001"; -- 0.08353430617830082
	pesos_i(17661) := b"1111111111111111_1111111111111111_1111001111100000_0100100001110001"; -- -0.04735896347843746
	pesos_i(17662) := b"1111111111111111_1111111111111111_1101110100101000_0010111110001100"; -- -0.13610556445170463
	pesos_i(17663) := b"1111111111111111_1111111111111111_1110100100110011_0110001001110110"; -- -0.08905968292863597
	pesos_i(17664) := b"0000000000000000_0000000000000000_0000001100001100_0101101011100101"; -- 0.011907273312060419
	pesos_i(17665) := b"0000000000000000_0000000000000000_0001010010000110_0010110011110110"; -- 0.08017235760312662
	pesos_i(17666) := b"0000000000000000_0000000000000000_0001110001100000_1010000011001001"; -- 0.11084942730692596
	pesos_i(17667) := b"0000000000000000_0000000000000000_0000011101110001_1101011001011111"; -- 0.029080770667825287
	pesos_i(17668) := b"0000000000000000_0000000000000000_0000001000000100_0010000101101111"; -- 0.007875528047125898
	pesos_i(17669) := b"0000000000000000_0000000000000000_0000110011101000_1110101010011111"; -- 0.050429023622712246
	pesos_i(17670) := b"0000000000000000_0000000000000000_0001101100101110_1100010100110010"; -- 0.1061824080609069
	pesos_i(17671) := b"1111111111111111_1111111111111111_1111011100100110_1101110100101100"; -- -0.034563233199076324
	pesos_i(17672) := b"0000000000000000_0000000000000000_0001100011000000_1011110000011100"; -- 0.09669089971538221
	pesos_i(17673) := b"0000000000000000_0000000000000000_0000100010011110_1100000001111101"; -- 0.033672361836577
	pesos_i(17674) := b"0000000000000000_0000000000000000_0000001100010100_1110100010000100"; -- 0.012037784818713477
	pesos_i(17675) := b"1111111111111111_1111111111111111_1110000000010110_1000110111110001"; -- -0.12465584638233858
	pesos_i(17676) := b"1111111111111111_1111111111111111_1111010000111001_0001110111011011"; -- -0.046003469399873695
	pesos_i(17677) := b"1111111111111111_1111111111111111_1111011001110000_0001100001010100"; -- -0.03735206564986624
	pesos_i(17678) := b"1111111111111111_1111111111111111_1111110100001011_0100101101000001"; -- -0.011546417764428746
	pesos_i(17679) := b"0000000000000000_0000000000000000_0000001101111111_1001000001100111"; -- 0.0136652233626037
	pesos_i(17680) := b"1111111111111111_1111111111111111_1110000101100011_1110011110111111"; -- -0.11956931669490402
	pesos_i(17681) := b"1111111111111111_1111111111111111_1111000010110101_0101000110010001"; -- -0.059733297344385525
	pesos_i(17682) := b"0000000000000000_0000000000000000_0000000110101011_1111010001101111"; -- 0.006530072386971741
	pesos_i(17683) := b"1111111111111111_1111111111111111_1110110010100101_1100111011101001"; -- -0.07559496703108447
	pesos_i(17684) := b"1111111111111111_1111111111111111_1111101111001001_0110011111110000"; -- -0.016458038305150288
	pesos_i(17685) := b"0000000000000000_0000000000000000_0000110000011100_0001001101010110"; -- 0.047303398514332524
	pesos_i(17686) := b"0000000000000000_0000000000000000_0001100001010101_0101100110111000"; -- 0.09505234466804394
	pesos_i(17687) := b"0000000000000000_0000000000000000_0001110110110010_1000001010101111"; -- 0.11600510376666874
	pesos_i(17688) := b"0000000000000000_0000000000000000_0000100001001010_1000010100011011"; -- 0.032387083997021664
	pesos_i(17689) := b"0000000000000000_0000000000000000_0010011000111111_1101010110111101"; -- 0.14941154358707576
	pesos_i(17690) := b"0000000000000000_0000000000000000_0001101000000110_0010011110001011"; -- 0.10165640965032596
	pesos_i(17691) := b"1111111111111111_1111111111111111_1110011110101000_0100011101100110"; -- -0.0950885177153004
	pesos_i(17692) := b"1111111111111111_1111111111111111_1110000110000101_0110100000111100"; -- -0.11905811820062456
	pesos_i(17693) := b"1111111111111111_1111111111111111_1110001111101111_0100011011100110"; -- -0.10963017353482445
	pesos_i(17694) := b"1111111111111111_1111111111111111_1110001001011110_1111001000101100"; -- -0.11573873923799391
	pesos_i(17695) := b"1111111111111111_1111111111111111_1111011001110010_1001011111000100"; -- -0.037313952002580905
	pesos_i(17696) := b"0000000000000000_0000000000000000_0001000010001100_1101000110101111"; -- 0.06464872861151708
	pesos_i(17697) := b"0000000000000000_0000000000000000_0001110010011011_1001011000011101"; -- 0.1117490597105054
	pesos_i(17698) := b"1111111111111111_1111111111111111_1111100011001111_1100100011010100"; -- -0.02807946042983304
	pesos_i(17699) := b"0000000000000000_0000000000000000_0001000100010000_1101000101000100"; -- 0.0666628639119648
	pesos_i(17700) := b"1111111111111111_1111111111111111_1110111101011001_0010011111000011"; -- -0.06504584785080512
	pesos_i(17701) := b"0000000000000000_0000000000000000_0000111000100011_0101000000010001"; -- 0.055226329844665675
	pesos_i(17702) := b"1111111111111111_1111111111111111_1101100100000111_0000111000010001"; -- -0.15223610016347408
	pesos_i(17703) := b"0000000000000000_0000000000000000_0001010010110100_0111101011111101"; -- 0.08087891267168175
	pesos_i(17704) := b"1111111111111111_1111111111111111_1110010110111000_0000000000010010"; -- -0.10266112856894553
	pesos_i(17705) := b"1111111111111111_1111111111111111_1111000001001010_1101011101111010"; -- -0.06135800612313222
	pesos_i(17706) := b"1111111111111111_1111111111111111_1111111111110100_0101100110001011"; -- -0.0001777682123431292
	pesos_i(17707) := b"0000000000000000_0000000000000000_0000101001010101_1100010010000000"; -- 0.04037120927021627
	pesos_i(17708) := b"1111111111111111_1111111111111111_1101101111000001_1101011001111001"; -- -0.1415735201071833
	pesos_i(17709) := b"1111111111111111_1111111111111111_1111110111101110_0000111111101110"; -- -0.008086208619026451
	pesos_i(17710) := b"0000000000000000_0000000000000000_0000100011000011_0101111100101110"; -- 0.03423113705926199
	pesos_i(17711) := b"0000000000000000_0000000000000000_0000100100010101_0000000011111011"; -- 0.0354767431118669
	pesos_i(17712) := b"1111111111111111_1111111111111111_1101101010000001_1001110001100100"; -- -0.1464597946609734
	pesos_i(17713) := b"0000000000000000_0000000000000000_0001101100100000_0100011001010000"; -- 0.10596122219577433
	pesos_i(17714) := b"1111111111111111_1111111111111111_1101101100000001_1100100111000011"; -- -0.14450396524891024
	pesos_i(17715) := b"0000000000000000_0000000000000000_0001010010100110_0100010101101111"; -- 0.0806620975191963
	pesos_i(17716) := b"1111111111111111_1111111111111111_1110010101000100_0000000111111100"; -- -0.10443103406619571
	pesos_i(17717) := b"1111111111111111_1111111111111111_1111101110110010_0110001100111000"; -- -0.016809271663980753
	pesos_i(17718) := b"0000000000000000_0000000000000000_0010000001010111_0110110100100010"; -- 0.12633401938193148
	pesos_i(17719) := b"0000000000000000_0000000000000000_0000100101111100_0000001110101100"; -- 0.03704855873108019
	pesos_i(17720) := b"0000000000000000_0000000000000000_0001001110010110_0001011101000000"; -- 0.07650895408896517
	pesos_i(17721) := b"1111111111111111_1111111111111111_1111000110100010_1000010111100110"; -- -0.056113845258880836
	pesos_i(17722) := b"1111111111111111_1111111111111111_1111000100110011_0010100100001101"; -- -0.05781310490965821
	pesos_i(17723) := b"0000000000000000_0000000000000000_0000110110110111_1010011001111110"; -- 0.0535835321821869
	pesos_i(17724) := b"0000000000000000_0000000000000000_0000010010111001_0100110010010011"; -- 0.018452440234157562
	pesos_i(17725) := b"1111111111111111_1111111111111111_1111011111010110_1011100110101000"; -- -0.03187980325874232
	pesos_i(17726) := b"1111111111111111_1111111111111111_1101111000010100_1111010110111001"; -- -0.13249267795957476
	pesos_i(17727) := b"0000000000000000_0000000000000000_0001011100011001_0111010011010110"; -- 0.09023218359508692
	pesos_i(17728) := b"1111111111111111_1111111111111111_1111111100000101_0100010110011111"; -- -0.0038258062296420018
	pesos_i(17729) := b"0000000000000000_0000000000000000_0001000011100000_1011001111000100"; -- 0.0659286835097244
	pesos_i(17730) := b"0000000000000000_0000000000000000_0010010010110111_0001111111111011"; -- 0.14341926456874293
	pesos_i(17731) := b"1111111111111111_1111111111111111_1110010100001110_1111110011101100"; -- -0.10524005168127713
	pesos_i(17732) := b"1111111111111111_1111111111111111_1110010000001000_0010001000111000"; -- -0.10925089020282858
	pesos_i(17733) := b"0000000000000000_0000000000000000_0000100101011001_0001000100110000"; -- 0.03651530673643753
	pesos_i(17734) := b"0000000000000000_0000000000000000_0000011100110110_1101000000001111"; -- 0.02818012584209413
	pesos_i(17735) := b"1111111111111111_1111111111111111_1111010110110101_0011001011110110"; -- -0.04020387157853893
	pesos_i(17736) := b"0000000000000000_0000000000000000_0001001011100010_1100010000000111"; -- 0.0737726704195436
	pesos_i(17737) := b"1111111111111111_1111111111111111_1110111101001111_1000010100010110"; -- -0.0651928730543973
	pesos_i(17738) := b"0000000000000000_0000000000000000_0001100101101110_0001101001001011"; -- 0.09933628406016719
	pesos_i(17739) := b"0000000000000000_0000000000000000_0001100001110000_0000100111101010"; -- 0.09545957518423531
	pesos_i(17740) := b"1111111111111111_1111111111111111_1110111111100100_0101100010110000"; -- -0.06292195990432116
	pesos_i(17741) := b"1111111111111111_1111111111111111_1110110000001101_0000101100001011"; -- -0.07792597742816343
	pesos_i(17742) := b"0000000000000000_0000000000000000_0001010110110001_0101000111000000"; -- 0.084736928316322
	pesos_i(17743) := b"0000000000000000_0000000000000000_0010001110101100_1011011100011011"; -- 0.13935417570664624
	pesos_i(17744) := b"1111111111111111_1111111111111111_1110010100110010_0010110010110110"; -- -0.10470314556276113
	pesos_i(17745) := b"0000000000000000_0000000000000000_0010001010110011_0111111111110111"; -- 0.1355514506144644
	pesos_i(17746) := b"0000000000000000_0000000000000000_0000001111101001_0011110101001101"; -- 0.015277701682436001
	pesos_i(17747) := b"1111111111111111_1111111111111111_1111111111011110_0001110101111001"; -- -0.0005170420769837707
	pesos_i(17748) := b"1111111111111111_1111111111111111_1111100101001010_1101110000101111"; -- -0.026201475615839104
	pesos_i(17749) := b"1111111111111111_1111111111111111_1111101001011100_1001100000001111"; -- -0.022024628011259654
	pesos_i(17750) := b"1111111111111111_1111111111111111_1110100111000100_0101100011001100"; -- -0.08684773463420098
	pesos_i(17751) := b"1111111111111111_1111111111111111_1101100110010100_1001100010010110"; -- -0.15007635431678482
	pesos_i(17752) := b"1111111111111111_1111111111111111_1111011010110010_1001101111010001"; -- -0.036337148148840225
	pesos_i(17753) := b"1111111111111111_1111111111111111_1101101110101011_0111011010001111"; -- -0.14191493037211542
	pesos_i(17754) := b"1111111111111111_1111111111111111_1110001001110000_1101110100010001"; -- -0.11546533913454286
	pesos_i(17755) := b"1111111111111111_1111111111111111_1101101010001011_0111110001000111"; -- -0.14630912092976395
	pesos_i(17756) := b"1111111111111111_1111111111111111_1111000010111010_1011111100101110"; -- -0.05965047006677669
	pesos_i(17757) := b"1111111111111111_1111111111111111_1110010101001011_0001110000111010"; -- -0.10432265844663842
	pesos_i(17758) := b"1111111111111111_1111111111111111_1101100111100011_0000100000010011"; -- -0.14887952352281808
	pesos_i(17759) := b"1111111111111111_1111111111111111_1111010011010100_0111111010111101"; -- -0.04363258251557352
	pesos_i(17760) := b"1111111111111111_1111111111111111_1111111000001101_1110011010010101"; -- -0.007600391904985342
	pesos_i(17761) := b"1111111111111111_1111111111111111_1110111000000010_1001111111011011"; -- -0.07027245418301288
	pesos_i(17762) := b"1111111111111111_1111111111111111_1110110000101000_0001100000101101"; -- -0.07751320737933173
	pesos_i(17763) := b"0000000000000000_0000000000000000_0010001100111100_0100001111001111"; -- 0.13763831910629615
	pesos_i(17764) := b"0000000000000000_0000000000000000_0000111101100101_1111110000101110"; -- 0.060149918713936476
	pesos_i(17765) := b"0000000000000000_0000000000000000_0001001000100001_0000110110010011"; -- 0.0708168490645536
	pesos_i(17766) := b"1111111111111111_1111111111111111_1101101101010100_1101101110111110"; -- -0.14323641399387319
	pesos_i(17767) := b"0000000000000000_0000000000000000_0000001011011001_0011011011001010"; -- 0.0111269229632399
	pesos_i(17768) := b"0000000000000000_0000000000000000_0000110110001010_1001101000001101"; -- 0.05289614492925398
	pesos_i(17769) := b"1111111111111111_1111111111111111_1111101011001100_1000000011001001"; -- -0.020317030755152687
	pesos_i(17770) := b"0000000000000000_0000000000000000_0010001101000010_0111000001010001"; -- 0.13773252464889224
	pesos_i(17771) := b"0000000000000000_0000000000000000_0010011110101010_1001110010001101"; -- 0.15494707521372267
	pesos_i(17772) := b"1111111111111111_1111111111111111_1110111110011011_0111110000101100"; -- -0.06403373656136875
	pesos_i(17773) := b"0000000000000000_0000000000000000_0010000001110011_1010100011000000"; -- 0.12676481905688988
	pesos_i(17774) := b"0000000000000000_0000000000000000_0010011100011110_1001010111100011"; -- 0.15281044770210842
	pesos_i(17775) := b"1111111111111111_1111111111111111_1110111101101110_0110000000000111"; -- -0.0647220594537153
	pesos_i(17776) := b"1111111111111111_1111111111111111_1110001011011111_1110010101000110"; -- -0.11377112428005351
	pesos_i(17777) := b"1111111111111111_1111111111111111_1111001110010011_1011011010101001"; -- -0.04852732071471415
	pesos_i(17778) := b"0000000000000000_0000000000000000_0010001001011000_1011010010000011"; -- 0.13416603284211898
	pesos_i(17779) := b"0000000000000000_0000000000000000_0001101111000101_1001010010001100"; -- 0.10848358554718492
	pesos_i(17780) := b"0000000000000000_0000000000000000_0000111100110000_0111000101100011"; -- 0.05933293030273884
	pesos_i(17781) := b"0000000000000000_0000000000000000_0000001010111111_0010110101111011"; -- 0.010729639503002411
	pesos_i(17782) := b"0000000000000000_0000000000000000_0000111110000010_1011010000011010"; -- 0.06058812741801551
	pesos_i(17783) := b"1111111111111111_1111111111111111_1111110011111000_0101101100000011"; -- -0.011835395683382644
	pesos_i(17784) := b"1111111111111111_1111111111111111_1111010111010110_1100010111000100"; -- -0.039691581428122985
	pesos_i(17785) := b"0000000000000000_0000000000000000_0000111111001101_0001001000000100"; -- 0.06172287557798392
	pesos_i(17786) := b"1111111111111111_1111111111111111_1110101110000100_1000011010101001"; -- -0.08000906345970561
	pesos_i(17787) := b"1111111111111111_1111111111111111_1111011000010011_0101011101100111"; -- -0.03876737352238819
	pesos_i(17788) := b"1111111111111111_1111111111111111_1110111100111101_1010010111001000"; -- -0.06546558252408381
	pesos_i(17789) := b"1111111111111111_1111111111111111_1111000100110111_1110011100110110"; -- -0.057740735332046295
	pesos_i(17790) := b"1111111111111111_1111111111111111_1111000011111100_1011011101010111"; -- -0.05864385713602134
	pesos_i(17791) := b"1111111111111111_1111111111111111_1111111011110100_0010101011101000"; -- -0.004086797941147298
	pesos_i(17792) := b"0000000000000000_0000000000000000_0001011001100101_0010110010011000"; -- 0.08748129557387697
	pesos_i(17793) := b"0000000000000000_0000000000000000_0001111100000111_1111111011100111"; -- 0.12121575490279941
	pesos_i(17794) := b"1111111111111111_1111111111111111_1111101100010000_0010011001101111"; -- -0.019284818659870223
	pesos_i(17795) := b"0000000000000000_0000000000000000_0001100011011111_0101000001011110"; -- 0.09715750018788771
	pesos_i(17796) := b"0000000000000000_0000000000000000_0000011111000010_1011000010011000"; -- 0.030314480771284607
	pesos_i(17797) := b"1111111111111111_1111111111111111_1110010000111011_1100110100011011"; -- -0.10846250617754115
	pesos_i(17798) := b"1111111111111111_1111111111111111_1110000010111100_0001110110101000"; -- -0.12212957998692767
	pesos_i(17799) := b"0000000000000000_0000000000000000_0001111000010010_0011100011101001"; -- 0.11746555030813635
	pesos_i(17800) := b"0000000000000000_0000000000000000_0001111001000100_0010011111010000"; -- 0.11822747069391525
	pesos_i(17801) := b"0000000000000000_0000000000000000_0000011000010110_0111010011010111"; -- 0.023780157546471708
	pesos_i(17802) := b"1111111111111111_1111111111111111_1110000110010011_1110101010110100"; -- -0.11883671862170549
	pesos_i(17803) := b"0000000000000000_0000000000000000_0000110100001011_1101011101100010"; -- 0.05096193440863193
	pesos_i(17804) := b"1111111111111111_1111111111111111_1110110100011010_0100011000010111"; -- -0.07381784388318156
	pesos_i(17805) := b"1111111111111111_1111111111111111_1111101000001000_0100100101001010"; -- -0.023311061285381393
	pesos_i(17806) := b"0000000000000000_0000000000000000_0001111010000101_1001101000111010"; -- 0.11922611155126026
	pesos_i(17807) := b"0000000000000000_0000000000000000_0000101111100000_1011011011101001"; -- 0.04639762109542577
	pesos_i(17808) := b"0000000000000000_0000000000000000_0000001101010101_0100110100000010"; -- 0.013020337198533651
	pesos_i(17809) := b"0000000000000000_0000000000000000_0001101101000011_1010111010011100"; -- 0.10650149648072002
	pesos_i(17810) := b"1111111111111111_1111111111111111_1110011111011101_1001000110110010"; -- -0.09427537347718729
	pesos_i(17811) := b"1111111111111111_1111111111111111_1111110010001000_1011010000101100"; -- -0.013539065551483442
	pesos_i(17812) := b"1111111111111111_1111111111111111_1111110101100101_1110100111010001"; -- -0.010163675853885572
	pesos_i(17813) := b"0000000000000000_0000000000000000_0001110110101111_1100100001011110"; -- 0.1159634809802793
	pesos_i(17814) := b"0000000000000000_0000000000000000_0000101010111110_1111101000011010"; -- 0.041976577091315935
	pesos_i(17815) := b"0000000000000000_0000000000000000_0001000010010110_1011000001100011"; -- 0.06479933176548244
	pesos_i(17816) := b"0000000000000000_0000000000000000_0010001001111011_1000100001001111"; -- 0.13469745562778213
	pesos_i(17817) := b"1111111111111111_1111111111111111_1110001100100001_1011010000000010"; -- -0.11276698058364573
	pesos_i(17818) := b"0000000000000000_0000000000000000_0000101010101100_0000100000111110"; -- 0.04168750295759362
	pesos_i(17819) := b"0000000000000000_0000000000000000_0001100101001001_1010111000001000"; -- 0.0987805146674831
	pesos_i(17820) := b"1111111111111111_1111111111111111_1110100101010111_0000111111111100"; -- -0.08851528269247017
	pesos_i(17821) := b"1111111111111111_1111111111111111_1110110110000010_1011011000111110"; -- -0.07222424495851006
	pesos_i(17822) := b"1111111111111111_1111111111111111_1111010101011101_1010111010111011"; -- -0.04153926790003913
	pesos_i(17823) := b"1111111111111111_1111111111111111_1110110110011011_0110101010011011"; -- -0.07184728362890239
	pesos_i(17824) := b"0000000000000000_0000000000000000_0001100010011011_1111000011000100"; -- 0.09612946304917902
	pesos_i(17825) := b"1111111111111111_1111111111111111_1110110101010101_0101000010111010"; -- -0.07291694132045233
	pesos_i(17826) := b"1111111111111111_1111111111111111_1110101010110011_1001110100101000"; -- -0.08319680947296984
	pesos_i(17827) := b"0000000000000000_0000000000000000_0000011011000110_0110000001000011"; -- 0.02646447778578043
	pesos_i(17828) := b"1111111111111111_1111111111111111_1111000111000111_0011101110101011"; -- -0.05555369449159547
	pesos_i(17829) := b"0000000000000000_0000000000000000_0001101111010100_1111110010111001"; -- 0.10871867669663961
	pesos_i(17830) := b"1111111111111111_1111111111111111_1111101100011000_0100111011111001"; -- -0.019160331826534167
	pesos_i(17831) := b"0000000000000000_0000000000000000_0010001000101111_0110000011110111"; -- 0.13353544261444839
	pesos_i(17832) := b"0000000000000000_0000000000000000_0000101100101010_1110011011000101"; -- 0.04362337418451445
	pesos_i(17833) := b"0000000000000000_0000000000000000_0000011000000111_0001110001001011"; -- 0.023545997958642338
	pesos_i(17834) := b"1111111111111111_1111111111111111_1110010111101111_0010001001001010"; -- -0.10181985556279728
	pesos_i(17835) := b"0000000000000000_0000000000000000_0001111111001100_0001010011001001"; -- 0.12420778176896277
	pesos_i(17836) := b"1111111111111111_1111111111111111_1110000001000011_0010100000100111"; -- -0.12397526793475314
	pesos_i(17837) := b"0000000000000000_0000000000000000_0000110010100101_1110000010011001"; -- 0.0494060872619095
	pesos_i(17838) := b"0000000000000000_0000000000000000_0010001000000101_1010000000011010"; -- 0.13289833676176663
	pesos_i(17839) := b"0000000000000000_0000000000000000_0001011101100110_1000110001110011"; -- 0.09140851783259085
	pesos_i(17840) := b"0000000000000000_0000000000000000_0010001101101110_0110110111100101"; -- 0.13840376709856242
	pesos_i(17841) := b"0000000000000000_0000000000000000_0001001001001110_1010010000010010"; -- 0.07151246498381011
	pesos_i(17842) := b"0000000000000000_0000000000000000_0000001101010111_1001100000000000"; -- 0.013055324466858712
	pesos_i(17843) := b"0000000000000000_0000000000000000_0001100001100010_0001001111100011"; -- 0.0952465467366918
	pesos_i(17844) := b"0000000000000000_0000000000000000_0001000110101001_0011110101010001"; -- 0.06898864016508888
	pesos_i(17845) := b"0000000000000000_0000000000000000_0000001111101110_1100000001100011"; -- 0.015361808919923161
	pesos_i(17846) := b"1111111111111111_1111111111111111_1111010010000010_0011000001001110"; -- -0.0448884782344507
	pesos_i(17847) := b"1111111111111111_1111111111111111_1111000010011111_0000100110010011"; -- -0.0600732819052724
	pesos_i(17848) := b"1111111111111111_1111111111111111_1101110101110010_1100100010011111"; -- -0.13496729005511637
	pesos_i(17849) := b"0000000000000000_0000000000000000_0000110111011110_0000010011110001"; -- 0.054168995644473916
	pesos_i(17850) := b"1111111111111111_1111111111111111_1111010000011101_1101001100100001"; -- -0.046419910814608854
	pesos_i(17851) := b"0000000000000000_0000000000000000_0000101011000001_1100010101111100"; -- 0.04201921723528174
	pesos_i(17852) := b"0000000000000000_0000000000000000_0000001010000001_0110110100010010"; -- 0.009787384839701749
	pesos_i(17853) := b"0000000000000000_0000000000000000_0001101100001111_1010001110000001"; -- 0.1057073774738402
	pesos_i(17854) := b"1111111111111111_1111111111111111_1110110101111001_1110011010101000"; -- -0.07235868828156039
	pesos_i(17855) := b"1111111111111111_1111111111111111_1111111001110001_1100000000101000"; -- -0.006076803346883191
	pesos_i(17856) := b"1111111111111111_1111111111111111_1111010110010010_0001110111001101"; -- -0.04073919059177261
	pesos_i(17857) := b"1111111111111111_1111111111111111_1110110001011000_1001010000011100"; -- -0.07677339847022456
	pesos_i(17858) := b"1111111111111111_1111111111111111_1111111100111000_0001111011001101"; -- -0.003049922017054317
	pesos_i(17859) := b"0000000000000000_0000000000000000_0000110111101011_0000001000100011"; -- 0.05436719276682413
	pesos_i(17860) := b"0000000000000000_0000000000000000_0000100101011001_0110110101100000"; -- 0.03652080156644192
	pesos_i(17861) := b"1111111111111111_1111111111111111_1110010001010111_1100011001111010"; -- -0.10803565524661739
	pesos_i(17862) := b"0000000000000000_0000000000000000_0001101111110101_0001000000111000"; -- 0.10920812014189127
	pesos_i(17863) := b"1111111111111111_1111111111111111_1111000100101110_1111100100010010"; -- -0.057876999885152554
	pesos_i(17864) := b"1111111111111111_1111111111111111_1110000000011011_1110000110110100"; -- -0.12457455981790294
	pesos_i(17865) := b"1111111111111111_1111111111111111_1111110101100100_0101000111000111"; -- -0.010187996740585513
	pesos_i(17866) := b"0000000000000000_0000000000000000_0001011100100110_1010111010110010"; -- 0.09043399672047447
	pesos_i(17867) := b"0000000000000000_0000000000000000_0001000010111101_1110010111100100"; -- 0.06539761376544573
	pesos_i(17868) := b"1111111111111111_1111111111111111_1111101010110110_0101010011011011"; -- -0.0206553426983796
	pesos_i(17869) := b"0000000000000000_0000000000000000_0010100100000000_0000110010110001"; -- 0.16015700638750208
	pesos_i(17870) := b"1111111111111111_1111111111111111_1110100010110100_0010010011100010"; -- -0.09100121954129353
	pesos_i(17871) := b"1111111111111111_1111111111111111_1111101010101000_0010110000101110"; -- -0.020871390115562907
	pesos_i(17872) := b"1111111111111111_1111111111111111_1110111101101000_0001000110000100"; -- -0.06481829185318182
	pesos_i(17873) := b"1111111111111111_1111111111111111_1110001111110111_1110100111000010"; -- -0.10949839608948819
	pesos_i(17874) := b"0000000000000000_0000000000000000_0000000000010010_1111001110001100"; -- 0.0002891747831114147
	pesos_i(17875) := b"1111111111111111_1111111111111111_1111010101000001_1001111100100110"; -- -0.04196744271916586
	pesos_i(17876) := b"1111111111111111_1111111111111111_1111111100011101_1111110000100110"; -- -0.0034487158316411633
	pesos_i(17877) := b"0000000000000000_0000000000000000_0010010001000011_1110011111011001"; -- 0.1416611581597958
	pesos_i(17878) := b"1111111111111111_1111111111111111_1101101010011011_0110100010010001"; -- -0.14606615499116465
	pesos_i(17879) := b"1111111111111111_1111111111111111_1101101110101100_1011100110000101"; -- -0.1418956804313066
	pesos_i(17880) := b"1111111111111111_1111111111111111_1101110010010001_1100000000011110"; -- -0.13840102455956355
	pesos_i(17881) := b"1111111111111111_1111111111111111_1110111111011010_1000110001010100"; -- -0.06307146987643804
	pesos_i(17882) := b"0000000000000000_0000000000000000_0001101010100100_1001010001010100"; -- 0.10407378238271306
	pesos_i(17883) := b"0000000000000000_0000000000000000_0001100010010000_1101010010101111"; -- 0.09595994259138307
	pesos_i(17884) := b"1111111111111111_1111111111111111_1111110100001001_0011111110000101"; -- -0.011577634816960893
	pesos_i(17885) := b"0000000000000000_0000000000000000_0010011011110110_0101001101111011"; -- 0.15219613803744214
	pesos_i(17886) := b"1111111111111111_1111111111111111_1110101100110101_0010000101001111"; -- -0.08122054888360705
	pesos_i(17887) := b"0000000000000000_0000000000000000_0000000011001111_0001011011001011"; -- 0.0031599278550478046
	pesos_i(17888) := b"1111111111111111_1111111111111111_1111101100110100_0000111010100110"; -- -0.0187369199195718
	pesos_i(17889) := b"0000000000000000_0000000000000000_0010010001010011_1000110000001101"; -- 0.14189982721898614
	pesos_i(17890) := b"1111111111111111_1111111111111111_1111100110010000_1101101100010101"; -- -0.025133426139057988
	pesos_i(17891) := b"1111111111111111_1111111111111111_1110111100010011_0011110110010011"; -- -0.06611266292788
	pesos_i(17892) := b"0000000000000000_0000000000000000_0000000000101010_0011110000101001"; -- 0.0006444550104517985
	pesos_i(17893) := b"1111111111111111_1111111111111111_1110110111100100_0010100001001001"; -- -0.07073734494182177
	pesos_i(17894) := b"0000000000000000_0000000000000000_0001100000110101_1100001011001010"; -- 0.09457032615171966
	pesos_i(17895) := b"1111111111111111_1111111111111111_1111011110001011_0100111001000100"; -- -0.033030613228364716
	pesos_i(17896) := b"0000000000000000_0000000000000000_0000101011101111_1110000011100100"; -- 0.04272275516142427
	pesos_i(17897) := b"0000000000000000_0000000000000000_0000010011001111_0111011011001011"; -- 0.01879065000140101
	pesos_i(17898) := b"1111111111111111_1111111111111111_1101101011001000_0110111011101001"; -- -0.1453791314631553
	pesos_i(17899) := b"0000000000000000_0000000000000000_0001101011100110_1001110100110101"; -- 0.1050813917942424
	pesos_i(17900) := b"0000000000000000_0000000000000000_0010001010100000_1000001111111111"; -- 0.13526177379187987
	pesos_i(17901) := b"1111111111111111_1111111111111111_1110101000001100_1101011110001000"; -- -0.08574154795832228
	pesos_i(17902) := b"0000000000000000_0000000000000000_0000011001000010_1101100001000001"; -- 0.02445746988354392
	pesos_i(17903) := b"1111111111111111_1111111111111111_1110000001000011_0011011001100101"; -- -0.1239744189101961
	pesos_i(17904) := b"0000000000000000_0000000000000000_0000100001000101_1011111101110110"; -- 0.032314268408027064
	pesos_i(17905) := b"0000000000000000_0000000000000000_0000011110001100_1101111100000011"; -- 0.029493273095199654
	pesos_i(17906) := b"0000000000000000_0000000000000000_0010000010001100_1010001011111111"; -- 0.12714594588639794
	pesos_i(17907) := b"0000000000000000_0000000000000000_0000001001000010_0101111011100100"; -- 0.008825235946039848
	pesos_i(17908) := b"1111111111111111_1111111111111111_1110111000110010_1100010110111010"; -- -0.06953777519110553
	pesos_i(17909) := b"0000000000000000_0000000000000000_0001001000011001_0100001110011011"; -- 0.07069799929088737
	pesos_i(17910) := b"1111111111111111_1111111111111111_1111111001111111_1111100001001111"; -- -0.005859833403494226
	pesos_i(17911) := b"0000000000000000_0000000000000000_0001010110011011_0010010000110101"; -- 0.08439852034192787
	pesos_i(17912) := b"1111111111111111_1111111111111111_1101110100111100_1100010101010100"; -- -0.13579146089659966
	pesos_i(17913) := b"0000000000000000_0000000000000000_0000100000101111_0001101101001010"; -- 0.031968789531905524
	pesos_i(17914) := b"1111111111111111_1111111111111111_1111000001010010_1100010111010010"; -- -0.0612369883480303
	pesos_i(17915) := b"0000000000000000_0000000000000000_0010101000110001_1110110100011001"; -- 0.16482431287175417
	pesos_i(17916) := b"1111111111111111_1111111111111111_1111010101111011_1010110011110000"; -- -0.041081610969733846
	pesos_i(17917) := b"1111111111111111_1111111111111111_1110000000110011_0000001010101110"; -- -0.12422164213740794
	pesos_i(17918) := b"1111111111111111_1111111111111111_1101100101111111_1000001010101101"; -- -0.15039809496600662
	pesos_i(17919) := b"1111111111111111_1111111111111111_1111010101110111_0000010101010111"; -- -0.04115263581174801
	pesos_i(17920) := b"1111111111111111_1111111111111111_1111010011101101_1110010110010111"; -- -0.04324498238690944
	pesos_i(17921) := b"1111111111111111_1111111111111111_1111111110110010_1000111110000110"; -- -0.0011816309814309152
	pesos_i(17922) := b"1111111111111111_1111111111111111_1111111010111011_1111110011010001"; -- -0.004944037346244727
	pesos_i(17923) := b"0000000000000000_0000000000000000_0010000111010110_1010010001100110"; -- 0.13218142981912126
	pesos_i(17924) := b"1111111111111111_1111111111111111_1111000100010010_1101011110111100"; -- -0.058306233107506385
	pesos_i(17925) := b"1111111111111111_1111111111111111_1111100010100001_1101011000010000"; -- -0.0287805759277856
	pesos_i(17926) := b"1111111111111111_1111111111111111_1111111000001011_1111111101110101"; -- -0.007629426818300195
	pesos_i(17927) := b"0000000000000000_0000000000000000_0000110100111111_1111101110100001"; -- 0.05175755189704061
	pesos_i(17928) := b"1111111111111111_1111111111111111_1111010001000010_0000101110010000"; -- -0.04586723082605335
	pesos_i(17929) := b"0000000000000000_0000000000000000_0010011000110110_0110100010101001"; -- 0.1492677129117376
	pesos_i(17930) := b"0000000000000000_0000000000000000_0010101001001010_1110100000011100"; -- 0.1652054853038164
	pesos_i(17931) := b"0000000000000000_0000000000000000_0000000000101000_0001011001011101"; -- 0.0006116844617773138
	pesos_i(17932) := b"1111111111111111_1111111111111111_1111101110010010_0111011000110000"; -- -0.017296422206230306
	pesos_i(17933) := b"0000000000000000_0000000000000000_0010010011111001_0011011011011000"; -- 0.14442770742644323
	pesos_i(17934) := b"1111111111111111_1111111111111111_1110111101100001_1011100110101111"; -- -0.06491507978019788
	pesos_i(17935) := b"0000000000000000_0000000000000000_0001100011100100_1001001100001010"; -- 0.09723776813585247
	pesos_i(17936) := b"0000000000000000_0000000000000000_0000001011010010_1101101001011010"; -- 0.011029860371190244
	pesos_i(17937) := b"0000000000000000_0000000000000000_0000000100000001_1001110001001010"; -- 0.00393082425953678
	pesos_i(17938) := b"0000000000000000_0000000000000000_0010010110010011_1000101001101011"; -- 0.1467825422791202
	pesos_i(17939) := b"1111111111111111_1111111111111111_1101110110111111_1000000110000111"; -- -0.1337966008540396
	pesos_i(17940) := b"0000000000000000_0000000000000000_0000000001110001_1001110100101101"; -- 0.0017336115664950396
	pesos_i(17941) := b"0000000000000000_0000000000000000_0000110100110110_1111011110010001"; -- 0.05161998077749029
	pesos_i(17942) := b"1111111111111111_1111111111111111_1110001011100110_1101100110110001"; -- -0.11366500301888363
	pesos_i(17943) := b"1111111111111111_1111111111111111_1111101000111011_0101000011001010"; -- -0.0225324160269867
	pesos_i(17944) := b"1111111111111111_1111111111111111_1110111011010100_0000001110000011"; -- -0.06707742740239614
	pesos_i(17945) := b"1111111111111111_1111111111111111_1111001001000001_1011101110011111"; -- -0.05368449564737194
	pesos_i(17946) := b"1111111111111111_1111111111111111_1111010101001010_0010000000111011"; -- -0.04183767859210968
	pesos_i(17947) := b"1111111111111111_1111111111111111_1110010111010010_1000010011101111"; -- -0.10225648088284628
	pesos_i(17948) := b"0000000000000000_0000000000000000_0000100001101000_1011110001100000"; -- 0.032848142080528414
	pesos_i(17949) := b"1111111111111111_1111111111111111_1101111000110111_1111101000101100"; -- -0.1319583552617255
	pesos_i(17950) := b"0000000000000000_0000000000000000_0001100001100010_1010001110001000"; -- 0.09525510863210941
	pesos_i(17951) := b"0000000000000000_0000000000000000_0010000111010110_1000001000011100"; -- 0.13217938594525358
	pesos_i(17952) := b"1111111111111111_1111111111111111_1110011001000001_1111110110101100"; -- -0.10055555860792129
	pesos_i(17953) := b"0000000000000000_0000000000000000_0000001011111001_1001011001011100"; -- 0.011620900680862316
	pesos_i(17954) := b"1111111111111111_1111111111111111_1111011110101011_0100101000110010"; -- -0.032542574764428754
	pesos_i(17955) := b"1111111111111111_1111111111111111_1111000001000000_0001001011100011"; -- -0.06152231180186595
	pesos_i(17956) := b"1111111111111111_1111111111111111_1110001111100011_1010010000000000"; -- -0.1098077296086965
	pesos_i(17957) := b"1111111111111111_1111111111111111_1110001011100000_1110000011000000"; -- -0.11375613520989072
	pesos_i(17958) := b"1111111111111111_1111111111111111_1111100110101010_1011101000000101"; -- -0.02473866822008005
	pesos_i(17959) := b"1111111111111111_1111111111111111_1101100100101100_1001100001000000"; -- -0.15166328851823793
	pesos_i(17960) := b"1111111111111111_1111111111111111_1110010101000101_0011101011101001"; -- -0.10441238228867233
	pesos_i(17961) := b"1111111111111111_1111111111111111_1111100010101011_1110100011100111"; -- -0.028626865094427908
	pesos_i(17962) := b"1111111111111111_1111111111111111_1110100010000111_0101100100011000"; -- -0.0916847530233903
	pesos_i(17963) := b"1111111111111111_1111111111111111_1111100010101110_1110001101100101"; -- -0.028581416922422727
	pesos_i(17964) := b"0000000000000000_0000000000000000_0000100110110000_0101100100111001"; -- 0.03784711493569538
	pesos_i(17965) := b"1111111111111111_1111111111111111_1111011100111111_0001011010000011"; -- -0.03419360448163474
	pesos_i(17966) := b"1111111111111111_1111111111111111_1111010111101110_1111110111010101"; -- -0.039322028647997526
	pesos_i(17967) := b"1111111111111111_1111111111111111_1111110010011110_0110101100100000"; -- -0.013207726266653796
	pesos_i(17968) := b"1111111111111111_1111111111111111_1110110001001011_1010101101101101"; -- -0.07697037309086087
	pesos_i(17969) := b"0000000000000000_0000000000000000_0010010010101101_1011010101010111"; -- 0.1432755791148949
	pesos_i(17970) := b"0000000000000000_0000000000000000_0000100000011000_0100010010001100"; -- 0.03162029659907124
	pesos_i(17971) := b"0000000000000000_0000000000000000_0010011100100100_0001111100101001"; -- 0.15289492368965468
	pesos_i(17972) := b"0000000000000000_0000000000000000_0010001100010111_1111100111000100"; -- 0.13708458923502054
	pesos_i(17973) := b"0000000000000000_0000000000000000_0000011001011111_1001100010101111"; -- 0.024896185572830003
	pesos_i(17974) := b"1111111111111111_1111111111111111_1110110110001001_0101001101010001"; -- -0.07212332977617458
	pesos_i(17975) := b"1111111111111111_1111111111111111_1111010011011011_1001011110111010"; -- -0.04352428153766549
	pesos_i(17976) := b"1111111111111111_1111111111111111_1110010110000010_1101001010001000"; -- -0.10347255868142963
	pesos_i(17977) := b"0000000000000000_0000000000000000_0000010011100000_0100011101000101"; -- 0.019047216782453927
	pesos_i(17978) := b"1111111111111111_1111111111111111_1111010101100101_0001110110110110"; -- -0.04142584144133741
	pesos_i(17979) := b"1111111111111111_1111111111111111_1101110000110011_1000101011000111"; -- -0.13983853001946
	pesos_i(17980) := b"0000000000000000_0000000000000000_0001111001010000_0111001011001101"; -- 0.11841504588352608
	pesos_i(17981) := b"0000000000000000_0000000000000000_0001000001000010_0010011101011011"; -- 0.06350942576654935
	pesos_i(17982) := b"0000000000000000_0000000000000000_0001000000000001_0001100010011000"; -- 0.06251672462475895
	pesos_i(17983) := b"1111111111111111_1111111111111111_1110001000010111_1110111101010100"; -- -0.11682228280371541
	pesos_i(17984) := b"0000000000000000_0000000000000000_0000100011010101_0110100110100010"; -- 0.03450641836782989
	pesos_i(17985) := b"0000000000000000_0000000000000000_0010001111101111_0001011000101100"; -- 0.14036692202375675
	pesos_i(17986) := b"0000000000000000_0000000000000000_0001011011111101_1110101111001011"; -- 0.08981202799368106
	pesos_i(17987) := b"0000000000000000_0000000000000000_0000001001010100_1000011111001000"; -- 0.009102331473811084
	pesos_i(17988) := b"1111111111111111_1111111111111111_1110101010110011_0110101000100000"; -- -0.08319985127227682
	pesos_i(17989) := b"0000000000000000_0000000000000000_0000111001111110_0011010010000101"; -- 0.05661323774920881
	pesos_i(17990) := b"1111111111111111_1111111111111111_1110110100000111_0100010010000011"; -- -0.07410785483242843
	pesos_i(17991) := b"0000000000000000_0000000000000000_0000000111001101_1111000010010000"; -- 0.007048640449589833
	pesos_i(17992) := b"0000000000000000_0000000000000000_0001110100011110_1001000101100001"; -- 0.11374767886886948
	pesos_i(17993) := b"1111111111111111_1111111111111111_1101101011000110_0001001101001001"; -- -0.14541511025037993
	pesos_i(17994) := b"1111111111111111_1111111111111111_1101110110100101_0101000010100100"; -- -0.13419624319697707
	pesos_i(17995) := b"1111111111111111_1111111111111111_1110100110111110_0000010010011111"; -- -0.08694430463613892
	pesos_i(17996) := b"0000000000000000_0000000000000000_0001000010010110_0010100101001111"; -- 0.06479128052445898
	pesos_i(17997) := b"1111111111111111_1111111111111111_1110101000101011_1101011011111011"; -- -0.08526855823084796
	pesos_i(17998) := b"0000000000000000_0000000000000000_0001111000000100_0111000100000111"; -- 0.11725527204026795
	pesos_i(17999) := b"0000000000000000_0000000000000000_0000001011011011_0101101011001000"; -- 0.01115958580308403
	pesos_i(18000) := b"1111111111111111_1111111111111111_1110010011010111_0100111011101000"; -- -0.10608965727552655
	pesos_i(18001) := b"0000000000000000_0000000000000000_0001011100100010_0110010001000110"; -- 0.09036852556568364
	pesos_i(18002) := b"0000000000000000_0000000000000000_0000011101001100_0100010011110111"; -- 0.028507528570939474
	pesos_i(18003) := b"0000000000000000_0000000000000000_0000111001000101_0001001100110001"; -- 0.05574150025027285
	pesos_i(18004) := b"0000000000000000_0000000000000000_0001000000100100_0001101000000110"; -- 0.06305086753445784
	pesos_i(18005) := b"0000000000000000_0000000000000000_0000010101111111_1101000101111100"; -- 0.021481602353257526
	pesos_i(18006) := b"1111111111111111_1111111111111111_1111101100011110_0011110000110111"; -- -0.01906989731497717
	pesos_i(18007) := b"0000000000000000_0000000000000000_0001111000101101_0101110101100010"; -- 0.11787971153018649
	pesos_i(18008) := b"1111111111111111_1111111111111111_1111001010001011_1010111110111110"; -- -0.05255605318218622
	pesos_i(18009) := b"0000000000000000_0000000000000000_0000011101011101_1011000001110111"; -- 0.02877333552588307
	pesos_i(18010) := b"0000000000000000_0000000000000000_0010001101101010_1001001110011011"; -- 0.1383449795375672
	pesos_i(18011) := b"1111111111111111_1111111111111111_1111110001111001_1000010100010110"; -- -0.013770753951513816
	pesos_i(18012) := b"0000000000000000_0000000000000000_0001101001100010_0001011110110011"; -- 0.10305927400585639
	pesos_i(18013) := b"0000000000000000_0000000000000000_0001011100011100_0111010110100100"; -- 0.0902780080272212
	pesos_i(18014) := b"1111111111111111_1111111111111111_1111101001001000_1011010111010001"; -- -0.022328029998601742
	pesos_i(18015) := b"0000000000000000_0000000000000000_0000000001001011_1011001011101010"; -- 0.0011550733060973527
	pesos_i(18016) := b"0000000000000000_0000000000000000_0001000111101010_0000101100111010"; -- 0.06997747589168925
	pesos_i(18017) := b"0000000000000000_0000000000000000_0001000101010000_1011100011000101"; -- 0.06763796634646109
	pesos_i(18018) := b"1111111111111111_1111111111111111_1111001111101100_1011110011010110"; -- -0.04716892035208508
	pesos_i(18019) := b"0000000000000000_0000000000000000_0010000110111100_0010110010011010"; -- 0.13177756075554714
	pesos_i(18020) := b"0000000000000000_0000000000000000_0001010110110101_0111011100001001"; -- 0.0848001859069309
	pesos_i(18021) := b"1111111111111111_1111111111111111_1111010101010001_0000100011001001"; -- -0.04173226437670573
	pesos_i(18022) := b"0000000000000000_0000000000000000_0000011001011000_1110100010101000"; -- 0.0247941408542457
	pesos_i(18023) := b"0000000000000000_0000000000000000_0010001100000101_1101010110111000"; -- 0.13680778247584788
	pesos_i(18024) := b"0000000000000000_0000000000000000_0001001111111110_1011010101100001"; -- 0.07810529348267256
	pesos_i(18025) := b"1111111111111111_1111111111111111_1111110000100000_1000110110111000"; -- -0.0151282717197054
	pesos_i(18026) := b"0000000000000000_0000000000000000_0000010100011101_1100110101010111"; -- 0.019985994149243305
	pesos_i(18027) := b"1111111111111111_1111111111111111_1111100111011011_1111011011100100"; -- -0.023987359400668273
	pesos_i(18028) := b"0000000000000000_0000000000000000_0000101110010110_0101110000111001"; -- 0.04526306534855083
	pesos_i(18029) := b"1111111111111111_1111111111111111_1111110100000101_0000111010101101"; -- -0.011641581388887228
	pesos_i(18030) := b"1111111111111111_1111111111111111_1111111010101000_1000011001001001"; -- -0.005241019492859704
	pesos_i(18031) := b"1111111111111111_1111111111111111_1111101011101110_0001100010110111"; -- -0.019804434973900945
	pesos_i(18032) := b"1111111111111111_1111111111111111_1111010110111011_1000011001111100"; -- -0.040107340640582474
	pesos_i(18033) := b"1111111111111111_1111111111111111_1111100001100000_0000110010000101"; -- -0.029784409999585305
	pesos_i(18034) := b"1111111111111111_1111111111111111_1111101110101101_0110101110111111"; -- -0.016885057379024463
	pesos_i(18035) := b"0000000000000000_0000000000000000_0001001001100100_0100110011000110"; -- 0.07184295499344491
	pesos_i(18036) := b"1111111111111111_1111111111111111_1101110101111101_0010101011000001"; -- -0.13480885296670925
	pesos_i(18037) := b"1111111111111111_1111111111111111_1110110011100101_1101010000111001"; -- -0.07461808782174517
	pesos_i(18038) := b"1111111111111111_1111111111111111_1110100010100011_0100101010101010"; -- -0.09125836711407039
	pesos_i(18039) := b"1111111111111111_1111111111111111_1111110011000110_1101101010111000"; -- -0.012590723024604731
	pesos_i(18040) := b"0000000000000000_0000000000000000_0000001100100100_1000110101101001"; -- 0.012276495102845402
	pesos_i(18041) := b"0000000000000000_0000000000000000_0000110100110010_1110100110001011"; -- 0.05155810959193252
	pesos_i(18042) := b"1111111111111111_1111111111111111_1110011111110111_1111110010110110"; -- -0.09387226639280863
	pesos_i(18043) := b"1111111111111111_1111111111111111_1110101100110010_0011011100101111"; -- -0.08126502124369392
	pesos_i(18044) := b"0000000000000000_0000000000000000_0000101001010001_1101111001100010"; -- 0.04031171693355565
	pesos_i(18045) := b"1111111111111111_1111111111111111_1111110001010110_1101011000110101"; -- -0.014299976297245715
	pesos_i(18046) := b"1111111111111111_1111111111111111_1101111010111110_0100011110111110"; -- -0.12990905392300073
	pesos_i(18047) := b"0000000000000000_0000000000000000_0001100010110001_0001111000100011"; -- 0.09645260198532227
	pesos_i(18048) := b"1111111111111111_1111111111111111_1110010111001010_0010011001110001"; -- -0.10238418341028371
	pesos_i(18049) := b"1111111111111111_1111111111111111_1111111010001010_0110010011001001"; -- -0.0057007798598298215
	pesos_i(18050) := b"0000000000000000_0000000000000000_0000010001011110_0110010101011011"; -- 0.017065367540537096
	pesos_i(18051) := b"0000000000000000_0000000000000000_0010011001100111_0110011000010011"; -- 0.15001523925473398
	pesos_i(18052) := b"0000000000000000_0000000000000000_0001110011110000_1001000000010010"; -- 0.11304569667702721
	pesos_i(18053) := b"1111111111111111_1111111111111111_1101101101101000_1101000011100001"; -- -0.14293188567583603
	pesos_i(18054) := b"1111111111111111_1111111111111111_1111111000111100_1010111000111111"; -- -0.006886586697932543
	pesos_i(18055) := b"0000000000000000_0000000000000000_0000011111011010_0111011111100100"; -- 0.03067731206269491
	pesos_i(18056) := b"1111111111111111_1111111111111111_1110111100010110_0001100110111110"; -- -0.06606902230379243
	pesos_i(18057) := b"0000000000000000_0000000000000000_0010010011101010_0000110011111100"; -- 0.14419633067902446
	pesos_i(18058) := b"0000000000000000_0000000000000000_0001000010001101_0010001101011000"; -- 0.06465359594717808
	pesos_i(18059) := b"1111111111111111_1111111111111111_1110100010101100_0011111100001011"; -- -0.0911217307367576
	pesos_i(18060) := b"1111111111111111_1111111111111111_1111001110000001_0011101111011010"; -- -0.0488092987648952
	pesos_i(18061) := b"1111111111111111_1111111111111111_1110000111011010_0011111100000010"; -- -0.11776357847355072
	pesos_i(18062) := b"1111111111111111_1111111111111111_1101111001001101_0000100010000011"; -- -0.13163706590994326
	pesos_i(18063) := b"0000000000000000_0000000000000000_0001000011010000_0100100110011101"; -- 0.06567821581161778
	pesos_i(18064) := b"0000000000000000_0000000000000000_0000100001001000_0000110000010110"; -- 0.03234935313530576
	pesos_i(18065) := b"1111111111111111_1111111111111111_1110001010111001_0110001100111100"; -- -0.11435870912364073
	pesos_i(18066) := b"0000000000000000_0000000000000000_0010010001011110_1111010100100001"; -- 0.142073936886769
	pesos_i(18067) := b"1111111111111111_1111111111111111_1111000001110110_1011000000101010"; -- -0.06068896269743044
	pesos_i(18068) := b"0000000000000000_0000000000000000_0000100110111101_0111011110011000"; -- 0.038047289471677265
	pesos_i(18069) := b"0000000000000000_0000000000000000_0001100011010111_0001110001000011"; -- 0.09703232417432008
	pesos_i(18070) := b"0000000000000000_0000000000000000_0001000100000010_1000111001011010"; -- 0.06644525248282038
	pesos_i(18071) := b"1111111111111111_1111111111111111_1101110001111111_0001100011010100"; -- -0.13868565392459334
	pesos_i(18072) := b"0000000000000000_0000000000000000_0010010001110001_1110101100011011"; -- 0.14236325661147137
	pesos_i(18073) := b"0000000000000000_0000000000000000_0001100011100101_0000110010011111"; -- 0.09724501506753215
	pesos_i(18074) := b"1111111111111111_1111111111111111_1111101111100101_1100000000010000"; -- -0.016025539463464328
	pesos_i(18075) := b"1111111111111111_1111111111111111_1111100110011101_0101101110101000"; -- -0.02494265688810841
	pesos_i(18076) := b"0000000000000000_0000000000000000_0001110110111101_1001000010110110"; -- 0.11617378650590555
	pesos_i(18077) := b"0000000000000000_0000000000000000_0001110101001110_0011011001110001"; -- 0.11447468044767138
	pesos_i(18078) := b"1111111111111111_1111111111111111_1111000101110111_0111000111001000"; -- -0.056771172220772936
	pesos_i(18079) := b"0000000000000000_0000000000000000_0001001101110010_0101100110110110"; -- 0.07596359909078991
	pesos_i(18080) := b"1111111111111111_1111111111111111_1110011010001011_1100100101001010"; -- -0.0994295304995959
	pesos_i(18081) := b"1111111111111111_1111111111111111_1110100011000011_1100011100100100"; -- -0.09076266643854755
	pesos_i(18082) := b"1111111111111111_1111111111111111_1111001000111000_0101100011111111"; -- -0.05382770332335289
	pesos_i(18083) := b"1111111111111111_1111111111111111_1111001110010000_1010111010001001"; -- -0.04857358131334488
	pesos_i(18084) := b"0000000000000000_0000000000000000_0010010011001110_0110100000010010"; -- 0.1437745136548478
	pesos_i(18085) := b"1111111111111111_1111111111111111_1101101101010100_0110001001000000"; -- -0.14324365546212955
	pesos_i(18086) := b"1111111111111111_1111111111111111_1110110001001101_0011110010000110"; -- -0.07694646583861678
	pesos_i(18087) := b"0000000000000000_0000000000000000_0010000011001101_0101011110001110"; -- 0.12813327033032107
	pesos_i(18088) := b"0000000000000000_0000000000000000_0000110010100001_0000101001001000"; -- 0.049332277742823206
	pesos_i(18089) := b"1111111111111111_1111111111111111_1111001111001111_1111011000101011"; -- -0.04760800787652948
	pesos_i(18090) := b"1111111111111111_1111111111111111_1110100110110110_1110101010101110"; -- -0.08705266238679193
	pesos_i(18091) := b"1111111111111111_1111111111111111_1110001101101110_0001001101001110"; -- -0.11160163248006816
	pesos_i(18092) := b"1111111111111111_1111111111111111_1111010001010000_0110110001010110"; -- -0.045647839571492786
	pesos_i(18093) := b"1111111111111111_1111111111111111_1101110000100010_1101110101001100"; -- -0.14009301078046904
	pesos_i(18094) := b"0000000000000000_0000000000000000_0000011010110111_1100110010111110"; -- 0.02624206191813986
	pesos_i(18095) := b"1111111111111111_1111111111111111_1110011001010101_1110111000000111"; -- -0.10025131541974809
	pesos_i(18096) := b"0000000000000000_0000000000000000_0001110011101110_0010000000010001"; -- 0.11300850308665303
	pesos_i(18097) := b"1111111111111111_1111111111111111_1111101001000000_0111011110010101"; -- -0.02245380983924015
	pesos_i(18098) := b"1111111111111111_1111111111111111_1110110100000001_0011110111001011"; -- -0.07419980808610106
	pesos_i(18099) := b"1111111111111111_1111111111111111_1111111111111001_0000000101000100"; -- -0.00010673599290808916
	pesos_i(18100) := b"1111111111111111_1111111111111111_1110101100100001_1111111000000011"; -- -0.08151256977883059
	pesos_i(18101) := b"0000000000000000_0000000000000000_0010010110000010_0010001101010011"; -- 0.14651699798516496
	pesos_i(18102) := b"1111111111111111_1111111111111111_1111110110010010_1011100001000110"; -- -0.009479983344723815
	pesos_i(18103) := b"1111111111111111_1111111111111111_1111101011010101_0010111001110111"; -- -0.020184608523771116
	pesos_i(18104) := b"0000000000000000_0000000000000000_0000000011011010_1001101111110001"; -- 0.0033357107525606743
	pesos_i(18105) := b"1111111111111111_1111111111111111_1101100111000110_0010101110000100"; -- -0.14931991604203654
	pesos_i(18106) := b"1111111111111111_1111111111111111_1111100001000110_0101011001000110"; -- -0.030176742509412227
	pesos_i(18107) := b"0000000000000000_0000000000000000_0000101001001010_1010111001111001"; -- 0.04020204986110323
	pesos_i(18108) := b"1111111111111111_1111111111111111_1110111011010011_1110111010011000"; -- -0.06707867432684393
	pesos_i(18109) := b"1111111111111111_1111111111111111_1110011000110010_0100111011111111"; -- -0.10079485212601508
	pesos_i(18110) := b"0000000000000000_0000000000000000_0010011000110110_1010101010010101"; -- 0.14927164220031838
	pesos_i(18111) := b"0000000000000000_0000000000000000_0001111001100000_0011001101001100"; -- 0.11865540134347585
	pesos_i(18112) := b"1111111111111111_1111111111111111_1110010010101001_1011111011001111"; -- -0.106784891481733
	pesos_i(18113) := b"1111111111111111_1111111111111111_1110000011010010_0010101100010101"; -- -0.12179308640391821
	pesos_i(18114) := b"0000000000000000_0000000000000000_0001100100110011_0010100101101000"; -- 0.09843691624908887
	pesos_i(18115) := b"0000000000000000_0000000000000000_0000010101101001_0110101001000110"; -- 0.021139757148204635
	pesos_i(18116) := b"1111111111111111_1111111111111111_1101111011100111_0110111011111100"; -- -0.1292811044390511
	pesos_i(18117) := b"0000000000000000_0000000000000000_0001000000010010_1001100001100111"; -- 0.06278374211233724
	pesos_i(18118) := b"0000000000000000_0000000000000000_0001001111101100_0101111100001001"; -- 0.07782548878903887
	pesos_i(18119) := b"1111111111111111_1111111111111111_1101100110101110_0110011011111101"; -- -0.1496825821601168
	pesos_i(18120) := b"0000000000000000_0000000000000000_0000100001111100_0111110010101101"; -- 0.033149521080551934
	pesos_i(18121) := b"1111111111111111_1111111111111111_1110110101101110_1110101111101011"; -- -0.07252622150991009
	pesos_i(18122) := b"0000000000000000_0000000000000000_0010000111010110_1100111111001110"; -- 0.13218401705552146
	pesos_i(18123) := b"0000000000000000_0000000000000000_0000100011001111_0100110000000010"; -- 0.034413099745776735
	pesos_i(18124) := b"0000000000000000_0000000000000000_0001101000000111_0101000010011010"; -- 0.10167411568240337
	pesos_i(18125) := b"0000000000000000_0000000000000000_0010001010001010_1001000111101100"; -- 0.13492691062403955
	pesos_i(18126) := b"1111111111111111_1111111111111111_1110011010110101_0000000011111101"; -- -0.09880060029691702
	pesos_i(18127) := b"0000000000000000_0000000000000000_0001011100100010_1000100100001100"; -- 0.09037071743272757
	pesos_i(18128) := b"1111111111111111_1111111111111111_1110110110000011_0100000011110011"; -- -0.07221597744745525
	pesos_i(18129) := b"1111111111111111_1111111111111111_1111010110110010_0111111110000110"; -- -0.04024508446620336
	pesos_i(18130) := b"1111111111111111_1111111111111111_1110010010001110_0001000101111001"; -- -0.10720721051357714
	pesos_i(18131) := b"1111111111111111_1111111111111111_1110011010101000_0101110001011000"; -- -0.09899351936824069
	pesos_i(18132) := b"0000000000000000_0000000000000000_0001100000000101_1001111111110100"; -- 0.09383582789143959
	pesos_i(18133) := b"0000000000000000_0000000000000000_0000101110100101_1001111000000101"; -- 0.04549586894700856
	pesos_i(18134) := b"0000000000000000_0000000000000000_0001101001010101_1000101001000100"; -- 0.10286773823535865
	pesos_i(18135) := b"1111111111111111_1111111111111111_1101100001000111_0111001011100100"; -- -0.15515977786673524
	pesos_i(18136) := b"1111111111111111_1111111111111111_1111010111100011_1010101111100111"; -- -0.03949475863220829
	pesos_i(18137) := b"0000000000000000_0000000000000000_0001000110111010_0111101010011100"; -- 0.06925169292866742
	pesos_i(18138) := b"0000000000000000_0000000000000000_0000010001111001_1010010001010011"; -- 0.017481107968387682
	pesos_i(18139) := b"1111111111111111_1111111111111111_1110000110111111_0010100011111101"; -- -0.11817687817263205
	pesos_i(18140) := b"0000000000000000_0000000000000000_0001010000111010_0100001110111011"; -- 0.07901404675112884
	pesos_i(18141) := b"0000000000000000_0000000000000000_0001000010111101_0001010011011110"; -- 0.06538515490478988
	pesos_i(18142) := b"0000000000000000_0000000000000000_0010000101010111_1011110101111100"; -- 0.13024505871322675
	pesos_i(18143) := b"1111111111111111_1111111111111111_1111111110110110_1101101011110101"; -- -0.0011160995056302902
	pesos_i(18144) := b"0000000000000000_0000000000000000_0001001110001001_0101111011100100"; -- 0.07631486004280028
	pesos_i(18145) := b"0000000000000000_0000000000000000_0001000011010110_1100011111010100"; -- 0.06577729150261782
	pesos_i(18146) := b"1111111111111111_1111111111111111_1110101101011010_1110010011000101"; -- -0.08064432333252523
	pesos_i(18147) := b"0000000000000000_0000000000000000_0001001010001001_0110100111011000"; -- 0.07240926284146922
	pesos_i(18148) := b"0000000000000000_0000000000000000_0000011110001010_1010111100001111"; -- 0.029459897165992004
	pesos_i(18149) := b"1111111111111111_1111111111111111_1111101111001111_0011001101001101"; -- -0.016369622971143145
	pesos_i(18150) := b"0000000000000000_0000000000000000_0000110001101011_1100010111101111"; -- 0.04851948810027387
	pesos_i(18151) := b"0000000000000000_0000000000000000_0010000001100001_0000100010101000"; -- 0.12648061845693978
	pesos_i(18152) := b"0000000000000000_0000000000000000_0010000001111111_0111111010011110"; -- 0.12694541317561547
	pesos_i(18153) := b"0000000000000000_0000000000000000_0000100110101000_0100100000110110"; -- 0.03772403073467053
	pesos_i(18154) := b"1111111111111111_1111111111111111_1111100011110001_0101000101110001"; -- -0.027567777483158473
	pesos_i(18155) := b"1111111111111111_1111111111111111_1111000001011010_0001111001101010"; -- -0.06112489624950908
	pesos_i(18156) := b"0000000000000000_0000000000000000_0010000110001111_1100101110111101"; -- 0.13110040065117792
	pesos_i(18157) := b"1111111111111111_1111111111111111_1111100000001100_1010000110110000"; -- -0.031057257176905176
	pesos_i(18158) := b"1111111111111111_1111111111111111_1111110100111010_0110011110100110"; -- -0.01082756219523334
	pesos_i(18159) := b"0000000000000000_0000000000000000_0000111110101000_0101110001111000"; -- 0.06116273811825353
	pesos_i(18160) := b"1111111111111111_1111111111111111_1111001010001010_0101001100000100"; -- -0.0525768390912892
	pesos_i(18161) := b"0000000000000000_0000000000000000_0000110010010010_1010010010010001"; -- 0.0491125921593786
	pesos_i(18162) := b"0000000000000000_0000000000000000_0001001010010000_1100111100011100"; -- 0.07252211034492916
	pesos_i(18163) := b"1111111111111111_1111111111111111_1110010111001000_1110100110100100"; -- -0.10240306613286901
	pesos_i(18164) := b"0000000000000000_0000000000000000_0001001100111110_0000000110111010"; -- 0.0751648979002172
	pesos_i(18165) := b"0000000000000000_0000000000000000_0000011100101111_0011111101000101"; -- 0.028064684353283076
	pesos_i(18166) := b"1111111111111111_1111111111111111_1110110010110010_0110000110011111"; -- -0.07540311682771497
	pesos_i(18167) := b"0000000000000000_0000000000000000_0000011010111101_1010010010001010"; -- 0.02633121831835473
	pesos_i(18168) := b"1111111111111111_1111111111111111_1111110000111101_0010110111010011"; -- -0.014691482627384057
	pesos_i(18169) := b"0000000000000000_0000000000000000_0000010001000001_1110101000001001"; -- 0.016630770841088497
	pesos_i(18170) := b"0000000000000000_0000000000000000_0000010010110100_0010100001111110"; -- 0.01837399566220975
	pesos_i(18171) := b"0000000000000000_0000000000000000_0000111110001101_1011101101110000"; -- 0.060756411435765156
	pesos_i(18172) := b"0000000000000000_0000000000000000_0000100110101111_1000011111000100"; -- 0.03783463043956056
	pesos_i(18173) := b"1111111111111111_1111111111111111_1101100100000101_1001100100111001"; -- -0.15225832334448083
	pesos_i(18174) := b"0000000000000000_0000000000000000_0000010011011001_1100111100010110"; -- 0.01894850045513013
	pesos_i(18175) := b"1111111111111111_1111111111111111_1110010001100110_0010111111000000"; -- -0.1078157573166004
	pesos_i(18176) := b"0000000000000000_0000000000000000_0001100100010111_0111010011111101"; -- 0.09801417527014404
	pesos_i(18177) := b"0000000000000000_0000000000000000_0000010110011001_1111001110110001"; -- 0.021880369817607652
	pesos_i(18178) := b"1111111111111111_1111111111111111_1110001000110000_0000001100100011"; -- -0.1164548910484826
	pesos_i(18179) := b"1111111111111111_1111111111111111_1110111010110011_0000011011001000"; -- -0.06758077250190767
	pesos_i(18180) := b"1111111111111111_1111111111111111_1101101000101001_1110100111100001"; -- -0.14779794935354934
	pesos_i(18181) := b"0000000000000000_0000000000000000_0001101000110000_1000000111000001"; -- 0.10230265571618233
	pesos_i(18182) := b"1111111111111111_1111111111111111_1110001111001001_1010111100010110"; -- -0.11020379738937515
	pesos_i(18183) := b"0000000000000000_0000000000000000_0010011111001111_1101100010111101"; -- 0.15551523793664918
	pesos_i(18184) := b"0000000000000000_0000000000000000_0001001011100000_1111000101001101"; -- 0.0737448514787681
	pesos_i(18185) := b"1111111111111111_1111111111111111_1111010011111011_1101110111100110"; -- -0.0430318177755893
	pesos_i(18186) := b"0000000000000000_0000000000000000_0001001001000011_1111100000000100"; -- 0.07134962166574815
	pesos_i(18187) := b"1111111111111111_1111111111111111_1101010111111111_1111101000000101"; -- -0.1640628564738433
	pesos_i(18188) := b"0000000000000000_0000000000000000_0001000010010110_0110111001101100"; -- 0.0647954001244557
	pesos_i(18189) := b"0000000000000000_0000000000000000_0000011100000001_1111111100011000"; -- 0.027374213584205373
	pesos_i(18190) := b"0000000000000000_0000000000000000_0001110001000011_1100111001100010"; -- 0.11040964033777854
	pesos_i(18191) := b"0000000000000000_0000000000000000_0010001001110100_0101010011110100"; -- 0.13458758308507962
	pesos_i(18192) := b"0000000000000000_0000000000000000_0001001001111011_0101111000111110"; -- 0.07219494822251235
	pesos_i(18193) := b"1111111111111111_1111111111111111_1101110000011111_0000111100010111"; -- -0.1401510781793772
	pesos_i(18194) := b"0000000000000000_0000000000000000_0001100000000011_0110111101100010"; -- 0.09380241540037977
	pesos_i(18195) := b"1111111111111111_1111111111111111_1111101001110010_1111111010010101"; -- -0.021682823804020947
	pesos_i(18196) := b"0000000000000000_0000000000000000_0000001000010110_0110011001000101"; -- 0.00815428899642154
	pesos_i(18197) := b"1111111111111111_1111111111111111_1101111100001011_0011000001100101"; -- -0.12873551876454217
	pesos_i(18198) := b"1111111111111111_1111111111111111_1111011111111001_0111001000101001"; -- -0.031350007113016276
	pesos_i(18199) := b"0000000000000000_0000000000000000_0000111000111001_1011111111001001"; -- 0.055568682225126224
	pesos_i(18200) := b"0000000000000000_0000000000000000_0010010000011101_1011101010100000"; -- 0.14107862854182865
	pesos_i(18201) := b"1111111111111111_1111111111111111_1110000111110100_1001100011011111"; -- -0.11736149360638849
	pesos_i(18202) := b"1111111111111111_1111111111111111_1101101110011110_1010101000100101"; -- -0.14211021997127934
	pesos_i(18203) := b"1111111111111111_1111111111111111_1111010101101010_0010110010110011"; -- -0.04134865398748827
	pesos_i(18204) := b"1111111111111111_1111111111111111_1111010100101001_0100101110100010"; -- -0.042338631524397395
	pesos_i(18205) := b"1111111111111111_1111111111111111_1111110001110101_0101000001101011"; -- -0.013834928416020074
	pesos_i(18206) := b"0000000000000000_0000000000000000_0001001111101011_1100001010000000"; -- 0.07781615859343201
	pesos_i(18207) := b"0000000000000000_0000000000000000_0001100000111000_1110000001111101"; -- 0.09461787278447102
	pesos_i(18208) := b"1111111111111111_1111111111111111_1101110100001110_0101001111001000"; -- -0.13650013321188384
	pesos_i(18209) := b"1111111111111111_1111111111111111_1110011101101111_1101000111001111"; -- -0.09595001887156787
	pesos_i(18210) := b"1111111111111111_1111111111111111_1110101110110110_1110010001101000"; -- -0.07924053631252632
	pesos_i(18211) := b"0000000000000000_0000000000000000_0000010101101111_1100001010101001"; -- 0.02123657825435822
	pesos_i(18212) := b"1111111111111111_1111111111111111_1110000111101010_1011001001100000"; -- -0.1175125612776915
	pesos_i(18213) := b"1111111111111111_1111111111111111_1111000100000101_0110011110011101"; -- -0.0585112801860246
	pesos_i(18214) := b"1111111111111111_1111111111111111_1110111111100110_1000001110100011"; -- -0.06288888228207717
	pesos_i(18215) := b"0000000000000000_0000000000000000_0010001001000000_0111001000000010"; -- 0.13379585798254442
	pesos_i(18216) := b"1111111111111111_1111111111111111_1111111010001111_0111010010011000"; -- -0.005623543734863396
	pesos_i(18217) := b"0000000000000000_0000000000000000_0010011000100000_0000100011110010"; -- 0.14892631449001567
	pesos_i(18218) := b"0000000000000000_0000000000000000_0010001110100101_0110010110001111"; -- 0.1392425035325958
	pesos_i(18219) := b"1111111111111111_1111111111111111_1110101000111011_1000010010100101"; -- -0.08502932528637737
	pesos_i(18220) := b"1111111111111111_1111111111111111_1111101001010110_0101100011111110"; -- -0.022119939684917485
	pesos_i(18221) := b"0000000000000000_0000000000000000_0000101111011100_1000001011000101"; -- 0.046333478075439104
	pesos_i(18222) := b"1111111111111111_1111111111111111_1101110000010010_1110000100000111"; -- -0.1403369291944474
	pesos_i(18223) := b"0000000000000000_0000000000000000_0001110111001001_0011111111110010"; -- 0.11635207809531015
	pesos_i(18224) := b"1111111111111111_1111111111111111_1101110111011100_1110111101011011"; -- -0.13334754972808457
	pesos_i(18225) := b"1111111111111111_1111111111111111_1110010100110101_1010110001110111"; -- -0.10464975441988252
	pesos_i(18226) := b"0000000000000000_0000000000000000_0001110000000000_0101011010111001"; -- 0.10938016912856928
	pesos_i(18227) := b"0000000000000000_0000000000000000_0000101101101111_1100000110001100"; -- 0.04467401196722976
	pesos_i(18228) := b"1111111111111111_1111111111111111_1111011010011100_1010101101011011"; -- -0.03667191525613475
	pesos_i(18229) := b"0000000000000000_0000000000000000_0001010000111111_0010100010101100"; -- 0.07908872784211049
	pesos_i(18230) := b"1111111111111111_1111111111111111_1111111000111110_1001011001011001"; -- -0.006857493549281558
	pesos_i(18231) := b"0000000000000000_0000000000000000_0000100110100100_1001011110010011"; -- 0.037667725911554845
	pesos_i(18232) := b"0000000000000000_0000000000000000_0001100100101001_0110011111010000"; -- 0.09828804800439424
	pesos_i(18233) := b"0000000000000000_0000000000000000_0001110101011001_1000011010111000"; -- 0.11464731214057185
	pesos_i(18234) := b"1111111111111111_1111111111111111_1110111010100110_1110111110000101"; -- -0.06776526444186347
	pesos_i(18235) := b"1111111111111111_1111111111111111_1111000011100110_1101111010111011"; -- -0.05897720266864914
	pesos_i(18236) := b"1111111111111111_1111111111111111_1111011100101010_0000011010100110"; -- -0.03451498451600332
	pesos_i(18237) := b"0000000000000000_0000000000000000_0000010010110001_0010111101011100"; -- 0.01832862853476965
	pesos_i(18238) := b"0000000000000000_0000000000000000_0010001111010110_0100101100010011"; -- 0.13998860565216628
	pesos_i(18239) := b"0000000000000000_0000000000000000_0001101011110001_0111100101110001"; -- 0.10524710663579072
	pesos_i(18240) := b"0000000000000000_0000000000000000_0000101010111011_1111010001001100"; -- 0.041930454773945545
	pesos_i(18241) := b"0000000000000000_0000000000000000_0000111100110111_1001001000010000"; -- 0.059441689445699455
	pesos_i(18242) := b"1111111111111111_1111111111111111_1110101101001011_0111001110000100"; -- -0.08087995554694748
	pesos_i(18243) := b"1111111111111111_1111111111111111_1111010000011010_0011010001111100"; -- -0.046475143126612065
	pesos_i(18244) := b"1111111111111111_1111111111111111_1110101101101001_0001011001110110"; -- -0.0804277383161773
	pesos_i(18245) := b"0000000000000000_0000000000000000_0001100000010010_1010010110011100"; -- 0.09403452938052125
	pesos_i(18246) := b"1111111111111111_1111111111111111_1101010000010111_0011111011110100"; -- -0.1715202954793232
	pesos_i(18247) := b"1111111111111111_1111111111111111_1110000100001111_1111110011110100"; -- -0.1208497910820845
	pesos_i(18248) := b"0000000000000000_0000000000000000_0010000010011110_1110100001010001"; -- 0.12742473584031763
	pesos_i(18249) := b"0000000000000000_0000000000000000_0001010101010100_0010110011001000"; -- 0.08331565747765493
	pesos_i(18250) := b"0000000000000000_0000000000000000_0001011000011000_1011101001010111"; -- 0.08631481769852169
	pesos_i(18251) := b"1111111111111111_1111111111111111_1111001111001100_1011001001100011"; -- -0.047657824248476546
	pesos_i(18252) := b"0000000000000000_0000000000000000_0000000010101001_0010111010000111"; -- 0.0025815085647790934
	pesos_i(18253) := b"1111111111111111_1111111111111111_1110011111001101_1110011010111001"; -- -0.09451444606076435
	pesos_i(18254) := b"0000000000000000_0000000000000000_0000000001100011_1010100000100101"; -- 0.0015206423546343638
	pesos_i(18255) := b"0000000000000000_0000000000000000_0001001010110010_0110101100100100"; -- 0.07303495053163862
	pesos_i(18256) := b"1111111111111111_1111111111111111_1110000011110100_1001110010100001"; -- -0.1212675197130393
	pesos_i(18257) := b"0000000000000000_0000000000000000_0001100011011100_1100110000111011"; -- 0.09711910672665496
	pesos_i(18258) := b"0000000000000000_0000000000000000_0010000110010011_1000100110001111"; -- 0.13115749122311537
	pesos_i(18259) := b"1111111111111111_1111111111111111_1101101100111010_0100110010010111"; -- -0.14364167501861
	pesos_i(18260) := b"1111111111111111_1111111111111111_1110110101010110_1100001001011010"; -- -0.07289490996157483
	pesos_i(18261) := b"1111111111111111_1111111111111111_1111101010001101_0110111011100001"; -- -0.02127940181735158
	pesos_i(18262) := b"1111111111111111_1111111111111111_1111101101001000_1101000100111010"; -- -0.018420146330063142
	pesos_i(18263) := b"1111111111111111_1111111111111111_1111111000010011_0111101011101101"; -- -0.007515256047337616
	pesos_i(18264) := b"0000000000000000_0000000000000000_0000110011001000_1010100001101101"; -- 0.0499367968346187
	pesos_i(18265) := b"0000000000000000_0000000000000000_0000011101101100_0010001010100010"; -- 0.02899376338883894
	pesos_i(18266) := b"0000000000000000_0000000000000000_0001110110101101_1111111100100100"; -- 0.11593622807152039
	pesos_i(18267) := b"0000000000000000_0000000000000000_0001011111110110_1000000101011101"; -- 0.09360512268819209
	pesos_i(18268) := b"0000000000000000_0000000000000000_0001101110001011_0101111111011101"; -- 0.10759543567499745
	pesos_i(18269) := b"0000000000000000_0000000000000000_0000000001111001_1110110101011001"; -- 0.0018604605438476169
	pesos_i(18270) := b"1111111111111111_1111111111111111_1111100000100001_0100110001100001"; -- -0.030741907418225783
	pesos_i(18271) := b"0000000000000000_0000000000000000_0001101010000110_0111111010000101"; -- 0.10361471899958884
	pesos_i(18272) := b"1111111111111111_1111111111111111_1101110110010010_0011111000100000"; -- -0.13448726395357008
	pesos_i(18273) := b"0000000000000000_0000000000000000_0001111000110000_0000000111011001"; -- 0.11792003194398147
	pesos_i(18274) := b"1111111111111111_1111111111111111_1111110101100111_1000100111011100"; -- -0.01013887767371482
	pesos_i(18275) := b"1111111111111111_1111111111111111_1101110000110000_1111100010000011"; -- -0.1398777657052725
	pesos_i(18276) := b"0000000000000000_0000000000000000_0001110001011101_1011010010000110"; -- 0.11080482743725963
	pesos_i(18277) := b"0000000000000000_0000000000000000_0000011111110000_1111110101100101"; -- 0.03102096279570633
	pesos_i(18278) := b"1111111111111111_1111111111111111_1111000101001111_1010011110010111"; -- -0.05737831652520319
	pesos_i(18279) := b"1111111111111111_1111111111111111_1111101111110101_0010100010011110"; -- -0.015790425813149458
	pesos_i(18280) := b"1111111111111111_1111111111111111_1110101110001001_1110101110010000"; -- -0.0799267552523511
	pesos_i(18281) := b"0000000000000000_0000000000000000_0000100010000001_1101011001010001"; -- 0.03323115801046554
	pesos_i(18282) := b"1111111111111111_1111111111111111_1111111011011000_0010110111010010"; -- -0.004513870451990224
	pesos_i(18283) := b"0000000000000000_0000000000000000_0000110001101010_1001010101100111"; -- 0.04850133671784909
	pesos_i(18284) := b"1111111111111111_1111111111111111_1110001100100100_0011010100101000"; -- -0.11272876529692683
	pesos_i(18285) := b"0000000000000000_0000000000000000_0001000000001000_1100001010000011"; -- 0.0626336640865637
	pesos_i(18286) := b"1111111111111111_1111111111111111_1110000101110001_0001111000000010"; -- -0.11936771821531736
	pesos_i(18287) := b"0000000000000000_0000000000000000_0000011010011110_1101100011000100"; -- 0.025861308846693985
	pesos_i(18288) := b"0000000000000000_0000000000000000_0000001101100101_0010011101110111"; -- 0.013262240070174142
	pesos_i(18289) := b"0000000000000000_0000000000000000_0001100101101001_0101000111110101"; -- 0.09926330779036709
	pesos_i(18290) := b"0000000000000000_0000000000000000_0001011010100011_1111110011101011"; -- 0.08843975774313924
	pesos_i(18291) := b"1111111111111111_1111111111111111_1111001001010001_0111111001011111"; -- -0.05344400572038285
	pesos_i(18292) := b"0000000000000000_0000000000000000_0010011100001011_1011010110011110"; -- 0.15252242184118606
	pesos_i(18293) := b"0000000000000000_0000000000000000_0001110101101101_1111010011111100"; -- 0.11495906013220461
	pesos_i(18294) := b"0000000000000000_0000000000000000_0000101101010111_1110101001111100"; -- 0.04431024091476005
	pesos_i(18295) := b"0000000000000000_0000000000000000_0000001101000011_1100010001010101"; -- 0.012752791096147357
	pesos_i(18296) := b"1111111111111111_1111111111111111_1111011011110101_1111011010011001"; -- -0.03530939821461026
	pesos_i(18297) := b"0000000000000000_0000000000000000_0000101100011101_0101101101000001"; -- 0.04341669411812063
	pesos_i(18298) := b"0000000000000000_0000000000000000_0001100111011110_0100100100000010"; -- 0.10104805279906509
	pesos_i(18299) := b"0000000000000000_0000000000000000_0001101011010110_0110001011111011"; -- 0.10483378054839255
	pesos_i(18300) := b"1111111111111111_1111111111111111_1111100111110011_1000010011101010"; -- -0.023627941999685424
	pesos_i(18301) := b"0000000000000000_0000000000000000_0001001110011000_0010111000110000"; -- 0.07654083886116222
	pesos_i(18302) := b"0000000000000000_0000000000000000_0010010100001000_0100000111010101"; -- 0.14465724414283052
	pesos_i(18303) := b"1111111111111111_1111111111111111_1101101011110111_0011010111011001"; -- -0.1446653695606237
	pesos_i(18304) := b"0000000000000000_0000000000000000_0000010011100000_0111000000000101"; -- 0.019049645604463265
	pesos_i(18305) := b"0000000000000000_0000000000000000_0001111110010010_0000010010010011"; -- 0.12332180584556512
	pesos_i(18306) := b"0000000000000000_0000000000000000_0001011100000001_0111101111101110"; -- 0.08986639567270888
	pesos_i(18307) := b"1111111111111111_1111111111111111_1110101110001000_1110100010110000"; -- -0.0799421853515681
	pesos_i(18308) := b"1111111111111111_1111111111111111_1110101010100100_1100110110001110"; -- -0.08342280660968401
	pesos_i(18309) := b"1111111111111111_1111111111111111_1111100110111011_0110011110011111"; -- -0.024484180167507596
	pesos_i(18310) := b"0000000000000000_0000000000000000_0001010100101101_1101011000101001"; -- 0.0827306605602374
	pesos_i(18311) := b"0000000000000000_0000000000000000_0000001011111001_0000011110001000"; -- 0.011612387466204334
	pesos_i(18312) := b"0000000000000000_0000000000000000_0001100000000100_1011100101000110"; -- 0.09382207831235718
	pesos_i(18313) := b"0000000000000000_0000000000000000_0001111010101011_0100110011001000"; -- 0.11980132944336741
	pesos_i(18314) := b"0000000000000000_0000000000000000_0000101010001111_1110010100100011"; -- 0.04125816435879317
	pesos_i(18315) := b"1111111111111111_1111111111111111_1101111101011100_0001001100000111"; -- -0.12750130727369086
	pesos_i(18316) := b"0000000000000000_0000000000000000_0000010100000000_0110001110001101"; -- 0.01953718379986885
	pesos_i(18317) := b"0000000000000000_0000000000000000_0001111001000010_1011000011110001"; -- 0.11820512659149734
	pesos_i(18318) := b"1111111111111111_1111111111111111_1110001000000001_0000011011111111"; -- -0.11717182417177822
	pesos_i(18319) := b"1111111111111111_1111111111111111_1101111110100001_0001110001110011"; -- -0.12644788931883763
	pesos_i(18320) := b"0000000000000000_0000000000000000_0010100101010101_0011111101011111"; -- 0.1614570243118146
	pesos_i(18321) := b"1111111111111111_1111111111111111_1111010110110011_1000110000100011"; -- -0.040229073877136846
	pesos_i(18322) := b"0000000000000000_0000000000000000_0000111000110111_1100000100010100"; -- 0.05553824165162162
	pesos_i(18323) := b"1111111111111111_1111111111111111_1110010100010110_0101000110110010"; -- -0.10512818730390396
	pesos_i(18324) := b"0000000000000000_0000000000000000_0001100100010001_1010010100011111"; -- 0.09792549146167655
	pesos_i(18325) := b"1111111111111111_1111111111111111_1101111100010111_0110100101100101"; -- -0.12854901580205974
	pesos_i(18326) := b"0000000000000000_0000000000000000_0001000010011000_0001110000110100"; -- 0.06482101699669068
	pesos_i(18327) := b"1111111111111111_1111111111111111_1111100101110101_1011100111011011"; -- -0.025547393924015845
	pesos_i(18328) := b"1111111111111111_1111111111111111_1111110110110100_1010001001111010"; -- -0.008962483611207505
	pesos_i(18329) := b"0000000000000000_0000000000000000_0000101111101111_1101110001111111"; -- 0.046628743212342866
	pesos_i(18330) := b"1111111111111111_1111111111111111_1110001011111110_1000100011010000"; -- -0.11330361300846357
	pesos_i(18331) := b"1111111111111111_1111111111111111_1110010011100010_1000010111111011"; -- -0.10591852775805012
	pesos_i(18332) := b"1111111111111111_1111111111111111_1110001010110000_1011101001111000"; -- -0.11449083870810958
	pesos_i(18333) := b"1111111111111111_1111111111111111_1110000010111111_0010110010110101"; -- -0.12208290646165418
	pesos_i(18334) := b"1111111111111111_1111111111111111_1110011110010000_1010100100101100"; -- -0.09544890088637972
	pesos_i(18335) := b"0000000000000000_0000000000000000_0001111001000111_1111001100111101"; -- 0.11828537212966365
	pesos_i(18336) := b"1111111111111111_1111111111111111_1111111101111100_0101001110110101"; -- -0.0020091708720706663
	pesos_i(18337) := b"0000000000000000_0000000000000000_0001010001100001_1011101001001010"; -- 0.07961620617944198
	pesos_i(18338) := b"1111111111111111_1111111111111111_1110111000010110_1101110000001001"; -- -0.0699636914413396
	pesos_i(18339) := b"1111111111111111_1111111111111111_1111100000010110_0110111100000001"; -- -0.03090769025504011
	pesos_i(18340) := b"1111111111111111_1111111111111111_1110101010100111_0100001101110000"; -- -0.08338526273669397
	pesos_i(18341) := b"0000000000000000_0000000000000000_0010100110100111_0000001001101010"; -- 0.16270461160357788
	pesos_i(18342) := b"0000000000000000_0000000000000000_0000100110101001_0001000011000101"; -- 0.03773598483282189
	pesos_i(18343) := b"1111111111111111_1111111111111111_1111000100111101_0001011000011101"; -- -0.05766164573459194
	pesos_i(18344) := b"1111111111111111_1111111111111111_1110010111110010_0010010010011100"; -- -0.10177394098461005
	pesos_i(18345) := b"0000000000000000_0000000000000000_0000101001101001_1001010001111110"; -- 0.04067352368765049
	pesos_i(18346) := b"1111111111111111_1111111111111111_1111101100011111_1011011011001000"; -- -0.019047332928570606
	pesos_i(18347) := b"1111111111111111_1111111111111111_1110000110110100_0101110011101000"; -- -0.11834163037388919
	pesos_i(18348) := b"0000000000000000_0000000000000000_0000101010110001_0010011100101111"; -- 0.041765641105229935
	pesos_i(18349) := b"1111111111111111_1111111111111111_1101110111111011_1001111000100011"; -- -0.13287936827035543
	pesos_i(18350) := b"1111111111111111_1111111111111111_1110010000000111_1101110010101001"; -- -0.10925503616935317
	pesos_i(18351) := b"0000000000000000_0000000000000000_0000111111001111_1110010100011110"; -- 0.061765975769677496
	pesos_i(18352) := b"0000000000000000_0000000000000000_0000100010111011_1001110011001001"; -- 0.034112738724982064
	pesos_i(18353) := b"1111111111111111_1111111111111111_1111000110111000_0101011011011111"; -- -0.055780954793654774
	pesos_i(18354) := b"0000000000000000_0000000000000000_0000001101111100_0101011100111101"; -- 0.013616039614156522
	pesos_i(18355) := b"1111111111111111_1111111111111111_1110111100111111_0110111001010111"; -- -0.06543836941675057
	pesos_i(18356) := b"1111111111111111_1111111111111111_1101111010000010_1110100101111111"; -- -0.1308149399270266
	pesos_i(18357) := b"1111111111111111_1111111111111111_1111101111101000_0001111111001011"; -- -0.015989315991325307
	pesos_i(18358) := b"1111111111111111_1111111111111111_1111110001100100_0100000110000100"; -- -0.014095216160517546
	pesos_i(18359) := b"1111111111111111_1111111111111111_1111110111110111_0101100100011111"; -- -0.007944517173667762
	pesos_i(18360) := b"0000000000000000_0000000000000000_0000110010010111_1010110000000010"; -- 0.04918932966870967
	pesos_i(18361) := b"0000000000000000_0000000000000000_0001110010010111_1111100111101000"; -- 0.1116939726404683
	pesos_i(18362) := b"0000000000000000_0000000000000000_0001001000100111_0000100100101011"; -- 0.07090813918481308
	pesos_i(18363) := b"1111111111111111_1111111111111111_1111101001000111_1110011001010100"; -- -0.022340397385616124
	pesos_i(18364) := b"1111111111111111_1111111111111111_1110101011111011_1010010001100000"; -- -0.08209774641181694
	pesos_i(18365) := b"1111111111111111_1111111111111111_1111111101010000_1101000011000100"; -- -0.0026731034497259705
	pesos_i(18366) := b"1111111111111111_1111111111111111_1110011111100111_1001011110011100"; -- -0.09412243307849531
	pesos_i(18367) := b"0000000000000000_0000000000000000_0000001001000101_1101010001110111"; -- 0.00887802041465915
	pesos_i(18368) := b"1111111111111111_1111111111111111_1111000111011111_1110111000011010"; -- -0.05517684796762688
	pesos_i(18369) := b"0000000000000000_0000000000000000_0001010110101100_0111111100011001"; -- 0.08466333734719961
	pesos_i(18370) := b"1111111111111111_1111111111111111_1111100111011000_1010011001101101"; -- -0.02403793190641062
	pesos_i(18371) := b"1111111111111111_1111111111111111_1110010001101111_0101001001100111"; -- -0.10767636296557948
	pesos_i(18372) := b"0000000000000000_0000000000000000_0001011011000100_0010011101001110"; -- 0.08893056537670842
	pesos_i(18373) := b"0000000000000000_0000000000000000_0000111111101101_0001001010100010"; -- 0.06221119372078535
	pesos_i(18374) := b"0000000000000000_0000000000000000_0010000011101111_1010101111100100"; -- 0.1286570961393055
	pesos_i(18375) := b"1111111111111111_1111111111111111_1111010101001011_0111101100001100"; -- -0.041817006597292344
	pesos_i(18376) := b"0000000000000000_0000000000000000_0010000010001110_1101110111101111"; -- 0.1271799762362115
	pesos_i(18377) := b"1111111111111111_1111111111111111_1101111011110101_1111001001000001"; -- -0.12905965719771112
	pesos_i(18378) := b"1111111111111111_1111111111111111_1111000100001000_1101000110000100"; -- -0.05845919156467102
	pesos_i(18379) := b"1111111111111111_1111111111111111_1101110000011101_1000001011110011"; -- -0.14017468989664428
	pesos_i(18380) := b"1111111111111111_1111111111111111_1110001101100011_1100111101111011"; -- -0.11175826307416555
	pesos_i(18381) := b"1111111111111111_1111111111111111_1111000111011110_0100111100001000"; -- -0.05520158825831692
	pesos_i(18382) := b"0000000000000000_0000000000000000_0010000011111111_0100111101100100"; -- 0.12889572323005052
	pesos_i(18383) := b"1111111111111111_1111111111111111_1111000000100010_1001011100001100"; -- -0.06197219815191762
	pesos_i(18384) := b"1111111111111111_1111111111111111_1101111110010000_1101100100110000"; -- -0.12669603894558884
	pesos_i(18385) := b"0000000000000000_0000000000000000_0001010100000101_0101011111101010"; -- 0.0821127841005208
	pesos_i(18386) := b"0000000000000000_0000000000000000_0001111110111000_1010010101000011"; -- 0.12391121760861956
	pesos_i(18387) := b"1111111111111111_1111111111111111_1111110100100110_1101100010101100"; -- -0.01112600136854015
	pesos_i(18388) := b"1111111111111111_1111111111111111_1111010101000001_1101100011010111"; -- -0.041964003956901995
	pesos_i(18389) := b"1111111111111111_1111111111111111_1110011111010001_1000001110100100"; -- -0.09445931670067921
	pesos_i(18390) := b"1111111111111111_1111111111111111_1110111001010101_0010000110011000"; -- -0.06901350069926458
	pesos_i(18391) := b"0000000000000000_0000000000000000_0010010111111101_1000110111010001"; -- 0.14840017644695183
	pesos_i(18392) := b"0000000000000000_0000000000000000_0000101101011111_0000001010000111"; -- 0.04441848550725874
	pesos_i(18393) := b"1111111111111111_1111111111111111_1110100010101001_1101000011000111"; -- -0.09115882050076411
	pesos_i(18394) := b"1111111111111111_1111111111111111_1101111100010011_0100111100111101"; -- -0.12861161001867594
	pesos_i(18395) := b"1111111111111111_1111111111111111_1111011010100000_0011111100011110"; -- -0.03661733171146398
	pesos_i(18396) := b"0000000000000000_0000000000000000_0001010101001001_1000110100100011"; -- 0.08315355404001781
	pesos_i(18397) := b"0000000000000000_0000000000000000_0000110011001001_1100100101010010"; -- 0.04995401623752335
	pesos_i(18398) := b"1111111111111111_1111111111111111_1111110111101010_1010010111001111"; -- -0.008138310361948665
	pesos_i(18399) := b"0000000000000000_0000000000000000_0000100101101000_0011011010110111"; -- 0.036746425296868016
	pesos_i(18400) := b"0000000000000000_0000000000000000_0000010000001001_1011010110110001"; -- 0.015773158744747398
	pesos_i(18401) := b"1111111111111111_1111111111111111_1101011011001110_0011100000101100"; -- -0.16091584131108527
	pesos_i(18402) := b"0000000000000000_0000000000000000_0000110010000010_0001100001100011"; -- 0.04886009607822663
	pesos_i(18403) := b"0000000000000000_0000000000000000_0000010110001001_0001110010001001"; -- 0.021623404814823062
	pesos_i(18404) := b"1111111111111111_1111111111111111_1110101010100110_0001010001010100"; -- -0.083403329349256
	pesos_i(18405) := b"1111111111111111_1111111111111111_1110011000111101_0011001010011010"; -- -0.10062869773716306
	pesos_i(18406) := b"0000000000000000_0000000000000000_0000101110100010_0111101111110110"; -- 0.04544806254515859
	pesos_i(18407) := b"1111111111111111_1111111111111111_1110010100001111_0010111001011011"; -- -0.10523710510044015
	pesos_i(18408) := b"1111111111111111_1111111111111111_1111100110101110_0110100100010010"; -- -0.02468245800861059
	pesos_i(18409) := b"1111111111111111_1111111111111111_1111101111001110_0100100011110101"; -- -0.016383590836960785
	pesos_i(18410) := b"0000000000000000_0000000000000000_0010000011101011_1101001010110100"; -- 0.12859837420118905
	pesos_i(18411) := b"1111111111111111_1111111111111111_1101010010001110_0011010100110001"; -- -0.16970508147889496
	pesos_i(18412) := b"1111111111111111_1111111111111111_1110100001101001_0100001110001000"; -- -0.09214380196257738
	pesos_i(18413) := b"0000000000000000_0000000000000000_0000100011010100_1001100011100110"; -- 0.03449397675644659
	pesos_i(18414) := b"1111111111111111_1111111111111111_1110011000101000_1011010110010010"; -- -0.10094132596468906
	pesos_i(18415) := b"0000000000000000_0000000000000000_0000010000111001_0111010001011111"; -- 0.016501687218165993
	pesos_i(18416) := b"0000000000000000_0000000000000000_0000110100101001_1011011111101111"; -- 0.05141782354400311
	pesos_i(18417) := b"0000000000000000_0000000000000000_0001001111110101_1011001001110101"; -- 0.077967790183229
	pesos_i(18418) := b"0000000000000000_0000000000000000_0001111110100101_1001000001100000"; -- 0.12362005561824777
	pesos_i(18419) := b"0000000000000000_0000000000000000_0010010110010000_0110100110010111"; -- 0.14673480930834293
	pesos_i(18420) := b"1111111111111111_1111111111111111_1111000001001101_1100010111111011"; -- -0.061313272671884515
	pesos_i(18421) := b"1111111111111111_1111111111111111_1111011000110001_0101001111110101"; -- -0.03830981500787464
	pesos_i(18422) := b"0000000000000000_0000000000000000_0000011000000110_1011101110001110"; -- 0.0235402318192165
	pesos_i(18423) := b"0000000000000000_0000000000000000_0001010101110110_1001000011011001"; -- 0.08384042070721288
	pesos_i(18424) := b"1111111111111111_1111111111111111_1111110110001001_1101001001001001"; -- -0.009615761945877294
	pesos_i(18425) := b"1111111111111111_1111111111111111_1110010100111001_0100011010000111"; -- -0.10459479530968255
	pesos_i(18426) := b"1111111111111111_1111111111111111_1111010010101010_1011100000001010"; -- -0.044270036363375904
	pesos_i(18427) := b"1111111111111111_1111111111111111_1111010101100001_0010111111000010"; -- -0.041485800946510186
	pesos_i(18428) := b"0000000000000000_0000000000000000_0000001011111111_1001001000001100"; -- 0.01171219632310492
	pesos_i(18429) := b"1111111111111111_1111111111111111_1111010100100111_1101110010101100"; -- -0.04236050404897659
	pesos_i(18430) := b"1111111111111111_1111111111111111_1111010000001110_1001011100000000"; -- -0.04665237665161222
	pesos_i(18431) := b"1111111111111111_1111111111111111_1111110100101110_0110001010101011"; -- -0.011010964590726115
	pesos_i(18432) := b"0000000000000000_0000000000000000_0001001111110110_0101100100010100"; -- 0.07797772151448328
	pesos_i(18433) := b"1111111111111111_1111111111111111_1111010111100101_0101000011010001"; -- -0.03946967018122351
	pesos_i(18434) := b"1111111111111111_1111111111111111_1111101010001111_0111010101001011"; -- -0.021248501889042058
	pesos_i(18435) := b"1111111111111111_1111111111111111_1110100110110111_0000101000110100"; -- -0.08705078353210821
	pesos_i(18436) := b"1111111111111111_1111111111111111_1111101010101010_0010111111100000"; -- -0.020840652231419066
	pesos_i(18437) := b"1111111111111111_1111111111111111_1110101011110100_1011100101010000"; -- -0.08220331003515689
	pesos_i(18438) := b"0000000000000000_0000000000000000_0001100111011100_0101111010010000"; -- 0.10101881995902814
	pesos_i(18439) := b"0000000000000000_0000000000000000_0000000000010111_0111111010000010"; -- 0.00035849265549935447
	pesos_i(18440) := b"0000000000000000_0000000000000000_0001111110000001_0100001011001100"; -- 0.12306611517498126
	pesos_i(18441) := b"0000000000000000_0000000000000000_0000111101011011_1011010101010110"; -- 0.059993108175162645
	pesos_i(18442) := b"0000000000000000_0000000000000000_0001101100010101_1111100100100101"; -- 0.10580403462531177
	pesos_i(18443) := b"0000000000000000_0000000000000000_0000000111000001_1101010101011001"; -- 0.006863912896232562
	pesos_i(18444) := b"1111111111111111_1111111111111111_1111000111000011_1001100011010100"; -- -0.055609176925500776
	pesos_i(18445) := b"1111111111111111_1111111111111111_1111111111010000_1000100110001010"; -- -0.000724223857460522
	pesos_i(18446) := b"1111111111111111_1111111111111111_1110110101010101_0011111111110111"; -- -0.07291794041547313
	pesos_i(18447) := b"0000000000000000_0000000000000000_0000100010011000_0110111111110010"; -- 0.033576008304046036
	pesos_i(18448) := b"0000000000000000_0000000000000000_0001111101000100_0000101100101111"; -- 0.12213201426745664
	pesos_i(18449) := b"0000000000000000_0000000000000000_0000011011101011_0001000101100001"; -- 0.027024351359040105
	pesos_i(18450) := b"0000000000000000_0000000000000000_0000010110011111_1111011001101100"; -- 0.02197208542353665
	pesos_i(18451) := b"0000000000000000_0000000000000000_0001101101101000_1010000000111110"; -- 0.10706521527541132
	pesos_i(18452) := b"0000000000000000_0000000000000000_0010000011101110_1111111110011010"; -- 0.12864682689338888
	pesos_i(18453) := b"1111111111111111_1111111111111111_1110000100000111_0110110010000011"; -- -0.12098047075795247
	pesos_i(18454) := b"1111111111111111_1111111111111111_1111000010110111_1010110010010110"; -- -0.05969735475294608
	pesos_i(18455) := b"1111111111111111_1111111111111111_1111000001001110_1000111110100000"; -- -0.061301253688339115
	pesos_i(18456) := b"0000000000000000_0000000000000000_0001111000001111_0111010001000000"; -- 0.11742331089339245
	pesos_i(18457) := b"1111111111111111_1111111111111111_1110001110100011_0111101001010001"; -- -0.1107867766550509
	pesos_i(18458) := b"1111111111111111_1111111111111111_1110000001100100_0001111001000001"; -- -0.1234723178720614
	pesos_i(18459) := b"0000000000000000_0000000000000000_0001110010001111_0000110100110110"; -- 0.11155779421877501
	pesos_i(18460) := b"0000000000000000_0000000000000000_0000000111100101_0011111100111001"; -- 0.00740428097538149
	pesos_i(18461) := b"1111111111111111_1111111111111111_1111011100001100_1000100010100000"; -- -0.03496500103769617
	pesos_i(18462) := b"0000000000000000_0000000000000000_0001101100011010_1110000011111001"; -- 0.10587888784536593
	pesos_i(18463) := b"1111111111111111_1111111111111111_1101101010010010_1101100110110001"; -- -0.1461967414016742
	pesos_i(18464) := b"0000000000000000_0000000000000000_0001101000100101_0000000101111010"; -- 0.10212716318753692
	pesos_i(18465) := b"1111111111111111_1111111111111111_1111000010010001_0000101110100110"; -- -0.060286781258554606
	pesos_i(18466) := b"1111111111111111_1111111111111111_1110100011011111_1100001011100010"; -- -0.09033567409640851
	pesos_i(18467) := b"1111111111111111_1111111111111111_1110101100111111_0000111001100010"; -- -0.08106908898366742
	pesos_i(18468) := b"0000000000000000_0000000000000000_0001011000110111_1000010111001011"; -- 0.08678470815348828
	pesos_i(18469) := b"0000000000000000_0000000000000000_0001101000000100_1001000110110111"; -- 0.1016322204228017
	pesos_i(18470) := b"0000000000000000_0000000000000000_0000011100001101_0010001000011001"; -- 0.027544146636574725
	pesos_i(18471) := b"1111111111111111_1111111111111111_1101111111011000_0100010010110001"; -- -0.1256062572928375
	pesos_i(18472) := b"0000000000000000_0000000000000000_0001110110011101_0111001111110100"; -- 0.1156837911617066
	pesos_i(18473) := b"0000000000000000_0000000000000000_0001010011100100_0100101110110110"; -- 0.08160851673465812
	pesos_i(18474) := b"0000000000000000_0000000000000000_0000101011000000_0100110001001001"; -- 0.04199673453279961
	pesos_i(18475) := b"0000000000000000_0000000000000000_0001111011010110_1001110000011101"; -- 0.12046218587372053
	pesos_i(18476) := b"1111111111111111_1111111111111111_1111000100011111_1001000110000101"; -- -0.058112053814081376
	pesos_i(18477) := b"0000000000000000_0000000000000000_0000101110110101_1010111011011011"; -- 0.045741013124291824
	pesos_i(18478) := b"1111111111111111_1111111111111111_1101100000111000_1110011111001000"; -- -0.1553816925996185
	pesos_i(18479) := b"0000000000000000_0000000000000000_0000010111010100_1000001110011001"; -- 0.02277395717052237
	pesos_i(18480) := b"0000000000000000_0000000000000000_0000111011101000_0111100010000110"; -- 0.058234722820508567
	pesos_i(18481) := b"1111111111111111_1111111111111111_1110010001100110_0001100010011111"; -- -0.10781713601320737
	pesos_i(18482) := b"0000000000000000_0000000000000000_0010001101101000_1000100001000101"; -- 0.1383137863585042
	pesos_i(18483) := b"0000000000000000_0000000000000000_0010001001010000_1000001011100011"; -- 0.13404100457070303
	pesos_i(18484) := b"0000000000000000_0000000000000000_0001100111000011_1101111000010010"; -- 0.10064495021439006
	pesos_i(18485) := b"0000000000000000_0000000000000000_0000110111110110_0101011110100010"; -- 0.05454013540425698
	pesos_i(18486) := b"0000000000000000_0000000000000000_0010001000011101_1011111100110111"; -- 0.13326640207387191
	pesos_i(18487) := b"1111111111111111_1111111111111111_1101111100000001_1011001001111100"; -- -0.12888035264080192
	pesos_i(18488) := b"1111111111111111_1111111111111111_1101101000110100_0110010010100100"; -- -0.14763804434420888
	pesos_i(18489) := b"0000000000000000_0000000000000000_0000000001001101_1011011010000010"; -- 0.0011858051035871767
	pesos_i(18490) := b"0000000000000000_0000000000000000_0000100111001000_1100000011111011"; -- 0.038219510322456185
	pesos_i(18491) := b"0000000000000000_0000000000000000_0001000000101111_1011110111110111"; -- 0.0632284859125213
	pesos_i(18492) := b"1111111111111111_1111111111111111_1111011111100100_0001100000001111"; -- -0.03167581205903844
	pesos_i(18493) := b"1111111111111111_1111111111111111_1111010011011110_0111000111011000"; -- -0.04348076317557338
	pesos_i(18494) := b"0000000000000000_0000000000000000_0000111110000001_1110100001111100"; -- 0.060575990880849466
	pesos_i(18495) := b"0000000000000000_0000000000000000_0000001011001011_0110100010111101"; -- 0.010916277066759725
	pesos_i(18496) := b"0000000000000000_0000000000000000_0010010110011110_1001100110111011"; -- 0.14695130179985474
	pesos_i(18497) := b"1111111111111111_1111111111111111_1111100000000011_1011110001011110"; -- -0.031192996114432624
	pesos_i(18498) := b"0000000000000000_0000000000000000_0001110000101101_0100110000100010"; -- 0.11006618333683336
	pesos_i(18499) := b"1111111111111111_1111111111111111_1110110011011001_0010111010010110"; -- -0.0748110659245411
	pesos_i(18500) := b"1111111111111111_1111111111111111_1101110100100011_0101111011110011"; -- -0.13617903292951986
	pesos_i(18501) := b"1111111111111111_1111111111111111_1111010001001011_1000110010111101"; -- -0.04572220226299013
	pesos_i(18502) := b"0000000000000000_0000000000000000_0000100111010100_0011100001001001"; -- 0.03839446807578312
	pesos_i(18503) := b"1111111111111111_1111111111111111_1111100100111010_1101010000101111"; -- -0.02644609311860555
	pesos_i(18504) := b"0000000000000000_0000000000000000_0000101110001100_0010110011000110"; -- 0.04510764914502127
	pesos_i(18505) := b"0000000000000000_0000000000000000_0000110100100001_1100111010010011"; -- 0.051297102785178295
	pesos_i(18506) := b"0000000000000000_0000000000000000_0000110011100011_0101011000101100"; -- 0.050343881460444696
	pesos_i(18507) := b"1111111111111111_1111111111111111_1111111010111101_0010100010101000"; -- -0.00492616553186024
	pesos_i(18508) := b"1111111111111111_1111111111111111_1110000000011110_0001111011110001"; -- -0.12454039211045591
	pesos_i(18509) := b"0000000000000000_0000000000000000_0000000100111001_0101111000100001"; -- 0.004781611425017751
	pesos_i(18510) := b"1111111111111111_1111111111111111_1110000010001101_0011000100110111"; -- -0.12284557734342266
	pesos_i(18511) := b"1111111111111111_1111111111111111_1110001000011010_0011010000110010"; -- -0.11678766043271131
	pesos_i(18512) := b"0000000000000000_0000000000000000_0000100011001010_0000001010000111"; -- 0.03433242593473512
	pesos_i(18513) := b"1111111111111111_1111111111111111_1111111011111100_0111010001110000"; -- -0.003960344930155835
	pesos_i(18514) := b"0000000000000000_0000000000000000_0001101100011101_1011000011101011"; -- 0.10592180007005185
	pesos_i(18515) := b"1111111111111111_1111111111111111_1110100011001000_1100001010101011"; -- -0.09068663902237953
	pesos_i(18516) := b"1111111111111111_1111111111111111_1111111000110010_0011111101010111"; -- -0.00704578511774993
	pesos_i(18517) := b"1111111111111111_1111111111111111_1110100010011000_1010000011001000"; -- -0.09142108068165225
	pesos_i(18518) := b"1111111111111111_1111111111111111_1101110100101110_1101010101000110"; -- -0.13600413365439018
	pesos_i(18519) := b"1111111111111111_1111111111111111_1110010000001010_1101110000111011"; -- -0.10920928524719312
	pesos_i(18520) := b"0000000000000000_0000000000000000_0001111110110111_1101101100101001"; -- 0.12389917129950073
	pesos_i(18521) := b"1111111111111111_1111111111111111_1111110100100011_0110111000100100"; -- -0.011178127603181546
	pesos_i(18522) := b"1111111111111111_1111111111111111_1101110010000011_1100110010010010"; -- -0.13861390536840734
	pesos_i(18523) := b"1111111111111111_1111111111111111_1101111101111101_1000110100001111"; -- -0.12699049366173232
	pesos_i(18524) := b"0000000000000000_0000000000000000_0000000011100101_1110010111101001"; -- 0.003507966424547322
	pesos_i(18525) := b"1111111111111111_1111111111111111_1110110100111011_0100011101000101"; -- -0.0733142333690878
	pesos_i(18526) := b"0000000000000000_0000000000000000_0001110011000000_0101000101110011"; -- 0.11230954219860838
	pesos_i(18527) := b"1111111111111111_1111111111111111_1110110100101110_0111011000000001"; -- -0.07350981203911143
	pesos_i(18528) := b"1111111111111111_1111111111111111_1110100110011100_0010011000110100"; -- -0.08746110173900175
	pesos_i(18529) := b"1111111111111111_1111111111111111_1111111011111011_0001101010001111"; -- -0.0039809608438244135
	pesos_i(18530) := b"0000000000000000_0000000000000000_0001000101011011_0011101001010010"; -- 0.06779827603068278
	pesos_i(18531) := b"1111111111111111_1111111111111111_1101100111010001_1111100101011110"; -- -0.14913979961624935
	pesos_i(18532) := b"0000000000000000_0000000000000000_0010001111101101_0111101011001101"; -- 0.1403424024519621
	pesos_i(18533) := b"1111111111111111_1111111111111111_1110100001010100_0111101010100111"; -- -0.09246095114934647
	pesos_i(18534) := b"0000000000000000_0000000000000000_0000011110111100_0001100000000100"; -- 0.030213833685365336
	pesos_i(18535) := b"1111111111111111_1111111111111111_1110100100001001_1010010100000111"; -- -0.08969658441566468
	pesos_i(18536) := b"1111111111111111_1111111111111111_1110001001001101_0000110010100010"; -- -0.11601182033811178
	pesos_i(18537) := b"0000000000000000_0000000000000000_0010000001111110_1000101110110101"; -- 0.12693093472504535
	pesos_i(18538) := b"1111111111111111_1111111111111111_1111010101001011_0111100001011011"; -- -0.04181716712049286
	pesos_i(18539) := b"0000000000000000_0000000000000000_0001101010011010_0010011001001001"; -- 0.10391463544151594
	pesos_i(18540) := b"0000000000000000_0000000000000000_0000010110010001_1001100001110000"; -- 0.021752860396945062
	pesos_i(18541) := b"0000000000000000_0000000000000000_0000011011101101_1000010010110011"; -- 0.027061742466045143
	pesos_i(18542) := b"1111111111111111_1111111111111111_1101101011110110_0111011001111100"; -- -0.14467677555543365
	pesos_i(18543) := b"1111111111111111_1111111111111111_1111100010100110_0111101001101101"; -- -0.02870974393025477
	pesos_i(18544) := b"0000000000000000_0000000000000000_0001101100001101_0011110110010110"; -- 0.10567078507792013
	pesos_i(18545) := b"0000000000000000_0000000000000000_0000101100010100_1010111000011111"; -- 0.0432843041723346
	pesos_i(18546) := b"1111111111111111_1111111111111111_1110111111011001_0111010010001010"; -- -0.06308814655514945
	pesos_i(18547) := b"0000000000000000_0000000000000000_0001100101110010_1011111100101111"; -- 0.09940714742435638
	pesos_i(18548) := b"1111111111111111_1111111111111111_1110111000111100_1101000100001101"; -- -0.06938451216128202
	pesos_i(18549) := b"1111111111111111_1111111111111111_1110110000011001_0001101101010000"; -- -0.0777419023912544
	pesos_i(18550) := b"1111111111111111_1111111111111111_1110100011100100_1011011001001101"; -- -0.09026013004877041
	pesos_i(18551) := b"1111111111111111_1111111111111111_1110011101000110_1110100110100001"; -- -0.09657420949827099
	pesos_i(18552) := b"0000000000000000_0000000000000000_0010001101111111_0101110011101110"; -- 0.1386621553005674
	pesos_i(18553) := b"1111111111111111_1111111111111111_1101111100001011_0101011110100010"; -- -0.12873317991577143
	pesos_i(18554) := b"0000000000000000_0000000000000000_0001100100001001_1101001100011111"; -- 0.09780616290817022
	pesos_i(18555) := b"0000000000000000_0000000000000000_0010101101001011_1000101001010000"; -- 0.16912140333783346
	pesos_i(18556) := b"0000000000000000_0000000000000000_0000111001001111_1000011010111000"; -- 0.05590097427280509
	pesos_i(18557) := b"1111111111111111_1111111111111111_1110110110101000_1011100010101111"; -- -0.07164426538550157
	pesos_i(18558) := b"0000000000000000_0000000000000000_0010000000110010_0000111111100011"; -- 0.12576388632732152
	pesos_i(18559) := b"1111111111111111_1111111111111111_1110101001010111_1110110101000010"; -- -0.0845958435823061
	pesos_i(18560) := b"1111111111111111_1111111111111111_1111111011000001_1010011111010001"; -- -0.004857551091294363
	pesos_i(18561) := b"0000000000000000_0000000000000000_0010010010011101_1101111001111001"; -- 0.14303389039271402
	pesos_i(18562) := b"1111111111111111_1111111111111111_1110011011101111_0000101001001111"; -- -0.09791503505797694
	pesos_i(18563) := b"0000000000000000_0000000000000000_0001011001001001_1010101010011111"; -- 0.08706156148893221
	pesos_i(18564) := b"0000000000000000_0000000000000000_0000000000001110_1001101001010011"; -- 0.00022282146659767226
	pesos_i(18565) := b"0000000000000000_0000000000000000_0001011010111001_0101011110111111"; -- 0.08876560600246552
	pesos_i(18566) := b"0000000000000000_0000000000000000_0001110010001111_0001000110011110"; -- 0.11155805695073816
	pesos_i(18567) := b"1111111111111111_1111111111111111_1111101010101101_0011001001100000"; -- -0.020794726887678812
	pesos_i(18568) := b"1111111111111111_1111111111111111_1111000010111001_1110010110011001"; -- -0.059663438942109785
	pesos_i(18569) := b"0000000000000000_0000000000000000_0001111110001100_1110111001111100"; -- 0.12324419526853682
	pesos_i(18570) := b"0000000000000000_0000000000000000_0000111111101110_1111001000011001"; -- 0.06223977185043302
	pesos_i(18571) := b"1111111111111111_1111111111111111_1111010011011011_1110110010011010"; -- -0.043519222652048946
	pesos_i(18572) := b"0000000000000000_0000000000000000_0001111001001000_1000100011100001"; -- 0.11829429134470879
	pesos_i(18573) := b"0000000000000000_0000000000000000_0000010010111001_0000100011011011"; -- 0.01844840380219286
	pesos_i(18574) := b"0000000000000000_0000000000000000_0001111110100001_0101111100011010"; -- 0.12355608360123771
	pesos_i(18575) := b"0000000000000000_0000000000000000_0000010101101101_1010000011101111"; -- 0.02120405050184183
	pesos_i(18576) := b"1111111111111111_1111111111111111_1110111011111000_1110000000010011"; -- -0.06651496456128012
	pesos_i(18577) := b"0000000000000000_0000000000000000_0000001001010001_1111001100100001"; -- 0.009062953559829997
	pesos_i(18578) := b"1111111111111111_1111111111111111_1111101100111110_1000000101011100"; -- -0.01857749468979692
	pesos_i(18579) := b"1111111111111111_1111111111111111_1111110111010010_0101111000111011"; -- -0.008508787615855037
	pesos_i(18580) := b"1111111111111111_1111111111111111_1110100111000001_1001001110010010"; -- -0.08689000794285405
	pesos_i(18581) := b"1111111111111111_1111111111111111_1111110111110001_1001010110110111"; -- -0.008032458220078668
	pesos_i(18582) := b"0000000000000000_0000000000000000_0000011001111010_0101110100010011"; -- 0.02530461986547119
	pesos_i(18583) := b"0000000000000000_0000000000000000_0001000001101101_1001101001101011"; -- 0.06417241195063199
	pesos_i(18584) := b"1111111111111111_1111111111111111_1111100101001010_0010010111111110"; -- -0.026212335121935538
	pesos_i(18585) := b"1111111111111111_1111111111111111_1111010101000000_1000100101010100"; -- -0.04198400220902646
	pesos_i(18586) := b"0000000000000000_0000000000000000_0001010001001101_0100001101001100"; -- 0.07930393799509318
	pesos_i(18587) := b"1111111111111111_1111111111111111_1111111000100001_1011111110101111"; -- -0.007297534811177864
	pesos_i(18588) := b"0000000000000000_0000000000000000_0010100001010101_1100110011001100"; -- 0.15755920391555422
	pesos_i(18589) := b"0000000000000000_0000000000000000_0001101000101000_0001101000100011"; -- 0.10217440952843079
	pesos_i(18590) := b"0000000000000000_0000000000000000_0001110000100011_1101111001111000"; -- 0.10992231785356017
	pesos_i(18591) := b"1111111111111111_1111111111111111_1110100111110111_0111100011011010"; -- -0.0860676256914235
	pesos_i(18592) := b"0000000000000000_0000000000000000_0010001011110001_1110010011001000"; -- 0.13650350451268184
	pesos_i(18593) := b"1111111111111111_1111111111111111_1111001100001111_0110010011001100"; -- -0.05054636029884617
	pesos_i(18594) := b"0000000000000000_0000000000000000_0000100110001001_1011101101100000"; -- 0.037257872628644925
	pesos_i(18595) := b"0000000000000000_0000000000000000_0000010101000110_0010000111101000"; -- 0.02060138620325356
	pesos_i(18596) := b"0000000000000000_0000000000000000_0001011110101110_1001011010000100"; -- 0.09250775083556308
	pesos_i(18597) := b"1111111111111111_1111111111111111_1110011110011001_1011001111000001"; -- -0.09531094103313895
	pesos_i(18598) := b"0000000000000000_0000000000000000_0000001100111000_0011001101000000"; -- 0.012576296869258945
	pesos_i(18599) := b"1111111111111111_1111111111111111_1110100100001001_1110010010001000"; -- -0.08969279931520961
	pesos_i(18600) := b"1111111111111111_1111111111111111_1110011100010111_0001000111010101"; -- -0.09730423505411841
	pesos_i(18601) := b"1111111111111111_1111111111111111_1110011111010100_0110011101010110"; -- -0.09441522732622984
	pesos_i(18602) := b"1111111111111111_1111111111111111_1110001011111100_1011100010110000"; -- -0.11333127699707392
	pesos_i(18603) := b"0000000000000000_0000000000000000_0001110110001110_0111110110111101"; -- 0.11545549266971133
	pesos_i(18604) := b"0000000000000000_0000000000000000_0000011001111101_1110101011011000"; -- 0.025358846525409345
	pesos_i(18605) := b"0000000000000000_0000000000000000_0000011011110001_1001111001011010"; -- 0.027124306621341118
	pesos_i(18606) := b"0000000000000000_0000000000000000_0010001011100011_0100100000100100"; -- 0.13628054503575623
	pesos_i(18607) := b"0000000000000000_0000000000000000_0000011101100000_0100101000100000"; -- 0.028813011895344638
	pesos_i(18608) := b"1111111111111111_1111111111111111_1111111101010000_0111011010111011"; -- -0.002678469886254332
	pesos_i(18609) := b"0000000000000000_0000000000000000_0010001011001111_0011010011110011"; -- 0.13597422537965043
	pesos_i(18610) := b"1111111111111111_1111111111111111_1110011101000100_0111011100000001"; -- -0.09661155906499465
	pesos_i(18611) := b"0000000000000000_0000000000000000_0001101010110100_1010111101001001"; -- 0.10431952982670664
	pesos_i(18612) := b"0000000000000000_0000000000000000_0001101101111011_1010011101011101"; -- 0.10735555668255248
	pesos_i(18613) := b"0000000000000000_0000000000000000_0001010000011000_0110001110110110"; -- 0.07849715411803465
	pesos_i(18614) := b"1111111111111111_1111111111111111_1111111001010010_0110101110110100"; -- -0.006554859680908675
	pesos_i(18615) := b"1111111111111111_1111111111111111_1111111101101011_1011100101101010"; -- -0.002262508077438762
	pesos_i(18616) := b"1111111111111111_1111111111111111_1111010110001010_1101011100111110"; -- -0.04085020762674212
	pesos_i(18617) := b"0000000000000000_0000000000000000_0001110011010100_0111101101110111"; -- 0.11261722235413416
	pesos_i(18618) := b"0000000000000000_0000000000000000_0010001101100111_0011111101100100"; -- 0.13829418361473497
	pesos_i(18619) := b"1111111111111111_1111111111111111_1111111001100011_0001011101000001"; -- -0.00630049377227351
	pesos_i(18620) := b"0000000000000000_0000000000000000_0010000011010011_1101010101110111"; -- 0.12823232808872276
	pesos_i(18621) := b"1111111111111111_1111111111111111_1111100000010001_0000110110110100"; -- -0.030989783924639445
	pesos_i(18622) := b"1111111111111111_1111111111111111_1111100000011101_0000111100000001"; -- -0.030806600745867142
	pesos_i(18623) := b"1111111111111111_1111111111111111_1110111100000000_0001111110000010"; -- -0.0664043719379919
	pesos_i(18624) := b"0000000000000000_0000000000000000_0000001111011101_0000100010000100"; -- 0.01509144993698448
	pesos_i(18625) := b"0000000000000000_0000000000000000_0000001011110011_0010011000111000"; -- 0.011522663696668408
	pesos_i(18626) := b"0000000000000000_0000000000000000_0000110101001001_1100111001110000"; -- 0.05190744613150877
	pesos_i(18627) := b"0000000000000000_0000000000000000_0001000010101011_0100110101110101"; -- 0.06511386964741865
	pesos_i(18628) := b"1111111111111111_1111111111111111_1110100111011000_1010111010100101"; -- -0.08653744193920716
	pesos_i(18629) := b"1111111111111111_1111111111111111_1111010111011111_1101100001110110"; -- -0.03955313803178741
	pesos_i(18630) := b"0000000000000000_0000000000000000_0000101111111011_1000001100000100"; -- 0.04680651520716886
	pesos_i(18631) := b"1111111111111111_1111111111111111_1101100101100000_0101110101101110"; -- -0.15087333742773154
	pesos_i(18632) := b"1111111111111111_1111111111111111_1111100100111110_0000001011100111"; -- -0.026397532080676384
	pesos_i(18633) := b"0000000000000000_0000000000000000_0001101011100011_0001000100010110"; -- 0.10502726341181054
	pesos_i(18634) := b"1111111111111111_1111111111111111_1110111110011101_1001110000010001"; -- -0.06400131784438852
	pesos_i(18635) := b"1111111111111111_1111111111111111_1111110110001100_1000011010011000"; -- -0.009574497220130112
	pesos_i(18636) := b"1111111111111111_1111111111111111_1110011110111011_0101011000001110"; -- -0.09479772718997614
	pesos_i(18637) := b"0000000000000000_0000000000000000_0010011010101100_0110111001100000"; -- 0.15106859052824795
	pesos_i(18638) := b"0000000000000000_0000000000000000_0010001011000111_0011000110001010"; -- 0.13585195178504214
	pesos_i(18639) := b"0000000000000000_0000000000000000_0001101000000000_1110001000011011"; -- 0.10157597689744566
	pesos_i(18640) := b"1111111111111111_1111111111111111_1101101011101010_0100100011011110"; -- -0.1448626000599221
	pesos_i(18641) := b"1111111111111111_1111111111111111_1111011110101111_1111000101000111"; -- -0.0324715806362047
	pesos_i(18642) := b"1111111111111111_1111111111111111_1110101100011111_0100000000011011"; -- -0.08155440666901448
	pesos_i(18643) := b"1111111111111111_1111111111111111_1110001101011001_1001101101110001"; -- -0.11191395276638846
	pesos_i(18644) := b"0000000000000000_0000000000000000_0000110001001000_0100100000100110"; -- 0.04797793311399626
	pesos_i(18645) := b"0000000000000000_0000000000000000_0000111111110100_1100110111000101"; -- 0.062329159423163895
	pesos_i(18646) := b"1111111111111111_1111111111111111_1111110101110001_1111111110010001"; -- -0.00997927392129287
	pesos_i(18647) := b"1111111111111111_1111111111111111_1110001111110101_1001100001000100"; -- -0.10953377096394636
	pesos_i(18648) := b"1111111111111111_1111111111111111_1110111011110100_0000100110011101"; -- -0.06658878237169673
	pesos_i(18649) := b"0000000000000000_0000000000000000_0000111010000110_0100001010001101"; -- 0.056736144420617515
	pesos_i(18650) := b"1111111111111111_1111111111111111_1111001011110011_1001100011111001"; -- -0.05097049645103526
	pesos_i(18651) := b"0000000000000000_0000000000000000_0001111111101001_1000001010101001"; -- 0.12465683578792802
	pesos_i(18652) := b"1111111111111111_1111111111111111_1101100111000101_1110000010111011"; -- -0.14932437361572987
	pesos_i(18653) := b"0000000000000000_0000000000000000_0001011011101100_1100100100100000"; -- 0.08955056224642205
	pesos_i(18654) := b"0000000000000000_0000000000000000_0010000000000111_1101000110010101"; -- 0.12511930364029678
	pesos_i(18655) := b"0000000000000000_0000000000000000_0000100001000110_0101100011010111"; -- 0.03232341048732262
	pesos_i(18656) := b"0000000000000000_0000000000000000_0001110011110101_0001010110111111"; -- 0.11311469957489889
	pesos_i(18657) := b"0000000000000000_0000000000000000_0001001010111110_1001000010011110"; -- 0.07322028966667483
	pesos_i(18658) := b"0000000000000000_0000000000000000_0010000000110001_1100100010101110"; -- 0.12575964208301108
	pesos_i(18659) := b"1111111111111111_1111111111111111_1111011101001110_0011000110111011"; -- -0.033963100186652787
	pesos_i(18660) := b"0000000000000000_0000000000000000_0001000111000011_1111011000011100"; -- 0.06939638304962077
	pesos_i(18661) := b"1111111111111111_1111111111111111_1101100111011111_0111111011010000"; -- -0.14893348131852452
	pesos_i(18662) := b"0000000000000000_0000000000000000_0000011110011100_1010010010100001"; -- 0.02973393370633027
	pesos_i(18663) := b"0000000000000000_0000000000000000_0001000100011001_0111000001011101"; -- 0.06679441707560453
	pesos_i(18664) := b"1111111111111111_1111111111111111_1111100010001001_1100011101010110"; -- -0.029147664634385083
	pesos_i(18665) := b"0000000000000000_0000000000000000_0001110000111000_1110110111011001"; -- 0.11024366910336317
	pesos_i(18666) := b"0000000000000000_0000000000000000_0000111101000011_1100010100110111"; -- 0.0596278438065338
	pesos_i(18667) := b"0000000000000000_0000000000000000_0000001001010001_1001001010001100"; -- 0.009057196691221991
	pesos_i(18668) := b"1111111111111111_1111111111111111_1110001100001111_0011011101000011"; -- -0.11304907427932741
	pesos_i(18669) := b"0000000000000000_0000000000000000_0010010101001111_0110101000111111"; -- 0.14574302707594936
	pesos_i(18670) := b"1111111111111111_1111111111111111_1111110000001000_0101110001010101"; -- -0.015497426202066159
	pesos_i(18671) := b"0000000000000000_0000000000000000_0000010011001100_0101101100000111"; -- 0.01874321867703324
	pesos_i(18672) := b"0000000000000000_0000000000000000_0010000111001110_1100101011111111"; -- 0.13206166005737652
	pesos_i(18673) := b"0000000000000000_0000000000000000_0010010100101110_0000000000001010"; -- 0.1452331565732203
	pesos_i(18674) := b"1111111111111111_1111111111111111_1111011000101111_1000001010100001"; -- -0.03833755084368358
	pesos_i(18675) := b"1111111111111111_1111111111111111_1110000111011100_0111000001110101"; -- -0.11773011355228138
	pesos_i(18676) := b"1111111111111111_1111111111111111_1110101000010010_1000110111001111"; -- -0.08565438934987264
	pesos_i(18677) := b"0000000000000000_0000000000000000_0000111111000110_0111010110000100"; -- 0.06162199463163845
	pesos_i(18678) := b"0000000000000000_0000000000000000_0001011101111110_1111110100011000"; -- 0.0917814429544339
	pesos_i(18679) := b"0000000000000000_0000000000000000_0001111000010110_1000001000110110"; -- 0.11753095461250994
	pesos_i(18680) := b"0000000000000000_0000000000000000_0001100110001011_1011101011101100"; -- 0.09978836303227442
	pesos_i(18681) := b"0000000000000000_0000000000000000_0000010101111000_1110100000110100"; -- 0.021376145081115554
	pesos_i(18682) := b"0000000000000000_0000000000000000_0001110011110011_0011001100010010"; -- 0.1130859298230756
	pesos_i(18683) := b"0000000000000000_0000000000000000_0000101111110111_0101000111011110"; -- 0.0467425504504925
	pesos_i(18684) := b"0000000000000000_0000000000000000_0010000111011000_0011110000010110"; -- 0.1322057298955749
	pesos_i(18685) := b"0000000000000000_0000000000000000_0000000100100000_0011110000000000"; -- 0.004398107437912682
	pesos_i(18686) := b"0000000000000000_0000000000000000_0001100100111100_0100110100111101"; -- 0.09857638107964242
	pesos_i(18687) := b"1111111111111111_1111111111111111_1110010100101010_0111101100110011"; -- -0.1048205376701647
	pesos_i(18688) := b"1111111111111111_1111111111111111_1111110011001011_1001000010101001"; -- -0.012518843446647984
	pesos_i(18689) := b"0000000000000000_0000000000000000_0001011001011011_1101000011101101"; -- 0.08733850284126787
	pesos_i(18690) := b"1111111111111111_1111111111111111_1111000110001011_1100011010001101"; -- -0.05646094383073437
	pesos_i(18691) := b"0000000000000000_0000000000000000_0001010001001100_0111010110001001"; -- 0.07929167364439908
	pesos_i(18692) := b"0000000000000000_0000000000000000_0000101101011011_0000000000100110"; -- 0.044357308766689627
	pesos_i(18693) := b"0000000000000000_0000000000000000_0001000110000000_1001100001000001"; -- 0.06836845015464574
	pesos_i(18694) := b"0000000000000000_0000000000000000_0001001110000010_0111101101001000"; -- 0.0762097408244954
	pesos_i(18695) := b"0000000000000000_0000000000000000_0000001100111000_1101100100101111"; -- 0.012586187225575328
	pesos_i(18696) := b"1111111111111111_1111111111111111_1101101010110110_1010000011110000"; -- -0.14565080769602326
	pesos_i(18697) := b"0000000000000000_0000000000000000_0000110001100100_0100100010110001"; -- 0.048405211665243204
	pesos_i(18698) := b"0000000000000000_0000000000000000_0010010000010111_0001010000011101"; -- 0.14097715107026584
	pesos_i(18699) := b"1111111111111111_1111111111111111_1111011001001011_1111101101000000"; -- -0.03790311523685715
	pesos_i(18700) := b"0000000000000000_0000000000000000_0001111000001000_1110000101111101"; -- 0.1173230105186926
	pesos_i(18701) := b"1111111111111111_1111111111111111_1110101000010011_1001100100001011"; -- -0.08563846097629078
	pesos_i(18702) := b"0000000000000000_0000000000000000_0000000110111110_0110100111000100"; -- 0.006811724003986571
	pesos_i(18703) := b"1111111111111111_1111111111111111_1101110010000110_0000101110110000"; -- -0.1385796255845961
	pesos_i(18704) := b"0000000000000000_0000000000000000_0000111101111110_1010001001000011"; -- 0.0605260290827075
	pesos_i(18705) := b"1111111111111111_1111111111111111_1111011100000011_1110101001101000"; -- -0.03509650196647263
	pesos_i(18706) := b"0000000000000000_0000000000000000_0000010010000110_1111111011001000"; -- 0.01768486393540687
	pesos_i(18707) := b"0000000000000000_0000000000000000_0010001111101101_0001011100011100"; -- 0.14033646038443984
	pesos_i(18708) := b"1111111111111111_1111111111111111_1111110001001000_1000010100110000"; -- -0.014518428662368387
	pesos_i(18709) := b"0000000000000000_0000000000000000_0001000000111010_1010101001010010"; -- 0.0633951617441997
	pesos_i(18710) := b"0000000000000000_0000000000000000_0000100001111101_1001100010011110"; -- 0.03316644525472487
	pesos_i(18711) := b"0000000000000000_0000000000000000_0000111111101010_1001001000111111"; -- 0.06217302347243892
	pesos_i(18712) := b"1111111111111111_1111111111111111_1111110011000100_1100111011100111"; -- -0.012621944907312428
	pesos_i(18713) := b"1111111111111111_1111111111111111_1110010110000111_1110111101100111"; -- -0.10339454409415072
	pesos_i(18714) := b"0000000000000000_0000000000000000_0000011010101010_1011111010001110"; -- 0.02604285208231266
	pesos_i(18715) := b"0000000000000000_0000000000000000_0000101111011011_0011000111011000"; -- 0.046313395618414625
	pesos_i(18716) := b"1111111111111111_1111111111111111_1110101110110010_1101100010111100"; -- -0.07930226724538583
	pesos_i(18717) := b"1111111111111111_1111111111111111_1101110011000101_0000110101010001"; -- -0.13761822474030114
	pesos_i(18718) := b"0000000000000000_0000000000000000_0001000011111011_0001001010110000"; -- 0.06633106991669015
	pesos_i(18719) := b"0000000000000000_0000000000000000_0010010110111011_0001100011011100"; -- 0.14738612535664916
	pesos_i(18720) := b"1111111111111111_1111111111111111_1111001000110110_1000100011000000"; -- -0.05385537442132408
	pesos_i(18721) := b"0000000000000000_0000000000000000_0001100001100111_0010100010000010"; -- 0.09532406979498359
	pesos_i(18722) := b"0000000000000000_0000000000000000_0010000011000100_0001011110001011"; -- 0.12799212596812007
	pesos_i(18723) := b"1111111111111111_1111111111111111_1110011110001111_1111110001111110"; -- -0.09545919349685915
	pesos_i(18724) := b"0000000000000000_0000000000000000_0001001100101111_0100011111001101"; -- 0.07494019284378355
	pesos_i(18725) := b"0000000000000000_0000000000000000_0000011111100010_1001100101000000"; -- 0.030801370671930013
	pesos_i(18726) := b"0000000000000000_0000000000000000_0000011111010001_1001101001000000"; -- 0.03054203095800047
	pesos_i(18727) := b"1111111111111111_1111111111111111_1101101000111100_1110000010110010"; -- -0.1475085797807893
	pesos_i(18728) := b"1111111111111111_1111111111111111_1111010111101110_0110110111000010"; -- -0.03933061622623886
	pesos_i(18729) := b"0000000000000000_0000000000000000_0000111010000111_1101110110011011"; -- 0.05676064529484793
	pesos_i(18730) := b"0000000000000000_0000000000000000_0001101100111010_0110011101111110"; -- 0.10635992849325841
	pesos_i(18731) := b"0000000000000000_0000000000000000_0000111001101101_1100001001001000"; -- 0.05636228798450132
	pesos_i(18732) := b"1111111111111111_1111111111111111_1111010001111100_0000101011011000"; -- -0.04498226374640301
	pesos_i(18733) := b"0000000000000000_0000000000000000_0000101000100000_0001011111000001"; -- 0.03955219697810586
	pesos_i(18734) := b"0000000000000000_0000000000000000_0001110111111111_1110101101011100"; -- 0.1171862697096897
	pesos_i(18735) := b"0000000000000000_0000000000000000_0001110101100010_0111101110001011"; -- 0.11478397497514893
	pesos_i(18736) := b"1111111111111111_1111111111111111_1111100011010101_1110110001100011"; -- -0.027985788238269575
	pesos_i(18737) := b"1111111111111111_1111111111111111_1110001001000101_1111000101001000"; -- -0.11612026200541853
	pesos_i(18738) := b"0000000000000000_0000000000000000_0001000010101101_1011101110011010"; -- 0.06515095239528658
	pesos_i(18739) := b"0000000000000000_0000000000000000_0010010010110010_1101011001010010"; -- 0.14335383903168283
	pesos_i(18740) := b"0000000000000000_0000000000000000_0001101110111111_0111110101100001"; -- 0.10839065187924754
	pesos_i(18741) := b"0000000000000000_0000000000000000_0000110100010011_0010001101101100"; -- 0.05107327832481373
	pesos_i(18742) := b"0000000000000000_0000000000000000_0001111010111111_1110011000000110"; -- 0.12011563916074001
	pesos_i(18743) := b"1111111111111111_1111111111111111_1111011000000000_0001011110100001"; -- -0.03906109169863832
	pesos_i(18744) := b"0000000000000000_0000000000000000_0000000001100110_0001000011100010"; -- 0.0015574027436206558
	pesos_i(18745) := b"0000000000000000_0000000000000000_0010110100101111_0100110101100001"; -- 0.1765030251271213
	pesos_i(18746) := b"1111111111111111_1111111111111111_1110010101010001_1110011011111010"; -- -0.10421902079671191
	pesos_i(18747) := b"1111111111111111_1111111111111111_1110111101110100_1001001011001010"; -- -0.06462748116455605
	pesos_i(18748) := b"1111111111111111_1111111111111111_1111000100001101_1100111100100100"; -- -0.05838303913118303
	pesos_i(18749) := b"0000000000000000_0000000000000000_0010000001110011_1100100000110000"; -- 0.12676669289912057
	pesos_i(18750) := b"1111111111111111_1111111111111111_1110000110000100_1100110010111011"; -- -0.11906738698384543
	pesos_i(18751) := b"1111111111111111_1111111111111111_1110011001000011_1010100110011100"; -- -0.1005300516365937
	pesos_i(18752) := b"0000000000000000_0000000000000000_0000101111001000_1110000101100110"; -- 0.046033942677622224
	pesos_i(18753) := b"0000000000000000_0000000000000000_0000000010010100_1001010101011001"; -- 0.0022672025134367426
	pesos_i(18754) := b"1111111111111111_1111111111111111_1101111011110011_1000010111011001"; -- -0.1290966362531979
	pesos_i(18755) := b"1111111111111111_1111111111111111_1111001100010101_1111011000001110"; -- -0.05044614939008672
	pesos_i(18756) := b"1111111111111111_1111111111111111_1111111111111100_1111011010001101"; -- -4.633960959027513e-05
	pesos_i(18757) := b"0000000000000000_0000000000000000_0000010110111000_1001010100011100"; -- 0.022347754907779058
	pesos_i(18758) := b"1111111111111111_1111111111111111_1110101110100111_0101000010101100"; -- -0.07947822379408788
	pesos_i(18759) := b"1111111111111111_1111111111111111_1111111000001001_0011110010110001"; -- -0.007671553378562619
	pesos_i(18760) := b"0000000000000000_0000000000000000_0001110100101101_0100100001000101"; -- 0.11397220313029359
	pesos_i(18761) := b"1111111111111111_1111111111111111_1101111100011111_1010111010011101"; -- -0.12842281988430437
	pesos_i(18762) := b"1111111111111111_1111111111111111_1101111111000100_1011110000001100"; -- -0.12590431880483033
	pesos_i(18763) := b"0000000000000000_0000000000000000_0000000011001000_1100111111111110"; -- 0.003064155214271848
	pesos_i(18764) := b"0000000000000000_0000000000000000_0000001110000110_1011111010001001"; -- 0.013774784463594736
	pesos_i(18765) := b"0000000000000000_0000000000000000_0000001010100011_1001110010010010"; -- 0.010309014929772792
	pesos_i(18766) := b"1111111111111111_1111111111111111_1110010111110111_1110011001000111"; -- -0.10168610357390596
	pesos_i(18767) := b"0000000000000000_0000000000000000_0001101111001001_0101101010000110"; -- 0.10854116231366386
	pesos_i(18768) := b"0000000000000000_0000000000000000_0010000010101100_0110000000101010"; -- 0.1276302436025674
	pesos_i(18769) := b"0000000000000000_0000000000000000_0001001001001111_0101111010011100"; -- 0.0715235835163744
	pesos_i(18770) := b"1111111111111111_1111111111111111_1111011101100011_1110110111100001"; -- -0.033631451296011014
	pesos_i(18771) := b"1111111111111111_1111111111111111_1111001010010001_0001000100011001"; -- -0.052473956373551366
	pesos_i(18772) := b"1111111111111111_1111111111111111_1111001100100111_1010011100011011"; -- -0.05017619706599245
	pesos_i(18773) := b"0000000000000000_0000000000000000_0000111010100010_1100010000001010"; -- 0.057171108612634955
	pesos_i(18774) := b"1111111111111111_1111111111111111_1111101000010110_1111001111111001"; -- -0.023087264687172107
	pesos_i(18775) := b"1111111111111111_1111111111111111_1110011110100110_0010110001100000"; -- -0.0951206460282721
	pesos_i(18776) := b"1111111111111111_1111111111111111_1111111001010101_0111010111000011"; -- -0.0065084838587742225
	pesos_i(18777) := b"1111111111111111_1111111111111111_1111110001110011_0001101001010011"; -- -0.013868670190961987
	pesos_i(18778) := b"1111111111111111_1111111111111111_1110001110001101_1110111110100101"; -- -0.1111154769194623
	pesos_i(18779) := b"1111111111111111_1111111111111111_1111100101011001_1101111101110100"; -- -0.025972398993769737
	pesos_i(18780) := b"1111111111111111_1111111111111111_1111101100111011_0011000011011001"; -- -0.01862806993474772
	pesos_i(18781) := b"0000000000000000_0000000000000000_0010000101000001_0011100111001001"; -- 0.12990151553458426
	pesos_i(18782) := b"1111111111111111_1111111111111111_1110001000101110_1101101101001111"; -- -0.11647252389305623
	pesos_i(18783) := b"1111111111111111_1111111111111111_1110111110010011_1110001111100100"; -- -0.06414962471127485
	pesos_i(18784) := b"0000000000000000_0000000000000000_0001011001001110_0001000100100011"; -- 0.0871287070672821
	pesos_i(18785) := b"0000000000000000_0000000000000000_0000001100101010_1001011011000101"; -- 0.012368605775269156
	pesos_i(18786) := b"0000000000000000_0000000000000000_0010000011001111_0111011011110001"; -- 0.12816565869167076
	pesos_i(18787) := b"0000000000000000_0000000000000000_0001001110011111_0010001110101110"; -- 0.07664702416178544
	pesos_i(18788) := b"1111111111111111_1111111111111111_1110110001111011_1100101010110101"; -- -0.07623608673123485
	pesos_i(18789) := b"1111111111111111_1111111111111111_1110001110010010_1101011101100111"; -- -0.11104062773775168
	pesos_i(18790) := b"1111111111111111_1111111111111111_1111011110101101_0011110010001111"; -- -0.032512869898234036
	pesos_i(18791) := b"1111111111111111_1111111111111111_1111100111000010_1001101111101111"; -- -0.024374250495905456
	pesos_i(18792) := b"1111111111111111_1111111111111111_1110001010101001_0001111001000111"; -- -0.11460695998812125
	pesos_i(18793) := b"0000000000000000_0000000000000000_0000001011010011_1011000101100001"; -- 0.011042677172287048
	pesos_i(18794) := b"1111111111111111_1111111111111111_1110100011001011_1001101111001101"; -- -0.0906431794561062
	pesos_i(18795) := b"0000000000000000_0000000000000000_0000010000011011_0111000110000000"; -- 0.016043752481351734
	pesos_i(18796) := b"0000000000000000_0000000000000000_0001100100000000_0111001101100110"; -- 0.09766312830045128
	pesos_i(18797) := b"0000000000000000_0000000000000000_0001100000111001_0001000100010110"; -- 0.09462076931845882
	pesos_i(18798) := b"1111111111111111_1111111111111111_1101000001111001_1111101101111010"; -- -0.18563869727030285
	pesos_i(18799) := b"0000000000000000_0000000000000000_0000000011101010_0101001011011100"; -- 0.003575495480351156
	pesos_i(18800) := b"0000000000000000_0000000000000000_0000000000000111_1101010011100010"; -- 0.00011950022152556345
	pesos_i(18801) := b"1111111111111111_1111111111111111_1110001000101110_1100011110111001"; -- -0.11647369131698358
	pesos_i(18802) := b"0000000000000000_0000000000000000_0000000011100011_1001111001111000"; -- 0.0034731904791786374
	pesos_i(18803) := b"1111111111111111_1111111111111111_1111011110010100_1001000111111100"; -- -0.03288924783589549
	pesos_i(18804) := b"1111111111111111_1111111111111111_1101110011110000_1110101101001011"; -- -0.13694886616703952
	pesos_i(18805) := b"0000000000000000_0000000000000000_0001011001011101_0111110111011111"; -- 0.0873640698702899
	pesos_i(18806) := b"0000000000000000_0000000000000000_0000011100001011_0000011011001011"; -- 0.02751200154012605
	pesos_i(18807) := b"1111111111111111_1111111111111111_1101101000100011_0010110010011010"; -- -0.14790078389693131
	pesos_i(18808) := b"0000000000000000_0000000000000000_0010011001010010_0011010000101101"; -- 0.14969183052022303
	pesos_i(18809) := b"0000000000000000_0000000000000000_0000010101101000_0111111100000011"; -- 0.02112573460060687
	pesos_i(18810) := b"1111111111111111_1111111111111111_1111011100110110_0100001011100000"; -- -0.03432828941083184
	pesos_i(18811) := b"1111111111111111_1111111111111111_1101001110011100_0011111000101100"; -- -0.1733971732174506
	pesos_i(18812) := b"1111111111111111_1111111111111111_1111011111010011_1110110000011010"; -- -0.031922572698688784
	pesos_i(18813) := b"1111111111111111_1111111111111111_1111101011000110_0000001000011110"; -- -0.02041613364131652
	pesos_i(18814) := b"1111111111111111_1111111111111111_1111101101110001_1001010001101101"; -- -0.017798159883624636
	pesos_i(18815) := b"1111111111111111_1111111111111111_1101101011111000_0000010111011101"; -- -0.14465297092598992
	pesos_i(18816) := b"0000000000000000_0000000000000000_0000101001001100_1111100000111101"; -- 0.040236964101955826
	pesos_i(18817) := b"1111111111111111_1111111111111111_1111111101110011_0001101110011000"; -- -0.002149844516376365
	pesos_i(18818) := b"0000000000000000_0000000000000000_0000110100101000_1111100010010101"; -- 0.05140641811521028
	pesos_i(18819) := b"1111111111111111_1111111111111111_1101100110011011_1110011000101010"; -- -0.14996491892310004
	pesos_i(18820) := b"1111111111111111_1111111111111111_1101110110101110_1111000101110010"; -- -0.13404932950060813
	pesos_i(18821) := b"1111111111111111_1111111111111111_1101100000101110_0111110010011100"; -- -0.1555406684145511
	pesos_i(18822) := b"1111111111111111_1111111111111111_1101100100110101_0010111001010100"; -- -0.15153227292456256
	pesos_i(18823) := b"0000000000000000_0000000000000000_0000010101000100_0010111111000111"; -- 0.020571695481441173
	pesos_i(18824) := b"1111111111111111_1111111111111111_1111010010010010_1101110101101101"; -- -0.044634018720741776
	pesos_i(18825) := b"0000000000000000_0000000000000000_0001110010000010_0001011101111001"; -- 0.11136004157097691
	pesos_i(18826) := b"1111111111111111_1111111111111111_1110001101011000_0000111000010000"; -- -0.1119376383378761
	pesos_i(18827) := b"0000000000000000_0000000000000000_0000111101000101_0001000011001111"; -- 0.059647608403025985
	pesos_i(18828) := b"1111111111111111_1111111111111111_1111101010011010_1111100001010000"; -- -0.021072845934899647
	pesos_i(18829) := b"0000000000000000_0000000000000000_0001101100111110_0010000100000101"; -- 0.10641676293699237
	pesos_i(18830) := b"0000000000000000_0000000000000000_0010010010000100_0101110010011110"; -- 0.14264468067449404
	pesos_i(18831) := b"1111111111111111_1111111111111111_1110011001101010_1011111101011010"; -- -0.09993366290732165
	pesos_i(18832) := b"1111111111111111_1111111111111111_1111110011001110_0100111011100111"; -- -0.012476986484642582
	pesos_i(18833) := b"1111111111111111_1111111111111111_1111111010101111_0111110000001101"; -- -0.005134817824117524
	pesos_i(18834) := b"1111111111111111_1111111111111111_1111101011111111_0010100111010001"; -- -0.01954401640918571
	pesos_i(18835) := b"0000000000000000_0000000000000000_0001111010101110_1101101000100101"; -- 0.11985553182176546
	pesos_i(18836) := b"1111111111111111_1111111111111111_1110011001111110_0001111011011010"; -- -0.09963805359017877
	pesos_i(18837) := b"0000000000000000_0000000000000000_0000010110001101_0010010010001111"; -- 0.021684918425851865
	pesos_i(18838) := b"0000000000000000_0000000000000000_0001100000011001_0010000111111000"; -- 0.09413349453062726
	pesos_i(18839) := b"1111111111111111_1111111111111111_1111001101111000_1110011001111001"; -- -0.04893645816204829
	pesos_i(18840) := b"1111111111111111_1111111111111111_1111100110111000_0010011010011110"; -- -0.02453383103495534
	pesos_i(18841) := b"0000000000000000_0000000000000000_0001000011001000_1010000100010110"; -- 0.06556135922925031
	pesos_i(18842) := b"0000000000000000_0000000000000000_0001111100101000_0000001101101000"; -- 0.12170430464373495
	pesos_i(18843) := b"1111111111111111_1111111111111111_1110010000100101_1110101011011110"; -- -0.10879642559815358
	pesos_i(18844) := b"0000000000000000_0000000000000000_0010000111010001_1110111010111101"; -- 0.1321095669329737
	pesos_i(18845) := b"0000000000000000_0000000000000000_0000110001100100_0111101100011111"; -- 0.048408217536529505
	pesos_i(18846) := b"1111111111111111_1111111111111111_1111001110010011_1011000101001110"; -- -0.04852763979280504
	pesos_i(18847) := b"0000000000000000_0000000000000000_0001000001101011_1011000111111010"; -- 0.06414329873226211
	pesos_i(18848) := b"1111111111111111_1111111111111111_1110001000110000_0000110100001010"; -- -0.11645430093621194
	pesos_i(18849) := b"0000000000000000_0000000000000000_0000110001000100_1001100001111000"; -- 0.047921685536107685
	pesos_i(18850) := b"1111111111111111_1111111111111111_1111100000100101_0001101011010000"; -- -0.03068382664752385
	pesos_i(18851) := b"0000000000000000_0000000000000000_0000001000011011_0001011011000011"; -- 0.008225843992106133
	pesos_i(18852) := b"1111111111111111_1111111111111111_1111111000001000_0010001111100010"; -- -0.007688290879220353
	pesos_i(18853) := b"1111111111111111_1111111111111111_1110101101111110_1100110100101011"; -- -0.08009641362878499
	pesos_i(18854) := b"1111111111111111_1111111111111111_1111011001101000_1111101111100111"; -- -0.03746057127998833
	pesos_i(18855) := b"0000000000000000_0000000000000000_0000110001000010_0011011010110010"; -- 0.04788534017844233
	pesos_i(18856) := b"1111111111111111_1111111111111111_1110100100010001_1110110111101101"; -- -0.08957016914596615
	pesos_i(18857) := b"0000000000000000_0000000000000000_0010010010011110_0111101101111011"; -- 0.14304324862728846
	pesos_i(18858) := b"1111111111111111_1111111111111111_1110011110100010_0000010111111001"; -- -0.09518397021962165
	pesos_i(18859) := b"1111111111111111_1111111111111111_1101111000101101_1001100011000111"; -- -0.13211674817504132
	pesos_i(18860) := b"0000000000000000_0000000000000000_0000110000111111_0011001010001001"; -- 0.047839315949656507
	pesos_i(18861) := b"1111111111111111_1111111111111111_1110011111111000_1111000110000110"; -- -0.09385767441190612
	pesos_i(18862) := b"0000000000000000_0000000000000000_0000010000110100_1110001001101111"; -- 0.016431953577062813
	pesos_i(18863) := b"1111111111111111_1111111111111111_1111101111001100_0101100110011000"; -- -0.016413116806102034
	pesos_i(18864) := b"1111111111111111_1111111111111111_1111000111100000_1000100111000000"; -- -0.05516757065160003
	pesos_i(18865) := b"0000000000000000_0000000000000000_0001000110100111_1101001010000100"; -- 0.06896701543762751
	pesos_i(18866) := b"1111111111111111_1111111111111111_1101101111000010_0111111101101110"; -- -0.1415634494207932
	pesos_i(18867) := b"1111111111111111_1111111111111111_1111110000000111_0100011011111010"; -- -0.0155139580544106
	pesos_i(18868) := b"0000000000000000_0000000000000000_0000100100101111_1010111000010001"; -- 0.03588378834142586
	pesos_i(18869) := b"0000000000000000_0000000000000000_0001001000101110_1001001010001011"; -- 0.07102313898523295
	pesos_i(18870) := b"1111111111111111_1111111111111111_1110000100001101_0101010011100111"; -- -0.12089032513996982
	pesos_i(18871) := b"1111111111111111_1111111111111111_1111010001010001_0001100010100111"; -- -0.04563756861898232
	pesos_i(18872) := b"0000000000000000_0000000000000000_0001111101010110_0011110111100101"; -- 0.12240969517669806
	pesos_i(18873) := b"1111111111111111_1111111111111111_1111011000100010_0010100101110010"; -- -0.038541230925636626
	pesos_i(18874) := b"1111111111111111_1111111111111111_1110001101101110_0000110101111110"; -- -0.11160197904523837
	pesos_i(18875) := b"0000000000000000_0000000000000000_0000110001010111_1110001011001011"; -- 0.048216032583543705
	pesos_i(18876) := b"0000000000000000_0000000000000000_0010000110011111_1011100110011110"; -- 0.1313434610607785
	pesos_i(18877) := b"0000000000000000_0000000000000000_0010000010000110_0010000100111101"; -- 0.1270466588383833
	pesos_i(18878) := b"1111111111111111_1111111111111111_1111110110111010_1110000001000011"; -- -0.00886724824242325
	pesos_i(18879) := b"0000000000000000_0000000000000000_0010011001100000_1110111001100110"; -- 0.14991655350844732
	pesos_i(18880) := b"0000000000000000_0000000000000000_0001011100100110_0110001000011101"; -- 0.09042943208342435
	pesos_i(18881) := b"0000000000000000_0000000000000000_0010100010100011_1111010100010000"; -- 0.1587517894906615
	pesos_i(18882) := b"1111111111111111_1111111111111111_1101110100000100_1100111010111011"; -- -0.1366453928082962
	pesos_i(18883) := b"0000000000000000_0000000000000000_0010000000101000_1111110010111010"; -- 0.12562541534170485
	pesos_i(18884) := b"0000000000000000_0000000000000000_0001101010000011_0010010101110010"; -- 0.10356363339755684
	pesos_i(18885) := b"0000000000000000_0000000000000000_0001011000110010_1000011111100001"; -- 0.08670853847967007
	pesos_i(18886) := b"1111111111111111_1111111111111111_1111011111101001_1101001100101100"; -- -0.03158836537576167
	pesos_i(18887) := b"0000000000000000_0000000000000000_0001111010110001_0100111001001010"; -- 0.11989297203735674
	pesos_i(18888) := b"1111111111111111_1111111111111111_1110001011001011_0111110111011110"; -- -0.11408246356218815
	pesos_i(18889) := b"0000000000000000_0000000000000000_0000011001010111_1100100111110000"; -- 0.02477705097023131
	pesos_i(18890) := b"1111111111111111_1111111111111111_1111000100101110_1110011110101000"; -- -0.05787803788621552
	pesos_i(18891) := b"0000000000000000_0000000000000000_0000010000001101_1011001100000000"; -- 0.01583403357500007
	pesos_i(18892) := b"1111111111111111_1111111111111111_1111010011110111_0111111011110100"; -- -0.04309851199351278
	pesos_i(18893) := b"0000000000000000_0000000000000000_0001000110110101_0011100110110111"; -- 0.06917153083889384
	pesos_i(18894) := b"0000000000000000_0000000000000000_0001001111010001_0000011101010011"; -- 0.07740827349149887
	pesos_i(18895) := b"1111111111111111_1111111111111111_1111011111101010_1101100110010110"; -- -0.03157272425843301
	pesos_i(18896) := b"1111111111111111_1111111111111111_1111011100000111_0110111110000100"; -- -0.03504279163762742
	pesos_i(18897) := b"1111111111111111_1111111111111111_1110110000110100_0001101000100011"; -- -0.07732998510950954
	pesos_i(18898) := b"1111111111111111_1111111111111111_1111101101101111_1110101010101010"; -- -0.017823537416829356
	pesos_i(18899) := b"1111111111111111_1111111111111111_1111011011011011_1101000100000111"; -- -0.035708366277133155
	pesos_i(18900) := b"1111111111111111_1111111111111111_1101111001110010_1000110101001000"; -- -0.1310645769808208
	pesos_i(18901) := b"0000000000000000_0000000000000000_0001110100101000_1101011111110011"; -- 0.11390447324950162
	pesos_i(18902) := b"1111111111111111_1111111111111111_1111110000111011_0000110011011111"; -- -0.014723964241493973
	pesos_i(18903) := b"1111111111111111_1111111111111111_1110110110011100_1010011001101101"; -- -0.07182845917762243
	pesos_i(18904) := b"0000000000000000_0000000000000000_0010011101111010_1011011101010111"; -- 0.1542162501244518
	pesos_i(18905) := b"1111111111111111_1111111111111111_1111000011010110_0011001111111000"; -- -0.059231521631167496
	pesos_i(18906) := b"1111111111111111_1111111111111111_1111000100010001_0011111100001000"; -- -0.05833059370489815
	pesos_i(18907) := b"1111111111111111_1111111111111111_1111010010100100_0001000010100000"; -- -0.044371567708906406
	pesos_i(18908) := b"1111111111111111_1111111111111111_1110101001001110_0000101010101100"; -- -0.08474667829561969
	pesos_i(18909) := b"1111111111111111_1111111111111111_1110011110100100_1100001011001100"; -- -0.09514219789368031
	pesos_i(18910) := b"1111111111111111_1111111111111111_1110101111000101_0100110101100010"; -- -0.07902065615843072
	pesos_i(18911) := b"1111111111111111_1111111111111111_1110100000000101_1100111111101100"; -- -0.09366131300091675
	pesos_i(18912) := b"1111111111111111_1111111111111111_1111000001010100_1010001010111010"; -- -0.06120856248138716
	pesos_i(18913) := b"1111111111111111_1111111111111111_1110001111000001_0011110101000100"; -- -0.11033265198076365
	pesos_i(18914) := b"0000000000000000_0000000000000000_0001111001000110_0111011010101011"; -- 0.1182626884470795
	pesos_i(18915) := b"0000000000000000_0000000000000000_0000011011111101_1110101100010010"; -- 0.02731198484315099
	pesos_i(18916) := b"0000000000000000_0000000000000000_0001111100011010_0100011111111001"; -- 0.12149476837281421
	pesos_i(18917) := b"0000000000000000_0000000000000000_0001111101110001_1010000110110101"; -- 0.12282763168535317
	pesos_i(18918) := b"0000000000000000_0000000000000000_0000101010111110_0010111010100011"; -- 0.041964449739142484
	pesos_i(18919) := b"1111111111111111_1111111111111111_1101110000011111_1001100101001111"; -- -0.14014283952017312
	pesos_i(18920) := b"1111111111111111_1111111111111111_1101101010111011_1000111000011010"; -- -0.14557563644866658
	pesos_i(18921) := b"1111111111111111_1111111111111111_1111110010000101_1000000101110011"; -- -0.013587865280999435
	pesos_i(18922) := b"1111111111111111_1111111111111111_1111100101101000_0011110110010101"; -- -0.025753165286755978
	pesos_i(18923) := b"0000000000000000_0000000000000000_0001010100001000_1100101011000000"; -- 0.08216540521483111
	pesos_i(18924) := b"1111111111111111_1111111111111111_1110010000100001_1011010001011110"; -- -0.10886070930202978
	pesos_i(18925) := b"0000000000000000_0000000000000000_0010010000111010_1010001101001110"; -- 0.14151974351154648
	pesos_i(18926) := b"0000000000000000_0000000000000000_0000101100110010_0101111100001001"; -- 0.04373735390397606
	pesos_i(18927) := b"1111111111111111_1111111111111111_1111110110011010_0100011001001110"; -- -0.009364705952857951
	pesos_i(18928) := b"0000000000000000_0000000000000000_0000010111101100_0000101110100111"; -- 0.023133018674747076
	pesos_i(18929) := b"1111111111111111_1111111111111111_1111100001011110_1111101110101010"; -- -0.02980067354395557
	pesos_i(18930) := b"1111111111111111_1111111111111111_1111001101100100_0011100011110000"; -- -0.049251977251143365
	pesos_i(18931) := b"1111111111111111_1111111111111111_1111001011000011_1101000110110010"; -- -0.05169953738824618
	pesos_i(18932) := b"0000000000000000_0000000000000000_0001101011011001_1101010000000100"; -- 0.10488629432415196
	pesos_i(18933) := b"1111111111111111_1111111111111111_1110100101010111_0010001110010000"; -- -0.08851411555344105
	pesos_i(18934) := b"0000000000000000_0000000000000000_0001001111010010_0010000101101111"; -- 0.07742508841169109
	pesos_i(18935) := b"1111111111111111_1111111111111111_1101101100101100_1000100001111100"; -- -0.14385172814460284
	pesos_i(18936) := b"0000000000000000_0000000000000000_0001100111011100_1110111010001001"; -- 0.10102740136737325
	pesos_i(18937) := b"1111111111111111_1111111111111111_1111001111000110_1011100100010001"; -- -0.04774897903692851
	pesos_i(18938) := b"0000000000000000_0000000000000000_0000011101010010_0001100011001111"; -- 0.028596449446090844
	pesos_i(18939) := b"0000000000000000_0000000000000000_0010100010011010_1001101001101000"; -- 0.1586090568869227
	pesos_i(18940) := b"0000000000000000_0000000000000000_0010000100101011_1011111111111011"; -- 0.12957382074654053
	pesos_i(18941) := b"0000000000000000_0000000000000000_0000001111101101_1001111111011101"; -- 0.015344611555338002
	pesos_i(18942) := b"1111111111111111_1111111111111111_1101110110011110_1010000100010100"; -- -0.13429826039144951
	pesos_i(18943) := b"1111111111111111_1111111111111111_1111011001110100_0010011111100001"; -- -0.03729010352695307
	pesos_i(18944) := b"1111111111111111_1111111111111111_1111111110101100_1000011111010000"; -- -0.00127364321601694
	pesos_i(18945) := b"0000000000000000_0000000000000000_0000000010110110_1110100101100000"; -- 0.0027910099080953343
	pesos_i(18946) := b"1111111111111111_1111111111111111_1110000000100011_0111101101001000"; -- -0.1244585941765386
	pesos_i(18947) := b"1111111111111111_1111111111111111_1111100011110011_0100101101110011"; -- -0.027537617022068726
	pesos_i(18948) := b"0000000000000000_0000000000000000_0001110100010000_1001100000100101"; -- 0.11353445926207453
	pesos_i(18949) := b"0000000000000000_0000000000000000_0010001111100010_1110010000011101"; -- 0.14018083299056472
	pesos_i(18950) := b"0000000000000000_0000000000000000_0000010001110000_0010110101001000"; -- 0.01733668340163071
	pesos_i(18951) := b"1111111111111111_1111111111111111_1111011000010111_0011101000011101"; -- -0.03870808413076686
	pesos_i(18952) := b"1111111111111111_1111111111111111_1110110010011000_1001111000010000"; -- -0.07579624290669863
	pesos_i(18953) := b"1111111111111111_1111111111111111_1111110101001100_1100111100101100"; -- -0.010546733543729757
	pesos_i(18954) := b"1111111111111111_1111111111111111_1111000101011000_1100000101101010"; -- -0.057239448286296686
	pesos_i(18955) := b"0000000000000000_0000000000000000_0000101110111010_1010101101100101"; -- 0.045817100729526904
	pesos_i(18956) := b"0000000000000000_0000000000000000_0001000000111011_0001100111101010"; -- 0.06340181322460521
	pesos_i(18957) := b"0000000000000000_0000000000000000_0001100000101011_0010100010110111"; -- 0.09440855474124533
	pesos_i(18958) := b"0000000000000000_0000000000000000_0001001001100010_0010010111010100"; -- 0.07181011599557909
	pesos_i(18959) := b"1111111111111111_1111111111111111_1111111100110110_0101101000110001"; -- -0.00307689960966668
	pesos_i(18960) := b"1111111111111111_1111111111111111_1110111101001000_1010011011011101"; -- -0.06529767139390615
	pesos_i(18961) := b"0000000000000000_0000000000000000_0001101000101000_0011100110110100"; -- 0.10217629092435865
	pesos_i(18962) := b"1111111111111111_1111111111111111_1110001011101011_0110101101001000"; -- -0.11359529020686893
	pesos_i(18963) := b"0000000000000000_0000000000000000_0001011000101000_0100101010011000"; -- 0.08655229771259865
	pesos_i(18964) := b"1111111111111111_1111111111111111_1110001001011010_1010001111000011"; -- -0.11580444802912608
	pesos_i(18965) := b"0000000000000000_0000000000000000_0000110000011110_0101010101101000"; -- 0.04733785427178212
	pesos_i(18966) := b"0000000000000000_0000000000000000_0000001100001100_1010001001000100"; -- 0.011911527139704817
	pesos_i(18967) := b"1111111111111111_1111111111111111_1110001011000000_0100010011111110"; -- -0.11425370030234923
	pesos_i(18968) := b"1111111111111111_1111111111111111_1111000011111110_1010100110111100"; -- -0.05861415060172817
	pesos_i(18969) := b"0000000000000000_0000000000000000_0000100001010111_1011110001100100"; -- 0.032588743679675916
	pesos_i(18970) := b"0000000000000000_0000000000000000_0000011001010100_0101110111101101"; -- 0.024724836716903186
	pesos_i(18971) := b"1111111111111111_1111111111111111_1110100000101000_0010110100010101"; -- -0.09313696125718061
	pesos_i(18972) := b"0000000000000000_0000000000000000_0000000101000101_1001000000111100"; -- 0.004967703381605559
	pesos_i(18973) := b"1111111111111111_1111111111111111_1111100001100001_1101101101111010"; -- -0.029756815715130808
	pesos_i(18974) := b"0000000000000000_0000000000000000_0010010000110000_0001110110111110"; -- 0.1413591946910431
	pesos_i(18975) := b"0000000000000000_0000000000000000_0000101001101010_0011010100111110"; -- 0.040683105028058275
	pesos_i(18976) := b"1111111111111111_1111111111111111_1110000010110011_0001000011110101"; -- -0.12226766594307745
	pesos_i(18977) := b"1111111111111111_1111111111111111_1111101101100000_0010110110100000"; -- -0.01806368680396867
	pesos_i(18978) := b"1111111111111111_1111111111111111_1111111101100011_0100011000111001"; -- -0.0023914442533226354
	pesos_i(18979) := b"0000000000000000_0000000000000000_0000111100100010_1001010100110010"; -- 0.05912144153624645
	pesos_i(18980) := b"0000000000000000_0000000000000000_0001111101111011_0010011001111110"; -- 0.12297287538579602
	pesos_i(18981) := b"1111111111111111_1111111111111111_1110000111010110_1000100011000011"; -- -0.11782021740971789
	pesos_i(18982) := b"1111111111111111_1111111111111111_1110111110100100_0000010011000001"; -- -0.06390352534788202
	pesos_i(18983) := b"0000000000000000_0000000000000000_0000110001010000_1010110001010001"; -- 0.04810597400392565
	pesos_i(18984) := b"1111111111111111_1111111111111111_1110110110111100_1111100011110110"; -- -0.07133525833908887
	pesos_i(18985) := b"0000000000000000_0000000000000000_0010000110111000_0101110101000011"; -- 0.13171942603278858
	pesos_i(18986) := b"0000000000000000_0000000000000000_0010000100100000_0111010001111101"; -- 0.12940147446655934
	pesos_i(18987) := b"1111111111111111_1111111111111111_1110010111100000_1010001100001111"; -- -0.10204106225804334
	pesos_i(18988) := b"1111111111111111_1111111111111111_1111110101111110_1110001100110011"; -- -0.009782600447559254
	pesos_i(18989) := b"0000000000000000_0000000000000000_0000100100001000_1110011110100100"; -- 0.03529212714050524
	pesos_i(18990) := b"0000000000000000_0000000000000000_0001100011001101_0111011000101110"; -- 0.09688509589746666
	pesos_i(18991) := b"1111111111111111_1111111111111111_1111101110010010_1010110001101010"; -- -0.017293190007438043
	pesos_i(18992) := b"1111111111111111_1111111111111111_1111110100011100_1101100010111110"; -- -0.011278585024970351
	pesos_i(18993) := b"1111111111111111_1111111111111111_1111011111010101_0110101110101111"; -- -0.031899709579011636
	pesos_i(18994) := b"0000000000000000_0000000000000000_0001001100001101_0110000010011011"; -- 0.07442287230892655
	pesos_i(18995) := b"1111111111111111_1111111111111111_1110100001000001_0111111111110100"; -- -0.09275055200805554
	pesos_i(18996) := b"0000000000000000_0000000000000000_0010000101100001_0111100111010011"; -- 0.13039361376350486
	pesos_i(18997) := b"0000000000000000_0000000000000000_0001001011001110_1101000010001101"; -- 0.07346824124239736
	pesos_i(18998) := b"1111111111111111_1111111111111111_1101110011110011_1011010010100100"; -- -0.13690634719942388
	pesos_i(18999) := b"1111111111111111_1111111111111111_1111001101110011_1010011110000100"; -- -0.04901650450653426
	pesos_i(19000) := b"0000000000000000_0000000000000000_0000100100100010_0111011010101101"; -- 0.03568212240389564
	pesos_i(19001) := b"1111111111111111_1111111111111111_1111101100001001_1101101001011111"; -- -0.019380904920223367
	pesos_i(19002) := b"0000000000000000_0000000000000000_0000101011100110_0111001100101101"; -- 0.04257888655183761
	pesos_i(19003) := b"1111111111111111_1111111111111111_1111010000001111_0111010001010101"; -- -0.04663918419423714
	pesos_i(19004) := b"1111111111111111_1111111111111111_1111011011000001_0101110100100110"; -- -0.03611200156273335
	pesos_i(19005) := b"1111111111111111_1111111111111111_1111111100001010_0101001000010100"; -- -0.0037487698134707065
	pesos_i(19006) := b"1111111111111111_1111111111111111_1111011001001000_1011110110011111"; -- -0.03795256477947552
	pesos_i(19007) := b"0000000000000000_0000000000000000_0000011010011000_1001101011000111"; -- 0.02576606135680772
	pesos_i(19008) := b"0000000000000000_0000000000000000_0001001110010111_0010110100101011"; -- 0.07652551943788224
	pesos_i(19009) := b"1111111111111111_1111111111111111_1101111001011110_0010011001000110"; -- -0.13137589264296295
	pesos_i(19010) := b"1111111111111111_1111111111111111_1101101000101111_1001101101101111"; -- -0.14771107232342012
	pesos_i(19011) := b"1111111111111111_1111111111111111_1110100101010011_0001001111110001"; -- -0.08857608179546485
	pesos_i(19012) := b"1111111111111111_1111111111111111_1111100101110110_0000101001011001"; -- -0.02554259607934509
	pesos_i(19013) := b"0000000000000000_0000000000000000_0001111110100100_1010001011000010"; -- 0.1236058924610431
	pesos_i(19014) := b"0000000000000000_0000000000000000_0000110011011111_1100110100011011"; -- 0.05028993520424573
	pesos_i(19015) := b"1111111111111111_1111111111111111_1111001010101100_0101110111110111"; -- -0.05205738748247797
	pesos_i(19016) := b"1111111111111111_1111111111111111_1101100110100100_1001011001101011"; -- -0.1498323429986637
	pesos_i(19017) := b"0000000000000000_0000000000000000_0000100000001100_1000100000110111"; -- 0.03144122460174048
	pesos_i(19018) := b"0000000000000000_0000000000000000_0001011101100101_1111101000001011"; -- 0.09139979132603025
	pesos_i(19019) := b"1111111111111111_1111111111111111_1111000111110110_1111101000011101"; -- -0.05482517993401543
	pesos_i(19020) := b"1111111111111111_1111111111111111_1111010110110000_1100111111001111"; -- -0.040270816822056646
	pesos_i(19021) := b"1111111111111111_1111111111111111_1101110111011111_1010101100010111"; -- -0.13330584221313987
	pesos_i(19022) := b"0000000000000000_0000000000000000_0010001110111011_1000001010111001"; -- 0.13957993517550876
	pesos_i(19023) := b"0000000000000000_0000000000000000_0001001001011110_1101001100110101"; -- 0.07175941511474736
	pesos_i(19024) := b"0000000000000000_0000000000000000_0000011110111110_0010100011101011"; -- 0.030245358800031215
	pesos_i(19025) := b"0000000000000000_0000000000000000_0000011000000000_1001001111101111"; -- 0.023446317621438097
	pesos_i(19026) := b"0000000000000000_0000000000000000_0010001100010100_0101110011111000"; -- 0.13702946703613053
	pesos_i(19027) := b"0000000000000000_0000000000000000_0001001011000011_1010001100001110"; -- 0.07329768274707073
	pesos_i(19028) := b"0000000000000000_0000000000000000_0000010110100010_0100001000110111"; -- 0.022007120484236736
	pesos_i(19029) := b"0000000000000000_0000000000000000_0001010000011110_0000001010000010"; -- 0.07858291318621471
	pesos_i(19030) := b"1111111111111111_1111111111111111_1101111001101100_0110100100000000"; -- -0.13115829240752452
	pesos_i(19031) := b"1111111111111111_1111111111111111_1110000110111011_1000110010011010"; -- -0.11823197582525916
	pesos_i(19032) := b"0000000000000000_0000000000000000_0010011000110010_1110101101000000"; -- 0.14921446144646003
	pesos_i(19033) := b"1111111111111111_1111111111111111_1110101111110011_1000101001000111"; -- -0.07831512238536253
	pesos_i(19034) := b"1111111111111111_1111111111111111_1110001100001011_0111000101101001"; -- -0.11310664350708872
	pesos_i(19035) := b"0000000000000000_0000000000000000_0001011001000101_0100110011000010"; -- 0.08699493156069654
	pesos_i(19036) := b"0000000000000000_0000000000000000_0010000110011001_0011010001011001"; -- 0.13124396486928283
	pesos_i(19037) := b"0000000000000000_0000000000000000_0000100000000111_0100000011101110"; -- 0.031360681544948754
	pesos_i(19038) := b"1111111111111111_1111111111111111_1110110000110110_1101001010101010"; -- -0.07728846874154618
	pesos_i(19039) := b"1111111111111111_1111111111111111_1111011110101100_1011111000001011"; -- -0.03252041087176697
	pesos_i(19040) := b"0000000000000000_0000000000000000_0001011100101011_0111011011110110"; -- 0.09050696864516755
	pesos_i(19041) := b"1111111111111111_1111111111111111_1101111100000111_1110111101011111"; -- -0.12878517088992603
	pesos_i(19042) := b"1111111111111111_1111111111111111_1110011001110100_1110001001111000"; -- -0.09977898197845049
	pesos_i(19043) := b"1111111111111111_1111111111111111_1110100101000101_1100011000010000"; -- -0.08877908819481241
	pesos_i(19044) := b"1111111111111111_1111111111111111_1111110011100110_0000111101000100"; -- -0.012114568690438006
	pesos_i(19045) := b"0000000000000000_0000000000000000_0010010101111110_0011110000100000"; -- 0.14645744109820877
	pesos_i(19046) := b"0000000000000000_0000000000000000_0000000011111001_0111011001100100"; -- 0.0038064951300258946
	pesos_i(19047) := b"1111111111111111_1111111111111111_1111011001000110_0110000111000100"; -- -0.03798855749115204
	pesos_i(19048) := b"1111111111111111_1111111111111111_1111110101000010_0011011110100100"; -- -0.010708353385048766
	pesos_i(19049) := b"0000000000000000_0000000000000000_0001100111001010_1010011000111001"; -- 0.1007484330273115
	pesos_i(19050) := b"1111111111111111_1111111111111111_1110101101101001_0010100011001100"; -- -0.08042664542503522
	pesos_i(19051) := b"1111111111111111_1111111111111111_1111010111101111_1010111101001010"; -- -0.03931145129645406
	pesos_i(19052) := b"1111111111111111_1111111111111111_1110011000000010_1101011100010010"; -- -0.10151916322642673
	pesos_i(19053) := b"0000000000000000_0000000000000000_0000111001000001_1111010111101000"; -- 0.055693978490414825
	pesos_i(19054) := b"1111111111111111_1111111111111111_1110100110000010_1011110110100000"; -- -0.08784880479719204
	pesos_i(19055) := b"0000000000000000_0000000000000000_0001101100001000_1111011100001110"; -- 0.10560554594917902
	pesos_i(19056) := b"0000000000000000_0000000000000000_0000110010100111_0110111101010010"; -- 0.04942985292292022
	pesos_i(19057) := b"0000000000000000_0000000000000000_0000111111100110_0011001111000010"; -- 0.06210635650680334
	pesos_i(19058) := b"1111111111111111_1111111111111111_1111111110011111_1001011111010100"; -- -0.0014710528406892283
	pesos_i(19059) := b"1111111111111111_1111111111111111_1110100100111001_0010011100101111"; -- -0.08897166348251634
	pesos_i(19060) := b"0000000000000000_0000000000000000_0000101100110100_1110100100101010"; -- 0.043776104672791395
	pesos_i(19061) := b"0000000000000000_0000000000000000_0000110101001001_0010001110001100"; -- 0.051897260439284554
	pesos_i(19062) := b"0000000000000000_0000000000000000_0000011101101110_0001100110001111"; -- 0.029023740206957183
	pesos_i(19063) := b"1111111111111111_1111111111111111_1110010100100000_0000010101000100"; -- -0.10498015499967159
	pesos_i(19064) := b"1111111111111111_1111111111111111_1111000110110110_0000101100101001"; -- -0.05581598519729757
	pesos_i(19065) := b"0000000000000000_0000000000000000_0001101000100111_1101001001100110"; -- 0.10217013351978857
	pesos_i(19066) := b"0000000000000000_0000000000000000_0000010100011000_1101001010101011"; -- 0.019910017781059566
	pesos_i(19067) := b"0000000000000000_0000000000000000_0001010111110010_0010110010110000"; -- 0.08572654052330396
	pesos_i(19068) := b"1111111111111111_1111111111111111_1101110000110111_0101100100100010"; -- -0.13978045379409726
	pesos_i(19069) := b"0000000000000000_0000000000000000_0000010011111101_0100001011011110"; -- 0.019489459181999784
	pesos_i(19070) := b"0000000000000000_0000000000000000_0001111010010011_0000001001111101"; -- 0.11943069035421565
	pesos_i(19071) := b"0000000000000000_0000000000000000_0010001100011000_0011111110010011"; -- 0.13708875015784747
	pesos_i(19072) := b"1111111111111111_1111111111111111_1111010110010100_1101000010101001"; -- -0.04069801208922773
	pesos_i(19073) := b"0000000000000000_0000000000000000_0000001001110001_0101111110011011"; -- 0.009542441613589263
	pesos_i(19074) := b"0000000000000000_0000000000000000_0000100001110111_0001001000010011"; -- 0.03306687312145503
	pesos_i(19075) := b"0000000000000000_0000000000000000_0001000001010010_1100100111011011"; -- 0.06376325218420942
	pesos_i(19076) := b"0000000000000000_0000000000000000_0001010100110010_1110001001110111"; -- 0.08280768773605292
	pesos_i(19077) := b"0000000000000000_0000000000000000_0001111001000110_0110101011011000"; -- 0.11826198370702402
	pesos_i(19078) := b"0000000000000000_0000000000000000_0001001011111011_0001000010001111"; -- 0.0741434429724015
	pesos_i(19079) := b"0000000000000000_0000000000000000_0000111011001111_1100110101111110"; -- 0.05785831757452986
	pesos_i(19080) := b"1111111111111111_1111111111111111_1111010001010011_1010000010111011"; -- -0.04559894022312108
	pesos_i(19081) := b"1111111111111111_1111111111111111_1110100100111100_1100111111010100"; -- -0.08891583507211542
	pesos_i(19082) := b"1111111111111111_1111111111111111_1110010100101000_1011110110110001"; -- -0.10484709188158747
	pesos_i(19083) := b"1111111111111111_1111111111111111_1110100011011000_0111100100111100"; -- -0.09044687532797621
	pesos_i(19084) := b"0000000000000000_0000000000000000_0001100100000010_0100111010100111"; -- 0.09769145563884417
	pesos_i(19085) := b"1111111111111111_1111111111111111_1110001111111101_0001011000010111"; -- -0.10941945963547106
	pesos_i(19086) := b"0000000000000000_0000000000000000_0000000001011110_0101100001001101"; -- 0.0014395892367548057
	pesos_i(19087) := b"1111111111111111_1111111111111111_1110111001011011_0010110110011111"; -- -0.06892123104153847
	pesos_i(19088) := b"0000000000000000_0000000000000000_0010001110001010_1100111011110111"; -- 0.13883679901230253
	pesos_i(19089) := b"1111111111111111_1111111111111111_1111010001111110_0101101001101000"; -- -0.04494700400707127
	pesos_i(19090) := b"1111111111111111_1111111111111111_1111100100111110_0011111010000101"; -- -0.026393978603624406
	pesos_i(19091) := b"0000000000000000_0000000000000000_0010011100101001_0101001001011001"; -- 0.15297426872383235
	pesos_i(19092) := b"0000000000000000_0000000000000000_0001011110101110_1001100001011111"; -- 0.0925078613793714
	pesos_i(19093) := b"1111111111111111_1111111111111111_1110000000010100_0110010100011110"; -- -0.1246887971257682
	pesos_i(19094) := b"1111111111111111_1111111111111111_1111110100010001_1101100101100011"; -- -0.011446393283389035
	pesos_i(19095) := b"1111111111111111_1111111111111111_1111000101111001_0111010010000000"; -- -0.05674049256749555
	pesos_i(19096) := b"0000000000000000_0000000000000000_0010011100001111_0010000110001011"; -- 0.1525746311065379
	pesos_i(19097) := b"0000000000000000_0000000000000000_0000001101000010_1101000011011111"; -- 0.012738279804630872
	pesos_i(19098) := b"0000000000000000_0000000000000000_0000000111101101_0001110011101010"; -- 0.007524306506589455
	pesos_i(19099) := b"1111111111111111_1111111111111111_1111111101111111_0010110101000001"; -- -0.001965686431531705
	pesos_i(19100) := b"1111111111111111_1111111111111111_1110001011010100_1000111101111110"; -- -0.11394408393773713
	pesos_i(19101) := b"1111111111111111_1111111111111111_1101110000110000_0101011111111101"; -- -0.13988733353068947
	pesos_i(19102) := b"0000000000000000_0000000000000000_0000010101001011_0100110111011111"; -- 0.02068030057187372
	pesos_i(19103) := b"1111111111111111_1111111111111111_1101001000110111_0111011101010010"; -- -0.17884115454325106
	pesos_i(19104) := b"0000000000000000_0000000000000000_0000010011101000_0001010011111110"; -- 0.01916629020607969
	pesos_i(19105) := b"1111111111111111_1111111111111111_1111100111000111_0011110000111001"; -- -0.02430366136793938
	pesos_i(19106) := b"1111111111111111_1111111111111111_1111001000001100_0011001010111011"; -- -0.05450137081938265
	pesos_i(19107) := b"1111111111111111_1111111111111111_1111001101110001_1101110011000101"; -- -0.049043847844642524
	pesos_i(19108) := b"1111111111111111_1111111111111111_1111010100001100_0100101110100100"; -- -0.042781135925081086
	pesos_i(19109) := b"1111111111111111_1111111111111111_1111100011111110_1010010111000101"; -- -0.027364387011304597
	pesos_i(19110) := b"1111111111111111_1111111111111111_1111000011001110_0011000000101100"; -- -0.05935381807108233
	pesos_i(19111) := b"0000000000000000_0000000000000000_0001110100111000_0100111111011001"; -- 0.11414050140282622
	pesos_i(19112) := b"1111111111111111_1111111111111111_1111111100101001_0010101001000000"; -- -0.0032781212944864207
	pesos_i(19113) := b"0000000000000000_0000000000000000_0001111011001110_1101110101000111"; -- 0.12034399964027682
	pesos_i(19114) := b"1111111111111111_1111111111111111_1101011001101010_0111010001101000"; -- -0.16243812989621387
	pesos_i(19115) := b"0000000000000000_0000000000000000_0001001011010011_1110010110000011"; -- 0.07354578454159505
	pesos_i(19116) := b"0000000000000000_0000000000000000_0000111001110000_1000100101101011"; -- 0.056404675172517564
	pesos_i(19117) := b"0000000000000000_0000000000000000_0000111001001111_0101101111101010"; -- 0.05589842278003892
	pesos_i(19118) := b"1111111111111111_1111111111111111_1110010000110101_1001011101001101"; -- -0.10855726585946636
	pesos_i(19119) := b"1111111111111111_1111111111111111_1111010111001101_0111111010110100"; -- -0.039833146196537675
	pesos_i(19120) := b"0000000000000000_0000000000000000_0001101101001010_0000110101010000"; -- 0.10659869388705526
	pesos_i(19121) := b"0000000000000000_0000000000000000_0001011111111000_0101010010001011"; -- 0.09363296873071529
	pesos_i(19122) := b"1111111111111111_1111111111111111_1111101100011111_0101110000100100"; -- -0.01905273557909136
	pesos_i(19123) := b"1111111111111111_1111111111111111_1111011010001110_1110001000000111"; -- -0.03688227963723173
	pesos_i(19124) := b"0000000000000000_0000000000000000_0000001101001000_1100100011011011"; -- 0.012829354632075579
	pesos_i(19125) := b"1111111111111111_1111111111111111_1101110110101101_1010000000001011"; -- -0.1340694402040511
	pesos_i(19126) := b"0000000000000000_0000000000000000_0001000100101100_1111001001010011"; -- 0.06709208032230173
	pesos_i(19127) := b"0000000000000000_0000000000000000_0001011101100100_0001011000011101"; -- 0.09137094694639249
	pesos_i(19128) := b"0000000000000000_0000000000000000_0000010010100110_1010100011111110"; -- 0.018168031625317247
	pesos_i(19129) := b"0000000000000000_0000000000000000_0000101111110100_0100100101111110"; -- 0.046696274945288954
	pesos_i(19130) := b"0000000000000000_0000000000000000_0000001001001101_0101110000101111"; -- 0.008992921302084858
	pesos_i(19131) := b"1111111111111111_1111111111111111_1110101001000011_1010001111100011"; -- -0.08490539281085888
	pesos_i(19132) := b"0000000000000000_0000000000000000_0001100011111101_1011001100001011"; -- 0.09762114536566173
	pesos_i(19133) := b"1111111111111111_1111111111111111_1110000001111000_0100001001000111"; -- -0.12316499480602314
	pesos_i(19134) := b"1111111111111111_1111111111111111_1111111110111000_0011011101101100"; -- -0.0010953294360485013
	pesos_i(19135) := b"0000000000000000_0000000000000000_0010101101011111_0000011011000110"; -- 0.1694187386059563
	pesos_i(19136) := b"0000000000000000_0000000000000000_0000011010101010_0111001011010100"; -- 0.02603833850605183
	pesos_i(19137) := b"0000000000000000_0000000000000000_0000111001011111_1001000100001100"; -- 0.05614573040394228
	pesos_i(19138) := b"0000000000000000_0000000000000000_0001101110011101_0011101011001011"; -- 0.10786788410956849
	pesos_i(19139) := b"0000000000000000_0000000000000000_0010000111101111_1100001101111011"; -- 0.13256475214153143
	pesos_i(19140) := b"1111111111111111_1111111111111111_1110001000001001_0010101000110001"; -- -0.11704765599913734
	pesos_i(19141) := b"0000000000000000_0000000000000000_0000000100100110_1101000110101001"; -- 0.004498580751055814
	pesos_i(19142) := b"1111111111111111_1111111111111111_1110101100001000_1111001101001011"; -- -0.08189467837828744
	pesos_i(19143) := b"1111111111111111_1111111111111111_1101011110001010_0011100010111100"; -- -0.15804715537240002
	pesos_i(19144) := b"1111111111111111_1111111111111111_1111101011111010_0101110011111110"; -- -0.019617259864596663
	pesos_i(19145) := b"1111111111111111_1111111111111111_1111100001010010_0010001000110010"; -- -0.02999674111153653
	pesos_i(19146) := b"0000000000000000_0000000000000000_0000011100100000_0010110010000110"; -- 0.027834684971385557
	pesos_i(19147) := b"0000000000000000_0000000000000000_0001110000101000_1011100000111101"; -- 0.10999633293480333
	pesos_i(19148) := b"0000000000000000_0000000000000000_0001000001101000_0110001111000111"; -- 0.06409286132072367
	pesos_i(19149) := b"0000000000000000_0000000000000000_0001101111001010_1001111011111011"; -- 0.10856050144449524
	pesos_i(19150) := b"1111111111111111_1111111111111111_1111001011001001_0110101100000010"; -- -0.05161410531742636
	pesos_i(19151) := b"1111111111111111_1111111111111111_1110101010011001_0010010011111101"; -- -0.08360070061151889
	pesos_i(19152) := b"1111111111111111_1111111111111111_1110110110000011_0101010000111101"; -- -0.0722148276547055
	pesos_i(19153) := b"1111111111111111_1111111111111111_1111010100000010_1101111100000110"; -- -0.04292493925766354
	pesos_i(19154) := b"1111111111111111_1111111111111111_1111101100001000_1001101110001101"; -- -0.019399908163188668
	pesos_i(19155) := b"0000000000000000_0000000000000000_0001110010010110_0011010100000110"; -- 0.11166697890409537
	pesos_i(19156) := b"1111111111111111_1111111111111111_1111100001000001_1101110100010011"; -- -0.030245001549520464
	pesos_i(19157) := b"1111111111111111_1111111111111111_1111101100100011_1010101101011011"; -- -0.018986978732342136
	pesos_i(19158) := b"1111111111111111_1111111111111111_1111101011111001_1110010010000011"; -- -0.019624441049445034
	pesos_i(19159) := b"0000000000000000_0000000000000000_0001110111111110_0000101101011101"; -- 0.11715765983338979
	pesos_i(19160) := b"1111111111111111_1111111111111111_1101101011110011_0011111010000111"; -- -0.144725887326542
	pesos_i(19161) := b"0000000000000000_0000000000000000_0010000001110011_1001111110011101"; -- 0.1267642744109965
	pesos_i(19162) := b"1111111111111111_1111111111111111_1111010011110000_1011100110011011"; -- -0.04320182774625158
	pesos_i(19163) := b"0000000000000000_0000000000000000_0001001001100011_0100110100001100"; -- 0.07182771243664098
	pesos_i(19164) := b"0000000000000000_0000000000000000_0001011011101001_1100000111101111"; -- 0.08950435726593524
	pesos_i(19165) := b"1111111111111111_1111111111111111_1111111111000011_1000001011011011"; -- -0.0009229866517536901
	pesos_i(19166) := b"0000000000000000_0000000000000000_0000011101101001_1110000000101101"; -- 0.02895928470314083
	pesos_i(19167) := b"0000000000000000_0000000000000000_0000101111000001_0100111100111011"; -- 0.04591841873144925
	pesos_i(19168) := b"1111111111111111_1111111111111111_1101101111111011_0101011010011011"; -- -0.1406961317961878
	pesos_i(19169) := b"1111111111111111_1111111111111111_1111011101101001_1011011111001100"; -- -0.033543122046428626
	pesos_i(19170) := b"1111111111111111_1111111111111111_1110000101111111_0011101100110101"; -- -0.11915235481995957
	pesos_i(19171) := b"0000000000000000_0000000000000000_0010001011111010_1001111110111010"; -- 0.13663671773393135
	pesos_i(19172) := b"1111111111111111_1111111111111111_1111001101010100_0010001001110100"; -- -0.049497458112679735
	pesos_i(19173) := b"0000000000000000_0000000000000000_0001111101101100_1010010001001100"; -- 0.12275149196332807
	pesos_i(19174) := b"1111111111111111_1111111111111111_1110101001000000_1011000111111111"; -- -0.0849503280713616
	pesos_i(19175) := b"1111111111111111_1111111111111111_1110100101101100_0000101010010011"; -- -0.08819517056195608
	pesos_i(19176) := b"0000000000000000_0000000000000000_0000111110101111_0001111010001011"; -- 0.06126585858835263
	pesos_i(19177) := b"0000000000000000_0000000000000000_0000101001010000_1001011100010110"; -- 0.040292208583931566
	pesos_i(19178) := b"1111111111111111_1111111111111111_1111110111101111_0000010000110001"; -- -0.008071649520790451
	pesos_i(19179) := b"0000000000000000_0000000000000000_0000110010011010_0110101111100100"; -- 0.04923128435828894
	pesos_i(19180) := b"1111111111111111_1111111111111111_1110110110001010_0001101011001010"; -- -0.07211144033011031
	pesos_i(19181) := b"0000000000000000_0000000000000000_0000011000010110_0000110000101100"; -- 0.02377391883326832
	pesos_i(19182) := b"1111111111111111_1111111111111111_1111101011010100_0100111001001011"; -- -0.020197969991425323
	pesos_i(19183) := b"0000000000000000_0000000000000000_0000011010100100_0001000000001010"; -- 0.025940897388720664
	pesos_i(19184) := b"1111111111111111_1111111111111111_1111101011100100_0100101011111000"; -- -0.01995402756122581
	pesos_i(19185) := b"0000000000000000_0000000000000000_0000011101001110_0100010101110110"; -- 0.028538075742828645
	pesos_i(19186) := b"0000000000000000_0000000000000000_0001111000100100_0010101001000110"; -- 0.11773933605076785
	pesos_i(19187) := b"0000000000000000_0000000000000000_0000010110011001_0010101011101110"; -- 0.021868403621745258
	pesos_i(19188) := b"0000000000000000_0000000000000000_0001111011001001_1100100010011111"; -- 0.12026647464575616
	pesos_i(19189) := b"1111111111111111_1111111111111111_1110011010010000_1110011100101001"; -- -0.0993514561590151
	pesos_i(19190) := b"0000000000000000_0000000000000000_0000001001101011_0000001101100000"; -- 0.009445391524463536
	pesos_i(19191) := b"1111111111111111_1111111111111111_1111100100000100_1010100000110010"; -- -0.027272689553684105
	pesos_i(19192) := b"1111111111111111_1111111111111111_1110001011110110_0000100101100111"; -- -0.11343327748248286
	pesos_i(19193) := b"1111111111111111_1111111111111111_1111100101100001_1000000001111111"; -- -0.025855988458575712
	pesos_i(19194) := b"1111111111111111_1111111111111111_1111101100100101_1110110110011000"; -- -0.018952513170212862
	pesos_i(19195) := b"0000000000000000_0000000000000000_0001100101100011_0110010110110001"; -- 0.09917293145209612
	pesos_i(19196) := b"0000000000000000_0000000000000000_0001001000111101_0011011011101100"; -- 0.07124655967999195
	pesos_i(19197) := b"1111111111111111_1111111111111111_1101100000100001_1011011100000100"; -- -0.15573555136784925
	pesos_i(19198) := b"0000000000000000_0000000000000000_0001001110110000_1010110111111011"; -- 0.0769146668752036
	pesos_i(19199) := b"1111111111111111_1111111111111111_1101111010010011_0010010110101110"; -- -0.1305672120806093
	pesos_i(19200) := b"1111111111111111_1111111111111111_1111001010000011_0001100010000001"; -- -0.052687138158434794
	pesos_i(19201) := b"0000000000000000_0000000000000000_0010010110100011_1111001111110011"; -- 0.14703297305213703
	pesos_i(19202) := b"1111111111111111_1111111111111111_1111110011101011_0000001101010111"; -- -0.012038985604838646
	pesos_i(19203) := b"0000000000000000_0000000000000000_0001000100111101_1111110010100110"; -- 0.06735209513070697
	pesos_i(19204) := b"1111111111111111_1111111111111111_1111110111011111_1010110111100001"; -- -0.008305676127147202
	pesos_i(19205) := b"0000000000000000_0000000000000000_0001110101110001_0110100000100111"; -- 0.11501170112479842
	pesos_i(19206) := b"0000000000000000_0000000000000000_0001001010101100_1010011101011011"; -- 0.07294698683501694
	pesos_i(19207) := b"0000000000000000_0000000000000000_0001011011110111_1011001001000001"; -- 0.08971704576465696
	pesos_i(19208) := b"1111111111111111_1111111111111111_1110010000000100_0111010001111111"; -- -0.10930702116286713
	pesos_i(19209) := b"1111111111111111_1111111111111111_1101111110101110_0110111101001011"; -- -0.12624458712616995
	pesos_i(19210) := b"1111111111111111_1111111111111111_1110111001001011_0100010110100111"; -- -0.06916393922168679
	pesos_i(19211) := b"1111111111111111_1111111111111111_1111110100001100_1101110011001000"; -- -0.011522484916542695
	pesos_i(19212) := b"1111111111111111_1111111111111111_1101111011110111_1110100111111000"; -- -0.12902963349723873
	pesos_i(19213) := b"0000000000000000_0000000000000000_0000010001001110_0101001001111100"; -- 0.01682010192043664
	pesos_i(19214) := b"0000000000000000_0000000000000000_0000101111100110_0111010001101001"; -- 0.04648520995419936
	pesos_i(19215) := b"1111111111111111_1111111111111111_1110111101111101_1110110001101110"; -- -0.06448480905619582
	pesos_i(19216) := b"0000000000000000_0000000000000000_0000100101110101_0010001001010111"; -- 0.03694357507403363
	pesos_i(19217) := b"0000000000000000_0000000000000000_0000101010011111_1001111100011000"; -- 0.04149813027375175
	pesos_i(19218) := b"1111111111111111_1111111111111111_1111101100010111_1011100001100000"; -- -0.01916930817077149
	pesos_i(19219) := b"1111111111111111_1111111111111111_1110101111110101_0010001000000000"; -- -0.07829082013515808
	pesos_i(19220) := b"0000000000000000_0000000000000000_0001100011101010_1000000100101010"; -- 0.0973282554371552
	pesos_i(19221) := b"0000000000000000_0000000000000000_0001110000010001_1110010100010000"; -- 0.10964805257924184
	pesos_i(19222) := b"1111111111111111_1111111111111111_1111000000000010_1110011000111001"; -- -0.06245576004113259
	pesos_i(19223) := b"0000000000000000_0000000000000000_0010010011101001_1000101001101011"; -- 0.14418854817815002
	pesos_i(19224) := b"1111111111111111_1111111111111111_1110110110110011_1000110101000101"; -- -0.0714790064708805
	pesos_i(19225) := b"1111111111111111_1111111111111111_1111100110101111_1110110111010111"; -- -0.024659285617484768
	pesos_i(19226) := b"1111111111111111_1111111111111111_1111010110010101_0110101001100010"; -- -0.04068884959084693
	pesos_i(19227) := b"0000000000000000_0000000000000000_0010010100001100_0101110001111000"; -- 0.14471986703876616
	pesos_i(19228) := b"0000000000000000_0000000000000000_0001110101110100_1101011111010001"; -- 0.11506413310129199
	pesos_i(19229) := b"0000000000000000_0000000000000000_0001100111000011_1011110010111001"; -- 0.10064296268992894
	pesos_i(19230) := b"1111111111111111_1111111111111111_1101110000110010_0010100101100001"; -- -0.13985959420007488
	pesos_i(19231) := b"1111111111111111_1111111111111111_1110011011011100_0001010010110110"; -- -0.09820433189111871
	pesos_i(19232) := b"0000000000000000_0000000000000000_0001110000000110_1011101001000110"; -- 0.1094776554239694
	pesos_i(19233) := b"0000000000000000_0000000000000000_0010011110000111_1011100101100111"; -- 0.1544147373460263
	pesos_i(19234) := b"0000000000000000_0000000000000000_0001011011100101_1100001100100101"; -- 0.08944339419158888
	pesos_i(19235) := b"1111111111111111_1111111111111111_1111110100110100_0010010010001110"; -- -0.0109231140680382
	pesos_i(19236) := b"1111111111111111_1111111111111111_1110001101011110_1010111100111000"; -- -0.11183648005222686
	pesos_i(19237) := b"1111111111111111_1111111111111111_1111110100101000_1110101001101000"; -- -0.011094426759285165
	pesos_i(19238) := b"1111111111111111_1111111111111111_1111100011011110_1110011001101100"; -- -0.0278488145745748
	pesos_i(19239) := b"0000000000000000_0000000000000000_0001010010011100_0000101011000110"; -- 0.08050601321798598
	pesos_i(19240) := b"1111111111111111_1111111111111111_1110000100111001_1010111100000111"; -- -0.12021356654601119
	pesos_i(19241) := b"0000000000000000_0000000000000000_0000000110100011_0001000110101010"; -- 0.0063944855882618
	pesos_i(19242) := b"1111111111111111_1111111111111111_1111111101011101_1010110101000110"; -- -0.0024768547473351253
	pesos_i(19243) := b"0000000000000000_0000000000000000_0000010101011100_1111100011000111"; -- 0.020949886866320554
	pesos_i(19244) := b"0000000000000000_0000000000000000_0000101000000000_1100010011001011"; -- 0.03907422970366109
	pesos_i(19245) := b"1111111111111111_1111111111111111_1110010011010001_1001100000101001"; -- -0.10617684366903536
	pesos_i(19246) := b"1111111111111111_1111111111111111_1101111011011110_0101010010100001"; -- -0.12942000455990907
	pesos_i(19247) := b"0000000000000000_0000000000000000_0001100100100001_0000100011000111"; -- 0.09816031313312795
	pesos_i(19248) := b"0000000000000000_0000000000000000_0000001100011011_1011101101001110"; -- 0.012141901574741341
	pesos_i(19249) := b"0000000000000000_0000000000000000_0001110000100110_0111110101000010"; -- 0.10996229993985328
	pesos_i(19250) := b"0000000000000000_0000000000000000_0000010010110000_1110111111101001"; -- 0.018324846648523168
	pesos_i(19251) := b"1111111111111111_1111111111111111_1111000000101011_1001101111011000"; -- -0.06183458310343271
	pesos_i(19252) := b"1111111111111111_1111111111111111_1101100011110010_0110000101101001"; -- -0.15255156695938563
	pesos_i(19253) := b"0000000000000000_0000000000000000_0000000010111101_1001101010000010"; -- 0.0028931205830683444
	pesos_i(19254) := b"1111111111111111_1111111111111111_1101111100011001_0001110000011100"; -- -0.128523104881904
	pesos_i(19255) := b"0000000000000000_0000000000000000_0000111001011101_1101010010001110"; -- 0.05611923662874553
	pesos_i(19256) := b"1111111111111111_1111111111111111_1110110101110100_0111010001111101"; -- -0.07244178713701827
	pesos_i(19257) := b"1111111111111111_1111111111111111_1111000010110101_0100011101111111"; -- -0.05973389771651917
	pesos_i(19258) := b"1111111111111111_1111111111111111_1111111110111001_0111101010010010"; -- -0.001076068164591545
	pesos_i(19259) := b"0000000000000000_0000000000000000_0000111000011111_1100111010101001"; -- 0.05517284036312007
	pesos_i(19260) := b"0000000000000000_0000000000000000_0010001101110001_0111011010011010"; -- 0.13845006228112208
	pesos_i(19261) := b"0000000000000000_0000000000000000_0001100110101011_1010111011111101"; -- 0.10027593311071212
	pesos_i(19262) := b"0000000000000000_0000000000000000_0000100000101000_0010111000011101"; -- 0.03186310002059333
	pesos_i(19263) := b"1111111111111111_1111111111111111_1111100001010111_1011000100011101"; -- -0.029911928542820952
	pesos_i(19264) := b"0000000000000000_0000000000000000_0001000011010011_0010000110010010"; -- 0.0657216053620883
	pesos_i(19265) := b"1111111111111111_1111111111111111_1111110011001010_0100111110111101"; -- -0.012537971947772278
	pesos_i(19266) := b"0000000000000000_0000000000000000_0001010110001011_1011101101110111"; -- 0.08416339555810472
	pesos_i(19267) := b"0000000000000000_0000000000000000_0000001110111100_1101010110010011"; -- 0.01460013225060039
	pesos_i(19268) := b"0000000000000000_0000000000000000_0001110100111000_0010011000011001"; -- 0.11413801302849254
	pesos_i(19269) := b"1111111111111111_1111111111111111_1110101001101010_1110000010010100"; -- -0.08430668250582465
	pesos_i(19270) := b"1111111111111111_1111111111111111_1101111011111001_1111010100000110"; -- -0.12899845693243064
	pesos_i(19271) := b"1111111111111111_1111111111111111_1110010111100100_0100001011111110"; -- -0.10198575302369206
	pesos_i(19272) := b"0000000000000000_0000000000000000_0001101000001100_0011011111000000"; -- 0.10174892836427289
	pesos_i(19273) := b"0000000000000000_0000000000000000_0001010101000001_1000111011011101"; -- 0.08303158667531073
	pesos_i(19274) := b"1111111111111111_1111111111111111_1111101100010001_0111111110010011"; -- -0.019264246663619606
	pesos_i(19275) := b"0000000000000000_0000000000000000_0001101011101110_1000011110111101"; -- 0.10520218239178171
	pesos_i(19276) := b"0000000000000000_0000000000000000_0001000100111110_1001110101100101"; -- 0.06736167640911012
	pesos_i(19277) := b"1111111111111111_1111111111111111_1110100101111011_1000010111111011"; -- -0.08795893316882594
	pesos_i(19278) := b"0000000000000000_0000000000000000_0000010100011100_1011011001011110"; -- 0.01996936596168062
	pesos_i(19279) := b"0000000000000000_0000000000000000_0000111011000000_1000000110001011"; -- 0.05762490894134323
	pesos_i(19280) := b"1111111111111111_1111111111111111_1101111011111010_1111011000000000"; -- -0.12898313988852012
	pesos_i(19281) := b"0000000000000000_0000000000000000_0010001111001100_0101011011000000"; -- 0.139836713696244
	pesos_i(19282) := b"0000000000000000_0000000000000000_0001110100101001_0000101100011111"; -- 0.11390752319756851
	pesos_i(19283) := b"0000000000000000_0000000000000000_0001101001010011_1011111011111110"; -- 0.10284036353689271
	pesos_i(19284) := b"0000000000000000_0000000000000000_0010000000110011_0100111111000000"; -- 0.12578295182846072
	pesos_i(19285) := b"0000000000000000_0000000000000000_0000100110100011_1000111011010010"; -- 0.03765194545769081
	pesos_i(19286) := b"0000000000000000_0000000000000000_0000010110110111_0111010010010100"; -- 0.022330556916986675
	pesos_i(19287) := b"1111111111111111_1111111111111111_1110110111001010_0011000101010010"; -- -0.07113353489587922
	pesos_i(19288) := b"0000000000000000_0000000000000000_0000010111101010_0101011110110111"; -- 0.02310703490399205
	pesos_i(19289) := b"1111111111111111_1111111111111111_1101011111011000_1010111000111110"; -- -0.15684996584616656
	pesos_i(19290) := b"1111111111111111_1111111111111111_1110011100111101_0110110110011011"; -- -0.09671893079451065
	pesos_i(19291) := b"0000000000000000_0000000000000000_0000000010101110_1010001011001010"; -- 0.0026647323675710716
	pesos_i(19292) := b"1111111111111111_1111111111111111_1111000000111010_0110110111010001"; -- -0.06160844456082941
	pesos_i(19293) := b"1111111111111111_1111111111111111_1111000000111110_0101011001011100"; -- -0.06154880756082779
	pesos_i(19294) := b"0000000000000000_0000000000000000_0001010001000101_1000001000110110"; -- 0.07918561755910283
	pesos_i(19295) := b"1111111111111111_1111111111111111_1110010100010010_1000010010101110"; -- -0.10518618352239474
	pesos_i(19296) := b"1111111111111111_1111111111111111_1111011100101101_0101101000000111"; -- -0.03446423834525009
	pesos_i(19297) := b"1111111111111111_1111111111111111_1111110010111101_0101000111000011"; -- -0.012736215449201244
	pesos_i(19298) := b"0000000000000000_0000000000000000_0001011011010101_0010101110100111"; -- 0.0891902240642432
	pesos_i(19299) := b"1111111111111111_1111111111111111_1111010010100111_0011110110111111"; -- -0.04432310180422742
	pesos_i(19300) := b"1111111111111111_1111111111111111_1110110100110100_0001000000100111"; -- -0.07342433018471083
	pesos_i(19301) := b"0000000000000000_0000000000000000_0000010010101001_1011110110111100"; -- 0.018215044482712488
	pesos_i(19302) := b"0000000000000000_0000000000000000_0010011010101101_1000011010001110"; -- 0.151085290637992
	pesos_i(19303) := b"0000000000000000_0000000000000000_0000010011110110_0111111111111101"; -- 0.019386290874414992
	pesos_i(19304) := b"0000000000000000_0000000000000000_0001001010000110_0001101001100001"; -- 0.07235875010381708
	pesos_i(19305) := b"1111111111111111_1111111111111111_1111110000111011_1111011010000011"; -- -0.014710038193489752
	pesos_i(19306) := b"1111111111111111_1111111111111111_1110000100101001_1000101010011000"; -- -0.12045987885202747
	pesos_i(19307) := b"0000000000000000_0000000000000000_0010000110001111_0110011011101011"; -- 0.13109439126020278
	pesos_i(19308) := b"0000000000000000_0000000000000000_0001011110101000_1001000011010110"; -- 0.0924158594635279
	pesos_i(19309) := b"1111111111111111_1111111111111111_1101111111001000_0010110110001101"; -- -0.1258517772622121
	pesos_i(19310) := b"1111111111111111_1111111111111111_1101110111011011_0101011001010100"; -- -0.13337192974583278
	pesos_i(19311) := b"1111111111111111_1111111111111111_1111110101000001_1010111101101000"; -- -0.010716473665248688
	pesos_i(19312) := b"1111111111111111_1111111111111111_1111000100101011_0010011000110111"; -- -0.05793534434184688
	pesos_i(19313) := b"1111111111111111_1111111111111111_1101110101111001_1000001101110011"; -- -0.13486460146582274
	pesos_i(19314) := b"0000000000000000_0000000000000000_0000110011000000_0111110101101111"; -- 0.049812163963188286
	pesos_i(19315) := b"0000000000000000_0000000000000000_0001010000000111_1011000000101000"; -- 0.07824231133636339
	pesos_i(19316) := b"0000000000000000_0000000000000000_0000011000111000_1101011010101000"; -- 0.024304786779160863
	pesos_i(19317) := b"1111111111111111_1111111111111111_1101111011110011_1100110001100110"; -- -0.12909243114198987
	pesos_i(19318) := b"1111111111111111_1111111111111111_1110101001101010_0011001001110110"; -- -0.08431706059531598
	pesos_i(19319) := b"1111111111111111_1111111111111111_1101101010011110_1011000110010100"; -- -0.14601602682224996
	pesos_i(19320) := b"1111111111111111_1111111111111111_1111010100000110_1011101110001110"; -- -0.0428660181970962
	pesos_i(19321) := b"1111111111111111_1111111111111111_1111000101111011_0101000001010000"; -- -0.05671213184964322
	pesos_i(19322) := b"1111111111111111_1111111111111111_1110001100100010_0111110000011010"; -- -0.11275505407353119
	pesos_i(19323) := b"0000000000000000_0000000000000000_0001101010101010_0100101110111110"; -- 0.10416100884306465
	pesos_i(19324) := b"1111111111111111_1111111111111111_1111111100000100_0000100111111101"; -- -0.003844619539777145
	pesos_i(19325) := b"0000000000000000_0000000000000000_0001111010110001_0001111101110010"; -- 0.11989017989632263
	pesos_i(19326) := b"1111111111111111_1111111111111111_1111110110101100_0010010011100000"; -- -0.009092040457483188
	pesos_i(19327) := b"0000000000000000_0000000000000000_0000001110010111_0010000101101011"; -- 0.014024819089799365
	pesos_i(19328) := b"0000000000000000_0000000000000000_0000100000010011_0111111011000000"; -- 0.03154747196541981
	pesos_i(19329) := b"0000000000000000_0000000000000000_0001011110111000_0011000010110001"; -- 0.09265426945804821
	pesos_i(19330) := b"1111111111111111_1111111111111111_1111100010010100_0000000101000010"; -- -0.028991624144706567
	pesos_i(19331) := b"1111111111111111_1111111111111111_1101101111110000_1100010010010001"; -- -0.14085742430345563
	pesos_i(19332) := b"1111111111111111_1111111111111111_1110010000110101_1011111000100111"; -- -0.10855495023757247
	pesos_i(19333) := b"0000000000000000_0000000000000000_0000000110011001_0000111100101111"; -- 0.0062417497577303424
	pesos_i(19334) := b"1111111111111111_1111111111111111_1101010111010000_0000010000011010"; -- -0.1647946774590684
	pesos_i(19335) := b"1111111111111111_1111111111111111_1111101110110100_1100110000010110"; -- -0.016772503416253044
	pesos_i(19336) := b"1111111111111111_1111111111111111_1110011011101101_0010110100001101"; -- -0.09794348176238789
	pesos_i(19337) := b"1111111111111111_1111111111111111_1111110100011100_1110011110000100"; -- -0.01127770444277919
	pesos_i(19338) := b"0000000000000000_0000000000000000_0001001110110100_1001010011111110"; -- 0.0769742126855437
	pesos_i(19339) := b"1111111111111111_1111111111111111_1111011011100101_0110110111000101"; -- -0.03556169443044933
	pesos_i(19340) := b"1111111111111111_1111111111111111_1110010110011001_0101101011000011"; -- -0.10312874537312963
	pesos_i(19341) := b"1111111111111111_1111111111111111_1110000010110101_0010010000100111"; -- -0.12223600435912975
	pesos_i(19342) := b"1111111111111111_1111111111111111_1110110111111011_0010000001100001"; -- -0.0703868640493077
	pesos_i(19343) := b"0000000000000000_0000000000000000_0010010010001011_0101110010011010"; -- 0.14275149125348366
	pesos_i(19344) := b"1111111111111111_1111111111111111_1110111010000001_0111111110101111"; -- -0.06833650563060538
	pesos_i(19345) := b"0000000000000000_0000000000000000_0000111101101000_1110000101111010"; -- 0.060194103409859694
	pesos_i(19346) := b"0000000000000000_0000000000000000_0010000011110111_1000000011110011"; -- 0.12877660694144494
	pesos_i(19347) := b"1111111111111111_1111111111111111_1111101100100110_1100100100101111"; -- -0.018939424556336733
	pesos_i(19348) := b"1111111111111111_1111111111111111_1101111011000110_1011011101011111"; -- -0.12978033010546378
	pesos_i(19349) := b"1111111111111111_1111111111111111_1110011100000111_0001101011110100"; -- -0.09754783200168182
	pesos_i(19350) := b"0000000000000000_0000000000000000_0001000000010100_0101000101110001"; -- 0.06281003016341485
	pesos_i(19351) := b"1111111111111111_1111111111111111_1111111111111111_0011100110011101"; -- -1.1824712306824807e-05
	pesos_i(19352) := b"0000000000000000_0000000000000000_0001101001001101_1010011110101000"; -- 0.10274741992402191
	pesos_i(19353) := b"0000000000000000_0000000000000000_0000101101010111_1001111101001011"; -- 0.04430575916802075
	pesos_i(19354) := b"1111111111111111_1111111111111111_1101101011011101_0000100011010010"; -- -0.14506478186289176
	pesos_i(19355) := b"0000000000000000_0000000000000000_0000110110100010_0100001110011110"; -- 0.053257204213636854
	pesos_i(19356) := b"1111111111111111_1111111111111111_1111111000110101_1011011101011110"; -- -0.006992854590568123
	pesos_i(19357) := b"1111111111111111_1111111111111111_1110100001111000_1111110111001110"; -- -0.09190381736581808
	pesos_i(19358) := b"1111111111111111_1111111111111111_1110111111111000_0111010111011000"; -- -0.06261504628984761
	pesos_i(19359) := b"0000000000000000_0000000000000000_0000011000110000_0000110011111000"; -- 0.02417069480646635
	pesos_i(19360) := b"1111111111111111_1111111111111111_1111001101000101_0010110110010010"; -- -0.049725677342093204
	pesos_i(19361) := b"1111111111111111_1111111111111111_1110101000000100_0010000111011011"; -- -0.0858744469228477
	pesos_i(19362) := b"0000000000000000_0000000000000000_0001110001000000_1110010001011110"; -- 0.11036517435111592
	pesos_i(19363) := b"0000000000000000_0000000000000000_0001011101001011_0101001001101010"; -- 0.09099307149729978
	pesos_i(19364) := b"1111111111111111_1111111111111111_1111111110101000_0110111010010001"; -- -0.0013361832676087929
	pesos_i(19365) := b"0000000000000000_0000000000000000_0001111000000000_1010110101111000"; -- 0.11719783945167693
	pesos_i(19366) := b"1111111111111111_1111111111111111_1111111010111011_1011010101000011"; -- -0.004948302441580564
	pesos_i(19367) := b"0000000000000000_0000000000000000_0001001100100111_1110001110000101"; -- 0.07482740392970931
	pesos_i(19368) := b"1111111111111111_1111111111111111_1110010010010111_1000110101100000"; -- -0.10706249620550284
	pesos_i(19369) := b"0000000000000000_0000000000000000_0010011000000100_1111101000000001"; -- 0.14851343662520702
	pesos_i(19370) := b"1111111111111111_1111111111111111_1101110111011010_0001011011011110"; -- -0.13339097102833464
	pesos_i(19371) := b"0000000000000000_0000000000000000_0001101101000010_1001110110001011"; -- 0.10648522037010683
	pesos_i(19372) := b"1111111111111111_1111111111111111_1111111100000100_0111101101001110"; -- -0.0038378652208860306
	pesos_i(19373) := b"1111111111111111_1111111111111111_1110110000010100_1000000011100111"; -- -0.07781214115102505
	pesos_i(19374) := b"1111111111111111_1111111111111111_1111101100000110_1000010101001101"; -- -0.019431752031585953
	pesos_i(19375) := b"0000000000000000_0000000000000000_0010001110001011_1001010100001010"; -- 0.13884860512375097
	pesos_i(19376) := b"1111111111111111_1111111111111111_1110001111101100_1010110010110000"; -- -0.10966988284140243
	pesos_i(19377) := b"0000000000000000_0000000000000000_0000111000001101_1100001010100111"; -- 0.05489746654363421
	pesos_i(19378) := b"0000000000000000_0000000000000000_0000011101011100_1110110000010010"; -- 0.028761629397119796
	pesos_i(19379) := b"1111111111111111_1111111111111111_1101111110111110_1100010011011100"; -- -0.12599534640958565
	pesos_i(19380) := b"0000000000000000_0000000000000000_0010001101111011_0001011001001111"; -- 0.13859691068521476
	pesos_i(19381) := b"0000000000000000_0000000000000000_0000010000001000_1101000010001100"; -- 0.01575950062403514
	pesos_i(19382) := b"1111111111111111_1111111111111111_1101111010000000_0110011001001111"; -- -0.1308532768280223
	pesos_i(19383) := b"0000000000000000_0000000000000000_0001101000110001_1001111000101101"; -- 0.10231960875600078
	pesos_i(19384) := b"1111111111111111_1111111111111111_1101111001100100_0100001001101110"; -- -0.13128266158973134
	pesos_i(19385) := b"1111111111111111_1111111111111111_1110101110110100_0101000001001101"; -- -0.07927988173243815
	pesos_i(19386) := b"0000000000000000_0000000000000000_0000101101110001_0110001001010101"; -- 0.044698854144803304
	pesos_i(19387) := b"1111111111111111_1111111111111111_1101101001001100_1010000011011010"; -- -0.14726824445017064
	pesos_i(19388) := b"0000000000000000_0000000000000000_0010010111100011_0001011010101110"; -- 0.14799634682649246
	pesos_i(19389) := b"1111111111111111_1111111111111111_1110100111100100_1000001001100011"; -- -0.08635697441089832
	pesos_i(19390) := b"1111111111111111_1111111111111111_1101101111001110_1111111000011110"; -- -0.1413727928995251
	pesos_i(19391) := b"1111111111111111_1111111111111111_1111000100011001_0011011100111001"; -- -0.058208988783435466
	pesos_i(19392) := b"0000000000000000_0000000000000000_0010001100100010_0000000101001111"; -- 0.13723762690310562
	pesos_i(19393) := b"0000000000000000_0000000000000000_0001101010100000_0111010010011001"; -- 0.1040108561237433
	pesos_i(19394) := b"0000000000000000_0000000000000000_0000011011011110_0110010010010000"; -- 0.026830945243973805
	pesos_i(19395) := b"1111111111111111_1111111111111111_1111000001010000_1011101111001000"; -- -0.0612681043099247
	pesos_i(19396) := b"0000000000000000_0000000000000000_0000011111101110_0010110110011110"; -- 0.030978060844887807
	pesos_i(19397) := b"0000000000000000_0000000000000000_0001110001100000_0011110110101100"; -- 0.11084351978372868
	pesos_i(19398) := b"0000000000000000_0000000000000000_0010001111101110_1010011001101000"; -- 0.14036026028464718
	pesos_i(19399) := b"1111111111111111_1111111111111111_1111101010001100_1110111110110010"; -- -0.021286982674778496
	pesos_i(19400) := b"1111111111111111_1111111111111111_1111111101010010_0001101110110111"; -- -0.0026533774218687523
	pesos_i(19401) := b"0000000000000000_0000000000000000_0010011010100000_0011110010101011"; -- 0.15088252238826352
	pesos_i(19402) := b"0000000000000000_0000000000000000_0001101111111010_0010000001110011"; -- 0.10928538134168686
	pesos_i(19403) := b"0000000000000000_0000000000000000_0010001100011110_1100111011001011"; -- 0.13718883955939873
	pesos_i(19404) := b"0000000000000000_0000000000000000_0000000110111001_0110011010001111"; -- 0.0067352389981345144
	pesos_i(19405) := b"1111111111111111_1111111111111111_1111010110001101_1001100100101100"; -- -0.040808130987574145
	pesos_i(19406) := b"1111111111111111_1111111111111111_1111010001111101_1111100110111100"; -- -0.04495276598684442
	pesos_i(19407) := b"1111111111111111_1111111111111111_1111111011010110_1011111101111111"; -- -0.004535705139742464
	pesos_i(19408) := b"1111111111111111_1111111111111111_1111101010110010_0111101000100000"; -- -0.020714156397780122
	pesos_i(19409) := b"1111111111111111_1111111111111111_1111000010000100_0100110011111101"; -- -0.06048125099609335
	pesos_i(19410) := b"0000000000000000_0000000000000000_0001101111111011_1001000010001110"; -- 0.10930732216279031
	pesos_i(19411) := b"1111111111111111_1111111111111111_1110000111110101_1001000110011010"; -- -0.1173466681673868
	pesos_i(19412) := b"1111111111111111_1111111111111111_1110110000100001_1110111011010011"; -- -0.07760722495788759
	pesos_i(19413) := b"1111111111111111_1111111111111111_1110011110110011_1011011001010110"; -- -0.0949140587844185
	pesos_i(19414) := b"0000000000000000_0000000000000000_0001011000101000_0100111011000110"; -- 0.08655254676591909
	pesos_i(19415) := b"0000000000000000_0000000000000000_0000010001110110_0101101000101000"; -- 0.01743091084700059
	pesos_i(19416) := b"0000000000000000_0000000000000000_0001111010011110_1001100110001010"; -- 0.11960754034056598
	pesos_i(19417) := b"1111111111111111_1111111111111111_1111101101101010_1111111000111111"; -- -0.01789866405124067
	pesos_i(19418) := b"1111111111111111_1111111111111111_1110011000100110_1100101000000011"; -- -0.1009706251652895
	pesos_i(19419) := b"1111111111111111_1111111111111111_1110110111011000_1100011001011110"; -- -0.070911027855097
	pesos_i(19420) := b"1111111111111111_1111111111111111_1110100010101110_1011001011001010"; -- -0.09108431401550635
	pesos_i(19421) := b"0000000000000000_0000000000000000_0010001110010010_0101100011001000"; -- 0.13895182497098182
	pesos_i(19422) := b"1111111111111111_1111111111111111_1110100011010110_1110010001001001"; -- -0.09047101231399071
	pesos_i(19423) := b"0000000000000000_0000000000000000_0001000100011101_0000010110011110"; -- 0.06684908979793934
	pesos_i(19424) := b"1111111111111111_1111111111111111_1110101000101101_1101000110010011"; -- -0.08523836299644139
	pesos_i(19425) := b"0000000000000000_0000000000000000_0000010110001101_1001110101111111"; -- 0.021692126751549436
	pesos_i(19426) := b"0000000000000000_0000000000000000_0000110011111100_0110010001001010"; -- 0.05072619261420444
	pesos_i(19427) := b"1111111111111111_1111111111111111_1101111000000101_1000011101110011"; -- -0.13272813274981107
	pesos_i(19428) := b"0000000000000000_0000000000000000_0001101100010001_0111100100101101"; -- 0.10573537203325128
	pesos_i(19429) := b"0000000000000000_0000000000000000_0001110011000111_0111110010001001"; -- 0.11241892195465866
	pesos_i(19430) := b"1111111111111111_1111111111111111_1110010101100010_1011001111000111"; -- -0.1039626730845835
	pesos_i(19431) := b"1111111111111111_1111111111111111_1101101110000110_0011110001010011"; -- -0.1424829767010306
	pesos_i(19432) := b"0000000000000000_0000000000000000_0010001100011100_0111000000111000"; -- 0.13715268495238378
	pesos_i(19433) := b"0000000000000000_0000000000000000_0000010110111111_1001011010111001"; -- 0.022454662487099614
	pesos_i(19434) := b"0000000000000000_0000000000000000_0001100101000111_1101100000010010"; -- 0.09875250276767294
	pesos_i(19435) := b"0000000000000000_0000000000000000_0001111011111011_1101100001010100"; -- 0.12103035012246859
	pesos_i(19436) := b"0000000000000000_0000000000000000_0001100110110011_1000010101110101"; -- 0.10039552779808233
	pesos_i(19437) := b"0000000000000000_0000000000000000_0000111110011001_1011001010010100"; -- 0.06093898872408669
	pesos_i(19438) := b"0000000000000000_0000000000000000_0000010001101100_0110110011100010"; -- 0.017279439166584542
	pesos_i(19439) := b"0000000000000000_0000000000000000_0001011010001100_0011010010010010"; -- 0.08807686387168269
	pesos_i(19440) := b"1111111111111111_1111111111111111_1111100111001011_1100111100100111"; -- -0.024233868472370572
	pesos_i(19441) := b"0000000000000000_0000000000000000_0010000101101011_0111111000101001"; -- 0.13054646011225027
	pesos_i(19442) := b"0000000000000000_0000000000000000_0000101000001000_1010100110111110"; -- 0.03919468766327067
	pesos_i(19443) := b"0000000000000000_0000000000000000_0001011000010111_0000000011001001"; -- 0.08628849900738099
	pesos_i(19444) := b"1111111111111111_1111111111111111_1110010000000001_0111010001000010"; -- -0.10935281159073719
	pesos_i(19445) := b"1111111111111111_1111111111111111_1111001100000101_1000101111000101"; -- -0.05069662506007434
	pesos_i(19446) := b"1111111111111111_1111111111111111_1101011111000000_1111111110000001"; -- -0.1572113332123111
	pesos_i(19447) := b"1111111111111111_1111111111111111_1111001000010111_1101010011011011"; -- -0.05432386056466776
	pesos_i(19448) := b"1111111111111111_1111111111111111_1110010111110110_0110011101100110"; -- -0.1017089248985707
	pesos_i(19449) := b"1111111111111111_1111111111111111_1111010110111110_1111011000110110"; -- -0.040054904788900954
	pesos_i(19450) := b"0000000000000000_0000000000000000_0000100111000110_1011010111100010"; -- 0.03818833137208089
	pesos_i(19451) := b"1111111111111111_1111111111111111_1111110111100100_1011010010111001"; -- -0.008228974241628608
	pesos_i(19452) := b"1111111111111111_1111111111111111_1111110011001011_1011100001111111"; -- -0.012516469075326225
	pesos_i(19453) := b"1111111111111111_1111111111111111_1101110010101101_1101011101101100"; -- -0.13797238929683225
	pesos_i(19454) := b"1111111111111111_1111111111111111_1101100001010011_1000101101010001"; -- -0.15497521656551314
	pesos_i(19455) := b"0000000000000000_0000000000000000_0000011001111100_0001000000000101"; -- 0.025330544612175748
	pesos_i(19456) := b"0000000000000000_0000000000000000_0001010011011111_0011011001111110"; -- 0.08153095802965271
	pesos_i(19457) := b"1111111111111111_1111111111111111_1110001011001100_0000011101000000"; -- -0.11407427485669115
	pesos_i(19458) := b"1111111111111111_1111111111111111_1110111111110101_1001001111011110"; -- -0.06265903321715452
	pesos_i(19459) := b"1111111111111111_1111111111111111_1111101011001101_1100011101101101"; -- -0.020297561536748374
	pesos_i(19460) := b"1111111111111111_1111111111111111_1101100000011011_1111101000011001"; -- -0.15582310578265743
	pesos_i(19461) := b"1111111111111111_1111111111111111_1111001000001111_1011101010001101"; -- -0.05444749890808099
	pesos_i(19462) := b"0000000000000000_0000000000000000_0001001000010011_0101101010000100"; -- 0.07060781223295173
	pesos_i(19463) := b"0000000000000000_0000000000000000_0001010110010010_1110001001000100"; -- 0.08427251959580126
	pesos_i(19464) := b"1111111111111111_1111111111111111_1110100000011110_0110000000001001"; -- -0.09328651214409583
	pesos_i(19465) := b"1111111111111111_1111111111111111_1111110000011100_0001100001111001"; -- -0.015196295289370956
	pesos_i(19466) := b"1111111111111111_1111111111111111_1110010010100110_1100111100011111"; -- -0.1068296955374813
	pesos_i(19467) := b"1111111111111111_1111111111111111_1111111111000101_1000111010001011"; -- -0.0008917722774172708
	pesos_i(19468) := b"1111111111111111_1111111111111111_1111100111000000_0001110000010110"; -- -0.024412388415514668
	pesos_i(19469) := b"1111111111111111_1111111111111111_1111011001100010_1101010111000111"; -- -0.037554396530188154
	pesos_i(19470) := b"0000000000000000_0000000000000000_0001101010101110_0010111011101110"; -- 0.10422032643176629
	pesos_i(19471) := b"1111111111111111_1111111111111111_1111001110000110_1100110011110011"; -- -0.04872435626470724
	pesos_i(19472) := b"0000000000000000_0000000000000000_0000000101011000_0001100010100111"; -- 0.005250492845885978
	pesos_i(19473) := b"0000000000000000_0000000000000000_0010001011110011_1100001111000110"; -- 0.13653205467373591
	pesos_i(19474) := b"1111111111111111_1111111111111111_1101110001010011_0000100101100011"; -- -0.13935796094688907
	pesos_i(19475) := b"0000000000000000_0000000000000000_0001111100111010_1011100101001000"; -- 0.12198980340606042
	pesos_i(19476) := b"1111111111111111_1111111111111111_1110101000100010_1010101110110010"; -- -0.08540846727170835
	pesos_i(19477) := b"1111111111111111_1111111111111111_1111110111010000_1111000010101010"; -- -0.008530577186304117
	pesos_i(19478) := b"1111111111111111_1111111111111111_1111010110011111_1110101010101111"; -- -0.040528614215371905
	pesos_i(19479) := b"0000000000000000_0000000000000000_0000000000001110_1001111111101101"; -- 0.00022315542658511307
	pesos_i(19480) := b"0000000000000000_0000000000000000_0001101110100001_0100011010111010"; -- 0.10792963078616388
	pesos_i(19481) := b"0000000000000000_0000000000000000_0001100001100010_1111000011100001"; -- 0.09525971882929639
	pesos_i(19482) := b"1111111111111111_1111111111111111_1111011000110100_1100111101001011"; -- -0.038256687425581984
	pesos_i(19483) := b"1111111111111111_1111111111111111_1101100111001001_1100101101110011"; -- -0.14926460695734448
	pesos_i(19484) := b"1111111111111111_1111111111111111_1111011100000001_1100110100000011"; -- -0.03512877165093399
	pesos_i(19485) := b"1111111111111111_1111111111111111_1111010000100110_1110110111110100"; -- -0.0462809830138662
	pesos_i(19486) := b"1111111111111111_1111111111111111_1111101110000010_1111110110010101"; -- -0.017532492747554043
	pesos_i(19487) := b"1111111111111111_1111111111111111_1111101101010111_1111010000101010"; -- -0.018189182076374252
	pesos_i(19488) := b"0000000000000000_0000000000000000_0000101001011010_1110110100001000"; -- 0.0404499191378997
	pesos_i(19489) := b"1111111111111111_1111111111111111_1111000011010000_0110111110001010"; -- -0.05931952366544723
	pesos_i(19490) := b"1111111111111111_1111111111111111_1110011100010110_1001100111000010"; -- -0.09731139195020246
	pesos_i(19491) := b"0000000000000000_0000000000000000_0000001010100001_1100000001111000"; -- 0.010280636995253311
	pesos_i(19492) := b"0000000000000000_0000000000000000_0010001101010100_0100011010100000"; -- 0.13800469779006622
	pesos_i(19493) := b"0000000000000000_0000000000000000_0000000100010100_0101010101001101"; -- 0.004216510044253366
	pesos_i(19494) := b"1111111111111111_1111111111111111_1110010010101110_0101000110110101"; -- -0.10671510061413175
	pesos_i(19495) := b"0000000000000000_0000000000000000_0001100110000100_1101011111001111"; -- 0.09968327343610252
	pesos_i(19496) := b"0000000000000000_0000000000000000_0000011110100111_1011101110110100"; -- 0.02990315578143109
	pesos_i(19497) := b"1111111111111111_1111111111111111_1101110011001100_1110100000010011"; -- -0.13749837422732739
	pesos_i(19498) := b"1111111111111111_1111111111111111_1110000111001110_0010100001000000"; -- -0.1179480403503964
	pesos_i(19499) := b"0000000000000000_0000000000000000_0001011011101010_1011001100110111"; -- 0.08951873876650109
	pesos_i(19500) := b"0000000000000000_0000000000000000_0000110010010110_1010001100001110"; -- 0.04917353717538998
	pesos_i(19501) := b"0000000000000000_0000000000000000_0001011000100111_0100011001000000"; -- 0.0865367799882523
	pesos_i(19502) := b"0000000000000000_0000000000000000_0001110110111110_0110011101101011"; -- 0.11618658422813209
	pesos_i(19503) := b"1111111111111111_1111111111111111_1111110100000011_1100001110111011"; -- -0.011661307207795058
	pesos_i(19504) := b"0000000000000000_0000000000000000_0000101010100001_0100001010010101"; -- 0.04152313353534933
	pesos_i(19505) := b"1111111111111111_1111111111111111_1111010111111100_1101101110101100"; -- -0.03911044178904035
	pesos_i(19506) := b"0000000000000000_0000000000000000_0000010001100000_0011100010001100"; -- 0.017093214252076407
	pesos_i(19507) := b"1111111111111111_1111111111111111_1111110101101010_0000010000101011"; -- -0.010101069893860216
	pesos_i(19508) := b"1111111111111111_1111111111111111_1110001010100000_0110001110011100"; -- -0.11474015660225753
	pesos_i(19509) := b"1111111111111111_1111111111111111_1110101110110001_1100110111110011"; -- -0.07931816870648578
	pesos_i(19510) := b"1111111111111111_1111111111111111_1111001100001010_1000111011110110"; -- -0.050620140867632495
	pesos_i(19511) := b"1111111111111111_1111111111111111_1110000010011011_1010101010100001"; -- -0.12262471753083623
	pesos_i(19512) := b"0000000000000000_0000000000000000_0010011010001010_1000010000010001"; -- 0.15055108473134196
	pesos_i(19513) := b"0000000000000000_0000000000000000_0001110001001001_1101010011010001"; -- 0.110501576444775
	pesos_i(19514) := b"0000000000000000_0000000000000000_0001110101010100_0111111100110101"; -- 0.11457057044594525
	pesos_i(19515) := b"0000000000000000_0000000000000000_0001000111001101_0110011100110100"; -- 0.06954045310534711
	pesos_i(19516) := b"1111111111111111_1111111111111111_1111011111011110_0101101101000000"; -- -0.03176335990820375
	pesos_i(19517) := b"0000000000000000_0000000000000000_0001110100000011_1011111010010011"; -- 0.11333838544323709
	pesos_i(19518) := b"0000000000000000_0000000000000000_0001100000000110_1101000101101000"; -- 0.09385403442261986
	pesos_i(19519) := b"1111111111111111_1111111111111111_1111010100010011_1010100100011001"; -- -0.04266875393807414
	pesos_i(19520) := b"1111111111111111_1111111111111111_1111110111101101_0010110010011011"; -- -0.008099758406408641
	pesos_i(19521) := b"1111111111111111_1111111111111111_1111110111100001_1111111000000001"; -- -0.008270382558180132
	pesos_i(19522) := b"0000000000000000_0000000000000000_0010001010001001_0111011011101101"; -- 0.13491004274678128
	pesos_i(19523) := b"1111111111111111_1111111111111111_1111001110111100_0100010110010101"; -- -0.04790845027181371
	pesos_i(19524) := b"0000000000000000_0000000000000000_0000011100100111_0010010101011001"; -- 0.027941068854291835
	pesos_i(19525) := b"1111111111111111_1111111111111111_1110011111111011_1000011000001100"; -- -0.09381830414047308
	pesos_i(19526) := b"1111111111111111_1111111111111111_1110110110000101_1110100100100001"; -- -0.07217543547010996
	pesos_i(19527) := b"0000000000000000_0000000000000000_0001010011011111_0111110001000100"; -- 0.08153511686065408
	pesos_i(19528) := b"1111111111111111_1111111111111111_1110001011010100_1001110101101011"; -- -0.11394325397028891
	pesos_i(19529) := b"0000000000000000_0000000000000000_0001010111110001_1010000011100111"; -- 0.08571820866669125
	pesos_i(19530) := b"0000000000000000_0000000000000000_0001000101101110_1110000000101001"; -- 0.06809807774178528
	pesos_i(19531) := b"1111111111111111_1111111111111111_1101111011010100_1110001011000100"; -- -0.1295641203604941
	pesos_i(19532) := b"0000000000000000_0000000000000000_0001011011000011_0011111100011010"; -- 0.08891672507479426
	pesos_i(19533) := b"1111111111111111_1111111111111111_1101110101111001_0100100100011000"; -- -0.13486807976807258
	pesos_i(19534) := b"0000000000000000_0000000000000000_0001111111111011_0001001111100110"; -- 0.1249248921784911
	pesos_i(19535) := b"1111111111111111_1111111111111111_1111111100100010_0101110010101000"; -- -0.003381928342680383
	pesos_i(19536) := b"1111111111111111_1111111111111111_1110110110010001_1010110111100101"; -- -0.07199586069868966
	pesos_i(19537) := b"1111111111111111_1111111111111111_1111000001000100_0000010010011100"; -- -0.06146212766522484
	pesos_i(19538) := b"1111111111111111_1111111111111111_1101011110000100_1010111011000011"; -- -0.15813167312002777
	pesos_i(19539) := b"0000000000000000_0000000000000000_0010011001010001_0101000000001111"; -- 0.14967823374064415
	pesos_i(19540) := b"0000000000000000_0000000000000000_0000000000000100_1110000011100001"; -- 7.443904469750707e-05
	pesos_i(19541) := b"0000000000000000_0000000000000000_0000010101011111_0101110111001100"; -- 0.020986425782361366
	pesos_i(19542) := b"1111111111111111_1111111111111111_1110111110011011_1001101000111110"; -- -0.06403194424047512
	pesos_i(19543) := b"1111111111111111_1111111111111111_1111101001001000_0000101000100011"; -- -0.022338262959963523
	pesos_i(19544) := b"1111111111111111_1111111111111111_1111010001000111_1111100010110000"; -- -0.045776802972350594
	pesos_i(19545) := b"1111111111111111_1111111111111111_1111010100111100_0100111100001101"; -- -0.04204851096311543
	pesos_i(19546) := b"0000000000000000_0000000000000000_0001101011011010_0110100000000000"; -- 0.10489511500371386
	pesos_i(19547) := b"1111111111111111_1111111111111111_1101110010101010_0110111001100011"; -- -0.13802442627830572
	pesos_i(19548) := b"0000000000000000_0000000000000000_0001101000011010_1101011101011011"; -- 0.10197206481645478
	pesos_i(19549) := b"1111111111111111_1111111111111111_1110011001010001_0110001110101101"; -- -0.10032059693499466
	pesos_i(19550) := b"1111111111111111_1111111111111111_1111100111101100_1100001001100010"; -- -0.023731089747701672
	pesos_i(19551) := b"1111111111111111_1111111111111111_1101100101101000_0001011110110010"; -- -0.15075542367922498
	pesos_i(19552) := b"0000000000000000_0000000000000000_0000101111100100_0001001100110110"; -- 0.046448899070225556
	pesos_i(19553) := b"0000000000000000_0000000000000000_0000000111100011_0011100010001010"; -- 0.007373365127756563
	pesos_i(19554) := b"0000000000000000_0000000000000000_0000101011000010_0100011000011111"; -- 0.042026884510248136
	pesos_i(19555) := b"0000000000000000_0000000000000000_0000010001111010_1010001011111100"; -- 0.017496286807117
	pesos_i(19556) := b"0000000000000000_0000000000000000_0000001100110001_0110110100010011"; -- 0.012472932100007016
	pesos_i(19557) := b"1111111111111111_1111111111111111_1110011111011011_1100111110000100"; -- -0.09430220639631884
	pesos_i(19558) := b"0000000000000000_0000000000000000_0000001001010100_1100000101000001"; -- 0.009105757143835224
	pesos_i(19559) := b"0000000000000000_0000000000000000_0000000001111100_0010000000010110"; -- 0.0018940022973882081
	pesos_i(19560) := b"1111111111111111_1111111111111111_1110000100110010_1110101100000110"; -- -0.12031680209794929
	pesos_i(19561) := b"1111111111111111_1111111111111111_1111111101010001_0101110000100110"; -- -0.0026647956746195817
	pesos_i(19562) := b"0000000000000000_0000000000000000_0000001100101101_1110101110111011"; -- 0.012419446082665455
	pesos_i(19563) := b"0000000000000000_0000000000000000_0000011011110100_1001011001010110"; -- 0.027169605138613526
	pesos_i(19564) := b"1111111111111111_1111111111111111_1111111100011101_1100001000101111"; -- -0.0034521708512991554
	pesos_i(19565) := b"1111111111111111_1111111111111111_1110111010010111_0100001101001010"; -- -0.06800441201349598
	pesos_i(19566) := b"0000000000000000_0000000000000000_0001110010100001_0000111111100101"; -- 0.11183261234433554
	pesos_i(19567) := b"0000000000000000_0000000000000000_0001010110011011_1010110010111000"; -- 0.08440665714106475
	pesos_i(19568) := b"0000000000000000_0000000000000000_0000110011101111_0000000010100100"; -- 0.05052188871027811
	pesos_i(19569) := b"1111111111111111_1111111111111111_1101110110000110_1110101010000011"; -- -0.1346600942883366
	pesos_i(19570) := b"0000000000000000_0000000000000000_0000001100000101_0010100000000000"; -- 0.011797428222911507
	pesos_i(19571) := b"0000000000000000_0000000000000000_0000011110000000_1011111010010100"; -- 0.029308234429132843
	pesos_i(19572) := b"0000000000000000_0000000000000000_0000101001111001_0101101111111100"; -- 0.04091429620351698
	pesos_i(19573) := b"0000000000000000_0000000000000000_0001101000101111_1111011001010001"; -- 0.10229434477290218
	pesos_i(19574) := b"1111111111111111_1111111111111111_1111010011010001_0000010110001100"; -- -0.043685582415540276
	pesos_i(19575) := b"1111111111111111_1111111111111111_1111100100011111_1101111011010000"; -- -0.02685744691528081
	pesos_i(19576) := b"1111111111111111_1111111111111111_1110110001101011_1010011100001000"; -- -0.07648235365091058
	pesos_i(19577) := b"1111111111111111_1111111111111111_1111111101001000_0110110011101001"; -- -0.0028011256366160925
	pesos_i(19578) := b"0000000000000000_0000000000000000_0001100011011000_0111011011001100"; -- 0.09705297917910367
	pesos_i(19579) := b"0000000000000000_0000000000000000_0001010100000110_1110110100011010"; -- 0.08213693519992665
	pesos_i(19580) := b"0000000000000000_0000000000000000_0001001110111000_1001110111000000"; -- 0.07703576971973897
	pesos_i(19581) := b"0000000000000000_0000000000000000_0000011111001001_1011111011100010"; -- 0.03042214400618443
	pesos_i(19582) := b"0000000000000000_0000000000000000_0010000110101001_0110000110011110"; -- 0.13149080372752286
	pesos_i(19583) := b"1111111111111111_1111111111111111_1110010100000000_1001110111011010"; -- -0.10545934132467014
	pesos_i(19584) := b"1111111111111111_1111111111111111_1111100000101110_1011110110101100"; -- -0.030536790355217176
	pesos_i(19585) := b"1111111111111111_1111111111111111_1101100011010101_0010111011101011"; -- -0.15299708151200203
	pesos_i(19586) := b"0000000000000000_0000000000000000_0010001111011101_1100111101010100"; -- 0.140103300007709
	pesos_i(19587) := b"1111111111111111_1111111111111111_1111111100101100_1111011110001011"; -- -0.003220108487342155
	pesos_i(19588) := b"1111111111111111_1111111111111111_1111110001110001_0100101101101011"; -- -0.01389626154604642
	pesos_i(19589) := b"0000000000000000_0000000000000000_0000111100100101_0000100010001001"; -- 0.059158833818634654
	pesos_i(19590) := b"0000000000000000_0000000000000000_0000001110101110_0010101111101011"; -- 0.0143763969526961
	pesos_i(19591) := b"1111111111111111_1111111111111111_1111011110111100_1000111011111111"; -- -0.03227907444103586
	pesos_i(19592) := b"0000000000000000_0000000000000000_0001000111111110_1111111010100111"; -- 0.07029716080753523
	pesos_i(19593) := b"0000000000000000_0000000000000000_0000101001010001_0101010101001111"; -- 0.04030354666140854
	pesos_i(19594) := b"0000000000000000_0000000000000000_0000000110101000_0000011010010100"; -- 0.0064701187611581595
	pesos_i(19595) := b"0000000000000000_0000000000000000_0010001000110111_0110001101111111"; -- 0.13365766393394857
	pesos_i(19596) := b"0000000000000000_0000000000000000_0001011011101000_1010001001011100"; -- 0.089487216446052
	pesos_i(19597) := b"1111111111111111_1111111111111111_1111111001111000_1011011111111111"; -- -0.005970478316077782
	pesos_i(19598) := b"1111111111111111_1111111111111111_1111001110100010_1010010101011111"; -- -0.04829946939641713
	pesos_i(19599) := b"0000000000000000_0000000000000000_0001000101111001_1101010000000101"; -- 0.06826520081385305
	pesos_i(19600) := b"0000000000000000_0000000000000000_0010000011000100_0111010000110000"; -- 0.12799764795585236
	pesos_i(19601) := b"1111111111111111_1111111111111111_1111010110100110_1101010011100000"; -- -0.040423102760329344
	pesos_i(19602) := b"1111111111111111_1111111111111111_1101101011101110_1011011100111010"; -- -0.1447949870882875
	pesos_i(19603) := b"0000000000000000_0000000000000000_0001000000101110_0101101000100111"; -- 0.06320727782476836
	pesos_i(19604) := b"1111111111111111_1111111111111111_1110010111111110_1100000010110100"; -- -0.10158153148222211
	pesos_i(19605) := b"1111111111111111_1111111111111111_1110011001011001_1100010001000010"; -- -0.10019276978156322
	pesos_i(19606) := b"0000000000000000_0000000000000000_0000000000110000_1101010101011001"; -- 0.0007451384683675271
	pesos_i(19607) := b"0000000000000000_0000000000000000_0001000101010010_1011101011101111"; -- 0.06766861283209867
	pesos_i(19608) := b"1111111111111111_1111111111111111_1110100011111111_1000010111100001"; -- -0.08985102908192547
	pesos_i(19609) := b"1111111111111111_1111111111111111_1110001110101001_1001110100101101"; -- -0.11069314633534577
	pesos_i(19610) := b"1111111111111111_1111111111111111_1111101011011011_0001011011011100"; -- -0.020094462680799705
	pesos_i(19611) := b"0000000000000000_0000000000000000_0000101001010001_1111010010100100"; -- 0.04031304357916695
	pesos_i(19612) := b"1111111111111111_1111111111111111_1110100111001110_1000001110100110"; -- -0.08669259260441824
	pesos_i(19613) := b"1111111111111111_1111111111111111_1111001111001101_1101010110000100"; -- -0.0476404717091387
	pesos_i(19614) := b"1111111111111111_1111111111111111_1101100111101010_0000010011000110"; -- -0.14877290881082245
	pesos_i(19615) := b"1111111111111111_1111111111111111_1111110011101000_0010011100101101"; -- -0.012082625770160924
	pesos_i(19616) := b"0000000000000000_0000000000000000_0001111000001011_1011101100110000"; -- 0.1173665038332253
	pesos_i(19617) := b"0000000000000000_0000000000000000_0001011100000111_0111011010010100"; -- 0.08995762926491228
	pesos_i(19618) := b"0000000000000000_0000000000000000_0001110101000001_0110100001011011"; -- 0.11427929137528262
	pesos_i(19619) := b"1111111111111111_1111111111111111_1111100101101101_1101011100110000"; -- -0.025667715797045444
	pesos_i(19620) := b"1111111111111111_1111111111111111_1111001000000001_1001101000101100"; -- -0.05466305185247461
	pesos_i(19621) := b"0000000000000000_0000000000000000_0000101101111101_1110011111100001"; -- 0.044889919786498964
	pesos_i(19622) := b"0000000000000000_0000000000000000_0001111110100010_0010100110111001"; -- 0.12356816071590146
	pesos_i(19623) := b"0000000000000000_0000000000000000_0001111010111110_0100010011001010"; -- 0.12009077014286419
	pesos_i(19624) := b"0000000000000000_0000000000000000_0010000100011011_1000100101010000"; -- 0.12932642184663676
	pesos_i(19625) := b"1111111111111111_1111111111111111_1110010111100101_0100101110001101"; -- -0.10196998409410647
	pesos_i(19626) := b"0000000000000000_0000000000000000_0001100101000111_0011010110000001"; -- 0.09874281315417235
	pesos_i(19627) := b"1111111111111111_1111111111111111_1111111111001101_1100010111101110"; -- -0.0007664006429791935
	pesos_i(19628) := b"0000000000000000_0000000000000000_0001011010000001_1100111011001111"; -- 0.08791821054081592
	pesos_i(19629) := b"1111111111111111_1111111111111111_1111000001010001_0001110000100101"; -- -0.06126236053870273
	pesos_i(19630) := b"1111111111111111_1111111111111111_1111001001101100_0110100101010100"; -- -0.05303327265135906
	pesos_i(19631) := b"1111111111111111_1111111111111111_1111111011111100_1000100101000010"; -- -0.0039591039449912765
	pesos_i(19632) := b"1111111111111111_1111111111111111_1110110011011111_0010010011001000"; -- -0.07472009778994211
	pesos_i(19633) := b"0000000000000000_0000000000000000_0000100001110101_0101110000001011"; -- 0.03304076449248049
	pesos_i(19634) := b"1111111111111111_1111111111111111_1110000010101010_0101011010110100"; -- -0.12240083784101355
	pesos_i(19635) := b"1111111111111111_1111111111111111_1110101010111010_1001101010010111"; -- -0.08309015101522267
	pesos_i(19636) := b"0000000000000000_0000000000000000_0001101011001011_0110111101101111"; -- 0.10466667612773935
	pesos_i(19637) := b"0000000000000000_0000000000000000_0000101101000101_0000010100010100"; -- 0.04402190902866972
	pesos_i(19638) := b"1111111111111111_1111111111111111_1111001100101010_1001100001110010"; -- -0.050131294330664766
	pesos_i(19639) := b"1111111111111111_1111111111111111_1110010110000101_0101000111110001"; -- -0.10343444692753441
	pesos_i(19640) := b"1111111111111111_1111111111111111_1110111100101010_0001010100001100"; -- -0.0657641263054588
	pesos_i(19641) := b"1111111111111111_1111111111111111_1110100100001001_1101000001101001"; -- -0.08969399868442432
	pesos_i(19642) := b"1111111111111111_1111111111111111_1110000100101011_0001001100100100"; -- -0.1204364812841586
	pesos_i(19643) := b"0000000000000000_0000000000000000_0000111001101111_1000100111001011"; -- 0.05638943878802258
	pesos_i(19644) := b"1111111111111111_1111111111111111_1111001111010011_1011011010010100"; -- -0.04755076297865573
	pesos_i(19645) := b"1111111111111111_1111111111111111_1111101010111011_0000010000100111"; -- -0.020583858932990886
	pesos_i(19646) := b"0000000000000000_0000000000000000_0000011110100011_1101011110100010"; -- 0.029843785315468017
	pesos_i(19647) := b"1111111111111111_1111111111111111_1110101011001010_0000110101100101"; -- -0.08285442620294452
	pesos_i(19648) := b"0000000000000000_0000000000000000_0000101110010010_1100000001110111"; -- 0.04520800497191667
	pesos_i(19649) := b"1111111111111111_1111111111111111_1101110001011111_0001000100101100"; -- -0.13917439151962172
	pesos_i(19650) := b"0000000000000000_0000000000000000_0001101001111100_1101111100101000"; -- 0.10346789095717886
	pesos_i(19651) := b"1111111111111111_1111111111111111_1111110000100101_0100001111000101"; -- -0.015056385496635485
	pesos_i(19652) := b"0000000000000000_0000000000000000_0000110100110111_0011011110001010"; -- 0.051623793892509824
	pesos_i(19653) := b"0000000000000000_0000000000000000_0000000011110101_1010010000000000"; -- 0.003748178365811089
	pesos_i(19654) := b"1111111111111111_1111111111111111_1111001111001010_0001001101010101"; -- -0.04769782234242874
	pesos_i(19655) := b"1111111111111111_1111111111111111_1101101001001101_0011111101110110"; -- -0.14725879064329084
	pesos_i(19656) := b"1111111111111111_1111111111111111_1111101000111001_1001001010001001"; -- -0.022559014835908234
	pesos_i(19657) := b"1111111111111111_1111111111111111_1111110000000111_0101101110101011"; -- -0.015512724749485994
	pesos_i(19658) := b"1111111111111111_1111111111111111_1110001011100110_0111011110000110"; -- -0.11367085447728635
	pesos_i(19659) := b"1111111111111111_1111111111111111_1111001011010001_1111100100000110"; -- -0.05148357012856189
	pesos_i(19660) := b"1111111111111111_1111111111111111_1111000100111100_0010010111110100"; -- -0.057675960390744394
	pesos_i(19661) := b"1111111111111111_1111111111111111_1111110101011000_0001011100110010"; -- -0.010374593932510626
	pesos_i(19662) := b"1111111111111111_1111111111111111_1110111110101101_1111001111000000"; -- -0.06375195095315904
	pesos_i(19663) := b"0000000000000000_0000000000000000_0000111011100011_0101100011101000"; -- 0.05815654438258185
	pesos_i(19664) := b"1111111111111111_1111111111111111_1101110101010001_1011100101000100"; -- -0.13547174548229501
	pesos_i(19665) := b"0000000000000000_0000000000000000_0001011001010001_1000011111111000"; -- 0.08718156630336607
	pesos_i(19666) := b"0000000000000000_0000000000000000_0001111110101010_0000000011101101"; -- 0.12368779936942731
	pesos_i(19667) := b"0000000000000000_0000000000000000_0001000010100000_1111001111011100"; -- 0.06495594148939608
	pesos_i(19668) := b"0000000000000000_0000000000000000_0000101101110110_0111010010000100"; -- 0.04477623208702816
	pesos_i(19669) := b"0000000000000000_0000000000000000_0001000110111100_0011011010101001"; -- 0.06927816033742178
	pesos_i(19670) := b"0000000000000000_0000000000000000_0000100100111101_0011101010011110"; -- 0.036090529970197516
	pesos_i(19671) := b"0000000000000000_0000000000000000_0000111001011001_1011010110111101"; -- 0.05605636464742265
	pesos_i(19672) := b"0000000000000000_0000000000000000_0000010011000101_0010000101011001"; -- 0.01863296912284369
	pesos_i(19673) := b"1111111111111111_1111111111111111_1101101001100010_0010000010110100"; -- -0.14694018936782255
	pesos_i(19674) := b"0000000000000000_0000000000000000_0001111101010111_1000100000011101"; -- 0.12242937758863827
	pesos_i(19675) := b"0000000000000000_0000000000000000_0001110101100010_0101111011001101"; -- 0.11478226191674598
	pesos_i(19676) := b"1111111111111111_1111111111111111_1111111001111000_1001001111010010"; -- -0.005972634498066417
	pesos_i(19677) := b"0000000000000000_0000000000000000_0000000111100001_1001110010100010"; -- 0.007348813502615414
	pesos_i(19678) := b"1111111111111111_1111111111111111_1110000000011011_1110111110111101"; -- -0.12457372326874293
	pesos_i(19679) := b"1111111111111111_1111111111111111_1110111010000111_1110011101011100"; -- -0.06823877342522935
	pesos_i(19680) := b"1111111111111111_1111111111111111_1110010000011001_0000100011011100"; -- -0.1089930022846571
	pesos_i(19681) := b"1111111111111111_1111111111111111_1101111100000010_1000011111100101"; -- -0.12886763256464837
	pesos_i(19682) := b"0000000000000000_0000000000000000_0000011010101011_1101011001100100"; -- 0.026059531700706583
	pesos_i(19683) := b"1111111111111111_1111111111111111_1111101011000111_1001000110000010"; -- -0.020392327966061722
	pesos_i(19684) := b"1111111111111111_1111111111111111_1101100110011000_1010110111100000"; -- -0.15001405035916743
	pesos_i(19685) := b"1111111111111111_1111111111111111_1110111111101000_1100000101000100"; -- -0.06285469137348619
	pesos_i(19686) := b"0000000000000000_0000000000000000_0001000011000010_0011101111100110"; -- 0.06546377518874955
	pesos_i(19687) := b"0000000000000000_0000000000000000_0000100101101100_0010000000001010"; -- 0.036806108957393856
	pesos_i(19688) := b"0000000000000000_0000000000000000_0010001101010101_0111001010001001"; -- 0.13802257397768256
	pesos_i(19689) := b"1111111111111111_1111111111111111_1111001110010010_0001101011101001"; -- -0.04855186286168427
	pesos_i(19690) := b"0000000000000000_0000000000000000_0000001111011011_0001011100100000"; -- 0.015061803264160118
	pesos_i(19691) := b"0000000000000000_0000000000000000_0000011111111010_0011001110100100"; -- 0.031161525277109612
	pesos_i(19692) := b"0000000000000000_0000000000000000_0000001111110101_0101110110010011"; -- 0.015462730750082771
	pesos_i(19693) := b"1111111111111111_1111111111111111_1101011011011011_1000010001110110"; -- -0.16071292993539166
	pesos_i(19694) := b"0000000000000000_0000000000000000_0000000101010100_1010010101111101"; -- 0.005197852055151678
	pesos_i(19695) := b"0000000000000000_0000000000000000_0000000101000101_1010011001110000"; -- 0.00496902682695615
	pesos_i(19696) := b"1111111111111111_1111111111111111_1110101100010111_0011111110001010"; -- -0.08167651061286338
	pesos_i(19697) := b"0000000000000000_0000000000000000_0001101110011111_1111110000110000"; -- 0.1079099291054884
	pesos_i(19698) := b"1111111111111111_1111111111111111_1110000010101000_0001001011101111"; -- -0.1224353949068029
	pesos_i(19699) := b"1111111111111111_1111111111111111_1111010110101010_1101011110100110"; -- -0.040361902099611484
	pesos_i(19700) := b"0000000000000000_0000000000000000_0001000011010110_1001010010011011"; -- 0.0657742384385595
	pesos_i(19701) := b"0000000000000000_0000000000000000_0000100111000011_1111111010101101"; -- 0.03814689377731092
	pesos_i(19702) := b"1111111111111111_1111111111111111_1111010011010101_1100110110011111"; -- -0.04361262195142285
	pesos_i(19703) := b"0000000000000000_0000000000000000_0000001001001100_1111100000011001"; -- 0.008986955710919207
	pesos_i(19704) := b"1111111111111111_1111111111111111_1101110000100000_1000000001110100"; -- -0.1401290624303028
	pesos_i(19705) := b"0000000000000000_0000000000000000_0010001010111011_0100001110111001"; -- 0.13566993016532938
	pesos_i(19706) := b"1111111111111111_1111111111111111_1110111010101100_1111001101101110"; -- -0.06767347885093952
	pesos_i(19707) := b"1111111111111111_1111111111111111_1101011001010001_0000110011111100"; -- -0.16282576410015065
	pesos_i(19708) := b"1111111111111111_1111111111111111_1110001000000100_1110101001011000"; -- -0.1171124968780761
	pesos_i(19709) := b"1111111111111111_1111111111111111_1110010100101111_0110010010111001"; -- -0.10474558339869537
	pesos_i(19710) := b"1111111111111111_1111111111111111_1110111111100000_1101110000001100"; -- -0.06297516548847917
	pesos_i(19711) := b"0000000000000000_0000000000000000_0000011110001000_0101001000100110"; -- 0.029423841737390728
	pesos_i(19712) := b"0000000000000000_0000000000000000_0000011001101011_1010010101000100"; -- 0.025080041060927868
	pesos_i(19713) := b"0000000000000000_0000000000000000_0000010011101000_1001101010000000"; -- 0.019174247995880866
	pesos_i(19714) := b"0000000000000000_0000000000000000_0001000001010000_0110111100110000"; -- 0.06372733051355024
	pesos_i(19715) := b"0000000000000000_0000000000000000_0001111110001110_1000011101101000"; -- 0.123268568851509
	pesos_i(19716) := b"1111111111111111_1111111111111111_1110011011010110_0111011110010000"; -- -0.09828999260968894
	pesos_i(19717) := b"0000000000000000_0000000000000000_0001011110101100_0110100101110101"; -- 0.09247454755660758
	pesos_i(19718) := b"1111111111111111_1111111111111111_1111000010011100_0100011010000111"; -- -0.060115425055539407
	pesos_i(19719) := b"1111111111111111_1111111111111111_1110110111010011_1011110010000010"; -- -0.07098790967344759
	pesos_i(19720) := b"1111111111111111_1111111111111111_1111101010110110_1100000100000101"; -- -0.02064889558109493
	pesos_i(19721) := b"1111111111111111_1111111111111111_1101101011011100_1010101001110110"; -- -0.1450704061901783
	pesos_i(19722) := b"1111111111111111_1111111111111111_1110010100011111_1110110100001000"; -- -0.10498159942290508
	pesos_i(19723) := b"0000000000000000_0000000000000000_0000001010111111_0011111100010000"; -- 0.010730687624339342
	pesos_i(19724) := b"1111111111111111_1111111111111111_1111111010001011_1000100100110011"; -- -0.0056833506839416015
	pesos_i(19725) := b"1111111111111111_1111111111111111_1110011011010010_0010111100100101"; -- -0.0983553443752731
	pesos_i(19726) := b"0000000000000000_0000000000000000_0010011000110110_1001001010001111"; -- 0.14927021027877832
	pesos_i(19727) := b"0000000000000000_0000000000000000_0001110111010111_0110010000111000"; -- 0.1165678631895559
	pesos_i(19728) := b"1111111111111111_1111111111111111_1111010111100001_0011100101001011"; -- -0.03953210744261301
	pesos_i(19729) := b"0000000000000000_0000000000000000_0001000011011110_1001111100101001"; -- 0.06589693786366513
	pesos_i(19730) := b"0000000000000000_0000000000000000_0000000111010001_0001001000101001"; -- 0.007096419244501199
	pesos_i(19731) := b"0000000000000000_0000000000000000_0000011111110101_1011011000001101"; -- 0.031093004452310682
	pesos_i(19732) := b"0000000000000000_0000000000000000_0000010000010000_0011010010010110"; -- 0.01587227501206907
	pesos_i(19733) := b"1111111111111111_1111111111111111_1101111010100110_1100001001101111"; -- -0.1302679518459227
	pesos_i(19734) := b"1111111111111111_1111111111111111_1111001000111001_1001010001100010"; -- -0.05380890461095819
	pesos_i(19735) := b"1111111111111111_1111111111111111_1110000010010100_1111101010000100"; -- -0.12272676731712225
	pesos_i(19736) := b"0000000000000000_0000000000000000_0001001011110100_1101111001001101"; -- 0.07404889461854537
	pesos_i(19737) := b"1111111111111111_1111111111111111_1110010111111000_1101111001100001"; -- -0.10167131542176687
	pesos_i(19738) := b"0000000000000000_0000000000000000_0001011111010110_0110110000111001"; -- 0.09311558135493953
	pesos_i(19739) := b"0000000000000000_0000000000000000_0010010011111100_0011101111011110"; -- 0.14447378330345437
	pesos_i(19740) := b"1111111111111111_1111111111111111_1111110010011101_0101100101101000"; -- -0.013224041189899264
	pesos_i(19741) := b"0000000000000000_0000000000000000_0000000101110000_0001000101100011"; -- 0.005616270674058075
	pesos_i(19742) := b"1111111111111111_1111111111111111_1110011010001101_1000110001110010"; -- -0.09940263965089426
	pesos_i(19743) := b"0000000000000000_0000000000000000_0001100111111101_1011110110101100"; -- 0.10152802899725565
	pesos_i(19744) := b"0000000000000000_0000000000000000_0001101011000111_1010010010100101"; -- 0.1046088126719043
	pesos_i(19745) := b"0000000000000000_0000000000000000_0000110101101101_1111011101000101"; -- 0.052459196342732814
	pesos_i(19746) := b"0000000000000000_0000000000000000_0000000000101100_0001101110000110"; -- 0.0006730272427004004
	pesos_i(19747) := b"0000000000000000_0000000000000000_0000001000100001_0011111111101100"; -- 0.008319850104327139
	pesos_i(19748) := b"1111111111111111_1111111111111111_1111100110111111_0010110000000010"; -- -0.02442669822441609
	pesos_i(19749) := b"0000000000000000_0000000000000000_0001000110110100_1010111011111101"; -- 0.06916326210657538
	pesos_i(19750) := b"1111111111111111_1111111111111111_1110100100101100_1101011110100101"; -- -0.08915950982645178
	pesos_i(19751) := b"1111111111111111_1111111111111111_1110111001100000_0111011111000000"; -- -0.06884051866722679
	pesos_i(19752) := b"0000000000000000_0000000000000000_0000010001110001_1000110110001010"; -- 0.017357679541545098
	pesos_i(19753) := b"0000000000000000_0000000000000000_0001101111011011_0110011000110100"; -- 0.10881651651992628
	pesos_i(19754) := b"1111111111111111_1111111111111111_1111010011110001_1001000101111111"; -- -0.04318895964739232
	pesos_i(19755) := b"0000000000000000_0000000000000000_0000010000011001_1100101000100100"; -- 0.016018518142731135
	pesos_i(19756) := b"1111111111111111_1111111111111111_1111100010011100_1010111100011111"; -- -0.028859190914115238
	pesos_i(19757) := b"0000000000000000_0000000000000000_0000011110011011_0010100100111001"; -- 0.029711319295314592
	pesos_i(19758) := b"0000000000000000_0000000000000000_0001010000101111_0100101000001101"; -- 0.07884657678913413
	pesos_i(19759) := b"1111111111111111_1111111111111111_1111100111101011_0000010111001000"; -- -0.02375759009517245
	pesos_i(19760) := b"0000000000000000_0000000000000000_0010011010001111_1100110101010001"; -- 0.15063174464959853
	pesos_i(19761) := b"0000000000000000_0000000000000000_0000101000111011_1000100011001010"; -- 0.03997092170320824
	pesos_i(19762) := b"0000000000000000_0000000000000000_0010010010000001_1101111100010100"; -- 0.14260668022656037
	pesos_i(19763) := b"0000000000000000_0000000000000000_0001000101001001_0010101010010100"; -- 0.06752267935730988
	pesos_i(19764) := b"0000000000000000_0000000000000000_0001110011110011_0000111011010000"; -- 0.1130837685601758
	pesos_i(19765) := b"1111111111111111_1111111111111111_1110010010111001_0011111011011111"; -- -0.10654837672668382
	pesos_i(19766) := b"1111111111111111_1111111111111111_1111101100111000_1010100110000100"; -- -0.01866665399453968
	pesos_i(19767) := b"0000000000000000_0000000000000000_0010010110111100_1000100101111101"; -- 0.1474080973075767
	pesos_i(19768) := b"1111111111111111_1111111111111111_1110011100011000_1001001111101010"; -- -0.09728122274319574
	pesos_i(19769) := b"1111111111111111_1111111111111111_1111100100110010_1011110101110001"; -- -0.02656951893617934
	pesos_i(19770) := b"0000000000000000_0000000000000000_0000000000111100_0111110111110110"; -- 0.0009230351443987908
	pesos_i(19771) := b"0000000000000000_0000000000000000_0001111101110100_0001000110001110"; -- 0.12286481592511707
	pesos_i(19772) := b"1111111111111111_1111111111111111_1110101101011001_0001001001110111"; -- -0.08067211715042573
	pesos_i(19773) := b"0000000000000000_0000000000000000_0010000101111001_1000101110101001"; -- 0.13076088794607957
	pesos_i(19774) := b"0000000000000000_0000000000000000_0001011001101010_0001110011101110"; -- 0.08755665596394276
	pesos_i(19775) := b"0000000000000000_0000000000000000_0000111001001100_1010110011010010"; -- 0.055857468888360545
	pesos_i(19776) := b"0000000000000000_0000000000000000_0000111101110000_0110110010011111"; -- 0.06030920877060159
	pesos_i(19777) := b"1111111111111111_1111111111111111_1111111100000010_1000000111111000"; -- -0.003867985625650596
	pesos_i(19778) := b"1111111111111111_1111111111111111_1111110010111111_0101000101110011"; -- -0.01270571662791687
	pesos_i(19779) := b"1111111111111111_1111111111111111_1101111011110011_0000001110000110"; -- -0.1291044043385333
	pesos_i(19780) := b"0000000000000000_0000000000000000_0001100011011001_0011001001101110"; -- 0.09706416305805908
	pesos_i(19781) := b"1111111111111111_1111111111111111_1110101111110000_1111110001010011"; -- -0.07835410104296205
	pesos_i(19782) := b"1111111111111111_1111111111111111_1110100010100010_0001011101000100"; -- -0.09127668940550958
	pesos_i(19783) := b"1111111111111111_1111111111111111_1110011111100001_1000110111000110"; -- -0.0942145721109327
	pesos_i(19784) := b"0000000000000000_0000000000000000_0000010100111000_1110101010000101"; -- 0.020399720565761545
	pesos_i(19785) := b"0000000000000000_0000000000000000_0001000101011000_1101010001000010"; -- 0.06776167498117615
	pesos_i(19786) := b"1111111111111111_1111111111111111_1101111000101000_1101001001010111"; -- -0.13218961111997576
	pesos_i(19787) := b"1111111111111111_1111111111111111_1110010000101000_1001101011000101"; -- -0.10875542341283138
	pesos_i(19788) := b"1111111111111111_1111111111111111_1110101100011100_1011010001101010"; -- -0.0815932504739673
	pesos_i(19789) := b"0000000000000000_0000000000000000_0000101101001001_1101111111000110"; -- 0.04409597955358139
	pesos_i(19790) := b"0000000000000000_0000000000000000_0001001010110110_0100100011111000"; -- 0.07309394898491926
	pesos_i(19791) := b"1111111111111111_1111111111111111_1111101100100001_0101111000001101"; -- -0.019022104069881984
	pesos_i(19792) := b"0000000000000000_0000000000000000_0001111001100011_1010011111101100"; -- 0.11870812915536735
	pesos_i(19793) := b"0000000000000000_0000000000000000_0001100011010110_1101001010011011"; -- 0.09702793384321831
	pesos_i(19794) := b"0000000000000000_0000000000000000_0000100011001111_0110000111100110"; -- 0.03441440455532145
	pesos_i(19795) := b"1111111111111111_1111111111111111_1111110011110100_0100000011100011"; -- -0.011897987808466142
	pesos_i(19796) := b"1111111111111111_1111111111111111_1101111011110011_0001110001101000"; -- -0.12910292109124513
	pesos_i(19797) := b"0000000000000000_0000000000000000_0000101011001100_1111000001011000"; -- 0.04218961854267168
	pesos_i(19798) := b"1111111111111111_1111111111111111_1101111110101110_1010000000000000"; -- -0.12624168402059416
	pesos_i(19799) := b"0000000000000000_0000000000000000_0001011100011010_0110001100010010"; -- 0.0902463835178528
	pesos_i(19800) := b"0000000000000000_0000000000000000_0000110111011100_0110100010000101"; -- 0.054144413398818377
	pesos_i(19801) := b"1111111111111111_1111111111111111_1111010000000010_0010111110110010"; -- -0.04684163966174922
	pesos_i(19802) := b"0000000000000000_0000000000000000_0000001111100111_1101010110001010"; -- 0.015256258077407615
	pesos_i(19803) := b"0000000000000000_0000000000000000_0001010101100110_1001011110101011"; -- 0.08359668663760039
	pesos_i(19804) := b"1111111111111111_1111111111111111_1110001010110101_0000101110110001"; -- -0.11442496240412901
	pesos_i(19805) := b"0000000000000000_0000000000000000_0010010001000100_1011000101110100"; -- 0.14167317458109716
	pesos_i(19806) := b"1111111111111111_1111111111111111_1101011111010011_0011001010001001"; -- -0.1569336333981362
	pesos_i(19807) := b"1111111111111111_1111111111111111_1111010110011110_0011010111110110"; -- -0.040554644890060595
	pesos_i(19808) := b"1111111111111111_1111111111111111_1111111111001110_0110111001111001"; -- -0.0007563547274684968
	pesos_i(19809) := b"1111111111111111_1111111111111111_1101111000000101_0011001110000011"; -- -0.13273313566437303
	pesos_i(19810) := b"0000000000000000_0000000000000000_0001110110001110_0110110010100010"; -- 0.11545447309548454
	pesos_i(19811) := b"0000000000000000_0000000000000000_0001000000111111_1100100001100101"; -- 0.06347324825280802
	pesos_i(19812) := b"0000000000000000_0000000000000000_0000110000111110_1110111011101110"; -- 0.04783528622224749
	pesos_i(19813) := b"1111111111111111_1111111111111111_1110100111111100_0100001011101100"; -- -0.08599454626000595
	pesos_i(19814) := b"1111111111111111_1111111111111111_1111010011111111_0111110101100010"; -- -0.042976535367325784
	pesos_i(19815) := b"1111111111111111_1111111111111111_1110111000011011_1001100000111011"; -- -0.06989143893676222
	pesos_i(19816) := b"0000000000000000_0000000000000000_0010001100000110_0101001011000110"; -- 0.1368152364274125
	pesos_i(19817) := b"1111111111111111_1111111111111111_1101011101101001_1100000110000010"; -- -0.15854254324383857
	pesos_i(19818) := b"1111111111111111_1111111111111111_1110000000001001_1110111011011101"; -- -0.12484843347332139
	pesos_i(19819) := b"1111111111111111_1111111111111111_1110111111101110_0001101111110111"; -- -0.06277299144486127
	pesos_i(19820) := b"0000000000000000_0000000000000000_0010101110001100_1000000100101011"; -- 0.17011267942553618
	pesos_i(19821) := b"0000000000000000_0000000000000000_0010000110101101_0001000010110100"; -- 0.13154701611882388
	pesos_i(19822) := b"1111111111111111_1111111111111111_1111011011110100_0001011101101110"; -- -0.03533795886902019
	pesos_i(19823) := b"1111111111111111_1111111111111111_1111001100101101_0110110001000100"; -- -0.05008815139961621
	pesos_i(19824) := b"1111111111111111_1111111111111111_1111001110110011_0001010101001111"; -- -0.048048656712823865
	pesos_i(19825) := b"1111111111111111_1111111111111111_1110100100100101_1000001101101011"; -- -0.08927134170860399
	pesos_i(19826) := b"1111111111111111_1111111111111111_1101100101111001_1111100101100000"; -- -0.15048257257177858
	pesos_i(19827) := b"1111111111111111_1111111111111111_1111111101111001_0001001001111001"; -- -0.0020588354829780887
	pesos_i(19828) := b"1111111111111111_1111111111111111_1101111011001000_0110101000110101"; -- -0.12975441178438477
	pesos_i(19829) := b"0000000000000000_0000000000000000_0000000000001001_1001101110100111"; -- 0.00014660675940678515
	pesos_i(19830) := b"0000000000000000_0000000000000000_0001111010010001_1100110100100100"; -- 0.11941225169778646
	pesos_i(19831) := b"1111111111111111_1111111111111111_1101101110101011_1111010010000011"; -- -0.14190742305467255
	pesos_i(19832) := b"1111111111111111_1111111111111111_1111110000010111_0111110011010000"; -- -0.015266608350792417
	pesos_i(19833) := b"0000000000000000_0000000000000000_0001100001000001_0011011101011110"; -- 0.09474512135276494
	pesos_i(19834) := b"1111111111111111_1111111111111111_1111011001001001_1001011001011101"; -- -0.037939646025760776
	pesos_i(19835) := b"1111111111111111_1111111111111111_1111001011000001_0101011000101000"; -- -0.05173741835124563
	pesos_i(19836) := b"0000000000000000_0000000000000000_0001100111011110_1010101001001111"; -- 0.10105385236114443
	pesos_i(19837) := b"0000000000000000_0000000000000000_0000100000011000_0000011000011100"; -- 0.03161657510276767
	pesos_i(19838) := b"1111111111111111_1111111111111111_1101111100110100_1000111101000001"; -- -0.12810425441509574
	pesos_i(19839) := b"0000000000000000_0000000000000000_0000101001001100_1110001101001010"; -- 0.04023571551843196
	pesos_i(19840) := b"1111111111111111_1111111111111111_1101010000100000_1100010011101111"; -- -0.17137498064677892
	pesos_i(19841) := b"1111111111111111_1111111111111111_1110001001001101_1100001101111110"; -- -0.11600092092402237
	pesos_i(19842) := b"1111111111111111_1111111111111111_1110001011001001_1001001000001100"; -- -0.11411177837167902
	pesos_i(19843) := b"1111111111111111_1111111111111111_1111111001111000_1000111001011000"; -- -0.00597296091195888
	pesos_i(19844) := b"0000000000000000_0000000000000000_0000011001110001_0010001010011101"; -- 0.025163806266591596
	pesos_i(19845) := b"0000000000000000_0000000000000000_0010000101100100_1100101010100001"; -- 0.1304442065455378
	pesos_i(19846) := b"1111111111111111_1111111111111111_1110000110000110_0110110100000011"; -- -0.11904257461467212
	pesos_i(19847) := b"0000000000000000_0000000000000000_0000100111100010_1101001000011111"; -- 0.038617260582313725
	pesos_i(19848) := b"0000000000000000_0000000000000000_0010001001111101_1001011011110001"; -- 0.13472884537247592
	pesos_i(19849) := b"1111111111111111_1111111111111111_1101100000101010_1111011110111000"; -- -0.15559436559176898
	pesos_i(19850) := b"0000000000000000_0000000000000000_0001001110000001_0101000100110100"; -- 0.07619197375913406
	pesos_i(19851) := b"0000000000000000_0000000000000000_0010100101011111_1101011100001100"; -- 0.16161865266384862
	pesos_i(19852) := b"1111111111111111_1111111111111111_1110001011001110_0001100111100000"; -- -0.11404264725726562
	pesos_i(19853) := b"1111111111111111_1111111111111111_1110011000100101_1000011000010011"; -- -0.10098993324961009
	pesos_i(19854) := b"1111111111111111_1111111111111111_1111001101101000_0001101111101011"; -- -0.04919267187558883
	pesos_i(19855) := b"0000000000000000_0000000000000000_0001011000001111_0101101001100110"; -- 0.08617177005986107
	pesos_i(19856) := b"0000000000000000_0000000000000000_0010100001110100_1110100100111111"; -- 0.15803392208964154
	pesos_i(19857) := b"0000000000000000_0000000000000000_0001001000000101_0111011000111100"; -- 0.07039584118344115
	pesos_i(19858) := b"0000000000000000_0000000000000000_0001011100000000_0001011100100010"; -- 0.089845128908549
	pesos_i(19859) := b"1111111111111111_1111111111111111_1110011111011101_0000111001001000"; -- -0.09428320636002031
	pesos_i(19860) := b"1111111111111111_1111111111111111_1101111111001011_1110100110100000"; -- -0.12579479066653687
	pesos_i(19861) := b"1111111111111111_1111111111111111_1110011100100111_1101001101100100"; -- -0.09704855736837538
	pesos_i(19862) := b"0000000000000000_0000000000000000_0001101111010100_0011011000010110"; -- 0.10870683698391213
	pesos_i(19863) := b"0000000000000000_0000000000000000_0000101001110000_1010110001101101"; -- 0.04078176165562326
	pesos_i(19864) := b"1111111111111111_1111111111111111_1111011111000001_1001001000101111"; -- -0.03220259048547135
	pesos_i(19865) := b"1111111111111111_1111111111111111_1111100101101110_0010001010101001"; -- -0.025663217334113874
	pesos_i(19866) := b"0000000000000000_0000000000000000_0000100110110010_0110010001101010"; -- 0.03787829948139739
	pesos_i(19867) := b"1111111111111111_1111111111111111_1110101011010010_0010111001011101"; -- -0.08273039089809028
	pesos_i(19868) := b"1111111111111111_1111111111111111_1111011010001110_1000110100111010"; -- -0.036887334180061425
	pesos_i(19869) := b"1111111111111111_1111111111111111_1110001101111100_1010100000001110"; -- -0.11137914325168193
	pesos_i(19870) := b"1111111111111111_1111111111111111_1111011110000001_0111110001100110"; -- -0.03318045150328569
	pesos_i(19871) := b"1111111111111111_1111111111111111_1110111111001010_0111010100100000"; -- -0.06331699342199539
	pesos_i(19872) := b"1111111111111111_1111111111111111_1110111010100111_1010110010001111"; -- -0.06775399689184082
	pesos_i(19873) := b"0000000000000000_0000000000000000_0000010000110101_1111010001110010"; -- 0.01644828589304404
	pesos_i(19874) := b"0000000000000000_0000000000000000_0001110101100111_0010101000110000"; -- 0.11485541978951687
	pesos_i(19875) := b"1111111111111111_1111111111111111_1110010100100011_1001010100011001"; -- -0.10492580541347439
	pesos_i(19876) := b"1111111111111111_1111111111111111_1110101010101011_1110101000100100"; -- -0.08331429130670169
	pesos_i(19877) := b"1111111111111111_1111111111111111_1101111010101011_0001011100100100"; -- -0.13020186782435228
	pesos_i(19878) := b"0000000000000000_0000000000000000_0001100001000101_1010111111111010"; -- 0.09481334541412016
	pesos_i(19879) := b"1111111111111111_1111111111111111_1110101001101101_0100011011111001"; -- -0.08427006162004283
	pesos_i(19880) := b"1111111111111111_1111111111111111_1111001010011001_0111101011111011"; -- -0.05234557504421568
	pesos_i(19881) := b"1111111111111111_1111111111111111_1111011010101110_0101010111001000"; -- -0.036402357712710665
	pesos_i(19882) := b"1111111111111111_1111111111111111_1111000001011101_1101110111010001"; -- -0.06106771123758869
	pesos_i(19883) := b"1111111111111111_1111111111111111_1111101000001001_0100101110101101"; -- -0.02329566015474565
	pesos_i(19884) := b"0000000000000000_0000000000000000_0001010100101101_0011000011000111"; -- 0.08272080292781826
	pesos_i(19885) := b"1111111111111111_1111111111111111_1110001001001000_0101100101110010"; -- -0.1160835357512459
	pesos_i(19886) := b"0000000000000000_0000000000000000_0010010011011110_1011110100101101"; -- 0.14402372695972462
	pesos_i(19887) := b"0000000000000000_0000000000000000_0001110110011001_0000010111001000"; -- 0.11561618926263849
	pesos_i(19888) := b"0000000000000000_0000000000000000_0000111100000011_1001000010011011"; -- 0.05864814541731201
	pesos_i(19889) := b"1111111111111111_1111111111111111_1111111011000011_0101110000011011"; -- -0.004831546217350453
	pesos_i(19890) := b"1111111111111111_1111111111111111_1110111001111100_1100000110001011"; -- -0.06840887420182028
	pesos_i(19891) := b"0000000000000000_0000000000000000_0001111100100010_1100000000101100"; -- 0.12162400318754932
	pesos_i(19892) := b"1111111111111111_1111111111111111_1111110001110010_0010000001111000"; -- -0.013883562840612103
	pesos_i(19893) := b"0000000000000000_0000000000000000_0001101101110101_0101100010100101"; -- 0.10725931194894069
	pesos_i(19894) := b"1111111111111111_1111111111111111_1111000001001101_0011011011010010"; -- -0.061321805651680564
	pesos_i(19895) := b"0000000000000000_0000000000000000_0000011101101101_0111110111110111"; -- 0.02901446611392192
	pesos_i(19896) := b"0000000000000000_0000000000000000_0000010111010100_0011001100110010"; -- 0.022769164705445318
	pesos_i(19897) := b"1111111111111111_1111111111111111_1110101010110111_0001001000111000"; -- -0.08314405577088717
	pesos_i(19898) := b"1111111111111111_1111111111111111_1111110010011111_0111001011000110"; -- -0.013192011425016279
	pesos_i(19899) := b"1111111111111111_1111111111111111_1110011010000010_1111011101001001"; -- -0.09956411802701624
	pesos_i(19900) := b"1111111111111111_1111111111111111_1110110001111100_0111011101001000"; -- -0.07622580047167107
	pesos_i(19901) := b"0000000000000000_0000000000000000_0010000000001101_1110110000011000"; -- 0.12521243650458067
	pesos_i(19902) := b"0000000000000000_0000000000000000_0000111110110010_0111010101010000"; -- 0.061316806709402996
	pesos_i(19903) := b"0000000000000000_0000000000000000_0000000111001100_1000111010001101"; -- 0.007027539623505256
	pesos_i(19904) := b"1111111111111111_1111111111111111_1111001101001001_1001111110100010"; -- -0.04965784358331026
	pesos_i(19905) := b"0000000000000000_0000000000000000_0001001101011110_1101011000000101"; -- 0.07566583271167616
	pesos_i(19906) := b"1111111111111111_1111111111111111_1111000000010001_1010100010000010"; -- -0.06223055683910772
	pesos_i(19907) := b"1111111111111111_1111111111111111_1110110111100101_1000111110010011"; -- -0.07071592950739128
	pesos_i(19908) := b"1111111111111111_1111111111111111_1101111100101101_1111000010010000"; -- -0.12820526591731923
	pesos_i(19909) := b"0000000000000000_0000000000000000_0001001110010100_1011111011000010"; -- 0.07648842089946219
	pesos_i(19910) := b"0000000000000000_0000000000000000_0001111010000000_1000110110011101"; -- 0.11914906588546702
	pesos_i(19911) := b"0000000000000000_0000000000000000_0010001100001101_1001111011000001"; -- 0.13692657679319709
	pesos_i(19912) := b"0000000000000000_0000000000000000_0000100011000111_0010000011111011"; -- 0.03428846484344254
	pesos_i(19913) := b"0000000000000000_0000000000000000_0000111110100100_1100111011111111"; -- 0.0611085293421347
	pesos_i(19914) := b"0000000000000000_0000000000000000_0000100001101100_0100101011010100"; -- 0.032902409414255325
	pesos_i(19915) := b"0000000000000000_0000000000000000_0000010001011000_0100010001000000"; -- 0.0169718414285455
	pesos_i(19916) := b"1111111111111111_1111111111111111_1110001001110110_1101000001011110"; -- -0.115374543284664
	pesos_i(19917) := b"0000000000000000_0000000000000000_0001011001101110_0110100110100111"; -- 0.08762226424261069
	pesos_i(19918) := b"0000000000000000_0000000000000000_0001010010101010_0101111010001011"; -- 0.08072462927032646
	pesos_i(19919) := b"1111111111111111_1111111111111111_1111010001011101_0101110000001110"; -- -0.045450445727984
	pesos_i(19920) := b"0000000000000000_0000000000000000_0001110110010100_0010011100010100"; -- 0.11554187998164665
	pesos_i(19921) := b"1111111111111111_1111111111111111_1110010110000110_1100100111101110"; -- -0.1034120363908495
	pesos_i(19922) := b"0000000000000000_0000000000000000_0000001011101111_0111010000100111"; -- 0.011466273825337913
	pesos_i(19923) := b"1111111111111111_1111111111111111_1111000110111010_0000001001111010"; -- -0.05575546752407868
	pesos_i(19924) := b"0000000000000000_0000000000000000_0001010110101100_0001111101001000"; -- 0.08465762622783281
	pesos_i(19925) := b"1111111111111111_1111111111111111_1110111010001001_0010110110100110"; -- -0.06821932499955309
	pesos_i(19926) := b"0000000000000000_0000000000000000_0000000011000010_0000011101111111"; -- 0.0029606519174041773
	pesos_i(19927) := b"0000000000000000_0000000000000000_0010000111101100_0101100011001100"; -- 0.13251261693782532
	pesos_i(19928) := b"0000000000000000_0000000000000000_0010000100110100_1000110100110110"; -- 0.12970812390952854
	pesos_i(19929) := b"0000000000000000_0000000000000000_0001111000011001_1011101011110100"; -- 0.11758011310300552
	pesos_i(19930) := b"0000000000000000_0000000000000000_0010100101100011_0011110000011110"; -- 0.16167045334728608
	pesos_i(19931) := b"0000000000000000_0000000000000000_0010010011011101_1010100011000101"; -- 0.14400725185295385
	pesos_i(19932) := b"1111111111111111_1111111111111111_1111011001111101_0010010011000100"; -- -0.037152959931546846
	pesos_i(19933) := b"1111111111111111_1111111111111111_1110010100101011_1111000010001100"; -- -0.10479828443406153
	pesos_i(19934) := b"0000000000000000_0000000000000000_0010011111001101_0011111110000110"; -- 0.15547558811211842
	pesos_i(19935) := b"0000000000000000_0000000000000000_0010000101100010_1101010100101011"; -- 0.13041431719877553
	pesos_i(19936) := b"0000000000000000_0000000000000000_0000100001010010_0100110101001011"; -- 0.03250582776110611
	pesos_i(19937) := b"0000000000000000_0000000000000000_0000001100011101_0001110111110000"; -- 0.01216303936342894
	pesos_i(19938) := b"0000000000000000_0000000000000000_0000000110111110_1110011000001110"; -- 0.006819132265433418
	pesos_i(19939) := b"1111111111111111_1111111111111111_1111000100000110_1111010010101001"; -- -0.0584876142822575
	pesos_i(19940) := b"0000000000000000_0000000000000000_0001111011110101_0000000110101000"; -- 0.12092600211339231
	pesos_i(19941) := b"0000000000000000_0000000000000000_0001110011110110_0010000110101011"; -- 0.11313066877136099
	pesos_i(19942) := b"1111111111111111_1111111111111111_1110110011010000_1111100100110110"; -- -0.07493631784574475
	pesos_i(19943) := b"1111111111111111_1111111111111111_1111111100011100_1010010101000100"; -- -0.003469153292017056
	pesos_i(19944) := b"1111111111111111_1111111111111111_1110110010000110_0111011001110011"; -- -0.07607326224611213
	pesos_i(19945) := b"0000000000000000_0000000000000000_0000000110101101_0000000011000110"; -- 0.006546066553240756
	pesos_i(19946) := b"1111111111111111_1111111111111111_1110001111100111_1100001101011011"; -- -0.1097448255751235
	pesos_i(19947) := b"0000000000000000_0000000000000000_0001001010010001_1100010000110101"; -- 0.07253671932587988
	pesos_i(19948) := b"1111111111111111_1111111111111111_1110011111111110_0000000010000110"; -- -0.09378048645189005
	pesos_i(19949) := b"1111111111111111_1111111111111111_1111011001010100_1110100001011001"; -- -0.03776691269305501
	pesos_i(19950) := b"0000000000000000_0000000000000000_0010000100101011_1000110101000101"; -- 0.12957079833844048
	pesos_i(19951) := b"1111111111111111_1111111111111111_1110001111000111_1101001001011111"; -- -0.11023221184501703
	pesos_i(19952) := b"1111111111111111_1111111111111111_1101111011110000_1101110000011100"; -- -0.12913727109050926
	pesos_i(19953) := b"1111111111111111_1111111111111111_1110000110010011_1000000101100110"; -- -0.11884299530985044
	pesos_i(19954) := b"1111111111111111_1111111111111111_1110111100011100_1100010111110110"; -- -0.06596720447047905
	pesos_i(19955) := b"0000000000000000_0000000000000000_0001011100000110_0110100000000010"; -- 0.08994150197822258
	pesos_i(19956) := b"0000000000000000_0000000000000000_0000011110100010_1111011010000110"; -- 0.02983036784037587
	pesos_i(19957) := b"1111111111111111_1111111111111111_1111001101110101_0101101101010011"; -- -0.0489905283922941
	pesos_i(19958) := b"1111111111111111_1111111111111111_1101101000111101_1011110110111011"; -- -0.14749540498374608
	pesos_i(19959) := b"1111111111111111_1111111111111111_1110111001011100_1010110111101010"; -- -0.06889832539204892
	pesos_i(19960) := b"1111111111111111_1111111111111111_1110110100001000_0001001001101111"; -- -0.07409558098695822
	pesos_i(19961) := b"0000000000000000_0000000000000000_0000101011011110_0100111000000001"; -- 0.042454600551246884
	pesos_i(19962) := b"1111111111111111_1111111111111111_1110001010110100_0011010111111000"; -- -0.11443770123462575
	pesos_i(19963) := b"0000000000000000_0000000000000000_0001110111011101_0000110010000111"; -- 0.1166541890024291
	pesos_i(19964) := b"1111111111111111_1111111111111111_1110011110101000_1101011001000101"; -- -0.09508000186347382
	pesos_i(19965) := b"1111111111111111_1111111111111111_1110101111011110_0101001111010001"; -- -0.07863880298052311
	pesos_i(19966) := b"0000000000000000_0000000000000000_0010001101011100_1111101101110011"; -- 0.13813754618098764
	pesos_i(19967) := b"0000000000000000_0000000000000000_0000101000110011_1000111010011000"; -- 0.03984919752830867
	pesos_i(19968) := b"1111111111111111_1111111111111111_1110110100010011_0001001011100110"; -- -0.07392770665503384
	pesos_i(19969) := b"1111111111111111_1111111111111111_1111100001010000_1111010100000110"; -- -0.03001469242143971
	pesos_i(19970) := b"1111111111111111_1111111111111111_1110011111000111_1001101011101100"; -- -0.09461051688804367
	pesos_i(19971) := b"0000000000000000_0000000000000000_0000111100101110_1000001100101011"; -- 0.05930347243292885
	pesos_i(19972) := b"0000000000000000_0000000000000000_0000110011100011_1101010100001100"; -- 0.05035144373553687
	pesos_i(19973) := b"1111111111111111_1111111111111111_1110010011001111_0000011110011000"; -- -0.10621597809554298
	pesos_i(19974) := b"0000000000000000_0000000000000000_0001000110101000_0110000101000001"; -- 0.06897552326600925
	pesos_i(19975) := b"0000000000000000_0000000000000000_0001001000010011_0110011000011110"; -- 0.07060850364291822
	pesos_i(19976) := b"0000000000000000_0000000000000000_0010001101110011_1110011110000100"; -- 0.1384873102607607
	pesos_i(19977) := b"1111111111111111_1111111111111111_1111000000011000_0110001001100101"; -- -0.06212792418996295
	pesos_i(19978) := b"0000000000000000_0000000000000000_0001010101011111_0001101011001110"; -- 0.08348243276065782
	pesos_i(19979) := b"1111111111111111_1111111111111111_1111001010100111_1110101101011110"; -- -0.05212525320585558
	pesos_i(19980) := b"1111111111111111_1111111111111111_1111000110010000_0100010111001100"; -- -0.056392324069637234
	pesos_i(19981) := b"1111111111111111_1111111111111111_1110110011110000_0000010000101011"; -- -0.07446264223479739
	pesos_i(19982) := b"1111111111111111_1111111111111111_1110001101000011_0010101100101010"; -- -0.11225633844226826
	pesos_i(19983) := b"1111111111111111_1111111111111111_1110111101010111_1101100011011010"; -- -0.06506580991447576
	pesos_i(19984) := b"1111111111111111_1111111111111111_1110010000111101_1001011010110010"; -- -0.10843523172300754
	pesos_i(19985) := b"0000000000000000_0000000000000000_0000100111011110_0001100001010010"; -- 0.038545150752136124
	pesos_i(19986) := b"0000000000000000_0000000000000000_0001001101100010_0100010111100111"; -- 0.07571827788367996
	pesos_i(19987) := b"0000000000000000_0000000000000000_0000101000000110_0101011111001001"; -- 0.039159285048732964
	pesos_i(19988) := b"1111111111111111_1111111111111111_1111000100110101_0010010000010111"; -- -0.05778288314386277
	pesos_i(19989) := b"0000000000000000_0000000000000000_0001110011101000_0111101110100100"; -- 0.11292240855049859
	pesos_i(19990) := b"0000000000000000_0000000000000000_0000111111011001_0000000000111011"; -- 0.061904921047099694
	pesos_i(19991) := b"1111111111111111_1111111111111111_1111000111001011_1111100000100001"; -- -0.05548142619152502
	pesos_i(19992) := b"1111111111111111_1111111111111111_1110111111010110_1011001010110010"; -- -0.06313021806050427
	pesos_i(19993) := b"0000000000000000_0000000000000000_0001100110110110_0110100010001100"; -- 0.10043958113618327
	pesos_i(19994) := b"0000000000000000_0000000000000000_0000011001101100_1110001100101001"; -- 0.025098988926989592
	pesos_i(19995) := b"1111111111111111_1111111111111111_1101111010001001_0101000101010101"; -- -0.13071719802272388
	pesos_i(19996) := b"1111111111111111_1111111111111111_1110101110100110_0000000100101101"; -- -0.07949822100866988
	pesos_i(19997) := b"0000000000000000_0000000000000000_0010001001000101_0000001010011010"; -- 0.13386551145566758
	pesos_i(19998) := b"1111111111111111_1111111111111111_1111010110001011_1111000111000010"; -- -0.040833368498003245
	pesos_i(19999) := b"1111111111111111_1111111111111111_1110110100100001_0110010001111011"; -- -0.07370922095320127
	pesos_i(20000) := b"0000000000000000_0000000000000000_0000000110110110_0110100110101011"; -- 0.006689647887875355
	pesos_i(20001) := b"1111111111111111_1111111111111111_1101101000010010_0101011111101010"; -- -0.14815760171593959
	pesos_i(20002) := b"1111111111111111_1111111111111111_1110000111110011_1011101000011111"; -- -0.11737477056366481
	pesos_i(20003) := b"1111111111111111_1111111111111111_1111011110100110_0001001111100110"; -- -0.03262210498764806
	pesos_i(20004) := b"0000000000000000_0000000000000000_0001100011110100_1101110011000101"; -- 0.09748630351563518
	pesos_i(20005) := b"0000000000000000_0000000000000000_0000001101011011_1101110110100110"; -- 0.013120511041623007
	pesos_i(20006) := b"1111111111111111_1111111111111111_1111100110000101_0101100101100010"; -- -0.02530900350552041
	pesos_i(20007) := b"1111111111111111_1111111111111111_1110111011011001_0000111000000010"; -- -0.06700050780955397
	pesos_i(20008) := b"1111111111111111_1111111111111111_1110010001111000_1101100001001101"; -- -0.107531052724309
	pesos_i(20009) := b"0000000000000000_0000000000000000_0001001101101011_0110100010011011"; -- 0.07585767531597037
	pesos_i(20010) := b"1111111111111111_1111111111111111_1111000001010010_1111001011010110"; -- -0.061234305043027216
	pesos_i(20011) := b"0000000000000000_0000000000000000_0001101101111111_0010101000010101"; -- 0.10740912448734045
	pesos_i(20012) := b"1111111111111111_1111111111111111_1101011111101111_1111101110010100"; -- -0.15649440409240678
	pesos_i(20013) := b"1111111111111111_1111111111111111_1110011011100110_1110011010010110"; -- -0.09803923451635488
	pesos_i(20014) := b"1111111111111111_1111111111111111_1111010111101001_1101010100011100"; -- -0.039400749776138576
	pesos_i(20015) := b"0000000000000000_0000000000000000_0010000100011111_1100000001110011"; -- 0.12939074338604584
	pesos_i(20016) := b"1111111111111111_1111111111111111_1111010111000110_1110111101100101"; -- -0.03993324084471828
	pesos_i(20017) := b"1111111111111111_1111111111111111_1110110000101111_1001110011111101"; -- -0.07739847962675428
	pesos_i(20018) := b"0000000000000000_0000000000000000_0000001110111011_0111011001100110"; -- 0.014579200600403533
	pesos_i(20019) := b"0000000000000000_0000000000000000_0000111001010011_1100101101010001"; -- 0.055966098039857
	pesos_i(20020) := b"1111111111111111_1111111111111111_1110001110010101_0111001000010010"; -- -0.11100089119556485
	pesos_i(20021) := b"0000000000000000_0000000000000000_0010010110110111_1111111010101000"; -- 0.14733878715934745
	pesos_i(20022) := b"0000000000000000_0000000000000000_0000100000111101_1110001101111110"; -- 0.03219434579689657
	pesos_i(20023) := b"0000000000000000_0000000000000000_0000011011110101_0011001111101010"; -- 0.027178997697808134
	pesos_i(20024) := b"1111111111111111_1111111111111111_1111111010010001_1100011001101001"; -- -0.005588149486405829
	pesos_i(20025) := b"0000000000000000_0000000000000000_0000010001010100_1010010111001110"; -- 0.016916621047801735
	pesos_i(20026) := b"0000000000000000_0000000000000000_0000101011001010_1010110000001001"; -- 0.042155029479680015
	pesos_i(20027) := b"0000000000000000_0000000000000000_0001111111010110_0011111010111100"; -- 0.12436287006277988
	pesos_i(20028) := b"1111111111111111_1111111111111111_1111100101010111_0010110000100110"; -- -0.026013603878200314
	pesos_i(20029) := b"0000000000000000_0000000000000000_0001010110111001_1101110100101010"; -- 0.08486730826582087
	pesos_i(20030) := b"0000000000000000_0000000000000000_0000001011001111_0111110010100011"; -- 0.010978498287221866
	pesos_i(20031) := b"0000000000000000_0000000000000000_0000011111010111_1001100101000100"; -- 0.030633525066809414
	pesos_i(20032) := b"1111111111111111_1111111111111111_1111001000000111_0100000101010110"; -- -0.054576794177604186
	pesos_i(20033) := b"0000000000000000_0000000000000000_0000000000110000_1111001101010101"; -- 0.0007469256909719506
	pesos_i(20034) := b"1111111111111111_1111111111111111_1111110000010110_1000010110111010"; -- -0.015281335834296087
	pesos_i(20035) := b"1111111111111111_1111111111111111_1110111001101110_1110100111111110"; -- -0.06862008615060847
	pesos_i(20036) := b"0000000000000000_0000000000000000_0001101010111111_0011010111001011"; -- 0.10448013492698617
	pesos_i(20037) := b"0000000000000000_0000000000000000_0010000100110100_1100001100110110"; -- 0.12971134251755545
	pesos_i(20038) := b"0000000000000000_0000000000000000_0001110011011000_0010111001011101"; -- 0.11267366187547877
	pesos_i(20039) := b"1111111111111111_1111111111111111_1110010110100101_1110010011101011"; -- -0.10293740517413201
	pesos_i(20040) := b"1111111111111111_1111111111111111_1110010101110000_0001111011100100"; -- -0.10375792448789346
	pesos_i(20041) := b"1111111111111111_1111111111111111_1111001010101001_0001100100011010"; -- -0.05210726838112803
	pesos_i(20042) := b"1111111111111111_1111111111111111_1101111111001101_0001011010011100"; -- -0.12577685073403688
	pesos_i(20043) := b"0000000000000000_0000000000000000_0001111011101101_1000001101110111"; -- 0.12081166882602751
	pesos_i(20044) := b"0000000000000000_0000000000000000_0010011010001000_1000000100010101"; -- 0.150520389189319
	pesos_i(20045) := b"0000000000000000_0000000000000000_0010010111011111_1110101000111001"; -- 0.1479479208206683
	pesos_i(20046) := b"1111111111111111_1111111111111111_1110000001101111_1110111110001011"; -- -0.12329199649186665
	pesos_i(20047) := b"0000000000000000_0000000000000000_0000110001100100_0000000000111100"; -- 0.04840089298049958
	pesos_i(20048) := b"1111111111111111_1111111111111111_1110100101011101_1001111100011001"; -- -0.08841519970914251
	pesos_i(20049) := b"0000000000000000_0000000000000000_0000011100011101_1110010011111011"; -- 0.027799903263407442
	pesos_i(20050) := b"1111111111111111_1111111111111111_1110110101001011_0110010100111101"; -- -0.07306830663086267
	pesos_i(20051) := b"1111111111111111_1111111111111111_1110010011001011_1000010011111100"; -- -0.10626953932113224
	pesos_i(20052) := b"1111111111111111_1111111111111111_1110100000011001_1001010101100000"; -- -0.093359626930556
	pesos_i(20053) := b"1111111111111111_1111111111111111_1110101100111101_0111101110111100"; -- -0.0810930887109476
	pesos_i(20054) := b"1111111111111111_1111111111111111_1111010001110101_1001100111110011"; -- -0.04508054547736012
	pesos_i(20055) := b"0000000000000000_0000000000000000_0000100000111001_1100111110000101"; -- 0.032132120031577414
	pesos_i(20056) := b"0000000000000000_0000000000000000_0000110100111011_1100010101101100"; -- 0.05169328580780815
	pesos_i(20057) := b"0000000000000000_0000000000000000_0001000111001101_0100001111111111"; -- 0.06953835467460731
	pesos_i(20058) := b"0000000000000000_0000000000000000_0001100100010110_1010000011100111"; -- 0.09800153387206832
	pesos_i(20059) := b"1111111111111111_1111111111111111_1110110111110001_1011100111110100"; -- -0.07053029824391882
	pesos_i(20060) := b"1111111111111111_1111111111111111_1111101000000011_1001100101010011"; -- -0.023382584714868027
	pesos_i(20061) := b"0000000000000000_0000000000000000_0001110000110100_1111110101101001"; -- 0.1101835613684617
	pesos_i(20062) := b"1111111111111111_1111111111111111_1110011111111011_0111000001101110"; -- -0.09381959252545863
	pesos_i(20063) := b"0000000000000000_0000000000000000_0010001000101100_1111001110011010"; -- 0.133498406517994
	pesos_i(20064) := b"0000000000000000_0000000000000000_0001110100100110_1011000110000001"; -- 0.11387166401503275
	pesos_i(20065) := b"0000000000000000_0000000000000000_0001001110010001_0000011001010110"; -- 0.07643165197506492
	pesos_i(20066) := b"0000000000000000_0000000000000000_0001100101111110_1111111111010100"; -- 0.09959410605221534
	pesos_i(20067) := b"1111111111111111_1111111111111111_1111001010010001_1011000111010111"; -- -0.05246437546501223
	pesos_i(20068) := b"0000000000000000_0000000000000000_0000110110111001_0110011101011110"; -- 0.05361028705291106
	pesos_i(20069) := b"1111111111111111_1111111111111111_1101101110100001_1101010011011110"; -- -0.14206189707670142
	pesos_i(20070) := b"1111111111111111_1111111111111111_1110101100101011_0011110010010101"; -- -0.08137151113757352
	pesos_i(20071) := b"0000000000000000_0000000000000000_0000001000000110_1011100111011011"; -- 0.007915130544601766
	pesos_i(20072) := b"1111111111111111_1111111111111111_1110111000000000_1001111111110000"; -- -0.07030296696126784
	pesos_i(20073) := b"1111111111111111_1111111111111111_1101111101100101_1110110110100100"; -- -0.12735094787674112
	pesos_i(20074) := b"1111111111111111_1111111111111111_1110011101111001_0111101110100000"; -- -0.09580256782265469
	pesos_i(20075) := b"1111111111111111_1111111111111111_1111010100111100_0000001001111101"; -- -0.042053074252195975
	pesos_i(20076) := b"0000000000000000_0000000000000000_0001101111000000_0010000101001111"; -- 0.10840042281027933
	pesos_i(20077) := b"0000000000000000_0000000000000000_0010001001001100_1000101101011001"; -- 0.1339804736435106
	pesos_i(20078) := b"0000000000000000_0000000000000000_0010001010011001_1001011111101111"; -- 0.13515615070038856
	pesos_i(20079) := b"1111111111111111_1111111111111111_1101100000101001_0101111100000100"; -- -0.1556187263103982
	pesos_i(20080) := b"1111111111111111_1111111111111111_1111010001100101_1011010001111101"; -- -0.04532310442478617
	pesos_i(20081) := b"0000000000000000_0000000000000000_0001101100100001_1100011001111111"; -- 0.10598412131879426
	pesos_i(20082) := b"0000000000000000_0000000000000000_0001100101100100_0110111010000100"; -- 0.09918871620374511
	pesos_i(20083) := b"1111111111111111_1111111111111111_1110000100111101_1011111100000111"; -- -0.12015157776870676
	pesos_i(20084) := b"0000000000000000_0000000000000000_0000101011011010_0011100011111111"; -- 0.04239231327859045
	pesos_i(20085) := b"1111111111111111_1111111111111111_1111011010000101_1111001010100110"; -- -0.037018618133854625
	pesos_i(20086) := b"1111111111111111_1111111111111111_1111110110101111_0100001011111000"; -- -0.009044470340380006
	pesos_i(20087) := b"1111111111111111_1111111111111111_1111000010001010_0001010100011010"; -- -0.06039302927753326
	pesos_i(20088) := b"0000000000000000_0000000000000000_0010111111100010_1000000111011100"; -- 0.18704997651270708
	pesos_i(20089) := b"1111111111111111_1111111111111111_1110100000001011_1011010101001000"; -- -0.09357134818350543
	pesos_i(20090) := b"0000000000000000_0000000000000000_0000011101011111_1110101100101111"; -- 0.028807353102413388
	pesos_i(20091) := b"1111111111111111_1111111111111111_1110011001000001_0000101011001101"; -- -0.10057003498788074
	pesos_i(20092) := b"0000000000000000_0000000000000000_0000111001000011_0101111111110111"; -- 0.05571555887180132
	pesos_i(20093) := b"0000000000000000_0000000000000000_0000110101000010_0000010001010000"; -- 0.05178858700947626
	pesos_i(20094) := b"0000000000000000_0000000000000000_0000011000001101_1111001011100000"; -- 0.0236503407803703
	pesos_i(20095) := b"0000000000000000_0000000000000000_0010001100101000_0010011001000000"; -- 0.13733138152006857
	pesos_i(20096) := b"1111111111111111_1111111111111111_1110101001111111_0101100011000100"; -- -0.08399434291540964
	pesos_i(20097) := b"1111111111111111_1111111111111111_1111101110000111_0101010110001001"; -- -0.01746621507521224
	pesos_i(20098) := b"1111111111111111_1111111111111111_1101110000001110_0101011101111111"; -- -0.1404061618681166
	pesos_i(20099) := b"0000000000000000_0000000000000000_0001110000001110_1001010111001110"; -- 0.10959755210334035
	pesos_i(20100) := b"1111111111111111_1111111111111111_1111111101001110_0111011100110101"; -- -0.002708959273644444
	pesos_i(20101) := b"1111111111111111_1111111111111111_1101111011101111_0111111011110110"; -- -0.1291580820217621
	pesos_i(20102) := b"0000000000000000_0000000000000000_0010000000100010_0111100010000011"; -- 0.1255259818415328
	pesos_i(20103) := b"0000000000000000_0000000000000000_0001110001100111_0000001011001010"; -- 0.11094682143282257
	pesos_i(20104) := b"1111111111111111_1111111111111111_1110111010110111_0000101101001000"; -- -0.06751946925069598
	pesos_i(20105) := b"1111111111111111_1111111111111111_1110001001010010_0101100010111011"; -- -0.11593099062568984
	pesos_i(20106) := b"0000000000000000_0000000000000000_0000000001110001_0001011010101100"; -- 0.001725594436140147
	pesos_i(20107) := b"1111111111111111_1111111111111111_1110110010011000_1011010011101110"; -- -0.07579487982523306
	pesos_i(20108) := b"1111111111111111_1111111111111111_1110101010011011_1101101101000110"; -- -0.0835593180708248
	pesos_i(20109) := b"1111111111111111_1111111111111111_1111011110111000_1111001000111100"; -- -0.03233419448071671
	pesos_i(20110) := b"0000000000000000_0000000000000000_0001100010110110_1010101000110011"; -- 0.096537244254524
	pesos_i(20111) := b"1111111111111111_1111111111111111_1111111001001100_1110010110011101"; -- -0.006639145903238029
	pesos_i(20112) := b"1111111111111111_1111111111111111_1111110010101000_1001010111000110"; -- -0.013052596354749639
	pesos_i(20113) := b"1111111111111111_1111111111111111_1110000011111011_0011110010011100"; -- -0.12116643138749375
	pesos_i(20114) := b"1111111111111111_1111111111111111_1110110010000110_1101011000011100"; -- -0.07606756034721902
	pesos_i(20115) := b"0000000000000000_0000000000000000_0001110101001101_1100010000101110"; -- 0.11446787008982708
	pesos_i(20116) := b"1111111111111111_1111111111111111_1111001000110101_1011100110111101"; -- -0.053867713329149636
	pesos_i(20117) := b"0000000000000000_0000000000000000_0000110100000100_1101010110010100"; -- 0.050855015372750334
	pesos_i(20118) := b"1111111111111111_1111111111111111_1111110110100010_1111100001100110"; -- -0.009232020519315784
	pesos_i(20119) := b"1111111111111111_1111111111111111_1110010110110110_1111101001110110"; -- -0.10267672183553568
	pesos_i(20120) := b"0000000000000000_0000000000000000_0000110010110111_1101101101000001"; -- 0.04968042703699741
	pesos_i(20121) := b"0000000000000000_0000000000000000_0000000111000110_0111110000111010"; -- 0.006934894687563438
	pesos_i(20122) := b"0000000000000000_0000000000000000_0001001011000111_0101101011100100"; -- 0.07335441657500058
	pesos_i(20123) := b"1111111111111111_1111111111111111_1111110011110010_1001010011110111"; -- -0.011923493970611557
	pesos_i(20124) := b"0000000000000000_0000000000000000_0001001100010110_1100011101011010"; -- 0.07456632571724463
	pesos_i(20125) := b"0000000000000000_0000000000000000_0001110011101000_0011010101010111"; -- 0.1129182182727439
	pesos_i(20126) := b"0000000000000000_0000000000000000_0000101101111000_1001011001010110"; -- 0.04480876547320128
	pesos_i(20127) := b"1111111111111111_1111111111111111_1110111110100011_1111101001001001"; -- -0.06390414932502862
	pesos_i(20128) := b"0000000000000000_0000000000000000_0001001001000001_1011011010100101"; -- 0.07131520779479551
	pesos_i(20129) := b"0000000000000000_0000000000000000_0001111001001010_0101100111010110"; -- 0.11832200507066937
	pesos_i(20130) := b"1111111111111111_1111111111111111_1101010111110010_1110100111000000"; -- -0.1642621903511398
	pesos_i(20131) := b"1111111111111111_1111111111111111_1110100011111001_1111010011100010"; -- -0.0899359654355288
	pesos_i(20132) := b"0000000000000000_0000000000000000_0000000110011011_0001000000100101"; -- 0.0062723245897593136
	pesos_i(20133) := b"1111111111111111_1111111111111111_1111000111011011_0100111011001001"; -- -0.05524737916954381
	pesos_i(20134) := b"0000000000000000_0000000000000000_0000001010001010_0100010101110001"; -- 0.009922351876237547
	pesos_i(20135) := b"0000000000000000_0000000000000000_0001100001111110_1101000111010000"; -- 0.0956851132565851
	pesos_i(20136) := b"1111111111111111_1111111111111111_1101110111010100_1001100101011011"; -- -0.13347474598008602
	pesos_i(20137) := b"1111111111111111_1111111111111111_1101111011100000_0101100011110001"; -- -0.12938923002463926
	pesos_i(20138) := b"1111111111111111_1111111111111111_1101110100111111_1110010100100001"; -- -0.13574378925567349
	pesos_i(20139) := b"0000000000000000_0000000000000000_0001111001001101_0111101010010011"; -- 0.118369732796402
	pesos_i(20140) := b"0000000000000000_0000000000000000_0000001110100000_0001100001011101"; -- 0.014161608315071262
	pesos_i(20141) := b"0000000000000000_0000000000000000_0001011011111110_0101010001011001"; -- 0.089818259851015
	pesos_i(20142) := b"0000000000000000_0000000000000000_0000111001110000_1010111101000010"; -- 0.05640693043930541
	pesos_i(20143) := b"1111111111111111_1111111111111111_1111011010010001_0101101011000100"; -- -0.03684456546606048
	pesos_i(20144) := b"1111111111111111_1111111111111111_1110111001100110_1001111010010010"; -- -0.06874665197209255
	pesos_i(20145) := b"1111111111111111_1111111111111111_1101111001000001_1111100010111111"; -- -0.13180585231649336
	pesos_i(20146) := b"1111111111111111_1111111111111111_1110001010000001_1000010011110110"; -- -0.11521119119419383
	pesos_i(20147) := b"1111111111111111_1111111111111111_1110101000001000_1000101110101110"; -- -0.08580710416553614
	pesos_i(20148) := b"0000000000000000_0000000000000000_0010011000100010_1101000110110100"; -- 0.14896879821689715
	pesos_i(20149) := b"0000000000000000_0000000000000000_0000001110000010_0001101111101111"; -- 0.013704057523486905
	pesos_i(20150) := b"0000000000000000_0000000000000000_0001100001111110_1110010101001111"; -- 0.09568627525522953
	pesos_i(20151) := b"1111111111111111_1111111111111111_1101111110010101_1000111001000110"; -- -0.12662421035226148
	pesos_i(20152) := b"0000000000000000_0000000000000000_0000111111001000_0110001111101101"; -- 0.06165146378210614
	pesos_i(20153) := b"0000000000000000_0000000000000000_0010010101000000_1011101101101001"; -- 0.14551898308943895
	pesos_i(20154) := b"1111111111111111_1111111111111111_1110100101001001_1111110001101100"; -- -0.08871481298672532
	pesos_i(20155) := b"0000000000000000_0000000000000000_0000001000011110_1111101000111111"; -- 0.008285179577517808
	pesos_i(20156) := b"1111111111111111_1111111111111111_1111101100100100_0001100011001110"; -- -0.01898045506841757
	pesos_i(20157) := b"0000000000000000_0000000000000000_0001100011111101_0000010011001000"; -- 0.09761075865939643
	pesos_i(20158) := b"0000000000000000_0000000000000000_0000110111100000_0000101001000110"; -- 0.054199831046709335
	pesos_i(20159) := b"0000000000000000_0000000000000000_0000010000001010_1001000110010111"; -- 0.015786265716333826
	pesos_i(20160) := b"1111111111111111_1111111111111111_1111001110111110_0010101010101011"; -- -0.047879536780266914
	pesos_i(20161) := b"0000000000000000_0000000000000000_0000100101001110_0010010100001010"; -- 0.03634864329359282
	pesos_i(20162) := b"0000000000000000_0000000000000000_0000110011000000_0000100111111110"; -- 0.04980528317906887
	pesos_i(20163) := b"1111111111111111_1111111111111111_1111000010011010_0001010111001111"; -- -0.06014884667415267
	pesos_i(20164) := b"0000000000000000_0000000000000000_0010001001011001_0101110001111110"; -- 0.1341760452844017
	pesos_i(20165) := b"1111111111111111_1111111111111111_1111010101001001_1011000000111111"; -- -0.04184435339429713
	pesos_i(20166) := b"1111111111111111_1111111111111111_1101111101111000_1111111010011110"; -- -0.1270600190100254
	pesos_i(20167) := b"1111111111111111_1111111111111111_1110110001111100_1100100100011101"; -- -0.07622092291622197
	pesos_i(20168) := b"0000000000000000_0000000000000000_0001010100110011_1100011100000010"; -- 0.08282130995189951
	pesos_i(20169) := b"1111111111111111_1111111111111111_1110101101110011_0101101000110110"; -- -0.08027111225066924
	pesos_i(20170) := b"1111111111111111_1111111111111111_1111110110000111_1100011011111000"; -- -0.009646953924755576
	pesos_i(20171) := b"1111111111111111_1111111111111111_1111001000111111_0000110001000011"; -- -0.053725465425549186
	pesos_i(20172) := b"0000000000000000_0000000000000000_0010001100110000_0111111011100000"; -- 0.1374587343183599
	pesos_i(20173) := b"1111111111111111_1111111111111111_1111010000010101_0000101101000010"; -- -0.046553894383982594
	pesos_i(20174) := b"0000000000000000_0000000000000000_0000011101110010_0101100110010010"; -- 0.029088590871284292
	pesos_i(20175) := b"0000000000000000_0000000000000000_0000110010011011_0011001100110000"; -- 0.04924316342373842
	pesos_i(20176) := b"0000000000000000_0000000000000000_0001101111010111_0011011000111100"; -- 0.10875262217996778
	pesos_i(20177) := b"1111111111111111_1111111111111111_1101110110101001_0010101000111101"; -- -0.1341374970454954
	pesos_i(20178) := b"1111111111111111_1111111111111111_1101101001101000_1011110011010000"; -- -0.1468393318091868
	pesos_i(20179) := b"0000000000000000_0000000000000000_0010001011100010_1111110101011010"; -- 0.13627608722541637
	pesos_i(20180) := b"0000000000000000_0000000000000000_0001110100100110_0100110001110111"; -- 0.11386564168556558
	pesos_i(20181) := b"0000000000000000_0000000000000000_0000110101110110_1000111101100001"; -- 0.052590333074408926
	pesos_i(20182) := b"1111111111111111_1111111111111111_1110001001010100_0000110001010011"; -- -0.11590502713394271
	pesos_i(20183) := b"0000000000000000_0000000000000000_0001000011000010_1010110111011111"; -- 0.06547056871063418
	pesos_i(20184) := b"1111111111111111_1111111111111111_1101111011001110_1010101011110110"; -- -0.12965899938867703
	pesos_i(20185) := b"0000000000000000_0000000000000000_0000111010101110_0001000101011101"; -- 0.057343564140091015
	pesos_i(20186) := b"0000000000000000_0000000000000000_0001010101110100_0011000011101010"; -- 0.08380418515248046
	pesos_i(20187) := b"0000000000000000_0000000000000000_0010100001010100_1111010111011101"; -- 0.15754639279131402
	pesos_i(20188) := b"0000000000000000_0000000000000000_0000000001101000_1010000101111011"; -- 0.0015965391516118493
	pesos_i(20189) := b"0000000000000000_0000000000000000_0000100110000111_0011110101111011"; -- 0.03721985115574974
	pesos_i(20190) := b"0000000000000000_0000000000000000_0001011000000000_1111111100101001"; -- 0.08595270871966494
	pesos_i(20191) := b"1111111111111111_1111111111111111_1111000000101101_1101101001111010"; -- -0.06180033217759975
	pesos_i(20192) := b"0000000000000000_0000000000000000_0000100110001001_1110011001000000"; -- 0.037260428092234746
	pesos_i(20193) := b"1111111111111111_1111111111111111_1111010100010010_0011111001101101"; -- -0.04269037092098519
	pesos_i(20194) := b"1111111111111111_1111111111111111_1111111100000001_1110101111000111"; -- -0.0038769377574919377
	pesos_i(20195) := b"1111111111111111_1111111111111111_1110111000001100_1111000010000010"; -- -0.07011505910411929
	pesos_i(20196) := b"1111111111111111_1111111111111111_1111011101010011_1010001100010011"; -- -0.03388005054446724
	pesos_i(20197) := b"1111111111111111_1111111111111111_1101100101101110_1001111011101010"; -- -0.15065581129528408
	pesos_i(20198) := b"0000000000000000_0000000000000000_0000001001001010_0110000111101011"; -- 0.008947486785310722
	pesos_i(20199) := b"1111111111111111_1111111111111111_1101100111110001_1101010001000111"; -- -0.14865372922099723
	pesos_i(20200) := b"0000000000000000_0000000000000000_0010011110110100_1101000100111110"; -- 0.15510280392523557
	pesos_i(20201) := b"1111111111111111_1111111111111111_1110100100001110_0010111110000010"; -- -0.08962729535793224
	pesos_i(20202) := b"0000000000000000_0000000000000000_0001001100101101_0010100011100111"; -- 0.07490783357657926
	pesos_i(20203) := b"0000000000000000_0000000000000000_0010000000010111_0110101000001110"; -- 0.1253572734286355
	pesos_i(20204) := b"0000000000000000_0000000000000000_0010011101010001_1100000111100011"; -- 0.1535912683683658
	pesos_i(20205) := b"0000000000000000_0000000000000000_0001111110011110_0011001000101111"; -- 0.12350762975509834
	pesos_i(20206) := b"1111111111111111_1111111111111111_1101101010011110_0110101011100010"; -- -0.1460202406890414
	pesos_i(20207) := b"0000000000000000_0000000000000000_0001000001000000_0001011110101010"; -- 0.06347797295409949
	pesos_i(20208) := b"1111111111111111_1111111111111111_1110111010111010_1001110110100111"; -- -0.06746496851476637
	pesos_i(20209) := b"0000000000000000_0000000000000000_0010011000011101_0000011100100111"; -- 0.14888043108355442
	pesos_i(20210) := b"1111111111111111_1111111111111111_1111000101000101_0100000111111111"; -- -0.05753695989183731
	pesos_i(20211) := b"0000000000000000_0000000000000000_0000000011100011_0001001100110001"; -- 0.0034648889949514144
	pesos_i(20212) := b"0000000000000000_0000000000000000_0000011000010010_1010101111101111"; -- 0.023722406190406768
	pesos_i(20213) := b"0000000000000000_0000000000000000_0000001010011101_1101111001111101"; -- 0.010221391235604867
	pesos_i(20214) := b"1111111111111111_1111111111111111_1111101010011011_0111110100100000"; -- -0.02106492955322418
	pesos_i(20215) := b"1111111111111111_1111111111111111_1110000101110011_1101111011111101"; -- -0.11932569808634143
	pesos_i(20216) := b"0000000000000000_0000000000000000_0000111100101000_0100111001110001"; -- 0.05920877699371746
	pesos_i(20217) := b"1111111111111111_1111111111111111_1111011011110000_1000001001010100"; -- -0.035392622512037376
	pesos_i(20218) := b"1111111111111111_1111111111111111_1110000111111011_1101100111101010"; -- -0.1172508052382069
	pesos_i(20219) := b"1111111111111111_1111111111111111_1111100001001010_0110010101100000"; -- -0.03011480728228515
	pesos_i(20220) := b"1111111111111111_1111111111111111_1110001111010100_0110001101010000"; -- -0.11004046716971981
	pesos_i(20221) := b"0000000000000000_0000000000000000_0000000111100010_0010010010100101"; -- 0.007356920619983224
	pesos_i(20222) := b"0000000000000000_0000000000000000_0000001101011011_1010110111110010"; -- 0.013117667704704952
	pesos_i(20223) := b"0000000000000000_0000000000000000_0001001100000001_0000100111001111"; -- 0.0742345935197926
	pesos_i(20224) := b"1111111111111111_1111111111111111_1101110001010111_0111101111010111"; -- -0.13929010381962997
	pesos_i(20225) := b"1111111111111111_1111111111111111_1111110010111001_0110011000100100"; -- -0.01279603591490686
	pesos_i(20226) := b"0000000000000000_0000000000000000_0010010111110001_1001010001100000"; -- 0.14821746193114194
	pesos_i(20227) := b"0000000000000000_0000000000000000_0000111101100110_1111111100111100"; -- 0.06016535962756017
	pesos_i(20228) := b"0000000000000000_0000000000000000_0001111010011011_1100001001011010"; -- 0.11956419659043509
	pesos_i(20229) := b"1111111111111111_1111111111111111_1110011101100111_0101111111001011"; -- -0.09607888497559801
	pesos_i(20230) := b"0000000000000000_0000000000000000_0000101011111010_0010011111000010"; -- 0.04287956702998573
	pesos_i(20231) := b"0000000000000000_0000000000000000_0000000010011000_0000000011011010"; -- 0.002319386659474727
	pesos_i(20232) := b"1111111111111111_1111111111111111_1110110100001111_1001011110100000"; -- -0.07398083055012226
	pesos_i(20233) := b"0000000000000000_0000000000000000_0000011000110111_1000011111100111"; -- 0.024284833911582145
	pesos_i(20234) := b"1111111111111111_1111111111111111_1110001100100110_0101010100000111"; -- -0.11269634789835091
	pesos_i(20235) := b"1111111111111111_1111111111111111_1111110100101011_1011011110001000"; -- -0.011051682711438688
	pesos_i(20236) := b"0000000000000000_0000000000000000_0000010001111001_1110001010111100"; -- 0.01748482794977443
	pesos_i(20237) := b"1111111111111111_1111111111111111_1111101010011010_1111100011100001"; -- -0.021072812130835603
	pesos_i(20238) := b"1111111111111111_1111111111111111_1110011010010101_0010101110101111"; -- -0.0992863366136257
	pesos_i(20239) := b"1111111111111111_1111111111111111_1101100100110110_1101111011011101"; -- -0.15150649161492535
	pesos_i(20240) := b"0000000000000000_0000000000000000_0010010011101010_0101001110001001"; -- 0.14420053565327878
	pesos_i(20241) := b"1111111111111111_1111111111111111_1111010111010110_1000101110011010"; -- -0.03969504835535005
	pesos_i(20242) := b"1111111111111111_1111111111111111_1111001110000110_1011101010000100"; -- -0.048725454964091135
	pesos_i(20243) := b"1111111111111111_1111111111111111_1111010100001110_0111111100110011"; -- -0.042747545247667044
	pesos_i(20244) := b"0000000000000000_0000000000000000_0001111001111010_0100010111010101"; -- 0.11905323455263146
	pesos_i(20245) := b"0000000000000000_0000000000000000_0001010000011101_1111000111010100"; -- 0.07858191901508405
	pesos_i(20246) := b"1111111111111111_1111111111111111_1111100001001001_1000100011010101"; -- -0.030127952671508706
	pesos_i(20247) := b"1111111111111111_1111111111111111_1111110000110010_0110100011100010"; -- -0.01485580903369803
	pesos_i(20248) := b"1111111111111111_1111111111111111_1111100011001011_0100011100101001"; -- -0.028148224242704932
	pesos_i(20249) := b"1111111111111111_1111111111111111_1110100001110110_0100101110101001"; -- -0.09194495323533601
	pesos_i(20250) := b"1111111111111111_1111111111111111_1111001101000101_0001111001011111"; -- -0.0497265832623545
	pesos_i(20251) := b"1111111111111111_1111111111111111_1110100000001110_0100111010101110"; -- -0.09353168725890722
	pesos_i(20252) := b"1111111111111111_1111111111111111_1111101101001001_0101011001111010"; -- -0.018412203955716508
	pesos_i(20253) := b"0000000000000000_0000000000000000_0001000100011110_1011110000110010"; -- 0.06687523108763097
	pesos_i(20254) := b"0000000000000000_0000000000000000_0000110010000111_1101111010100110"; -- 0.04894820736150084
	pesos_i(20255) := b"0000000000000000_0000000000000000_0001111011100010_1101010111000000"; -- 0.12064872677072061
	pesos_i(20256) := b"1111111111111111_1111111111111111_1111010010101100_1001010100100010"; -- -0.044241599361254894
	pesos_i(20257) := b"1111111111111111_1111111111111111_1110001011011101_1110111001001111"; -- -0.11380110342257177
	pesos_i(20258) := b"0000000000000000_0000000000000000_0000100011100110_0000100000010011"; -- 0.03476000274045191
	pesos_i(20259) := b"1111111111111111_1111111111111111_1111001101000101_1001001011111101"; -- -0.04971963228714959
	pesos_i(20260) := b"1111111111111111_1111111111111111_1111100001001110_0010110101001100"; -- -0.03005711460096789
	pesos_i(20261) := b"0000000000000000_0000000000000000_0000100001010011_0100001111011001"; -- 0.03252052362396011
	pesos_i(20262) := b"1111111111111111_1111111111111111_1110000011100010_0101011110000111"; -- -0.12154629660200844
	pesos_i(20263) := b"1111111111111111_1111111111111111_1110110011100100_0001000110000110"; -- -0.07464495150379538
	pesos_i(20264) := b"1111111111111111_1111111111111111_1110001010011010_1000000111010001"; -- -0.11482990893341564
	pesos_i(20265) := b"1111111111111111_1111111111111111_1110000000101010_0001100000010101"; -- -0.12435769545406314
	pesos_i(20266) := b"1111111111111111_1111111111111111_1101111011001000_1010101011110111"; -- -0.12975055193635
	pesos_i(20267) := b"1111111111111111_1111111111111111_1110110100111001_0111100001001010"; -- -0.07334182931572251
	pesos_i(20268) := b"1111111111111111_1111111111111111_1111110101110011_0100001010110001"; -- -0.009960014201401133
	pesos_i(20269) := b"0000000000000000_0000000000000000_0010011111110101_0011001111001010"; -- 0.1560852401283342
	pesos_i(20270) := b"0000000000000000_0000000000000000_0000100110110100_0000111001011111"; -- 0.03790368855580414
	pesos_i(20271) := b"1111111111111111_1111111111111111_1110101111111001_1000101001010111"; -- -0.07822356586146254
	pesos_i(20272) := b"1111111111111111_1111111111111111_1110010010001011_0101100001110101"; -- -0.1072487559526399
	pesos_i(20273) := b"1111111111111111_1111111111111111_1110001111101010_0001001101110000"; -- -0.10970953486060996
	pesos_i(20274) := b"0000000000000000_0000000000000000_0000111110011010_0101111001101001"; -- 0.060949230705590794
	pesos_i(20275) := b"0000000000000000_0000000000000000_0001010011001000_0010111111110000"; -- 0.08117961514933049
	pesos_i(20276) := b"1111111111111111_1111111111111111_1101111010000011_0111000011101111"; -- -0.1308068672219929
	pesos_i(20277) := b"0000000000000000_0000000000000000_0001001000111001_0100110101010111"; -- 0.07118686085582637
	pesos_i(20278) := b"0000000000000000_0000000000000000_0000111000010000_1101001110110111"; -- 0.05494425978766673
	pesos_i(20279) := b"1111111111111111_1111111111111111_1101111011100101_0111101011011111"; -- -0.12931091354096735
	pesos_i(20280) := b"1111111111111111_1111111111111111_1111101111100100_1111001110101110"; -- -0.01603772163671189
	pesos_i(20281) := b"0000000000000000_0000000000000000_0000010010000110_0010011111011110"; -- 0.01767205399475134
	pesos_i(20282) := b"1111111111111111_1111111111111111_1110111101001000_0001010011101100"; -- -0.06530637022221897
	pesos_i(20283) := b"1111111111111111_1111111111111111_1111000000011000_1001110100000010"; -- -0.06212443076593865
	pesos_i(20284) := b"0000000000000000_0000000000000000_0001110011110011_0000110100110111"; -- 0.11308367345947591
	pesos_i(20285) := b"1111111111111111_1111111111111111_1110011000110111_1111010010111111"; -- -0.10070867854410485
	pesos_i(20286) := b"1111111111111111_1111111111111111_1111100101011100_1101100111111110"; -- -0.025926948073756836
	pesos_i(20287) := b"1111111111111111_1111111111111111_1111110101011000_1100101110011101"; -- -0.010363840270058223
	pesos_i(20288) := b"1111111111111111_1111111111111111_1111000000111001_0010100100011010"; -- -0.061627799228163735
	pesos_i(20289) := b"0000000000000000_0000000000000000_0000010100110111_0100100110101110"; -- 0.02037487510178461
	pesos_i(20290) := b"0000000000000000_0000000000000000_0000000011110000_0001110111111000"; -- 0.003663895661113211
	pesos_i(20291) := b"0000000000000000_0000000000000000_0000000000110011_0111110101011110"; -- 0.0007856706379126546
	pesos_i(20292) := b"1111111111111111_1111111111111111_1110101010110110_0001111000111101"; -- -0.08315859814809225
	pesos_i(20293) := b"0000000000000000_0000000000000000_0010010100111010_0011000100101110"; -- 0.14541919103695378
	pesos_i(20294) := b"1111111111111111_1111111111111111_1110011101011011_0110000101000000"; -- -0.09626190368092138
	pesos_i(20295) := b"0000000000000000_0000000000000000_0010011101001011_1101011100000101"; -- 0.15350097527537082
	pesos_i(20296) := b"1111111111111111_1111111111111111_1111111001011011_1100111101000000"; -- -0.006411597146509715
	pesos_i(20297) := b"0000000000000000_0000000000000000_0001101101101000_1111101111001011"; -- 0.10707067204481001
	pesos_i(20298) := b"1111111111111111_1111111111111111_1101101010001010_1111110011011001"; -- -0.14631671613823063
	pesos_i(20299) := b"1111111111111111_1111111111111111_1101111000101110_1111000010101001"; -- -0.1320962512797472
	pesos_i(20300) := b"0000000000000000_0000000000000000_0000110101111000_1101001111000110"; -- 0.05262492741504896
	pesos_i(20301) := b"0000000000000000_0000000000000000_0010011011000010_0110000100110110"; -- 0.15140349933685582
	pesos_i(20302) := b"0000000000000000_0000000000000000_0001000101000111_0001000111011101"; -- 0.06749068878628363
	pesos_i(20303) := b"1111111111111111_1111111111111111_1111110010001100_1010110110001001"; -- -0.013478426063839928
	pesos_i(20304) := b"1111111111111111_1111111111111111_1110110100100001_1101011101011101"; -- -0.07370237320091552
	pesos_i(20305) := b"0000000000000000_0000000000000000_0001100111101000_0001010101001100"; -- 0.10119755849718436
	pesos_i(20306) := b"1111111111111111_1111111111111111_1110111001000010_1101110011011111"; -- -0.06929225506880335
	pesos_i(20307) := b"0000000000000000_0000000000000000_0001010111101000_1111101111100100"; -- 0.085586302852636
	pesos_i(20308) := b"1111111111111111_1111111111111111_1101101101110101_1100110000101010"; -- -0.14273380255203436
	pesos_i(20309) := b"0000000000000000_0000000000000000_0000111010110000_0001010100111001"; -- 0.05737431180625914
	pesos_i(20310) := b"1111111111111111_1111111111111111_1111110111011101_1011111111001010"; -- -0.008335126182717404
	pesos_i(20311) := b"0000000000000000_0000000000000000_0000000110111101_0110100010001100"; -- 0.00679639259159377
	pesos_i(20312) := b"1111111111111111_1111111111111111_1110010011010000_0011100000101111"; -- -0.10619782311153565
	pesos_i(20313) := b"0000000000000000_0000000000000000_0001101101110111_1111000011011001"; -- 0.10729890143139924
	pesos_i(20314) := b"1111111111111111_1111111111111111_1110100110111111_1010010000011011"; -- -0.08691953980991297
	pesos_i(20315) := b"0000000000000000_0000000000000000_0000100101101001_0000110111010000"; -- 0.036759246199072344
	pesos_i(20316) := b"0000000000000000_0000000000000000_0000011100101000_0101001010110101"; -- 0.027959031216468422
	pesos_i(20317) := b"0000000000000000_0000000000000000_0001111010111001_0110001001010100"; -- 0.12001623680399617
	pesos_i(20318) := b"1111111111111111_1111111111111111_1111001000010010_1111101100001100"; -- -0.05439787824527727
	pesos_i(20319) := b"1111111111111111_1111111111111111_1110101111001111_0011100101000101"; -- -0.07886926708946865
	pesos_i(20320) := b"0000000000000000_0000000000000000_0000110000010011_0010101111100001"; -- 0.047167532283200794
	pesos_i(20321) := b"1111111111111111_1111111111111111_1101101011101110_0000011001000101"; -- -0.1448055344865929
	pesos_i(20322) := b"0000000000000000_0000000000000000_0000101010000110_0101101101100001"; -- 0.04111262432592742
	pesos_i(20323) := b"1111111111111111_1111111111111111_1111011011101001_0000110000001010"; -- -0.035506484513330695
	pesos_i(20324) := b"0000000000000000_0000000000000000_0010010110110110_1101011010111110"; -- 0.14732114923396383
	pesos_i(20325) := b"0000000000000000_0000000000000000_0000111111011010_0000111000010001"; -- 0.061921004348578335
	pesos_i(20326) := b"0000000000000000_0000000000000000_0010000111110001_1010000100000100"; -- 0.13259321542253402
	pesos_i(20327) := b"0000000000000000_0000000000000000_0000010111100011_0101011110111010"; -- 0.023000224054859943
	pesos_i(20328) := b"0000000000000000_0000000000000000_0001110101100011_0111010101111110"; -- 0.11479887329974724
	pesos_i(20329) := b"1111111111111111_1111111111111111_1110101010000001_1010111001000011"; -- -0.08395872933948155
	pesos_i(20330) := b"0000000000000000_0000000000000000_0000110110110111_0011010000101001"; -- 0.053576717443080416
	pesos_i(20331) := b"0000000000000000_0000000000000000_0001000100001010_0100100110111010"; -- 0.06656323243680913
	pesos_i(20332) := b"0000000000000000_0000000000000000_0001110101101111_0111100111110100"; -- 0.11498224466909035
	pesos_i(20333) := b"1111111111111111_1111111111111111_1110101110011111_0001111001000101"; -- -0.07960329833130568
	pesos_i(20334) := b"1111111111111111_1111111111111111_1101110110000110_0000111111010101"; -- -0.13467312856008107
	pesos_i(20335) := b"0000000000000000_0000000000000000_0001100011001111_0001110010000100"; -- 0.09691026890252
	pesos_i(20336) := b"1111111111111111_1111111111111111_1110100010011000_0000100100101111"; -- -0.09143011678485877
	pesos_i(20337) := b"0000000000000000_0000000000000000_0001110110001011_1000100001101101"; -- 0.11541035326676606
	pesos_i(20338) := b"0000000000000000_0000000000000000_0001000011011101_1010100010101000"; -- 0.06588224497868359
	pesos_i(20339) := b"1111111111111111_1111111111111111_1110111010100101_1100111001000100"; -- -0.06778250545765895
	pesos_i(20340) := b"0000000000000000_0000000000000000_0010000110001101_1101000100000101"; -- 0.13107019770074388
	pesos_i(20341) := b"0000000000000000_0000000000000000_0000011010101110_1000010101111000"; -- 0.026100484600042866
	pesos_i(20342) := b"0000000000000000_0000000000000000_0001001010111111_1101100000000110"; -- 0.07323980462906829
	pesos_i(20343) := b"0000000000000000_0000000000000000_0000010100011100_1011110010011100"; -- 0.019969738169894134
	pesos_i(20344) := b"1111111111111111_1111111111111111_1111111101100110_0110101011010001"; -- -0.0023434867042919877
	pesos_i(20345) := b"1111111111111111_1111111111111111_1110100001010111_0100110111100000"; -- -0.09241784375145445
	pesos_i(20346) := b"1111111111111111_1111111111111111_1111101000010111_0110101010100011"; -- -0.023080191750958972
	pesos_i(20347) := b"0000000000000000_0000000000000000_0001111100001000_0011110010111011"; -- 0.12121944023957724
	pesos_i(20348) := b"0000000000000000_0000000000000000_0000001101111000_0101010011100011"; -- 0.01355486443335801
	pesos_i(20349) := b"1111111111111111_1111111111111111_1111101101000110_0101110000010101"; -- -0.01845764629404439
	pesos_i(20350) := b"1111111111111111_1111111111111111_1110100011101101_0100010000001111"; -- -0.09012961035241415
	pesos_i(20351) := b"1111111111111111_1111111111111111_1110100001100110_0100111001101110"; -- -0.09218892865767786
	pesos_i(20352) := b"1111111111111111_1111111111111111_1111111111000110_0010000100111000"; -- -0.000883029685890461
	pesos_i(20353) := b"0000000000000000_0000000000000000_0000011111110000_1110111101011110"; -- 0.03102012687652733
	pesos_i(20354) := b"0000000000000000_0000000000000000_0000001100000001_0000110011010010"; -- 0.01173477290125657
	pesos_i(20355) := b"1111111111111111_1111111111111111_1110100001001000_0010101111011100"; -- -0.09264875297744633
	pesos_i(20356) := b"0000000000000000_0000000000000000_0000110011110010_1011111010001011"; -- 0.05057898423932883
	pesos_i(20357) := b"0000000000000000_0000000000000000_0010001001101111_0101011010001101"; -- 0.13451138443164906
	pesos_i(20358) := b"1111111111111111_1111111111111111_1110100001001010_0001011100110001"; -- -0.0926194672275297
	pesos_i(20359) := b"1111111111111111_1111111111111111_1110100001010100_0110000000000000"; -- -0.09246253978165418
	pesos_i(20360) := b"0000000000000000_0000000000000000_0000101001010100_0111101000101001"; -- 0.04035151962768977
	pesos_i(20361) := b"1111111111111111_1111111111111111_1110011110110001_0100001111000000"; -- -0.09495140607438948
	pesos_i(20362) := b"0000000000000000_0000000000000000_0001000110100011_1011111001100101"; -- 0.0689047809706491
	pesos_i(20363) := b"1111111111111111_1111111111111111_1101111010101111_1001011111011110"; -- -0.13013316003755773
	pesos_i(20364) := b"1111111111111111_1111111111111111_1110100100011111_1010101100100101"; -- -0.0893605266329569
	pesos_i(20365) := b"0000000000000000_0000000000000000_0001111010010110_1110101010000010"; -- 0.11949029621411575
	pesos_i(20366) := b"1111111111111111_1111111111111111_1111011100000001_0110110100100001"; -- -0.03513448651155843
	pesos_i(20367) := b"1111111111111111_1111111111111111_1110100100111111_1011011101100101"; -- -0.08887151511518523
	pesos_i(20368) := b"1111111111111111_1111111111111111_1110001110101001_1000101000011100"; -- -0.11069428275733818
	pesos_i(20369) := b"0000000000000000_0000000000000000_0001000111000011_0011000011111101"; -- 0.06938463370814978
	pesos_i(20370) := b"0000000000000000_0000000000000000_0001111100110000_1100100100101010"; -- 0.12183816224082036
	pesos_i(20371) := b"0000000000000000_0000000000000000_0000110100110100_0010110100110000"; -- 0.05157740036551992
	pesos_i(20372) := b"0000000000000000_0000000000000000_0001011110011000_1101010011110101"; -- 0.09217577916185381
	pesos_i(20373) := b"1111111111111111_1111111111111111_1111110100011000_1011010001011001"; -- -0.011341789539068142
	pesos_i(20374) := b"0000000000000000_0000000000000000_0001010000011010_1010011101100000"; -- 0.07853170482441613
	pesos_i(20375) := b"1111111111111111_1111111111111111_1110011001001100_0101100001001010"; -- -0.10039756964107112
	pesos_i(20376) := b"0000000000000000_0000000000000000_0001101110101101_1100110000100001"; -- 0.10812068753946048
	pesos_i(20377) := b"1111111111111111_1111111111111111_1110110100111100_1100010011001000"; -- -0.07329149354029235
	pesos_i(20378) := b"1111111111111111_1111111111111111_1111100110010110_1010000101101100"; -- -0.025045310068097203
	pesos_i(20379) := b"0000000000000000_0000000000000000_0010000010100010_1111110001010100"; -- 0.12748696370178425
	pesos_i(20380) := b"1111111111111111_1111111111111111_1111101101000011_0000010100110001"; -- -0.018508601814437833
	pesos_i(20381) := b"1111111111111111_1111111111111111_1110011110111111_0111011100000100"; -- -0.09473472737893951
	pesos_i(20382) := b"0000000000000000_0000000000000000_0000001111111101_1011110010111010"; -- 0.015590472728288294
	pesos_i(20383) := b"0000000000000000_0000000000000000_0010001000010010_1101000110011110"; -- 0.13309965235527288
	pesos_i(20384) := b"0000000000000000_0000000000000000_0010010001001110_0100000110000011"; -- 0.14181909033751383
	pesos_i(20385) := b"1111111111111111_1111111111111111_1111110011111010_0101011011011100"; -- -0.011805125453988102
	pesos_i(20386) := b"1111111111111111_1111111111111111_1110110110000011_0111101010100110"; -- -0.07221253826768559
	pesos_i(20387) := b"1111111111111111_1111111111111111_1111010100101000_0110110110011010"; -- -0.04235186558423368
	pesos_i(20388) := b"1111111111111111_1111111111111111_1110010011111011_1001111001011010"; -- -0.10553560540679377
	pesos_i(20389) := b"1111111111111111_1111111111111111_1101101110010111_1010001110001101"; -- -0.14221742448065758
	pesos_i(20390) := b"1111111111111111_1111111111111111_1111010101100100_0110100110010010"; -- -0.04143657860409897
	pesos_i(20391) := b"0000000000000000_0000000000000000_0000100000100010_1100100111011101"; -- 0.03178083088381882
	pesos_i(20392) := b"0000000000000000_0000000000000000_0010000101011000_1000000011010000"; -- 0.1302567011865894
	pesos_i(20393) := b"1111111111111111_1111111111111111_1110011000110001_1010000000101100"; -- -0.10080527241936622
	pesos_i(20394) := b"0000000000000000_0000000000000000_0000000011101010_0101011111100000"; -- 0.00357579438327653
	pesos_i(20395) := b"1111111111111111_1111111111111111_1111110111011101_0101111110100111"; -- -0.008340856241776079
	pesos_i(20396) := b"1111111111111111_1111111111111111_1110111000111101_0101010100001000"; -- -0.06937664572379375
	pesos_i(20397) := b"1111111111111111_1111111111111111_1111110100011001_1011001001010010"; -- -0.011326651640684957
	pesos_i(20398) := b"0000000000000000_0000000000000000_0000100010111101_1111100011010100"; -- 0.034148742550123574
	pesos_i(20399) := b"0000000000000000_0000000000000000_0010010101001100_1010101111111110"; -- 0.14570116946657832
	pesos_i(20400) := b"0000000000000000_0000000000000000_0010010011010011_1101010110000001"; -- 0.1438573304131274
	pesos_i(20401) := b"0000000000000000_0000000000000000_0010001010011010_1111100111100111"; -- 0.13517724895607655
	pesos_i(20402) := b"0000000000000000_0000000000000000_0010000110010010_0001111010001011"; -- 0.13113585361800337
	pesos_i(20403) := b"0000000000000000_0000000000000000_0001101110001110_0100010001011111"; -- 0.10763957316683816
	pesos_i(20404) := b"0000000000000000_0000000000000000_0000111111011100_1000111110001000"; -- 0.061959238619635544
	pesos_i(20405) := b"0000000000000000_0000000000000000_0001010111001101_1111110011101100"; -- 0.08517437707596598
	pesos_i(20406) := b"1111111111111111_1111111111111111_1110101100000000_1110001111011011"; -- -0.08201766880556541
	pesos_i(20407) := b"0000000000000000_0000000000000000_0001111111101011_1011111111000110"; -- 0.12469099611489319
	pesos_i(20408) := b"0000000000000000_0000000000000000_0000000101010101_1010011010100110"; -- 0.005213180034136081
	pesos_i(20409) := b"0000000000000000_0000000000000000_0001111101110101_0010100110110010"; -- 0.12288151354919029
	pesos_i(20410) := b"0000000000000000_0000000000000000_0001100101011011_0110101101101101"; -- 0.09905120294810599
	pesos_i(20411) := b"1111111111111111_1111111111111111_1111011010000011_1010101111110010"; -- -0.03705334984195525
	pesos_i(20412) := b"1111111111111111_1111111111111111_1110111001001111_0011100110111100"; -- -0.06910361443029508
	pesos_i(20413) := b"1111111111111111_1111111111111111_1101110100001011_1100010110100010"; -- -0.13653912358263146
	pesos_i(20414) := b"0000000000000000_0000000000000000_0000011000000010_0000011100100111"; -- 0.02346844381316397
	pesos_i(20415) := b"0000000000000000_0000000000000000_0010010100100011_0101010011100001"; -- 0.14507036689526534
	pesos_i(20416) := b"0000000000000000_0000000000000000_0000010100000000_1101100010101101"; -- 0.019544164942572356
	pesos_i(20417) := b"1111111111111111_1111111111111111_1110001101001111_1111011011010111"; -- -0.11206109295654945
	pesos_i(20418) := b"0000000000000000_0000000000000000_0000100001010001_1010011100010111"; -- 0.03249592121985266
	pesos_i(20419) := b"0000000000000000_0000000000000000_0010010100011101_0100111100011101"; -- 0.14497847035192374
	pesos_i(20420) := b"0000000000000000_0000000000000000_0010011100000101_1110100101100000"; -- 0.1524339542289894
	pesos_i(20421) := b"0000000000000000_0000000000000000_0000011001111100_1001100111111011"; -- 0.025338767772098692
	pesos_i(20422) := b"1111111111111111_1111111111111111_1110010010111100_1111111101101011"; -- -0.10649112349764933
	pesos_i(20423) := b"1111111111111111_1111111111111111_1101110101100101_0010111000010001"; -- -0.13517486661143124
	pesos_i(20424) := b"1111111111111111_1111111111111111_1111100111101111_1010010110011000"; -- -0.02368702917417109
	pesos_i(20425) := b"0000000000000000_0000000000000000_0001001000101010_0011000110111001"; -- 0.07095633292661319
	pesos_i(20426) := b"1111111111111111_1111111111111111_1111100010100001_0100100111100001"; -- -0.028788931391395347
	pesos_i(20427) := b"0000000000000000_0000000000000000_0010011000110010_0100100011000101"; -- 0.14920477682790992
	pesos_i(20428) := b"1111111111111111_1111111111111111_1111110110001010_1011111001000000"; -- -0.009601697299122627
	pesos_i(20429) := b"1111111111111111_1111111111111111_1111101001110111_0000100110100101"; -- -0.02162112931989218
	pesos_i(20430) := b"1111111111111111_1111111111111111_1111110100011100_1011110101000011"; -- -0.011280222986993469
	pesos_i(20431) := b"0000000000000000_0000000000000000_0010000110001011_0110110001010001"; -- 0.13103367794968748
	pesos_i(20432) := b"0000000000000000_0000000000000000_0000001100111001_0111001111001010"; -- 0.01259540262540608
	pesos_i(20433) := b"0000000000000000_0000000000000000_0001110011001110_1011111000111110"; -- 0.11252964988402803
	pesos_i(20434) := b"1111111111111111_1111111111111111_1111110001100101_0111110001001111"; -- -0.01407645293244973
	pesos_i(20435) := b"1111111111111111_1111111111111111_1111100011010110_1100101011111111"; -- -0.02797251968688095
	pesos_i(20436) := b"0000000000000000_0000000000000000_0010011011111011_0110011010011010"; -- 0.1522735716838682
	pesos_i(20437) := b"1111111111111111_1111111111111111_1110010011010110_1111010000010010"; -- -0.10609507142100827
	pesos_i(20438) := b"0000000000000000_0000000000000000_0010000111110011_0110100010010101"; -- 0.13262036924151763
	pesos_i(20439) := b"1111111111111111_1111111111111111_1110000000100110_1000110010000110"; -- -0.12441179014292568
	pesos_i(20440) := b"1111111111111111_1111111111111111_1110000111101100_1001111011100010"; -- -0.11748320572764442
	pesos_i(20441) := b"0000000000000000_0000000000000000_0010010100100000_0001011110110011"; -- 0.14502094380854752
	pesos_i(20442) := b"1111111111111111_1111111111111111_1101101100101111_0110001110101011"; -- -0.14380814631599353
	pesos_i(20443) := b"1111111111111111_1111111111111111_1110101101101100_0001001000001001"; -- -0.08038222574245583
	pesos_i(20444) := b"1111111111111111_1111111111111111_1110111100111000_1001010111000000"; -- -0.06554283205403312
	pesos_i(20445) := b"0000000000000000_0000000000000000_0000001011100011_1000001010001111"; -- 0.01128402700918243
	pesos_i(20446) := b"0000000000000000_0000000000000000_0000110001100110_1001001011100000"; -- 0.048440150938245295
	pesos_i(20447) := b"0000000000000000_0000000000000000_0000010101100101_0110001101110110"; -- 0.021078316117729274
	pesos_i(20448) := b"1111111111111111_1111111111111111_1101110101101011_0000110011000001"; -- -0.13508529935422614
	pesos_i(20449) := b"0000000000000000_0000000000000000_0010001001100101_0101100011101100"; -- 0.13435893774315638
	pesos_i(20450) := b"1111111111111111_1111111111111111_1111000000010010_1000010000000010"; -- -0.06221747344135856
	pesos_i(20451) := b"1111111111111111_1111111111111111_1110101111010001_0010111110110101"; -- -0.07883931954736938
	pesos_i(20452) := b"1111111111111111_1111111111111111_1110001100101010_1101110011110001"; -- -0.11262721166900691
	pesos_i(20453) := b"1111111111111111_1111111111111111_1111101000011001_0010011100110011"; -- -0.02305369376373865
	pesos_i(20454) := b"1111111111111111_1111111111111111_1101110101001110_1001100100001011"; -- -0.13551944242882855
	pesos_i(20455) := b"0000000000000000_0000000000000000_0001101010100011_1010100000100001"; -- 0.10405970396485446
	pesos_i(20456) := b"0000000000000000_0000000000000000_0000100010111001_1011100000101010"; -- 0.03408385304581448
	pesos_i(20457) := b"0000000000000000_0000000000000000_0010010110100110_0100000111111110"; -- 0.14706814246516522
	pesos_i(20458) := b"0000000000000000_0000000000000000_0000011101111100_1001000111111001"; -- 0.029244540565281706
	pesos_i(20459) := b"1111111111111111_1111111111111111_1101011110110011_0011000100001111"; -- -0.15742200259307174
	pesos_i(20460) := b"1111111111111111_1111111111111111_1110111111000100_1110111000110010"; -- -0.06340132989895654
	pesos_i(20461) := b"1111111111111111_1111111111111111_1111010000010101_0000001000000110"; -- -0.046554444737038646
	pesos_i(20462) := b"1111111111111111_1111111111111111_1110110000001100_1100110101000010"; -- -0.07792966010945797
	pesos_i(20463) := b"1111111111111111_1111111111111111_1101110010011100_1000010010011111"; -- -0.1382367240028045
	pesos_i(20464) := b"0000000000000000_0000000000000000_0001100011101111_1011000110100000"; -- 0.09740743796259102
	pesos_i(20465) := b"0000000000000000_0000000000000000_0010011000100010_1110111101001111"; -- 0.14897056274855647
	pesos_i(20466) := b"0000000000000000_0000000000000000_0001111110011001_1101010011100111"; -- 0.12344103469977705
	pesos_i(20467) := b"1111111111111111_1111111111111111_1111000010000010_0010110110010011"; -- -0.06051364105317999
	pesos_i(20468) := b"1111111111111111_1111111111111111_1101111110111101_0001100010011101"; -- -0.12602087185382335
	pesos_i(20469) := b"0000000000000000_0000000000000000_0001001000011111_0111010010110111"; -- 0.07079247923030978
	pesos_i(20470) := b"1111111111111111_1111111111111111_1101110110110010_1011001000110110"; -- -0.13399206329120666
	pesos_i(20471) := b"0000000000000000_0000000000000000_0000011110011000_1100010000110010"; -- 0.029674780105624885
	pesos_i(20472) := b"1111111111111111_1111111111111111_1110111000101001_1011110000001000"; -- -0.06967568209281162
	pesos_i(20473) := b"0000000000000000_0000000000000000_0001100100000001_1110101000101001"; -- 0.0976854658351871
	pesos_i(20474) := b"0000000000000000_0000000000000000_0001101000001111_1101111010101111"; -- 0.10180465470036668
	pesos_i(20475) := b"1111111111111111_1111111111111111_1111110111110111_0000101010010010"; -- -0.007949199155203477
	pesos_i(20476) := b"1111111111111111_1111111111111111_1111111001001100_0110000011000011"; -- -0.006647064488535288
	pesos_i(20477) := b"1111111111111111_1111111111111111_1111100001010011_0011111010101001"; -- -0.029979785707951536
	pesos_i(20478) := b"0000000000000000_0000000000000000_0001110000010110_0111011101001000"; -- 0.10971780306351427
	pesos_i(20479) := b"0000000000000000_0000000000000000_0000010100001011_1010011010001101"; -- 0.019709023869295513
	pesos_i(20480) := b"0000000000000000_0000000000000000_0001011101011101_1101100101111110"; -- 0.09127578093114072
	pesos_i(20481) := b"0000000000000000_0000000000000000_0001111001101100_0111110111110000"; -- 0.11884295569697122
	pesos_i(20482) := b"0000000000000000_0000000000000000_0000010101011000_0111001101000110"; -- 0.02088089434146579
	pesos_i(20483) := b"1111111111111111_1111111111111111_1101101001111010_0010010110100010"; -- -0.1465736846313333
	pesos_i(20484) := b"1111111111111111_1111111111111111_1111000110111000_0100110100000100"; -- -0.05578154231104147
	pesos_i(20485) := b"0000000000000000_0000000000000000_0000110001110000_1011010101100100"; -- 0.04859479605154777
	pesos_i(20486) := b"1111111111111111_1111111111111111_1110011100000011_0110001110010000"; -- -0.09760453914488211
	pesos_i(20487) := b"1111111111111111_1111111111111111_1111101011001001_0010010111011011"; -- -0.020368227071689907
	pesos_i(20488) := b"1111111111111111_1111111111111111_1101101001111110_1000000101110000"; -- -0.146507177447435
	pesos_i(20489) := b"1111111111111111_1111111111111111_1110001011000110_0100100011010010"; -- -0.11416191941747213
	pesos_i(20490) := b"1111111111111111_1111111111111111_1101010110101001_0001110011010110"; -- -0.165388295917796
	pesos_i(20491) := b"0000000000000000_0000000000000000_0000110110010111_1100001010111110"; -- 0.05309693469145133
	pesos_i(20492) := b"1111111111111111_1111111111111111_1110010011000001_1110101100000011"; -- -0.1064160458304935
	pesos_i(20493) := b"0000000000000000_0000000000000000_0001101011100000_0111000111101000"; -- 0.10498725819723156
	pesos_i(20494) := b"1111111111111111_1111111111111111_1101101010001011_1111110111101110"; -- -0.14630139285900337
	pesos_i(20495) := b"0000000000000000_0000000000000000_0001010110111001_0110011111101001"; -- 0.08486031941455364
	pesos_i(20496) := b"0000000000000000_0000000000000000_0000101001001000_1010110010111000"; -- 0.040171427569730335
	pesos_i(20497) := b"1111111111111111_1111111111111111_1111111110100110_0000011101011010"; -- -0.0013728527373664274
	pesos_i(20498) := b"0000000000000000_0000000000000000_0010001001011101_0010010101000110"; -- 0.13423378916224368
	pesos_i(20499) := b"0000000000000000_0000000000000000_0010001001011110_1001011000011100"; -- 0.13425577342930833
	pesos_i(20500) := b"0000000000000000_0000000000000000_0000011011000111_1110111010111011"; -- 0.0264882284564692
	pesos_i(20501) := b"1111111111111111_1111111111111111_1101101000010010_1010111010001001"; -- -0.14815243865473104
	pesos_i(20502) := b"0000000000000000_0000000000000000_0001010001100011_1111011011010100"; -- 0.07965033224282504
	pesos_i(20503) := b"0000000000000000_0000000000000000_0000011010010001_1111110000101111"; -- 0.025665055736334083
	pesos_i(20504) := b"0000000000000000_0000000000000000_0000111001001001_1001101110110011"; -- 0.05581067201244515
	pesos_i(20505) := b"0000000000000000_0000000000000000_0000010100101110_1011111100101100"; -- 0.02024454894876563
	pesos_i(20506) := b"0000000000000000_0000000000000000_0001011101001100_1000001000110010"; -- 0.09101117819859156
	pesos_i(20507) := b"0000000000000000_0000000000000000_0000101110101010_1000111111010010"; -- 0.04557131643494988
	pesos_i(20508) := b"1111111111111111_1111111111111111_1110111001100000_1001000001100010"; -- -0.06883905036685378
	pesos_i(20509) := b"0000000000000000_0000000000000000_0001110111001001_1110101110111000"; -- 0.11636231644150938
	pesos_i(20510) := b"0000000000000000_0000000000000000_0010000000011001_1111101001100000"; -- 0.12539639334465624
	pesos_i(20511) := b"1111111111111111_1111111111111111_1111110010100100_1001110110101001"; -- -0.013113161225994707
	pesos_i(20512) := b"1111111111111111_1111111111111111_1110000100110011_1000101111001000"; -- -0.12030722021402256
	pesos_i(20513) := b"1111111111111111_1111111111111111_1111010010010001_0100001000000110"; -- -0.04465854019607078
	pesos_i(20514) := b"0000000000000000_0000000000000000_0001100011101011_0001000100011000"; -- 0.0973368341881254
	pesos_i(20515) := b"0000000000000000_0000000000000000_0000100110101011_0010000011100001"; -- 0.037767462741220635
	pesos_i(20516) := b"1111111111111111_1111111111111111_1101100110100001_0011011010011001"; -- -0.14988383063103855
	pesos_i(20517) := b"0000000000000000_0000000000000000_0010000011110010_0101001001101000"; -- 0.1286975387598276
	pesos_i(20518) := b"1111111111111111_1111111111111111_1110101000111100_1011101000010110"; -- -0.08501088098197472
	pesos_i(20519) := b"1111111111111111_1111111111111111_1110110101110001_0010011110100011"; -- -0.07249214441439267
	pesos_i(20520) := b"1111111111111111_1111111111111111_1110011000101011_0000101110010010"; -- -0.1009056823320826
	pesos_i(20521) := b"1111111111111111_1111111111111111_1110011100010100_1001110100111001"; -- -0.09734170309454836
	pesos_i(20522) := b"0000000000000000_0000000000000000_0000011100100110_1000100010100100"; -- 0.027931728416873417
	pesos_i(20523) := b"0000000000000000_0000000000000000_0000010001100011_1001100001110110"; -- 0.017144707540482647
	pesos_i(20524) := b"0000000000000000_0000000000000000_0000000100110101_1111101111010000"; -- 0.004729974971731299
	pesos_i(20525) := b"0000000000000000_0000000000000000_0001011111001001_1111110001111110"; -- 0.09292581622531208
	pesos_i(20526) := b"1111111111111111_1111111111111111_1110001110101110_0001100000111010"; -- -0.11062477671583941
	pesos_i(20527) := b"1111111111111111_1111111111111111_1101101110000010_0000101010100001"; -- -0.14254697397223703
	pesos_i(20528) := b"0000000000000000_0000000000000000_0001111010011111_1110001101111011"; -- 0.11962720639335238
	pesos_i(20529) := b"1111111111111111_1111111111111111_1110001110011100_0001000010101000"; -- -0.11089988608698158
	pesos_i(20530) := b"0000000000000000_0000000000000000_0000110101111000_0001100101010000"; -- 0.052613813527548646
	pesos_i(20531) := b"1111111111111111_1111111111111111_1101111100100100_1111101111111011"; -- -0.12834191435714298
	pesos_i(20532) := b"0000000000000000_0000000000000000_0010000000000110_1011110010011110"; -- 0.12510279522800752
	pesos_i(20533) := b"0000000000000000_0000000000000000_0000010100010010_1011111001011000"; -- 0.01981725357588445
	pesos_i(20534) := b"0000000000000000_0000000000000000_0001011011110100_1001101100111011"; -- 0.08966989698935018
	pesos_i(20535) := b"0000000000000000_0000000000000000_0001101101010100_1011001110100101"; -- 0.1067611959584385
	pesos_i(20536) := b"0000000000000000_0000000000000000_0010000111011000_1011111010101011"; -- 0.1322135131290996
	pesos_i(20537) := b"1111111111111111_1111111111111111_1110011010111100_0101101001010001"; -- -0.0986884643664621
	pesos_i(20538) := b"1111111111111111_1111111111111111_1110100110000100_0001000001110111"; -- -0.0878286085383027
	pesos_i(20539) := b"0000000000000000_0000000000000000_0010000100100110_1010111111101111"; -- 0.12949657038213153
	pesos_i(20540) := b"1111111111111111_1111111111111111_1110101100101010_1101110001000101"; -- -0.0813772518521917
	pesos_i(20541) := b"0000000000000000_0000000000000000_0010011100011101_0010101110001000"; -- 0.1527888496258551
	pesos_i(20542) := b"0000000000000000_0000000000000000_0001001001100001_0011011110111101"; -- 0.07179592471482223
	pesos_i(20543) := b"0000000000000000_0000000000000000_0001001110000110_1010000001000000"; -- 0.0762729794141598
	pesos_i(20544) := b"0000000000000000_0000000000000000_0000111010110000_1011100011100110"; -- 0.05738406775197704
	pesos_i(20545) := b"1111111111111111_1111111111111111_1110100110101100_1000100111100111"; -- -0.08721101869220732
	pesos_i(20546) := b"0000000000000000_0000000000000000_0001001101100100_0010001100110100"; -- 0.07574672723423738
	pesos_i(20547) := b"1111111111111111_1111111111111111_1111111110000111_0000000000111101"; -- -0.0018462991715746892
	pesos_i(20548) := b"1111111111111111_1111111111111111_1111001101001101_0010100110111110"; -- -0.04960383523756658
	pesos_i(20549) := b"1111111111111111_1111111111111111_1101101001110011_0111001101111000"; -- -0.14667585686461043
	pesos_i(20550) := b"0000000000000000_0000000000000000_0000111000100110_1111100010101111"; -- 0.05528215660758881
	pesos_i(20551) := b"1111111111111111_1111111111111111_1110101100001011_0001001111101010"; -- -0.0818622162345934
	pesos_i(20552) := b"0000000000000000_0000000000000000_0001010101100111_0110001110000101"; -- 0.08360883712116902
	pesos_i(20553) := b"1111111111111111_1111111111111111_1111000101101100_1100001110000100"; -- -0.05693414716057961
	pesos_i(20554) := b"1111111111111111_1111111111111111_1101111111000101_0001010000011000"; -- -0.12589907082079932
	pesos_i(20555) := b"1111111111111111_1111111111111111_1101110101000101_0010111100110101"; -- -0.1356630797404207
	pesos_i(20556) := b"0000000000000000_0000000000000000_0001000100111110_1010001110001111"; -- 0.06736204376924382
	pesos_i(20557) := b"1111111111111111_1111111111111111_1111001111111110_1100111010100010"; -- -0.046893201380625534
	pesos_i(20558) := b"1111111111111111_1111111111111111_1110010100110100_1111000110011110"; -- -0.10466089146973417
	pesos_i(20559) := b"0000000000000000_0000000000000000_0001100110000101_1000000111000000"; -- 0.09969340273853808
	pesos_i(20560) := b"0000000000000000_0000000000000000_0001111000111011_0000101100001100"; -- 0.11808842707495944
	pesos_i(20561) := b"1111111111111111_1111111111111111_1110110101101101_0010111101000110"; -- -0.07255272433015407
	pesos_i(20562) := b"0000000000000000_0000000000000000_0001011100010001_1100110101101000"; -- 0.09011539261852562
	pesos_i(20563) := b"1111111111111111_1111111111111111_1101111000000101_1001101111110010"; -- -0.13272691090095995
	pesos_i(20564) := b"0000000000000000_0000000000000000_0001101111000010_0111111100100110"; -- 0.10843653376431528
	pesos_i(20565) := b"1111111111111111_1111111111111111_1110110000000101_1111000001010101"; -- -0.07803438119796385
	pesos_i(20566) := b"1111111111111111_1111111111111111_1101110000101010_0010110001000101"; -- -0.1399814923051762
	pesos_i(20567) := b"0000000000000000_0000000000000000_0001000110010001_1111110101001111"; -- 0.06863387270879028
	pesos_i(20568) := b"1111111111111111_1111111111111111_1111001100110011_1010010100000100"; -- -0.0499932160567156
	pesos_i(20569) := b"0000000000000000_0000000000000000_0000110001101010_0100111101100111"; -- 0.04849716442750325
	pesos_i(20570) := b"0000000000000000_0000000000000000_0010001101001100_1100000001001010"; -- 0.13788987932018176
	pesos_i(20571) := b"0000000000000000_0000000000000000_0010000011000111_1011010011100011"; -- 0.12804728071240754
	pesos_i(20572) := b"0000000000000000_0000000000000000_0001000010001001_1111001010010111"; -- 0.06460491357831906
	pesos_i(20573) := b"0000000000000000_0000000000000000_0001111000000011_1110110100011101"; -- 0.11724740950304756
	pesos_i(20574) := b"0000000000000000_0000000000000000_0001100111011110_1011011010001001"; -- 0.10105458113002079
	pesos_i(20575) := b"1111111111111111_1111111111111111_1111011011110101_0001000110001100"; -- -0.0353230507098927
	pesos_i(20576) := b"1111111111111111_1111111111111111_1111010100010111_1001011101010011"; -- -0.042608778253623934
	pesos_i(20577) := b"0000000000000000_0000000000000000_0001110111111101_0101001001111000"; -- 0.11714663910166892
	pesos_i(20578) := b"1111111111111111_1111111111111111_1110001011101111_1100000110000000"; -- -0.1135291159842102
	pesos_i(20579) := b"1111111111111111_1111111111111111_1111110101011100_0011010101100001"; -- -0.010311759769196285
	pesos_i(20580) := b"0000000000000000_0000000000000000_0001101101001011_1110001110101001"; -- 0.10662672887772114
	pesos_i(20581) := b"1111111111111111_1111111111111111_1110000010011101_0111011101001010"; -- -0.12259725994093627
	pesos_i(20582) := b"0000000000000000_0000000000000000_0000100111000001_1010001001010000"; -- 0.03811087081478805
	pesos_i(20583) := b"1111111111111111_1111111111111111_1101110101100000_0010101000111001"; -- -0.13525138965491268
	pesos_i(20584) := b"0000000000000000_0000000000000000_0001011010110101_1100001001001011"; -- 0.08871092161249726
	pesos_i(20585) := b"0000000000000000_0000000000000000_0000000101000000_1011001010010111"; -- 0.004893457399403408
	pesos_i(20586) := b"0000000000000000_0000000000000000_0010000110101000_1001011111010001"; -- 0.13147877554950935
	pesos_i(20587) := b"1111111111111111_1111111111111111_1110100100100000_0110000000001001"; -- -0.08934974456181687
	pesos_i(20588) := b"1111111111111111_1111111111111111_1110111011001110_1110000010110001"; -- -0.06715579685917397
	pesos_i(20589) := b"1111111111111111_1111111111111111_1111100111111001_1111000011010100"; -- -0.023529956974740186
	pesos_i(20590) := b"0000000000000000_0000000000000000_0001100111101010_0110101110001000"; -- 0.10123321605054812
	pesos_i(20591) := b"1111111111111111_1111111111111111_1110110100100101_0001110100110010"; -- -0.07365243455492904
	pesos_i(20592) := b"0000000000000000_0000000000000000_0000101111011111_0101010111010111"; -- 0.04637657644427833
	pesos_i(20593) := b"1111111111111111_1111111111111111_1110101110000000_1100110010001101"; -- -0.08006593272023155
	pesos_i(20594) := b"1111111111111111_1111111111111111_1111101011111101_1001100000010011"; -- -0.019567962057447468
	pesos_i(20595) := b"1111111111111111_1111111111111111_1110111000111011_1001001110111011"; -- -0.06940342592295562
	pesos_i(20596) := b"1111111111111111_1111111111111111_1101111101100111_0100100100011010"; -- -0.12733023741816743
	pesos_i(20597) := b"1111111111111111_1111111111111111_1110011001111011_0101110010010101"; -- -0.09968015064140058
	pesos_i(20598) := b"1111111111111111_1111111111111111_1111101101001000_0000110000000101"; -- -0.018431900768223097
	pesos_i(20599) := b"1111111111111111_1111111111111111_1110001000110110_1110111100111011"; -- -0.11634926607955773
	pesos_i(20600) := b"1111111111111111_1111111111111111_1110000111010111_1100100000011010"; -- -0.11780118343332388
	pesos_i(20601) := b"1111111111111111_1111111111111111_1110110101111010_0101110000100110"; -- -0.07235168520613892
	pesos_i(20602) := b"1111111111111111_1111111111111111_1110111010010101_1100010111010000"; -- -0.06802714983132359
	pesos_i(20603) := b"1111111111111111_1111111111111111_1110101100111100_1101101111100110"; -- -0.08110261559482651
	pesos_i(20604) := b"1111111111111111_1111111111111111_1110011101001111_1110011000011011"; -- -0.09643709039615166
	pesos_i(20605) := b"0000000000000000_0000000000000000_0001110111010100_1101111011110010"; -- 0.1165294017754486
	pesos_i(20606) := b"1111111111111111_1111111111111111_1111001010101011_0011111111010101"; -- -0.05207444230122775
	pesos_i(20607) := b"0000000000000000_0000000000000000_0000111101001000_0101010110000011"; -- 0.059697479654779645
	pesos_i(20608) := b"0000000000000000_0000000000000000_0001110101010111_0010000011110110"; -- 0.1146107292268982
	pesos_i(20609) := b"1111111111111111_1111111111111111_1110101001101011_0111100100101011"; -- -0.08429758742038153
	pesos_i(20610) := b"0000000000000000_0000000000000000_0001111110110101_0001001000000010"; -- 0.12385666420842377
	pesos_i(20611) := b"1111111111111111_1111111111111111_1111010111111111_1010001110000111"; -- -0.03906801176688708
	pesos_i(20612) := b"1111111111111111_1111111111111111_1110101001011001_0001010001001100"; -- -0.08457825800008638
	pesos_i(20613) := b"1111111111111111_1111111111111111_1111101110101011_1001010000101100"; -- -0.01691316530486797
	pesos_i(20614) := b"0000000000000000_0000000000000000_0010000000011010_1101110110110011"; -- 0.1254099428499129
	pesos_i(20615) := b"1111111111111111_1111111111111111_1110010001100111_0100010110100001"; -- -0.10779919460628977
	pesos_i(20616) := b"1111111111111111_1111111111111111_1111010110111010_0000111010010111"; -- -0.04012974571799069
	pesos_i(20617) := b"0000000000000000_0000000000000000_0000000011100101_1110001111010110"; -- 0.003507842730151399
	pesos_i(20618) := b"0000000000000000_0000000000000000_0001001011100011_1010000101110011"; -- 0.07378586833554439
	pesos_i(20619) := b"1111111111111111_1111111111111111_1111110100000111_1100111001101011"; -- -0.011599634995104347
	pesos_i(20620) := b"1111111111111111_1111111111111111_1110000011000000_0111101111101111"; -- -0.12206292559175742
	pesos_i(20621) := b"1111111111111111_1111111111111111_1110010011100100_0010111100101001"; -- -0.10589318522504267
	pesos_i(20622) := b"0000000000000000_0000000000000000_0000101010011001_1111001110011000"; -- 0.041411613958857174
	pesos_i(20623) := b"0000000000000000_0000000000000000_0001011111001101_0000100111100001"; -- 0.09297239060122015
	pesos_i(20624) := b"0000000000000000_0000000000000000_0001110001110101_1100010111001010"; -- 0.11117206745671904
	pesos_i(20625) := b"0000000000000000_0000000000000000_0000110001001010_0000001011001100"; -- 0.04800431703721344
	pesos_i(20626) := b"1111111111111111_1111111111111111_1110000101100101_1000110000111100"; -- -0.11954425363611335
	pesos_i(20627) := b"0000000000000000_0000000000000000_0000100111101100_1001001001010001"; -- 0.038766045372305206
	pesos_i(20628) := b"0000000000000000_0000000000000000_0001100100001011_0010101100001010"; -- 0.09782666194472883
	pesos_i(20629) := b"0000000000000000_0000000000000000_0000010011001010_0000100011101100"; -- 0.01870780719637214
	pesos_i(20630) := b"0000000000000000_0000000000000000_0000111010011011_0010010001011011"; -- 0.057054779313202464
	pesos_i(20631) := b"0000000000000000_0000000000000000_0001110010001111_1110100011110101"; -- 0.11157089207991136
	pesos_i(20632) := b"0000000000000000_0000000000000000_0001010111101111_1100111011110001"; -- 0.0856904353494112
	pesos_i(20633) := b"0000000000000000_0000000000000000_0000101001100110_1110011010011001"; -- 0.04063264107860933
	pesos_i(20634) := b"0000000000000000_0000000000000000_0001000101111011_0010010001011110"; -- 0.0682852487521049
	pesos_i(20635) := b"1111111111111111_1111111111111111_1110000000011011_1001011000000011"; -- -0.12457907133386163
	pesos_i(20636) := b"0000000000000000_0000000000000000_0001011001111000_0100110101101111"; -- 0.08777317011577217
	pesos_i(20637) := b"1111111111111111_1111111111111111_1110010101000001_0011101010001001"; -- -0.10447343967774245
	pesos_i(20638) := b"1111111111111111_1111111111111111_1111011100001001_1100110000111110"; -- -0.035006747186032146
	pesos_i(20639) := b"1111111111111111_1111111111111111_1110111110010011_1101100100011111"; -- -0.06415026646653943
	pesos_i(20640) := b"0000000000000000_0000000000000000_0000000101100010_1011101110010111"; -- 0.005412792621603348
	pesos_i(20641) := b"1111111111111111_1111111111111111_1110000100001001_0000111000001101"; -- -0.12095558331587328
	pesos_i(20642) := b"1111111111111111_1111111111111111_1110000011100100_0100111010101101"; -- -0.12151630655905574
	pesos_i(20643) := b"0000000000000000_0000000000000000_0001000010001011_0111100100000001"; -- 0.06462818404621978
	pesos_i(20644) := b"0000000000000000_0000000000000000_0001001010111010_1110011110010010"; -- 0.0731644374762357
	pesos_i(20645) := b"0000000000000000_0000000000000000_0000101010100100_0111110111100010"; -- 0.04157244459265187
	pesos_i(20646) := b"1111111111111111_1111111111111111_1110010010111000_0001111010111111"; -- -0.10656555013786548
	pesos_i(20647) := b"1111111111111111_1111111111111111_1110101100111111_1101011000001010"; -- -0.08105718860395052
	pesos_i(20648) := b"0000000000000000_0000000000000000_0001001101011100_1111111011110010"; -- 0.07563775443709135
	pesos_i(20649) := b"1111111111111111_1111111111111111_1111100101000011_0111001000010101"; -- -0.02631461129079088
	pesos_i(20650) := b"1111111111111111_1111111111111111_1110011011011110_1101010010010000"; -- -0.09816237915296572
	pesos_i(20651) := b"0000000000000000_0000000000000000_0000001101110000_0001110010000010"; -- 0.013429433598167933
	pesos_i(20652) := b"1111111111111111_1111111111111111_1111010001010111_0111100100111010"; -- -0.04554025961522085
	pesos_i(20653) := b"1111111111111111_1111111111111111_1110001110101011_1000001001110100"; -- -0.1106642215497852
	pesos_i(20654) := b"1111111111111111_1111111111111111_1110100111101000_1010010000001011"; -- -0.08629393315448952
	pesos_i(20655) := b"0000000000000000_0000000000000000_0001011011100000_0011110011111001"; -- 0.08935910301876893
	pesos_i(20656) := b"0000000000000000_0000000000000000_0000111110011100_0000111001110011"; -- 0.06097498225712958
	pesos_i(20657) := b"0000000000000000_0000000000000000_0010001011011111_0011111111010001"; -- 0.13621901368867623
	pesos_i(20658) := b"0000000000000000_0000000000000000_0001001101100100_1001111011001111"; -- 0.0757540947367616
	pesos_i(20659) := b"0000000000000000_0000000000000000_0010001101110011_1110001100011011"; -- 0.13848704729990427
	pesos_i(20660) := b"0000000000000000_0000000000000000_0010001001100001_1101100001011011"; -- 0.1343054982348152
	pesos_i(20661) := b"1111111111111111_1111111111111111_1111001100101001_1000101011101101"; -- -0.05014735896856348
	pesos_i(20662) := b"0000000000000000_0000000000000000_0001000000101110_1110100110100000"; -- 0.06321582935612775
	pesos_i(20663) := b"0000000000000000_0000000000000000_0000111110111101_1110011011100100"; -- 0.061491423264349275
	pesos_i(20664) := b"0000000000000000_0000000000000000_0001001100000010_1010101110010110"; -- 0.07425949487623432
	pesos_i(20665) := b"0000000000000000_0000000000000000_0010010010001110_0101111100111001"; -- 0.1427974237608761
	pesos_i(20666) := b"1111111111111111_1111111111111111_1110000010010101_0011011010010111"; -- -0.12272318668489829
	pesos_i(20667) := b"0000000000000000_0000000000000000_0010001011100101_1101100011100000"; -- 0.13631968954750512
	pesos_i(20668) := b"0000000000000000_0000000000000000_0000110100010101_0111010010110001"; -- 0.051108639840826905
	pesos_i(20669) := b"0000000000000000_0000000000000000_0000100011100010_0000110011110100"; -- 0.034699258464447935
	pesos_i(20670) := b"1111111111111111_1111111111111111_1110011010011011_1011111000010111"; -- -0.0991860575350411
	pesos_i(20671) := b"1111111111111111_1111111111111111_1110011100001010_0100010010111010"; -- -0.09749956571564133
	pesos_i(20672) := b"1111111111111111_1111111111111111_1110000000011011_0010001100001001"; -- -0.12458592442717709
	pesos_i(20673) := b"0000000000000000_0000000000000000_0001000100000111_1010110101000111"; -- 0.06652338970005764
	pesos_i(20674) := b"0000000000000000_0000000000000000_0000001011111001_0111010100100110"; -- 0.011618921082271545
	pesos_i(20675) := b"0000000000000000_0000000000000000_0001000000110111_0111010110111001"; -- 0.06334625027760839
	pesos_i(20676) := b"0000000000000000_0000000000000000_0000110010010100_1001000110000101"; -- 0.049141974474768445
	pesos_i(20677) := b"0000000000000000_0000000000000000_0000001101001111_1011101100111010"; -- 0.012935353841602854
	pesos_i(20678) := b"1111111111111111_1111111111111111_1111011000110100_0010110100011110"; -- -0.038266353707052364
	pesos_i(20679) := b"0000000000000000_0000000000000000_0001110011101010_1001010100001000"; -- 0.11295443964608803
	pesos_i(20680) := b"0000000000000000_0000000000000000_0001001111011010_1100111001100111"; -- 0.07755746846802908
	pesos_i(20681) := b"0000000000000000_0000000000000000_0001100101100010_0111010110110010"; -- 0.09915862654948275
	pesos_i(20682) := b"1111111111111111_1111111111111111_1101111111101101_1010001010000111"; -- -0.12528022952783485
	pesos_i(20683) := b"1111111111111111_1111111111111111_1111000111101100_1011110010101100"; -- -0.054981430098149986
	pesos_i(20684) := b"1111111111111111_1111111111111111_1110001100100100_0001011110101000"; -- -0.11273052348838193
	pesos_i(20685) := b"1111111111111111_1111111111111111_1111101101101001_0110100010111100"; -- -0.017922834476487667
	pesos_i(20686) := b"0000000000000000_0000000000000000_0001110011000111_0100111101010001"; -- 0.11241622671143374
	pesos_i(20687) := b"0000000000000000_0000000000000000_0001001100111010_1111110110110100"; -- 0.07511888172154034
	pesos_i(20688) := b"0000000000000000_0000000000000000_0001111100100110_1110011001110110"; -- 0.12168732046394193
	pesos_i(20689) := b"1111111111111111_1111111111111111_1110100000110000_1101101101011010"; -- -0.0930045036830523
	pesos_i(20690) := b"1111111111111111_1111111111111111_1111100111100101_0111110110011101"; -- -0.023842000058494895
	pesos_i(20691) := b"0000000000000000_0000000000000000_0001010010000111_0110110010000100"; -- 0.08019140458459274
	pesos_i(20692) := b"1111111111111111_1111111111111111_1110110001001001_0010110100010100"; -- -0.07700842143493421
	pesos_i(20693) := b"0000000000000000_0000000000000000_0000110111111110_1010000011011100"; -- 0.05466657034755097
	pesos_i(20694) := b"1111111111111111_1111111111111111_1110001111100001_1101000110001000"; -- -0.10983553331643589
	pesos_i(20695) := b"1111111111111111_1111111111111111_1111110100001010_1001000110101101"; -- -0.011557479129335286
	pesos_i(20696) := b"0000000000000000_0000000000000000_0000100001011110_0111110010010100"; -- 0.03269175169269532
	pesos_i(20697) := b"0000000000000000_0000000000000000_0000000101111110_0110110000100010"; -- 0.005835302572249473
	pesos_i(20698) := b"0000000000000000_0000000000000000_0000110100001100_1101101110010011"; -- 0.05097744309558768
	pesos_i(20699) := b"1111111111111111_1111111111111111_1110011111101101_1100011110010000"; -- -0.09402802220580928
	pesos_i(20700) := b"1111111111111111_1111111111111111_1110101011100001_1101001110101101"; -- -0.0824916555842392
	pesos_i(20701) := b"1111111111111111_1111111111111111_1101110111010100_1010111000001101"; -- -0.13347351257758763
	pesos_i(20702) := b"1111111111111111_1111111111111111_1110100000111101_1011100011101100"; -- -0.09280819175953776
	pesos_i(20703) := b"1111111111111111_1111111111111111_1101101100111110_1101101100010101"; -- -0.14357214681434666
	pesos_i(20704) := b"0000000000000000_0000000000000000_0000001000111111_0101000111111111"; -- 0.008778691125929067
	pesos_i(20705) := b"0000000000000000_0000000000000000_0000101011001111_0110011110010000"; -- 0.04222724212369065
	pesos_i(20706) := b"1111111111111111_1111111111111111_1101111110110000_1001101011110001"; -- -0.1262114679558064
	pesos_i(20707) := b"0000000000000000_0000000000000000_0001110110001000_1001010000000111"; -- 0.11536526836306135
	pesos_i(20708) := b"0000000000000000_0000000000000000_0000001011101110_1111110101011000"; -- 0.011459192365971534
	pesos_i(20709) := b"0000000000000000_0000000000000000_0000100001010001_1101010010110011"; -- 0.03249863979340963
	pesos_i(20710) := b"0000000000000000_0000000000000000_0000100010011101_0101001110110110"; -- 0.03365061950695047
	pesos_i(20711) := b"0000000000000000_0000000000000000_0000101110100011_1011010101100000"; -- 0.0454667433167437
	pesos_i(20712) := b"1111111111111111_1111111111111111_1110101011010101_1010110111010010"; -- -0.08267701734425748
	pesos_i(20713) := b"0000000000000000_0000000000000000_0010010110101010_1011000001000111"; -- 0.14713575106907553
	pesos_i(20714) := b"0000000000000000_0000000000000000_0001111001001000_0100111101000111"; -- 0.11829085816371729
	pesos_i(20715) := b"1111111111111111_1111111111111111_1110000010110010_1011001001010010"; -- -0.12227330677297495
	pesos_i(20716) := b"1111111111111111_1111111111111111_1101101000101000_1101001101111101"; -- -0.14781454270515376
	pesos_i(20717) := b"0000000000000000_0000000000000000_0000011011000101_0001011100101101"; -- 0.026444862810457836
	pesos_i(20718) := b"0000000000000000_0000000000000000_0001011001011000_1101010011010100"; -- 0.08729295908382975
	pesos_i(20719) := b"0000000000000000_0000000000000000_0010001110010101_0110101001010010"; -- 0.13899864675008794
	pesos_i(20720) := b"1111111111111111_1111111111111111_1111010010110011_0001100110100101"; -- -0.04414214829462405
	pesos_i(20721) := b"1111111111111111_1111111111111111_1110001010110000_1100111100011001"; -- -0.11448960918262995
	pesos_i(20722) := b"1111111111111111_1111111111111111_1111110011011001_1010010011110101"; -- -0.012304010591308496
	pesos_i(20723) := b"0000000000000000_0000000000000000_0000011001001111_0011010010110100"; -- 0.02464608571646913
	pesos_i(20724) := b"1111111111111111_1111111111111111_1110111111111001_1101011101110101"; -- -0.06259396929771072
	pesos_i(20725) := b"0000000000000000_0000000000000000_0000010001000001_1010011010100010"; -- 0.016626753383219825
	pesos_i(20726) := b"0000000000000000_0000000000000000_0010000101110100_1100100111001110"; -- 0.13068829809557128
	pesos_i(20727) := b"1111111111111111_1111111111111111_1111111001000111_0101101010110111"; -- -0.006723718968929261
	pesos_i(20728) := b"0000000000000000_0000000000000000_0001111111010100_1101101010000110"; -- 0.12434163825330308
	pesos_i(20729) := b"1111111111111111_1111111111111111_1110101001101010_1011111011100111"; -- -0.08430868972451129
	pesos_i(20730) := b"1111111111111111_1111111111111111_1111010001011001_1111100110011011"; -- -0.045502090152248154
	pesos_i(20731) := b"0000000000000000_0000000000000000_0000000011110000_0000101110111001"; -- 0.0036628081248885613
	pesos_i(20732) := b"0000000000000000_0000000000000000_0000100010010000_1101100001000000"; -- 0.03346015509587752
	pesos_i(20733) := b"1111111111111111_1111111111111111_1111101110010100_0111111110011011"; -- -0.01726534332969988
	pesos_i(20734) := b"1111111111111111_1111111111111111_1110110011011101_1110100010101100"; -- -0.07473893936947891
	pesos_i(20735) := b"0000000000000000_0000000000000000_0010011001010010_1000110110101100"; -- 0.1496971650570182
	pesos_i(20736) := b"0000000000000000_0000000000000000_0000101110001110_1010101111001001"; -- 0.045145737167352464
	pesos_i(20737) := b"1111111111111111_1111111111111111_1101111100010000_1010111111110001"; -- -0.1286516225087603
	pesos_i(20738) := b"1111111111111111_1111111111111111_1110110111100000_0000100000010101"; -- -0.07080029952631739
	pesos_i(20739) := b"0000000000000000_0000000000000000_0000010011110010_1010111111000110"; -- 0.01932810396266322
	pesos_i(20740) := b"1111111111111111_1111111111111111_1110101001010110_1111110001001001"; -- -0.08461020672328404
	pesos_i(20741) := b"1111111111111111_1111111111111111_1101010101101101_1000011011010110"; -- -0.1662975052356636
	pesos_i(20742) := b"1111111111111111_1111111111111111_1110001111011000_1010001000010010"; -- -0.10997569151239914
	pesos_i(20743) := b"0000000000000000_0000000000000000_0000111001001110_1011100100010100"; -- 0.05588871700584282
	pesos_i(20744) := b"1111111111111111_1111111111111111_1101110111001110_0010000000110000"; -- -0.13357352090093486
	pesos_i(20745) := b"1111111111111111_1111111111111111_1111100101111000_0011011000111010"; -- -0.025509463078278706
	pesos_i(20746) := b"0000000000000000_0000000000000000_0000000010111011_0000011000001111"; -- 0.0028537547166724592
	pesos_i(20747) := b"1111111111111111_1111111111111111_1111100101010011_0100011011011100"; -- -0.026073047014782597
	pesos_i(20748) := b"1111111111111111_1111111111111111_1110100101111111_1010001111011100"; -- -0.0878961170828543
	pesos_i(20749) := b"1111111111111111_1111111111111111_1111010111111100_1100011010111111"; -- -0.03911168885167815
	pesos_i(20750) := b"1111111111111111_1111111111111111_1110111000001001_1110111000010100"; -- -0.07016098026322079
	pesos_i(20751) := b"1111111111111111_1111111111111111_1110000011100001_1001011110000111"; -- -0.12155774075424548
	pesos_i(20752) := b"1111111111111111_1111111111111111_1110111100011001_1001001011010010"; -- -0.06601602900668943
	pesos_i(20753) := b"0000000000000000_0000000000000000_0000111111110000_0100000101101011"; -- 0.062259758492041954
	pesos_i(20754) := b"0000000000000000_0000000000000000_0001101101010010_1001001000111100"; -- 0.10672868697693204
	pesos_i(20755) := b"0000000000000000_0000000000000000_0000100111011111_0110011011100111"; -- 0.038565093453999104
	pesos_i(20756) := b"0000000000000000_0000000000000000_0000110101010001_0000011100011110"; -- 0.052017636092376265
	pesos_i(20757) := b"1111111111111111_1111111111111111_1111110010000001_0010001101010001"; -- -0.013654511272998819
	pesos_i(20758) := b"1111111111111111_1111111111111111_1111000001010011_1111111110010100"; -- -0.061218286959778545
	pesos_i(20759) := b"0000000000000000_0000000000000000_0010010100000010_0100000010011011"; -- 0.14456561826984768
	pesos_i(20760) := b"1111111111111111_1111111111111111_1111101011000111_1100111101110010"; -- -0.020388636183008034
	pesos_i(20761) := b"1111111111111111_1111111111111111_1110111011001110_0101000110000110"; -- -0.06716433033122031
	pesos_i(20762) := b"0000000000000000_0000000000000000_0001101111100100_0000101011000010"; -- 0.10894839520097777
	pesos_i(20763) := b"0000000000000000_0000000000000000_0000001010110011_0110001011001000"; -- 0.01054971113356443
	pesos_i(20764) := b"1111111111111111_1111111111111111_1111101110000000_1010010011100011"; -- -0.01756829701357364
	pesos_i(20765) := b"1111111111111111_1111111111111111_1110111000110111_0000011100111011"; -- -0.06947283563426417
	pesos_i(20766) := b"0000000000000000_0000000000000000_0001010100001001_1001011110101110"; -- 0.08217761989236881
	pesos_i(20767) := b"0000000000000000_0000000000000000_0010011110101100_0000011100010001"; -- 0.15496868301106465
	pesos_i(20768) := b"1111111111111111_1111111111111111_1111110111111110_1000101100011111"; -- -0.007834725389464996
	pesos_i(20769) := b"1111111111111111_1111111111111111_1101110001101101_1001010001110100"; -- -0.13895294357293367
	pesos_i(20770) := b"0000000000000000_0000000000000000_0000010101111111_0100011100100111"; -- 0.021473357249486055
	pesos_i(20771) := b"1111111111111111_1111111111111111_1111001100000010_0100000100111000"; -- -0.05074684514925602
	pesos_i(20772) := b"1111111111111111_1111111111111111_1110101100001101_0001010010110001"; -- -0.08183165247720382
	pesos_i(20773) := b"1111111111111111_1111111111111111_1111111101111011_1001111010111010"; -- -0.0020199581453360176
	pesos_i(20774) := b"1111111111111111_1111111111111111_1111110010010011_0110111101110010"; -- -0.013375315464489399
	pesos_i(20775) := b"0000000000000000_0000000000000000_0000110100100011_1000110000111110"; -- 0.05132366664039975
	pesos_i(20776) := b"1111111111111111_1111111111111111_1111110100110010_1111100100001010"; -- -0.010940966688999099
	pesos_i(20777) := b"0000000000000000_0000000000000000_0001101100010000_1001101100001011"; -- 0.1057221318531206
	pesos_i(20778) := b"1111111111111111_1111111111111111_1110011010100110_1111101101000001"; -- -0.09901456520879126
	pesos_i(20779) := b"0000000000000000_0000000000000000_0001011101110001_1000100001110110"; -- 0.09157612692404608
	pesos_i(20780) := b"1111111111111111_1111111111111111_1101100100100001_0011110001100110"; -- -0.1518366100132087
	pesos_i(20781) := b"1111111111111111_1111111111111111_1110111100010100_1101111010000010"; -- -0.06608781181811692
	pesos_i(20782) := b"1111111111111111_1111111111111111_1111111001001010_1110110001011101"; -- -0.006669261330754338
	pesos_i(20783) := b"1111111111111111_1111111111111111_1111011100101111_1111110100000100"; -- -0.03442400611010432
	pesos_i(20784) := b"1111111111111111_1111111111111111_1101100110101010_1010001110000001"; -- -0.14974001036561585
	pesos_i(20785) := b"1111111111111111_1111111111111111_1110000001010100_0101110100100101"; -- -0.1237127098877029
	pesos_i(20786) := b"0000000000000000_0000000000000000_0001101111101100_0001101101000101"; -- 0.10907144952314757
	pesos_i(20787) := b"1111111111111111_1111111111111111_1110100010100011_0011100011100111"; -- -0.09125942567067002
	pesos_i(20788) := b"1111111111111111_1111111111111111_1110100011010011_0000010111101011"; -- -0.09053004283490647
	pesos_i(20789) := b"0000000000000000_0000000000000000_0000111110101011_0001111111110010"; -- 0.06120490712328714
	pesos_i(20790) := b"1111111111111111_1111111111111111_1111011100000100_1110011101001100"; -- -0.03508142837751618
	pesos_i(20791) := b"1111111111111111_1111111111111111_1111110101011010_0101111011100001"; -- -0.010339803841369235
	pesos_i(20792) := b"0000000000000000_0000000000000000_0000010010011010_0110101000110011"; -- 0.01798118350716002
	pesos_i(20793) := b"0000000000000000_0000000000000000_0000111000100011_0110001001001100"; -- 0.0552274166076738
	pesos_i(20794) := b"0000000000000000_0000000000000000_0001001111100101_0110010101010010"; -- 0.07771905180164704
	pesos_i(20795) := b"1111111111111111_1111111111111111_1110101010010101_1011110110100001"; -- -0.083652637581047
	pesos_i(20796) := b"0000000000000000_0000000000000000_0001010010111010_1100011010001100"; -- 0.08097496908486555
	pesos_i(20797) := b"0000000000000000_0000000000000000_0001000100110100_1101111101100100"; -- 0.06721302208821679
	pesos_i(20798) := b"0000000000000000_0000000000000000_0000101100011011_1001111101110000"; -- 0.043390240605957094
	pesos_i(20799) := b"1111111111111111_1111111111111111_1110100000101011_1011010010101111"; -- -0.09308310259046164
	pesos_i(20800) := b"1111111111111111_1111111111111111_1110001110010100_1100100110101101"; -- -0.11101092835317693
	pesos_i(20801) := b"1111111111111111_1111111111111111_1111001110001001_0101011100011010"; -- -0.04868560414420237
	pesos_i(20802) := b"0000000000000000_0000000000000000_0000111110010011_0010001110111000"; -- 0.06083892104252264
	pesos_i(20803) := b"0000000000000000_0000000000000000_0001101111011001_0101001101010011"; -- 0.10878487369029212
	pesos_i(20804) := b"0000000000000000_0000000000000000_0001010111011110_1100010010010100"; -- 0.08543041804752151
	pesos_i(20805) := b"0000000000000000_0000000000000000_0010011000001101_0111100001101010"; -- 0.1486430415424264
	pesos_i(20806) := b"0000000000000000_0000000000000000_0010001111110000_0000111000101000"; -- 0.1403817031135012
	pesos_i(20807) := b"0000000000000000_0000000000000000_0001001100101011_1011010100101110"; -- 0.07488567717524965
	pesos_i(20808) := b"0000000000000000_0000000000000000_0000010001000111_1010111011010101"; -- 0.016718794757113332
	pesos_i(20809) := b"1111111111111111_1111111111111111_1110111111011111_1001110111110000"; -- -0.0629941262648144
	pesos_i(20810) := b"1111111111111111_1111111111111111_1110000110001001_0001011101011100"; -- -0.11900190346282846
	pesos_i(20811) := b"1111111111111111_1111111111111111_1111110100101001_0000001110000110"; -- -0.011092929657359822
	pesos_i(20812) := b"0000000000000000_0000000000000000_0001011000101011_1111011100100100"; -- 0.08660835858889555
	pesos_i(20813) := b"0000000000000000_0000000000000000_0001001100111101_1000001111001101"; -- 0.07515739210280842
	pesos_i(20814) := b"1111111111111111_1111111111111111_1110000111100001_0101100101110111"; -- -0.11765518999888937
	pesos_i(20815) := b"1111111111111111_1111111111111111_1110101001000101_1010001010100101"; -- -0.08487494912181048
	pesos_i(20816) := b"0000000000000000_0000000000000000_0001010001111111_0111101100011001"; -- 0.08007020346889433
	pesos_i(20817) := b"1111111111111111_1111111111111111_1111000110011000_1101011101100011"; -- -0.056261576040020154
	pesos_i(20818) := b"0000000000000000_0000000000000000_0000000101001011_0100000001001111"; -- 0.005054492214038975
	pesos_i(20819) := b"1111111111111111_1111111111111111_1111000011001010_0001111110000110"; -- -0.059415845679062794
	pesos_i(20820) := b"0000000000000000_0000000000000000_0000101110111001_0111010011110000"; -- 0.04579859602034659
	pesos_i(20821) := b"1111111111111111_1111111111111111_1111100011010101_1110001110011111"; -- -0.02798631056932149
	pesos_i(20822) := b"1111111111111111_1111111111111111_1110001110001010_0011000101011100"; -- -0.11117259515266993
	pesos_i(20823) := b"1111111111111111_1111111111111111_1110110111011100_0100101100110010"; -- -0.07085733439970385
	pesos_i(20824) := b"1111111111111111_1111111111111111_1111010101110110_1111011001001011"; -- -0.04115353273784955
	pesos_i(20825) := b"1111111111111111_1111111111111111_1111110010001110_0101000111100001"; -- -0.013453371580520164
	pesos_i(20826) := b"0000000000000000_0000000000000000_0001100111011000_0010111001101011"; -- 0.1009549152456685
	pesos_i(20827) := b"0000000000000000_0000000000000000_0001100001111010_0101101000000010"; -- 0.09561693707570837
	pesos_i(20828) := b"0000000000000000_0000000000000000_0001000011110111_0111001110100111"; -- 0.06627581439487154
	pesos_i(20829) := b"0000000000000000_0000000000000000_0000110110001001_0110001000100110"; -- 0.05287755419453287
	pesos_i(20830) := b"1111111111111111_1111111111111111_1110011100110011_1010110001000110"; -- -0.09686778342793656
	pesos_i(20831) := b"1111111111111111_1111111111111111_1101110001101101_0110110100110111"; -- -0.1389552823166804
	pesos_i(20832) := b"1111111111111111_1111111111111111_1111111010010011_0000110011111010"; -- -0.005568684495000864
	pesos_i(20833) := b"0000000000000000_0000000000000000_0000010110110010_1111100011001111"; -- 0.022262144528541587
	pesos_i(20834) := b"0000000000000000_0000000000000000_0000110111111010_1100001101101101"; -- 0.054607595475997105
	pesos_i(20835) := b"1111111111111111_1111111111111111_1111101011001100_1011011101011010"; -- -0.020313778482333577
	pesos_i(20836) := b"0000000000000000_0000000000000000_0001011110111111_0111101110100111"; -- 0.09276554905674649
	pesos_i(20837) := b"1111111111111111_1111111111111111_1101110110001010_1010000100110111"; -- -0.1346034280527304
	pesos_i(20838) := b"1111111111111111_1111111111111111_1111010100110001_1101101111110110"; -- -0.04220795854156269
	pesos_i(20839) := b"0000000000000000_0000000000000000_0001100010001001_1001111101001001"; -- 0.09584994819334293
	pesos_i(20840) := b"1111111111111111_1111111111111111_1111101001011010_1000000101110100"; -- -0.022056493004102663
	pesos_i(20841) := b"0000000000000000_0000000000000000_0000100000110001_1110001000000010"; -- 0.03201115168974735
	pesos_i(20842) := b"1111111111111111_1111111111111111_1111010011100000_1101001001011010"; -- -0.04344449325473451
	pesos_i(20843) := b"0000000000000000_0000000000000000_0010001001000010_1111000101100101"; -- 0.13383396835537453
	pesos_i(20844) := b"1111111111111111_1111111111111111_1111011011100110_1001010111001111"; -- -0.03554404931635367
	pesos_i(20845) := b"1111111111111111_1111111111111111_1111010010110001_1010010101010010"; -- -0.044164340480896964
	pesos_i(20846) := b"0000000000000000_0000000000000000_0000110110101011_0000010100000000"; -- 0.05339080100480553
	pesos_i(20847) := b"1111111111111111_1111111111111111_1101111010011101_0000011000111100"; -- -0.13041649841341643
	pesos_i(20848) := b"0000000000000000_0000000000000000_0001111010101000_0111001101011000"; -- 0.11975785162216025
	pesos_i(20849) := b"0000000000000000_0000000000000000_0000110110000000_1010011111011000"; -- 0.05274437921296624
	pesos_i(20850) := b"0000000000000000_0000000000000000_0000111111000010_0011111111101110"; -- 0.061557765647749285
	pesos_i(20851) := b"0000000000000000_0000000000000000_0001011001110111_1011110100010101"; -- 0.08776456610275414
	pesos_i(20852) := b"1111111111111111_1111111111111111_1110011011110010_1101110011101101"; -- -0.09785670490799535
	pesos_i(20853) := b"0000000000000000_0000000000000000_0001000101110000_1100111100110111"; -- 0.06812758542584549
	pesos_i(20854) := b"0000000000000000_0000000000000000_0010001101101001_1110111000010011"; -- 0.13833511309168547
	pesos_i(20855) := b"0000000000000000_0000000000000000_0000010000110001_0101110000111100"; -- 0.01637817820406522
	pesos_i(20856) := b"1111111111111111_1111111111111111_1111001000010111_0011101100001111"; -- -0.05433302760244409
	pesos_i(20857) := b"1111111111111111_1111111111111111_1101111111110101_0101110011001001"; -- -0.1251623162517721
	pesos_i(20858) := b"0000000000000000_0000000000000000_0010001101110111_0001010000111101"; -- 0.13853575219613598
	pesos_i(20859) := b"1111111111111111_1111111111111111_1111101100011110_1111100001010101"; -- -0.019058684631250267
	pesos_i(20860) := b"1111111111111111_1111111111111111_1110000011101001_0101011100010000"; -- -0.12143951282305261
	pesos_i(20861) := b"0000000000000000_0000000000000000_0010010101000011_1011110101010000"; -- 0.14556487267814916
	pesos_i(20862) := b"1111111111111111_1111111111111111_1110010011101001_0011110101010111"; -- -0.10581604601413515
	pesos_i(20863) := b"0000000000000000_0000000000000000_0001101111111011_1110110000000101"; -- 0.10931277398484454
	pesos_i(20864) := b"0000000000000000_0000000000000000_0000101101111111_0101101011000000"; -- 0.04491202521633324
	pesos_i(20865) := b"0000000000000000_0000000000000000_0001011011000111_0011000110011011"; -- 0.08897695564517978
	pesos_i(20866) := b"1111111111111111_1111111111111111_1110010011100111_0100101100100110"; -- -0.10584574049372136
	pesos_i(20867) := b"1111111111111111_1111111111111111_1110010101100100_0100011001001000"; -- -0.10393868188861098
	pesos_i(20868) := b"1111111111111111_1111111111111111_1111100000100011_1000010001011000"; -- -0.03070805415693293
	pesos_i(20869) := b"1111111111111111_1111111111111111_1110101110000010_0001101100011101"; -- -0.08004599131528627
	pesos_i(20870) := b"0000000000000000_0000000000000000_0001110001000001_1111110101001010"; -- 0.11038191845679106
	pesos_i(20871) := b"0000000000000000_0000000000000000_0000000000011111_1001101101101101"; -- 0.00048228656568238316
	pesos_i(20872) := b"0000000000000000_0000000000000000_0001010110001111_1100000110010110"; -- 0.08422479542762216
	pesos_i(20873) := b"1111111111111111_1111111111111111_1110100100100011_1011100100110000"; -- -0.08929865428250987
	pesos_i(20874) := b"0000000000000000_0000000000000000_0001100100001010_1111000000010101"; -- 0.09782314794327064
	pesos_i(20875) := b"1111111111111111_1111111111111111_1111010101010010_1110110111101110"; -- -0.041703347615572546
	pesos_i(20876) := b"1111111111111111_1111111111111111_1110010011001010_1000000100101011"; -- -0.10628502563316523
	pesos_i(20877) := b"1111111111111111_1111111111111111_1101100111000100_1000001000011111"; -- -0.14934527156273789
	pesos_i(20878) := b"1111111111111111_1111111111111111_1101100111111101_0001011001000001"; -- -0.14848194983423518
	pesos_i(20879) := b"1111111111111111_1111111111111111_1101111111101101_0010011011110010"; -- -0.12528759569792117
	pesos_i(20880) := b"1111111111111111_1111111111111111_1110110101001110_1000001101000111"; -- -0.07302073967951853
	pesos_i(20881) := b"1111111111111111_1111111111111111_1110110000101101_0000010001110101"; -- -0.07743808877169495
	pesos_i(20882) := b"0000000000000000_0000000000000000_0001111000001010_0001011000000000"; -- 0.11734139913018893
	pesos_i(20883) := b"0000000000000000_0000000000000000_0000111000000100_1010011000001101"; -- 0.05475843259550634
	pesos_i(20884) := b"0000000000000000_0000000000000000_0000001000110011_0011110000010101"; -- 0.008594279363857933
	pesos_i(20885) := b"1111111111111111_1111111111111111_1111011000110011_1010100000101001"; -- -0.03827427873515892
	pesos_i(20886) := b"0000000000000000_0000000000000000_0000110100101111_0010101111011010"; -- 0.05150102676721275
	pesos_i(20887) := b"1111111111111111_1111111111111111_1101110100110011_1000010011010111"; -- -0.1359326338142818
	pesos_i(20888) := b"1111111111111111_1111111111111111_1101101100011110_0101110001011110"; -- -0.1440679807622394
	pesos_i(20889) := b"1111111111111111_1111111111111111_1111000010110011_0101010101000000"; -- -0.05976359546957227
	pesos_i(20890) := b"0000000000000000_0000000000000000_0010001100011010_1110111010001100"; -- 0.1371296971191319
	pesos_i(20891) := b"0000000000000000_0000000000000000_0000100010000011_1101110110000011"; -- 0.03326210439074442
	pesos_i(20892) := b"1111111111111111_1111111111111111_1111101100001001_1100110101000001"; -- -0.019381686843106167
	pesos_i(20893) := b"1111111111111111_1111111111111111_1101111100101010_1110111010001000"; -- -0.1282511632975256
	pesos_i(20894) := b"0000000000000000_0000000000000000_0000011010101100_1111011011010101"; -- 0.026076724150635965
	pesos_i(20895) := b"1111111111111111_1111111111111111_1111101111010101_0101110001100011"; -- -0.01627562126659242
	pesos_i(20896) := b"0000000000000000_0000000000000000_0000001011101110_0100110010100101"; -- 0.011448660157174533
	pesos_i(20897) := b"1111111111111111_1111111111111111_1110010110001101_1000101010100010"; -- -0.10330899751604
	pesos_i(20898) := b"1111111111111111_1111111111111111_1111011010001111_0101000100100101"; -- -0.036875656492656686
	pesos_i(20899) := b"0000000000000000_0000000000000000_0000111011100111_1011000010100010"; -- 0.05822280851592841
	pesos_i(20900) := b"0000000000000000_0000000000000000_0000110001001010_1001110011000101"; -- 0.04801349452764382
	pesos_i(20901) := b"1111111111111111_1111111111111111_1101101101110001_1110110011010100"; -- -0.14279289084000618
	pesos_i(20902) := b"1111111111111111_1111111111111111_1110010011111110_0111111110111010"; -- -0.10549165458733929
	pesos_i(20903) := b"1111111111111111_1111111111111111_1110111100111100_1111101000101010"; -- -0.06547581162758553
	pesos_i(20904) := b"1111111111111111_1111111111111111_1101010010000110_1100001101000110"; -- -0.16981868311305623
	pesos_i(20905) := b"0000000000000000_0000000000000000_0010011010101000_0111001010110111"; -- 0.15100781419710743
	pesos_i(20906) := b"0000000000000000_0000000000000000_0001100110011001_0101111010101011"; -- 0.0999964873211186
	pesos_i(20907) := b"0000000000000000_0000000000000000_0001000100101011_1100010101111110"; -- 0.06707414934846957
	pesos_i(20908) := b"1111111111111111_1111111111111111_1110100000111011_0001101010110111"; -- -0.09284813916347205
	pesos_i(20909) := b"0000000000000000_0000000000000000_0000010101000110_1100110011001111"; -- 0.02061157271184445
	pesos_i(20910) := b"1111111111111111_1111111111111111_1111111100011110_1011110110010010"; -- -0.003437187143856737
	pesos_i(20911) := b"0000000000000000_0000000000000000_0000101001011000_0111011111010011"; -- 0.040412415474878956
	pesos_i(20912) := b"0000000000000000_0000000000000000_0000111100100110_1011000001011101"; -- 0.05918409614067386
	pesos_i(20913) := b"1111111111111111_1111111111111111_1110101110001111_0101001111111011"; -- -0.07984423753058853
	pesos_i(20914) := b"0000000000000000_0000000000000000_0000010111111111_0111111111010100"; -- 0.023429860288011375
	pesos_i(20915) := b"0000000000000000_0000000000000000_0001000010000000_0101100101110000"; -- 0.06445845590549944
	pesos_i(20916) := b"1111111111111111_1111111111111111_1111100100100111_1100011101111101"; -- -0.02673676679512993
	pesos_i(20917) := b"1111111111111111_1111111111111111_1111100010011100_1100010000001111"; -- -0.028857942828246743
	pesos_i(20918) := b"1111111111111111_1111111111111111_1101110101101101_0110010111110100"; -- -0.13504946501088516
	pesos_i(20919) := b"1111111111111111_1111111111111111_1111000010001010_0111101001100000"; -- -0.06038699294444339
	pesos_i(20920) := b"0000000000000000_0000000000000000_0000101101100111_1011001001000010"; -- 0.04455103037759617
	pesos_i(20921) := b"0000000000000000_0000000000000000_0000110011011011_0000100001000010"; -- 0.05021716707578952
	pesos_i(20922) := b"1111111111111111_1111111111111111_1101100111000101_0101000011001111"; -- -0.1493329519964363
	pesos_i(20923) := b"1111111111111111_1111111111111111_1111001011101110_1011010011110000"; -- -0.051045123378114066
	pesos_i(20924) := b"0000000000000000_0000000000000000_0000100111011000_0010110101000110"; -- 0.03845484691256628
	pesos_i(20925) := b"0000000000000000_0000000000000000_0010001111000010_0100110110011010"; -- 0.1396835804967908
	pesos_i(20926) := b"1111111111111111_1111111111111111_1101111001011101_1000001110110011"; -- -0.13138558278338816
	pesos_i(20927) := b"0000000000000000_0000000000000000_0000111100000000_0100111100011011"; -- 0.05859846511925762
	pesos_i(20928) := b"1111111111111111_1111111111111111_1101111010100010_1001010101000110"; -- -0.13033167867745252
	pesos_i(20929) := b"0000000000000000_0000000000000000_0000110110110010_1101110001001110"; -- 0.053510445526312664
	pesos_i(20930) := b"0000000000000000_0000000000000000_0000011011110001_1101101111011010"; -- 0.02712797243064328
	pesos_i(20931) := b"0000000000000000_0000000000000000_0001000110100110_0011100101010111"; -- 0.06894262661780946
	pesos_i(20932) := b"0000000000000000_0000000000000000_0001001000100111_1110101010001101"; -- 0.0709215731031034
	pesos_i(20933) := b"0000000000000000_0000000000000000_0001010101010000_0101111001010000"; -- 0.08325757447880917
	pesos_i(20934) := b"0000000000000000_0000000000000000_0001101000100111_0110000111101111"; -- 0.10216342996028106
	pesos_i(20935) := b"0000000000000000_0000000000000000_0000101001111101_1000111010000001"; -- 0.04097834259187632
	pesos_i(20936) := b"1111111111111111_1111111111111111_1111001010110010_1101110111001110"; -- -0.051958215049511536
	pesos_i(20937) := b"1111111111111111_1111111111111111_1110100111100000_0111101111011010"; -- -0.08641839905737156
	pesos_i(20938) := b"0000000000000000_0000000000000000_0001000000010110_1010000101011000"; -- 0.06284531027287252
	pesos_i(20939) := b"1111111111111111_1111111111111111_1110110010011101_1100011101011000"; -- -0.07571748835638052
	pesos_i(20940) := b"1111111111111111_1111111111111111_1110110000111101_1011010101010100"; -- -0.07718340583519692
	pesos_i(20941) := b"1111111111111111_1111111111111111_1111001111001110_0011111101011110"; -- -0.047634162549172805
	pesos_i(20942) := b"0000000000000000_0000000000000000_0000001100000110_0100110011011111"; -- 0.011814884573849925
	pesos_i(20943) := b"0000000000000000_0000000000000000_0010011010110110_1001010011011000"; -- 0.15122347133880287
	pesos_i(20944) := b"0000000000000000_0000000000000000_0000111010010101_1010100010011011"; -- 0.05697110925108429
	pesos_i(20945) := b"1111111111111111_1111111111111111_1111111111001111_1000011110000111"; -- -0.0007396025006434983
	pesos_i(20946) := b"0000000000000000_0000000000000000_0001111001111110_0110000001110010"; -- 0.11911585591986551
	pesos_i(20947) := b"0000000000000000_0000000000000000_0001010010010111_0111110000100011"; -- 0.08043647635504185
	pesos_i(20948) := b"1111111111111111_1111111111111111_1110110100101111_1101101101111010"; -- -0.0734885051787193
	pesos_i(20949) := b"1111111111111111_1111111111111111_1101110111100100_1100011111101101"; -- -0.13322782955879098
	pesos_i(20950) := b"0000000000000000_0000000000000000_0001011111011011_0111101101001001"; -- 0.0931927732806538
	pesos_i(20951) := b"0000000000000000_0000000000000000_0010001000110010_1110111101011000"; -- 0.13358970555792282
	pesos_i(20952) := b"1111111111111111_1111111111111111_1101111101110001_1111101100100110"; -- -0.12716703726432474
	pesos_i(20953) := b"1111111111111111_1111111111111111_1111010000100101_0111101010001001"; -- -0.046303121150034404
	pesos_i(20954) := b"1111111111111111_1111111111111111_1110110010100110_1000001101010110"; -- -0.07558421280438885
	pesos_i(20955) := b"1111111111111111_1111111111111111_1110101011010101_1010110101000000"; -- -0.0826770514862267
	pesos_i(20956) := b"0000000000000000_0000000000000000_0001100101101000_0110000110111001"; -- 0.09924898882622005
	pesos_i(20957) := b"0000000000000000_0000000000000000_0000110101111110_1010110101110101"; -- 0.05271419638147475
	pesos_i(20958) := b"0000000000000000_0000000000000000_0000000100110111_1100101111010001"; -- 0.004757631820969904
	pesos_i(20959) := b"1111111111111111_1111111111111111_1111000100000110_0000100101010000"; -- -0.05850164218421553
	pesos_i(20960) := b"0000000000000000_0000000000000000_0001001001110101_0100111000110010"; -- 0.07210243913458234
	pesos_i(20961) := b"1111111111111111_1111111111111111_1110011001111010_1010000011101001"; -- -0.09969133681865952
	pesos_i(20962) := b"1111111111111111_1111111111111111_1111001000101111_0000101111110011"; -- -0.05396962475599868
	pesos_i(20963) := b"0000000000000000_0000000000000000_0000011000010010_0110111100011111"; -- 0.023718781487087608
	pesos_i(20964) := b"1111111111111111_1111111111111111_1111110101010011_0001000001110001"; -- -0.01045129063634122
	pesos_i(20965) := b"0000000000000000_0000000000000000_0001111100101101_1101100010000101"; -- 0.1217933011119999
	pesos_i(20966) := b"0000000000000000_0000000000000000_0001110010011001_0010101100110000"; -- 0.11171216892156823
	pesos_i(20967) := b"1111111111111111_1111111111111111_1111111111111001_0111111100101101"; -- -9.923118887786044e-05
	pesos_i(20968) := b"1111111111111111_1111111111111111_1111101101110111_0011010011001001"; -- -0.017712307749738875
	pesos_i(20969) := b"0000000000000000_0000000000000000_0001011110101011_0111100000110111"; -- 0.09246016833204897
	pesos_i(20970) := b"0000000000000000_0000000000000000_0001011111101101_0011011001010101"; -- 0.09346332153559792
	pesos_i(20971) := b"0000000000000000_0000000000000000_0001100001100100_0111000100001010"; -- 0.09528261650450291
	pesos_i(20972) := b"1111111111111111_1111111111111111_1111000011011110_0101100000001111"; -- -0.05910730018453266
	pesos_i(20973) := b"0000000000000000_0000000000000000_0000010110110010_0110100010101011"; -- 0.022253553157560457
	pesos_i(20974) := b"0000000000000000_0000000000000000_0001011000101001_1111110110010000"; -- 0.0865782239570061
	pesos_i(20975) := b"1111111111111111_1111111111111111_1111101101000000_1010010000011000"; -- -0.018544906706866995
	pesos_i(20976) := b"1111111111111111_1111111111111111_1111101110001011_0001101111111111"; -- -0.017408609626873933
	pesos_i(20977) := b"0000000000000000_0000000000000000_0001010111001010_0101010100001011"; -- 0.08511859428298593
	pesos_i(20978) := b"1111111111111111_1111111111111111_1111000000110001_0111001100001101"; -- -0.06174546169985227
	pesos_i(20979) := b"0000000000000000_0000000000000000_0000111111111101_0001001011000110"; -- 0.06245534266706811
	pesos_i(20980) := b"1111111111111111_1111111111111111_1110111110110001_1011110111010000"; -- -0.06369413068911355
	pesos_i(20981) := b"1111111111111111_1111111111111111_1101110111110000_1000001000011000"; -- -0.13304888633625606
	pesos_i(20982) := b"0000000000000000_0000000000000000_0010001101011000_1101010101111110"; -- 0.13807424859635184
	pesos_i(20983) := b"1111111111111111_1111111111111111_1111011011011101_1110110001000001"; -- -0.03567622571442673
	pesos_i(20984) := b"1111111111111111_1111111111111111_1110010110101111_1001100011100010"; -- -0.10278934931673188
	pesos_i(20985) := b"0000000000000000_0000000000000000_0001000010010001_0010101000111101"; -- 0.06471504196361395
	pesos_i(20986) := b"1111111111111111_1111111111111111_1110010111000000_1111111101101000"; -- -0.10252383909833247
	pesos_i(20987) := b"1111111111111111_1111111111111111_1110110111100001_1110001001011101"; -- -0.07077203005730275
	pesos_i(20988) := b"1111111111111111_1111111111111111_1110010111101110_0000010101011011"; -- -0.10183683895522307
	pesos_i(20989) := b"0000000000000000_0000000000000000_0010001001100010_1111010000111011"; -- 0.1343224185652767
	pesos_i(20990) := b"1111111111111111_1111111111111111_1111110010110010_1110111100010101"; -- -0.012894685194071564
	pesos_i(20991) := b"0000000000000000_0000000000000000_0010000111001100_0001011110010100"; -- 0.13202044827497372
	pesos_i(20992) := b"0000000000000000_0000000000000000_0000111010011101_1100010100001001"; -- 0.05709487415143888
	pesos_i(20993) := b"0000000000000000_0000000000000000_0001011011100011_0100000101111010"; -- 0.08940514782736873
	pesos_i(20994) := b"0000000000000000_0000000000000000_0010000000101100_1111101000010000"; -- 0.12568629160034342
	pesos_i(20995) := b"1111111111111111_1111111111111111_1101110110001001_1111110011111010"; -- -0.13461321731413242
	pesos_i(20996) := b"1111111111111111_1111111111111111_1110011111100000_0000110011111110"; -- -0.09423750695715782
	pesos_i(20997) := b"0000000000000000_0000000000000000_0000110000111100_1010011101101010"; -- 0.047800506013720566
	pesos_i(20998) := b"1111111111111111_1111111111111111_1110011101111000_1010111010011111"; -- -0.09581478700871933
	pesos_i(20999) := b"0000000000000000_0000000000000000_0000011110110101_1110010110111000"; -- 0.030119283103139893
	pesos_i(21000) := b"1111111111111111_1111111111111111_1110101000000110_0101110010100000"; -- -0.08584042642750715
	pesos_i(21001) := b"0000000000000000_0000000000000000_0001110100101001_1000000011000010"; -- 0.1139145349778774
	pesos_i(21002) := b"1111111111111111_1111111111111111_1110000111011011_1000001100010010"; -- -0.11774426271216143
	pesos_i(21003) := b"0000000000000000_0000000000000000_0001100000000100_1101110111010110"; -- 0.09382425762451371
	pesos_i(21004) := b"1111111111111111_1111111111111111_1111010100010000_0100101111110101"; -- -0.04272008186871426
	pesos_i(21005) := b"0000000000000000_0000000000000000_0010010011010110_1010110001000001"; -- 0.143900648001816
	pesos_i(21006) := b"0000000000000000_0000000000000000_0000000011100110_1000011111000011"; -- 0.0035176135200684997
	pesos_i(21007) := b"0000000000000000_0000000000000000_0000100110010001_1101110001001000"; -- 0.03738190426018916
	pesos_i(21008) := b"1111111111111111_1111111111111111_1101100001111111_1111100101100101"; -- -0.1542972687796827
	pesos_i(21009) := b"1111111111111111_1111111111111111_1101111011101010_0111010011110111"; -- -0.1292349718156501
	pesos_i(21010) := b"0000000000000000_0000000000000000_0001010011100100_1011000101100101"; -- 0.08161457735406426
	pesos_i(21011) := b"1111111111111111_1111111111111111_1111100000000110_0111001101110100"; -- -0.031151565649351953
	pesos_i(21012) := b"0000000000000000_0000000000000000_0001111100110011_0110011010011100"; -- 0.12187806432349978
	pesos_i(21013) := b"0000000000000000_0000000000000000_0000100110110101_0000110101100001"; -- 0.03791888818371321
	pesos_i(21014) := b"1111111111111111_1111111111111111_1110000101100000_0000011001101011"; -- -0.11962852368491458
	pesos_i(21015) := b"1111111111111111_1111111111111111_1111010111010100_1111100100111001"; -- -0.0397190319390667
	pesos_i(21016) := b"1111111111111111_1111111111111111_1110000001010100_1101101011000111"; -- -0.12370522145895894
	pesos_i(21017) := b"1111111111111111_1111111111111111_1110001111100010_0101101001000011"; -- -0.1098273837068147
	pesos_i(21018) := b"1111111111111111_1111111111111111_1101110100010000_0111010001110001"; -- -0.13646766883780437
	pesos_i(21019) := b"0000000000000000_0000000000000000_0001111111010110_1110100011111100"; -- 0.12437301770290077
	pesos_i(21020) := b"1111111111111111_1111111111111111_1101100011111101_0111100111001011"; -- -0.15238226696698717
	pesos_i(21021) := b"1111111111111111_1111111111111111_1110000111011011_1110001000101111"; -- -0.11773859357652877
	pesos_i(21022) := b"1111111111111111_1111111111111111_1111100111100000_0100001001100101"; -- -0.02392182381394815
	pesos_i(21023) := b"0000000000000000_0000000000000000_0001101010111011_1010000010011110"; -- 0.10442546707197652
	pesos_i(21024) := b"0000000000000000_0000000000000000_0000111111111101_0001100100011101"; -- 0.06245572045410275
	pesos_i(21025) := b"1111111111111111_1111111111111111_1111001011010111_0100100100100010"; -- -0.051402501239871216
	pesos_i(21026) := b"1111111111111111_1111111111111111_1101111001100111_0000010000100111"; -- -0.13124059722667358
	pesos_i(21027) := b"1111111111111111_1111111111111111_1111101100010011_0011010010001111"; -- -0.019238200272704904
	pesos_i(21028) := b"1111111111111111_1111111111111111_1111011110000110_1011001001100111"; -- -0.03310093865137824
	pesos_i(21029) := b"1111111111111111_1111111111111111_1101101111110000_1000101101100101"; -- -0.14086083210475517
	pesos_i(21030) := b"0000000000000000_0000000000000000_0001101010110000_1110000001111001"; -- 0.10426142651038334
	pesos_i(21031) := b"0000000000000000_0000000000000000_0000111110110101_1111010000111010"; -- 0.06137014795937988
	pesos_i(21032) := b"0000000000000000_0000000000000000_0001001100110100_1011111000101111"; -- 0.07502354284921214
	pesos_i(21033) := b"0000000000000000_0000000000000000_0001111110101110_1101100001000110"; -- 0.1237616701903143
	pesos_i(21034) := b"0000000000000000_0000000000000000_0001101001110101_0101110100000101"; -- 0.10335332273852466
	pesos_i(21035) := b"0000000000000000_0000000000000000_0010110000000001_1101001100010111"; -- 0.17190284082708737
	pesos_i(21036) := b"0000000000000000_0000000000000000_0010000010111001_1100100101100100"; -- 0.1278348797257761
	pesos_i(21037) := b"0000000000000000_0000000000000000_0001111101010011_0001011111010101"; -- 0.12236164990735046
	pesos_i(21038) := b"1111111111111111_1111111111111111_1110101110000101_0111100101110101"; -- -0.07999459175076704
	pesos_i(21039) := b"1111111111111111_1111111111111111_1111111110000011_1010110010000010"; -- -0.0018970662618874132
	pesos_i(21040) := b"1111111111111111_1111111111111111_1110010011000010_1100011100100101"; -- -0.10640292497255703
	pesos_i(21041) := b"1111111111111111_1111111111111111_1111000010011001_1011111110010110"; -- -0.06015398588564482
	pesos_i(21042) := b"1111111111111111_1111111111111111_1110110011100011_0101110111001011"; -- -0.07465566443207368
	pesos_i(21043) := b"0000000000000000_0000000000000000_0000000110010110_0111110101100101"; -- 0.006202542349065545
	pesos_i(21044) := b"0000000000000000_0000000000000000_0010001100001001_0010010110100111"; -- 0.1368583233907964
	pesos_i(21045) := b"0000000000000000_0000000000000000_0000110000111011_1011001000011011"; -- 0.04778588441888123
	pesos_i(21046) := b"1111111111111111_1111111111111111_1110110101011100_0111110000000111"; -- -0.07280754887072306
	pesos_i(21047) := b"0000000000000000_0000000000000000_0000000001111010_0001001111100100"; -- 0.001862757758134418
	pesos_i(21048) := b"1111111111111111_1111111111111111_1111000100001101_1000000101100110"; -- -0.05838767300959165
	pesos_i(21049) := b"1111111111111111_1111111111111111_1111011101100100_1111111101111010"; -- -0.03361514358237793
	pesos_i(21050) := b"0000000000000000_0000000000000000_0001100011110111_0011100001111001"; -- 0.09752228685821945
	pesos_i(21051) := b"0000000000000000_0000000000000000_0001110110111101_1101110001100011"; -- 0.11617829730124588
	pesos_i(21052) := b"1111111111111111_1111111111111111_1111111010000110_0100000100011101"; -- -0.005763941262087745
	pesos_i(21053) := b"1111111111111111_1111111111111111_1110010111011011_0011100010010011"; -- -0.10212370305860746
	pesos_i(21054) := b"0000000000000000_0000000000000000_0010001111101011_1110011101110110"; -- 0.14031836154939747
	pesos_i(21055) := b"0000000000000000_0000000000000000_0000001011111100_0111111001011001"; -- 0.011665245697253183
	pesos_i(21056) := b"0000000000000000_0000000000000000_0001011101100010_0010111111110000"; -- 0.09134196865649544
	pesos_i(21057) := b"0000000000000000_0000000000000000_0001011001100011_0101000011001000"; -- 0.08745293509975217
	pesos_i(21058) := b"0000000000000000_0000000000000000_0010010111010101_1010010100001100"; -- 0.14779120971914744
	pesos_i(21059) := b"1111111111111111_1111111111111111_1110111101111001_1011110001001011"; -- -0.06454871328984708
	pesos_i(21060) := b"1111111111111111_1111111111111111_1110000010110101_0111101101110110"; -- -0.12223080032595969
	pesos_i(21061) := b"1111111111111111_1111111111111111_1110110001111101_0101011101010011"; -- -0.0762124464850382
	pesos_i(21062) := b"0000000000000000_0000000000000000_0000100001110011_0111111110001000"; -- 0.033012362216814854
	pesos_i(21063) := b"0000000000000000_0000000000000000_0001011011110100_0000001011001100"; -- 0.0896608112625231
	pesos_i(21064) := b"0000000000000000_0000000000000000_0001000001010110_1001101001001001"; -- 0.06382145188481853
	pesos_i(21065) := b"0000000000000000_0000000000000000_0001111111101011_0100001010101011"; -- 0.12468353917728489
	pesos_i(21066) := b"1111111111111111_1111111111111111_1110101101011101_1000011101001110"; -- -0.08060411771977125
	pesos_i(21067) := b"1111111111111111_1111111111111111_1101110111010101_1111101001100000"; -- -0.1334537043132836
	pesos_i(21068) := b"0000000000000000_0000000000000000_0001010000101100_1110001111111110"; -- 0.07880997621472367
	pesos_i(21069) := b"0000000000000000_0000000000000000_0000111011001000_1000000011010101"; -- 0.0577469369110528
	pesos_i(21070) := b"0000000000000000_0000000000000000_0000010001101001_0111010000011011"; -- 0.01723409320931535
	pesos_i(21071) := b"1111111111111111_1111111111111111_1111100111101111_1001000010011111"; -- -0.023688279240885457
	pesos_i(21072) := b"1111111111111111_1111111111111111_1110000001110011_0001001000010011"; -- -0.12324416185109704
	pesos_i(21073) := b"0000000000000000_0000000000000000_0000001010101110_1110110101001100"; -- 0.01048167339209266
	pesos_i(21074) := b"0000000000000000_0000000000000000_0000000010100001_1011000111010111"; -- 0.002467265197193146
	pesos_i(21075) := b"1111111111111111_1111111111111111_1110001001100000_0100001101000001"; -- -0.11571864769200801
	pesos_i(21076) := b"1111111111111111_1111111111111111_1101101000110001_0111010000000001"; -- -0.14768290504081613
	pesos_i(21077) := b"1111111111111111_1111111111111111_1111000010100011_1110001000110111"; -- -0.05999933404186057
	pesos_i(21078) := b"1111111111111111_1111111111111111_1111001000111001_0011111100000101"; -- -0.053813992820401835
	pesos_i(21079) := b"1111111111111111_1111111111111111_1111110001010100_0001100111010111"; -- -0.014341721501653892
	pesos_i(21080) := b"0000000000000000_0000000000000000_0000100100010110_0101101000001001"; -- 0.0354973097779659
	pesos_i(21081) := b"1111111111111111_1111111111111111_1110001010011000_0001000010000111"; -- -0.11486717899271809
	pesos_i(21082) := b"1111111111111111_1111111111111111_1110100011000010_1001001101111000"; -- -0.09078100505032258
	pesos_i(21083) := b"0000000000000000_0000000000000000_0010000010111100_1111110110011011"; -- 0.12788376835482038
	pesos_i(21084) := b"1111111111111111_1111111111111111_1110011110101111_1111011110110101"; -- -0.09497119735987676
	pesos_i(21085) := b"0000000000000000_0000000000000000_0001110100101110_1011110011110000"; -- 0.11399441590498695
	pesos_i(21086) := b"1111111111111111_1111111111111111_1110011100000000_0111111001010100"; -- -0.0976487203361384
	pesos_i(21087) := b"0000000000000000_0000000000000000_0001100000000000_1000000000110101"; -- 0.09375764181572216
	pesos_i(21088) := b"1111111111111111_1111111111111111_1101111101101011_0010011111001111"; -- -0.12727118684195474
	pesos_i(21089) := b"1111111111111111_1111111111111111_1101110101100001_1001001101101011"; -- -0.13522986069671003
	pesos_i(21090) := b"1111111111111111_1111111111111111_1110011110010110_0101100000010011"; -- -0.09536218191993591
	pesos_i(21091) := b"1111111111111111_1111111111111111_1101110011101111_1100111000100011"; -- -0.1369658628084176
	pesos_i(21092) := b"1111111111111111_1111111111111111_1110100010010001_0011101001011101"; -- -0.09153399677013531
	pesos_i(21093) := b"1111111111111111_1111111111111111_1111011111001010_1001011110000000"; -- -0.03206494460871554
	pesos_i(21094) := b"1111111111111111_1111111111111111_1110100101000101_0001000100101011"; -- -0.08878987018681789
	pesos_i(21095) := b"0000000000000000_0000000000000000_0000100001001110_0110100101101010"; -- 0.03244646862685945
	pesos_i(21096) := b"1111111111111111_1111111111111111_1110111010011100_0000000111011010"; -- -0.06793201853522071
	pesos_i(21097) := b"0000000000000000_0000000000000000_0001010001100011_1110101111000011"; -- 0.0796496725598331
	pesos_i(21098) := b"0000000000000000_0000000000000000_0001011000000100_0011101011110011"; -- 0.08600204872508717
	pesos_i(21099) := b"0000000000000000_0000000000000000_0000101001101011_0010000110100101"; -- 0.04069719569254768
	pesos_i(21100) := b"0000000000000000_0000000000000000_0010000100010111_1110101111000100"; -- 0.1292712548847068
	pesos_i(21101) := b"0000000000000000_0000000000000000_0000011101001100_0011100101101110"; -- 0.028506840993037307
	pesos_i(21102) := b"1111111111111111_1111111111111111_1110111001000111_0110000111000001"; -- -0.06922329931081425
	pesos_i(21103) := b"0000000000000000_0000000000000000_0000110011011110_0011100100000000"; -- 0.05026584874751232
	pesos_i(21104) := b"0000000000000000_0000000000000000_0000111000110111_0000010100111111"; -- 0.05552704609842319
	pesos_i(21105) := b"1111111111111111_1111111111111111_1110101111101101_0001100111101011"; -- -0.07841337217512731
	pesos_i(21106) := b"0000000000000000_0000000000000000_0000001110010000_1000111111000010"; -- 0.013924584307906801
	pesos_i(21107) := b"0000000000000000_0000000000000000_0001000010101101_0111010001110001"; -- 0.06514671103037042
	pesos_i(21108) := b"1111111111111111_1111111111111111_1110010010000000_0011011110010101"; -- -0.1074185620047032
	pesos_i(21109) := b"0000000000000000_0000000000000000_0000101001000001_0111101101110011"; -- 0.04006167939289448
	pesos_i(21110) := b"0000000000000000_0000000000000000_0001000101111000_0000000111100011"; -- 0.06823741715273199
	pesos_i(21111) := b"0000000000000000_0000000000000000_0000100001111010_1101100110100010"; -- 0.03312454423149683
	pesos_i(21112) := b"0000000000000000_0000000000000000_0010010001001000_0001010001011110"; -- 0.14172484679460315
	pesos_i(21113) := b"1111111111111111_1111111111111111_1110101100111001_0000100000011011"; -- -0.08116101592923837
	pesos_i(21114) := b"0000000000000000_0000000000000000_0000011001010000_1110010010011110"; -- 0.02467182986336257
	pesos_i(21115) := b"1111111111111111_1111111111111111_1111110011000010_1110010001101001"; -- -0.012651180513578358
	pesos_i(21116) := b"1111111111111111_1111111111111111_1110110010110101_0011101111001110"; -- -0.07535959444819372
	pesos_i(21117) := b"1111111111111111_1111111111111111_1111000110101001_1001000110011110"; -- -0.05600633512543011
	pesos_i(21118) := b"1111111111111111_1111111111111111_1110001001010000_0101110111011100"; -- -0.1159612024843477
	pesos_i(21119) := b"1111111111111111_1111111111111111_1111110011110100_1010110000011100"; -- -0.011891597046458827
	pesos_i(21120) := b"0000000000000000_0000000000000000_0001000110000111_1001000001111010"; -- 0.06847479805802235
	pesos_i(21121) := b"0000000000000000_0000000000000000_0001000000101100_1000111111100100"; -- 0.06317996323868096
	pesos_i(21122) := b"1111111111111111_1111111111111111_1101110010010001_0100100000011100"; -- -0.13840817748333367
	pesos_i(21123) := b"1111111111111111_1111111111111111_1111101010110111_0111111100101011"; -- -0.020637561891838376
	pesos_i(21124) := b"1111111111111111_1111111111111111_1110010010101110_0101100101101111"; -- -0.10671463997201344
	pesos_i(21125) := b"1111111111111111_1111111111111111_1111000100011110_0100100111011100"; -- -0.05813158403594332
	pesos_i(21126) := b"1111111111111111_1111111111111111_1110000011110111_1000010000111110"; -- -0.12122319688626762
	pesos_i(21127) := b"1111111111111111_1111111111111111_1110010111001100_1010001100101010"; -- -0.10234623167265736
	pesos_i(21128) := b"1111111111111111_1111111111111111_1101100011110101_1010010101010011"; -- -0.15250174263142047
	pesos_i(21129) := b"1111111111111111_1111111111111111_1110100111000001_1111101110110110"; -- -0.0868838005044035
	pesos_i(21130) := b"0000000000000000_0000000000000000_0001111101000000_0010110000000010"; -- 0.12207293550020352
	pesos_i(21131) := b"1111111111111111_1111111111111111_1110100010000011_0110101011001101"; -- -0.09174473278977041
	pesos_i(21132) := b"1111111111111111_1111111111111111_1111001010011011_1110001110111010"; -- -0.05230881422126162
	pesos_i(21133) := b"1111111111111111_1111111111111111_1110100111110011_0001101010101110"; -- -0.08613427392775348
	pesos_i(21134) := b"0000000000000000_0000000000000000_0001000000110100_0110000100100000"; -- 0.0632992461980697
	pesos_i(21135) := b"1111111111111111_1111111111111111_1101111101011101_1111111001110011"; -- -0.12747201631098562
	pesos_i(21136) := b"0000000000000000_0000000000000000_0001110100010110_0101100010110001"; -- 0.11362222979599852
	pesos_i(21137) := b"0000000000000000_0000000000000000_0000111111001111_0100111100011010"; -- 0.06175703404729808
	pesos_i(21138) := b"1111111111111111_1111111111111111_1111000101110000_1100100011101011"; -- -0.05687278996357413
	pesos_i(21139) := b"0000000000000000_0000000000000000_0001111100101011_0001010111100111"; -- 0.12175118351762454
	pesos_i(21140) := b"0000000000000000_0000000000000000_0000110001000111_1011100101010101"; -- 0.04796942078303988
	pesos_i(21141) := b"0000000000000000_0000000000000000_0001100100101010_0101000000010000"; -- 0.09830189121384292
	pesos_i(21142) := b"1111111111111111_1111111111111111_1111110111111010_1011001100101001"; -- -0.007893373927526324
	pesos_i(21143) := b"0000000000000000_0000000000000000_0001110111111110_0100101010011101"; -- 0.11716142974498377
	pesos_i(21144) := b"1111111111111111_1111111111111111_1110111001010001_0101110001011001"; -- -0.06907103378179737
	pesos_i(21145) := b"0000000000000000_0000000000000000_0000101110001110_0011110000111010"; -- 0.045139087766323506
	pesos_i(21146) := b"0000000000000000_0000000000000000_0001000111110110_0110101010011101"; -- 0.07016626681495647
	pesos_i(21147) := b"0000000000000000_0000000000000000_0001100000011100_0110111011101100"; -- 0.09418385751511203
	pesos_i(21148) := b"0000000000000000_0000000000000000_0000100001110100_0000011110111100"; -- 0.03302048047506713
	pesos_i(21149) := b"0000000000000000_0000000000000000_0010000001010101_0010101001101010"; -- 0.1262995250428909
	pesos_i(21150) := b"1111111111111111_1111111111111111_1111101101011001_0110010001001011"; -- -0.018167239914414282
	pesos_i(21151) := b"0000000000000000_0000000000000000_0001110010100111_1011000110111011"; -- 0.11193381125947552
	pesos_i(21152) := b"0000000000000000_0000000000000000_0001101111011001_1010100000110101"; -- 0.10878993305350595
	pesos_i(21153) := b"0000000000000000_0000000000000000_0001011011000100_1100101100101001"; -- 0.08894033192990738
	pesos_i(21154) := b"1111111111111111_1111111111111111_1110000011100000_1100110010011011"; -- -0.12156983579879732
	pesos_i(21155) := b"1111111111111111_1111111111111111_1111110110111000_0011110111010111"; -- -0.008907446950404161
	pesos_i(21156) := b"1111111111111111_1111111111111111_1111111100000101_0011100001110101"; -- -0.0038265908662940547
	pesos_i(21157) := b"0000000000000000_0000000000000000_0001101000101001_1110110110001001"; -- 0.10220226847246316
	pesos_i(21158) := b"0000000000000000_0000000000000000_0000111001000010_0111110110001101"; -- 0.055702063486133234
	pesos_i(21159) := b"0000000000000000_0000000000000000_0001011000101111_0011011000000010"; -- 0.08665788211073233
	pesos_i(21160) := b"0000000000000000_0000000000000000_0000000001110110_0010100101000101"; -- 0.001802996907373466
	pesos_i(21161) := b"0000000000000000_0000000000000000_0010001000101111_0000111101010110"; -- 0.13353057716580316
	pesos_i(21162) := b"0000000000000000_0000000000000000_0001010101010101_1100000110111011"; -- 0.08333979432331678
	pesos_i(21163) := b"1111111111111111_1111111111111111_1110101011100000_1001000111011001"; -- -0.08251083815863808
	pesos_i(21164) := b"0000000000000000_0000000000000000_0000110011010110_1000101000110000"; -- 0.05014861739825297
	pesos_i(21165) := b"1111111111111111_1111111111111111_1110001011100000_1010001001110101"; -- -0.1137598480782603
	pesos_i(21166) := b"1111111111111111_1111111111111111_1110001100101001_1000110000101110"; -- -0.11264728429660016
	pesos_i(21167) := b"0000000000000000_0000000000000000_0010001100101110_1010111100001001"; -- 0.1374310872858224
	pesos_i(21168) := b"1111111111111111_1111111111111111_1110101000000011_0110011011010001"; -- -0.08588559538367817
	pesos_i(21169) := b"0000000000000000_0000000000000000_0010010110100100_1001010110111100"; -- 0.14704261628542745
	pesos_i(21170) := b"1111111111111111_1111111111111111_1111100011011110_0101100100010011"; -- -0.02785723948993854
	pesos_i(21171) := b"0000000000000000_0000000000000000_0000100101010000_1110101111100100"; -- 0.03639101340456067
	pesos_i(21172) := b"0000000000000000_0000000000000000_0000110111010101_1111000001111000"; -- 0.05404570519059269
	pesos_i(21173) := b"1111111111111111_1111111111111111_1111011101111010_1010000010000100"; -- -0.03328511018577774
	pesos_i(21174) := b"0000000000000000_0000000000000000_0001001011000110_1001111011000110"; -- 0.07334320393520805
	pesos_i(21175) := b"0000000000000000_0000000000000000_0000010011011110_0101011101011001"; -- 0.019017657561742424
	pesos_i(21176) := b"1111111111111111_1111111111111111_1110100100111001_1110011001110010"; -- -0.0889602633322126
	pesos_i(21177) := b"1111111111111111_1111111111111111_1110111110000110_0001100100111101"; -- -0.06436006783732
	pesos_i(21178) := b"0000000000000000_0000000000000000_0001101111001001_1111101000001111"; -- 0.10855067120855683
	pesos_i(21179) := b"0000000000000000_0000000000000000_0000101011001010_1111001010010100"; -- 0.0421592341722262
	pesos_i(21180) := b"1111111111111111_1111111111111111_1110001011010010_0100011011100001"; -- -0.11397892951890413
	pesos_i(21181) := b"1111111111111111_1111111111111111_1111010111000011_1011111100100111"; -- -0.03998189246838852
	pesos_i(21182) := b"0000000000000000_0000000000000000_0000000000101100_0110010011110011"; -- 0.0006774038274855485
	pesos_i(21183) := b"1111111111111111_1111111111111111_1101101111111111_1101001101001010"; -- -0.14062766499204904
	pesos_i(21184) := b"0000000000000000_0000000000000000_0000101110100111_1111100100011000"; -- 0.045531814900301164
	pesos_i(21185) := b"0000000000000000_0000000000000000_0000011001110011_0000011101000011"; -- 0.025192693640905376
	pesos_i(21186) := b"0000000000000000_0000000000000000_0000010110010111_0001000010110001"; -- 0.021836321934772574
	pesos_i(21187) := b"0000000000000000_0000000000000000_0000011111010000_0010011001011000"; -- 0.030519863663857744
	pesos_i(21188) := b"0000000000000000_0000000000000000_0000011001010100_1100000001111001"; -- 0.02473071054729154
	pesos_i(21189) := b"1111111111111111_1111111111111111_1110011111110010_0001101111001001"; -- -0.09396196686679015
	pesos_i(21190) := b"0000000000000000_0000000000000000_0001001110100010_1001000001100010"; -- 0.07669927981961588
	pesos_i(21191) := b"0000000000000000_0000000000000000_0000111110100110_0101011101101010"; -- 0.061131919187219164
	pesos_i(21192) := b"1111111111111111_1111111111111111_1110011011000110_1110110001100000"; -- -0.09852717062095423
	pesos_i(21193) := b"1111111111111111_1111111111111111_1110001000101110_1100000100110110"; -- -0.11647407946363636
	pesos_i(21194) := b"0000000000000000_0000000000000000_0000000100001110_0000101110010001"; -- 0.004120562494299843
	pesos_i(21195) := b"0000000000000000_0000000000000000_0001010011100110_0010100001011101"; -- 0.08163692723494884
	pesos_i(21196) := b"1111111111111111_1111111111111111_1111111110011010_1001011111101001"; -- -0.001547341895552272
	pesos_i(21197) := b"1111111111111111_1111111111111111_1110101001000010_0011001001001100"; -- -0.08492742203266745
	pesos_i(21198) := b"1111111111111111_1111111111111111_1101101010110001_1000100011101111"; -- -0.1457285325523822
	pesos_i(21199) := b"0000000000000000_0000000000000000_0000110100111101_0110011010111100"; -- 0.05171815952616141
	pesos_i(21200) := b"1111111111111111_1111111111111111_1110010010100111_0110110000111110"; -- -0.10682033055370026
	pesos_i(21201) := b"0000000000000000_0000000000000000_0001001101010011_1110000101101100"; -- 0.07549866568412535
	pesos_i(21202) := b"0000000000000000_0000000000000000_0001010001110101_1011110001011110"; -- 0.07992150593575126
	pesos_i(21203) := b"0000000000000000_0000000000000000_0000000101101111_0000011101101111"; -- 0.005600418597760028
	pesos_i(21204) := b"0000000000000000_0000000000000000_0001011001111000_0100000101111111"; -- 0.08777245845849248
	pesos_i(21205) := b"0000000000000000_0000000000000000_0000011000011000_0111110010110101"; -- 0.023811143982506014
	pesos_i(21206) := b"0000000000000000_0000000000000000_0001101000111110_1001000100101100"; -- 0.10251719784534664
	pesos_i(21207) := b"1111111111111111_1111111111111111_1111000000000100_0000000111000011"; -- -0.062438859864009266
	pesos_i(21208) := b"1111111111111111_1111111111111111_1110011111101001_1111101111010110"; -- -0.09408594152296386
	pesos_i(21209) := b"0000000000000000_0000000000000000_0001101000100001_0111001101111110"; -- 0.10207292389279225
	pesos_i(21210) := b"1111111111111111_1111111111111111_1110000101100110_1000001101010101"; -- -0.11952952541319263
	pesos_i(21211) := b"0000000000000000_0000000000000000_0000001010000011_1011100110111011"; -- 0.009822471855876065
	pesos_i(21212) := b"1111111111111111_1111111111111111_1111101011110010_1011001001001011"; -- -0.01973424601335251
	pesos_i(21213) := b"0000000000000000_0000000000000000_0001111010010001_0110100001101010"; -- 0.11940624805033544
	pesos_i(21214) := b"0000000000000000_0000000000000000_0001100100100011_1111010010010001"; -- 0.098204884823711
	pesos_i(21215) := b"0000000000000000_0000000000000000_0000110000000100_1001010010011001"; -- 0.04694489229471705
	pesos_i(21216) := b"0000000000000000_0000000000000000_0001011011011100_0110101001100111"; -- 0.08930077560419268
	pesos_i(21217) := b"0000000000000000_0000000000000000_0000001001110011_0010001100001011"; -- 0.009569349458722613
	pesos_i(21218) := b"1111111111111111_1111111111111111_1111011011000110_0100101100011111"; -- -0.03603678209146574
	pesos_i(21219) := b"1111111111111111_1111111111111111_1111011100000101_1010000110010101"; -- -0.035070325055118964
	pesos_i(21220) := b"1111111111111111_1111111111111111_1101100111111000_1001001101110110"; -- -0.14855078096490504
	pesos_i(21221) := b"0000000000000000_0000000000000000_0000110110000001_0000110011001000"; -- 0.052750395671466326
	pesos_i(21222) := b"1111111111111111_1111111111111111_1111100101011010_1010000001101111"; -- -0.025960896392082728
	pesos_i(21223) := b"1111111111111111_1111111111111111_1111011110001101_1010101011100001"; -- -0.03299457550047555
	pesos_i(21224) := b"0000000000000000_0000000000000000_0001000000010100_0011000010111010"; -- 0.06280807999710356
	pesos_i(21225) := b"1111111111111111_1111111111111111_1110100100010001_0110111101011110"; -- -0.08957771257306557
	pesos_i(21226) := b"0000000000000000_0000000000000000_0000010000000010_1111001110110011"; -- 0.01567004321451426
	pesos_i(21227) := b"1111111111111111_1111111111111111_1111110001110100_1111110101011010"; -- -0.013839879608725217
	pesos_i(21228) := b"1111111111111111_1111111111111111_1111101011010010_0110001001101101"; -- -0.020227287593516344
	pesos_i(21229) := b"0000000000000000_0000000000000000_0000010111111110_0111000111011100"; -- 0.023413769013477866
	pesos_i(21230) := b"1111111111111111_1111111111111111_1111001001111101_0100001010001000"; -- -0.05277618584683177
	pesos_i(21231) := b"0000000000000000_0000000000000000_0001000011000110_0000101011001010"; -- 0.06552188330242403
	pesos_i(21232) := b"0000000000000000_0000000000000000_0001001010100000_1001001011010111"; -- 0.07276265859525434
	pesos_i(21233) := b"0000000000000000_0000000000000000_0000001100110100_0100011001100011"; -- 0.012516402517928543
	pesos_i(21234) := b"0000000000000000_0000000000000000_0000111010101000_1100111101000100"; -- 0.05726333065218138
	pesos_i(21235) := b"0000000000000000_0000000000000000_0010010101010101_1100111100001001"; -- 0.14584058732823274
	pesos_i(21236) := b"1111111111111111_1111111111111111_1110110101100111_0111000001001000"; -- -0.07264040222554599
	pesos_i(21237) := b"0000000000000000_0000000000000000_0000101101101001_0100011110101001"; -- 0.04457519410411797
	pesos_i(21238) := b"1111111111111111_1111111111111111_1101110110011000_1100000110011101"; -- -0.13438787381585565
	pesos_i(21239) := b"0000000000000000_0000000000000000_0010010011100001_0110001110000110"; -- 0.14406415951005366
	pesos_i(21240) := b"0000000000000000_0000000000000000_0000000001110111_0111001100110100"; -- 0.0018226625733866126
	pesos_i(21241) := b"0000000000000000_0000000000000000_0001001100001110_1101001101001111"; -- 0.07444496792476012
	pesos_i(21242) := b"1111111111111111_1111111111111111_1110000101110111_1001000000010011"; -- -0.11926936656985904
	pesos_i(21243) := b"1111111111111111_1111111111111111_1110011110110110_0110101101100000"; -- -0.09487275028759472
	pesos_i(21244) := b"1111111111111111_1111111111111111_1111101110110001_0101111000000010"; -- -0.016824840928930454
	pesos_i(21245) := b"0000000000000000_0000000000000000_0001100011111111_0000110111111100"; -- 0.09764182463375089
	pesos_i(21246) := b"0000000000000000_0000000000000000_0000000100110111_1011100011010111"; -- 0.0047565005960567616
	pesos_i(21247) := b"1111111111111111_1111111111111111_1110110101101010_0111100000000001"; -- -0.07259416554282053
	pesos_i(21248) := b"0000000000000000_0000000000000000_0000110111100111_1100001001011100"; -- 0.05431761504677906
	pesos_i(21249) := b"0000000000000000_0000000000000000_0000110001000110_1000011111000100"; -- 0.04795120740815189
	pesos_i(21250) := b"0000000000000000_0000000000000000_0001010011111100_0010001010110010"; -- 0.08197228274603909
	pesos_i(21251) := b"1111111111111111_1111111111111111_1110100111001010_0111000100100101"; -- -0.08675473062448423
	pesos_i(21252) := b"1111111111111111_1111111111111111_1110101100100101_0010010010001100"; -- -0.08146449646226815
	pesos_i(21253) := b"0000000000000000_0000000000000000_0001110101100001_0010001111100101"; -- 0.11476349194683824
	pesos_i(21254) := b"0000000000000000_0000000000000000_0001101010100101_0100011000101010"; -- 0.10408438229108578
	pesos_i(21255) := b"0000000000000000_0000000000000000_0010001101010010_1000110000111111"; -- 0.1379783300574549
	pesos_i(21256) := b"1111111111111111_1111111111111111_1111100001100011_0110101001000101"; -- -0.029733045609654913
	pesos_i(21257) := b"0000000000000000_0000000000000000_0000101110100100_0110000011101010"; -- 0.04547696782750959
	pesos_i(21258) := b"0000000000000000_0000000000000000_0010001011110000_1100100011000011"; -- 0.13648657576625117
	pesos_i(21259) := b"0000000000000000_0000000000000000_0000000010010111_0010011100010001"; -- 0.0023064057105323804
	pesos_i(21260) := b"1111111111111111_1111111111111111_1110110100101011_0010010000011100"; -- -0.07356046983819843
	pesos_i(21261) := b"0000000000000000_0000000000000000_0000010111010110_0001001011011000"; -- 0.02279775409411757
	pesos_i(21262) := b"1111111111111111_1111111111111111_1111110011110011_1000100001110100"; -- -0.011908980915608559
	pesos_i(21263) := b"1111111111111111_1111111111111111_1111000001000001_0101010001101100"; -- -0.06150314669769738
	pesos_i(21264) := b"1111111111111111_1111111111111111_1101110110100010_1100001011001011"; -- -0.13423521562978646
	pesos_i(21265) := b"0000000000000000_0000000000000000_0001101011010101_0000011010010111"; -- 0.10481301478192141
	pesos_i(21266) := b"0000000000000000_0000000000000000_0000010001101001_1010110111011001"; -- 0.017237535026553393
	pesos_i(21267) := b"1111111111111111_1111111111111111_1110010101010000_0000010110000000"; -- -0.1042477189649167
	pesos_i(21268) := b"0000000000000000_0000000000000000_0000000001010100_1011001000001111"; -- 0.0012923514246040034
	pesos_i(21269) := b"1111111111111111_1111111111111111_1110011111111010_0101011010000101"; -- -0.09383639578753691
	pesos_i(21270) := b"1111111111111111_1111111111111111_1110100100011100_1001101001111011"; -- -0.08940729620397987
	pesos_i(21271) := b"0000000000000000_0000000000000000_0000001110001001_0000100010010111"; -- 0.013809716010877233
	pesos_i(21272) := b"1111111111111111_1111111111111111_1110100001001000_1011101111110010"; -- -0.09264016467074317
	pesos_i(21273) := b"0000000000000000_0000000000000000_0001100001100001_0010101011001111"; -- 0.09523265422238204
	pesos_i(21274) := b"1111111111111111_1111111111111111_1111011011101111_1001100100000110"; -- -0.03540652861228417
	pesos_i(21275) := b"0000000000000000_0000000000000000_0000000101110010_0001011111110001"; -- 0.005647178884278952
	pesos_i(21276) := b"1111111111111111_1111111111111111_1110011000111011_0100000000100010"; -- -0.10065840876095652
	pesos_i(21277) := b"1111111111111111_1111111111111111_1101101001001110_1101100110101011"; -- -0.14723434049764597
	pesos_i(21278) := b"0000000000000000_0000000000000000_0001111100101101_0011111011110110"; -- 0.1217841483043449
	pesos_i(21279) := b"1111111111111111_1111111111111111_1111100010100100_0101100111100100"; -- -0.028742200687249638
	pesos_i(21280) := b"0000000000000000_0000000000000000_0001011000100101_0110111001110011"; -- 0.0865086585581552
	pesos_i(21281) := b"1111111111111111_1111111111111111_1110011010010010_1111000011100000"; -- -0.09932035956145906
	pesos_i(21282) := b"0000000000000000_0000000000000000_0001000100110110_1100001110001011"; -- 0.0672418799200448
	pesos_i(21283) := b"0000000000000000_0000000000000000_0000111000101001_1101111111000111"; -- 0.0553264485640655
	pesos_i(21284) := b"0000000000000000_0000000000000000_0001101100010011_1001001111010111"; -- 0.10576747895071306
	pesos_i(21285) := b"0000000000000000_0000000000000000_0001100110011111_0000100101000100"; -- 0.1000829496621273
	pesos_i(21286) := b"0000000000000000_0000000000000000_0000101010001011_0000000001001010"; -- 0.04118348888306997
	pesos_i(21287) := b"1111111111111111_1111111111111111_1101100100100011_1001101110100110"; -- -0.15180041493887056
	pesos_i(21288) := b"0000000000000000_0000000000000000_0000101111100111_0001010101010001"; -- 0.046494800833224444
	pesos_i(21289) := b"0000000000000000_0000000000000000_0010000011010010_1110010101010111"; -- 0.12821801540552147
	pesos_i(21290) := b"1111111111111111_1111111111111111_1111100110101000_0100011001010110"; -- -0.024776081175004627
	pesos_i(21291) := b"0000000000000000_0000000000000000_0001101000000101_1011011001001100"; -- 0.1016496596624429
	pesos_i(21292) := b"0000000000000000_0000000000000000_0010011001011010_1011111011100011"; -- 0.14982216866331843
	pesos_i(21293) := b"0000000000000000_0000000000000000_0000011100001001_0011110000111101"; -- 0.027484669633604037
	pesos_i(21294) := b"1111111111111111_1111111111111111_1111010110111100_0111111101111110"; -- -0.04009249844985805
	pesos_i(21295) := b"0000000000000000_0000000000000000_0000100000110011_0000000010011001"; -- 0.032028233780266195
	pesos_i(21296) := b"1111111111111111_1111111111111111_1101110000110000_0101110100101100"; -- -0.13988702469068218
	pesos_i(21297) := b"0000000000000000_0000000000000000_0000001010011001_0100111010111000"; -- 0.010151786667759772
	pesos_i(21298) := b"1111111111111111_1111111111111111_1101110111011011_1001010011000100"; -- -0.1333682080209318
	pesos_i(21299) := b"1111111111111111_1111111111111111_1111011000100000_1100111110000010"; -- -0.03856185033346144
	pesos_i(21300) := b"0000000000000000_0000000000000000_0000000111011101_0101101101101110"; -- 0.007283891934485957
	pesos_i(21301) := b"1111111111111111_1111111111111111_1111100010010010_1001010011101011"; -- -0.029013340652158888
	pesos_i(21302) := b"0000000000000000_0000000000000000_0001111001111011_1100111010001100"; -- 0.11907664219821132
	pesos_i(21303) := b"0000000000000000_0000000000000000_0010001111111011_0111111001010010"; -- 0.14055623541747966
	pesos_i(21304) := b"0000000000000000_0000000000000000_0000110001110011_1010100000011011"; -- 0.0486397806701896
	pesos_i(21305) := b"0000000000000000_0000000000000000_0000111111101111_0000110011011000"; -- 0.06224136612216373
	pesos_i(21306) := b"0000000000000000_0000000000000000_0000101001110100_1011111110100101"; -- 0.040843942397723
	pesos_i(21307) := b"0000000000000000_0000000000000000_0001100100010001_1000100111111000"; -- 0.09792387298884044
	pesos_i(21308) := b"1111111111111111_1111111111111111_1111000101100111_0100111000111010"; -- -0.057017432105329495
	pesos_i(21309) := b"0000000000000000_0000000000000000_0000110000110111_0000111011101100"; -- 0.04771512289781587
	pesos_i(21310) := b"0000000000000000_0000000000000000_0000000111111101_1100001111010110"; -- 0.007778396273282055
	pesos_i(21311) := b"1111111111111111_1111111111111111_1111110100100111_1001110010101110"; -- -0.011114318335737379
	pesos_i(21312) := b"0000000000000000_0000000000000000_0010000001100100_0111101110100010"; -- 0.12653324804847957
	pesos_i(21313) := b"0000000000000000_0000000000000000_0001011100101100_0111110010011111"; -- 0.09052256465377206
	pesos_i(21314) := b"0000000000000000_0000000000000000_0001111010100011_1111000010110100"; -- 0.11968902952562359
	pesos_i(21315) := b"1111111111111111_1111111111111111_1110100001011101_0010010110111111"; -- -0.0923286828185683
	pesos_i(21316) := b"0000000000000000_0000000000000000_0001111010001001_1101101001110011"; -- 0.11929097478058284
	pesos_i(21317) := b"0000000000000000_0000000000000000_0001011000111010_1110110101110000"; -- 0.08683666203121042
	pesos_i(21318) := b"0000000000000000_0000000000000000_0010001010101011_0100101011011010"; -- 0.1354262144804884
	pesos_i(21319) := b"0000000000000000_0000000000000000_0010001101000110_0011000010110101"; -- 0.13778976829406425
	pesos_i(21320) := b"1111111111111111_1111111111111111_1111000001011010_1100010111011000"; -- -0.06111491664093261
	pesos_i(21321) := b"0000000000000000_0000000000000000_0000110010011111_0000011111001010"; -- 0.04930161183539842
	pesos_i(21322) := b"1111111111111111_1111111111111111_1111001111110011_0111011111110111"; -- -0.04706621390384919
	pesos_i(21323) := b"0000000000000000_0000000000000000_0001101100111110_1000101111000010"; -- 0.10642312513512998
	pesos_i(21324) := b"1111111111111111_1111111111111111_1110100010101000_0111101011110100"; -- -0.0911791949535947
	pesos_i(21325) := b"1111111111111111_1111111111111111_1111110010110010_0010000001000010"; -- -0.012907012923599805
	pesos_i(21326) := b"0000000000000000_0000000000000000_0001010001100111_1011111100001111"; -- 0.07970804319428396
	pesos_i(21327) := b"1111111111111111_1111111111111111_1110101010110101_1100010001100000"; -- -0.08316395424958883
	pesos_i(21328) := b"1111111111111111_1111111111111111_1101110010011110_0101111000111100"; -- -0.13820849461639179
	pesos_i(21329) := b"1111111111111111_1111111111111111_1101100100001100_0101110111011101"; -- -0.15215504984542438
	pesos_i(21330) := b"0000000000000000_0000000000000000_0000000011101011_1011110110100000"; -- 0.0035971178468707007
	pesos_i(21331) := b"1111111111111111_1111111111111111_1110110101110011_0111111110001011"; -- -0.0724563870599195
	pesos_i(21332) := b"0000000000000000_0000000000000000_0000000101001000_1110100100010101"; -- 0.005018775679722711
	pesos_i(21333) := b"0000000000000000_0000000000000000_0001010010001001_0001110111100010"; -- 0.08021723527306834
	pesos_i(21334) := b"1111111111111111_1111111111111111_1101111100000100_0001001000001001"; -- -0.12884413991204932
	pesos_i(21335) := b"0000000000000000_0000000000000000_0001011100101100_0111101111001101"; -- 0.09052251587296144
	pesos_i(21336) := b"1111111111111111_1111111111111111_1101110001001100_0010111000011011"; -- -0.1394625839193535
	pesos_i(21337) := b"1111111111111111_1111111111111111_1111111011101011_0010011100010110"; -- -0.0042243547764988666
	pesos_i(21338) := b"0000000000000000_0000000000000000_0000111110010000_0000000001101100"; -- 0.06079104087283045
	pesos_i(21339) := b"0000000000000000_0000000000000000_0001110110100011_1001010001101101"; -- 0.11577727957106093
	pesos_i(21340) := b"0000000000000000_0000000000000000_0000100000001111_0011101001010101"; -- 0.03148235876872258
	pesos_i(21341) := b"0000000000000000_0000000000000000_0001110010011010_1100000010101100"; -- 0.1117363376547923
	pesos_i(21342) := b"0000000000000000_0000000000000000_0000000010100101_1011010001000111"; -- 0.002528445616525877
	pesos_i(21343) := b"1111111111111111_1111111111111111_1111000011111001_0101000001010011"; -- -0.05869577378850578
	pesos_i(21344) := b"1111111111111111_1111111111111111_1111101001011011_0001111000001111"; -- -0.022047158569972043
	pesos_i(21345) := b"1111111111111111_1111111111111111_1111101010001111_0110001001000010"; -- -0.021249636517971897
	pesos_i(21346) := b"0000000000000000_0000000000000000_0000110010100011_0110111100000010"; -- 0.04936879910551225
	pesos_i(21347) := b"1111111111111111_1111111111111111_1110011000011110_0101101010111001"; -- -0.10109932889853812
	pesos_i(21348) := b"0000000000000000_0000000000000000_0000100010101010_1000100110111011"; -- 0.03385220352037984
	pesos_i(21349) := b"1111111111111111_1111111111111111_1111101111111011_1001000001100101"; -- -0.015692687337462582
	pesos_i(21350) := b"0000000000000000_0000000000000000_0001101010101101_0110011101010010"; -- 0.10420842890219799
	pesos_i(21351) := b"1111111111111111_1111111111111111_1110011011111110_0001010001100110"; -- -0.09768555168114168
	pesos_i(21352) := b"1111111111111111_1111111111111111_1111110101101110_1010110110001101"; -- -0.010029938811059121
	pesos_i(21353) := b"1111111111111111_1111111111111111_1110010001000001_0000101011110100"; -- -0.10838252594291749
	pesos_i(21354) := b"1111111111111111_1111111111111111_1110100000011101_0000110010101111"; -- -0.09330673915576862
	pesos_i(21355) := b"0000000000000000_0000000000000000_0001101001010111_1010111010001100"; -- 0.10290041853939956
	pesos_i(21356) := b"1111111111111111_1111111111111111_1111110011110110_0011111101000101"; -- -0.01186756674665732
	pesos_i(21357) := b"0000000000000000_0000000000000000_0001001111011111_1100100101100100"; -- 0.07763346386912284
	pesos_i(21358) := b"1111111111111111_1111111111111111_1111001101011111_1010010001001100"; -- -0.04932187210077389
	pesos_i(21359) := b"1111111111111111_1111111111111111_1110100101100000_1000110111001101"; -- -0.08837045415540337
	pesos_i(21360) := b"1111111111111111_1111111111111111_1111011001001100_1001101011110010"; -- -0.03789359658419198
	pesos_i(21361) := b"0000000000000000_0000000000000000_0010010111100011_0011000001001001"; -- 0.14799787323668212
	pesos_i(21362) := b"0000000000000000_0000000000000000_0001010110010111_0101011010110110"; -- 0.08434049545654922
	pesos_i(21363) := b"1111111111111111_1111111111111111_1111111011000110_0110100100001111"; -- -0.004784997708826291
	pesos_i(21364) := b"1111111111111111_1111111111111111_1110010110110111_1010001110101010"; -- -0.10266663651092374
	pesos_i(21365) := b"0000000000000000_0000000000000000_0010000110110011_1011100100010111"; -- 0.13164860546469745
	pesos_i(21366) := b"0000000000000000_0000000000000000_0010010101101101_1011111001110001"; -- 0.14620580925360188
	pesos_i(21367) := b"0000000000000000_0000000000000000_0000101010011100_1010011000100101"; -- 0.04145277402138036
	pesos_i(21368) := b"0000000000000000_0000000000000000_0000011111101111_0011100010011111"; -- 0.030993975471195638
	pesos_i(21369) := b"1111111111111111_1111111111111111_1110101100101011_1011111110101110"; -- -0.08136369709396264
	pesos_i(21370) := b"1111111111111111_1111111111111111_1111001101010110_1100101011101000"; -- -0.04945689988493585
	pesos_i(21371) := b"0000000000000000_0000000000000000_0010011110100110_0001110001000000"; -- 0.1548783928834127
	pesos_i(21372) := b"0000000000000000_0000000000000000_0001110111011101_1000001110111110"; -- 0.11666129492710864
	pesos_i(21373) := b"1111111111111111_1111111111111111_1110111101101110_0000111000100111"; -- -0.06472693965765204
	pesos_i(21374) := b"0000000000000000_0000000000000000_0000101001010011_0100110001110111"; -- 0.040333537218124035
	pesos_i(21375) := b"0000000000000000_0000000000000000_0001100000001001_1110110110000101"; -- 0.09390148638591998
	pesos_i(21376) := b"1111111111111111_1111111111111111_1110000101010101_1110001001110100"; -- -0.1197832553873368
	pesos_i(21377) := b"1111111111111111_1111111111111111_1111001010100001_1011110100000100"; -- -0.05221956882125085
	pesos_i(21378) := b"0000000000000000_0000000000000000_0000100100011011_1110110100010101"; -- 0.035582368537983675
	pesos_i(21379) := b"1111111111111111_1111111111111111_1110011100011010_1011110100000010"; -- -0.09724825583234031
	pesos_i(21380) := b"0000000000000000_0000000000000000_0010010100100111_1010000000001010"; -- 0.14513588183683174
	pesos_i(21381) := b"1111111111111111_1111111111111111_1110111101011111_0101011010100111"; -- -0.06495150010278762
	pesos_i(21382) := b"1111111111111111_1111111111111111_1110001001110101_0011011000111101"; -- -0.11539898885779452
	pesos_i(21383) := b"1111111111111111_1111111111111111_1111001000011010_0001011010011000"; -- -0.05428942473656753
	pesos_i(21384) := b"1111111111111111_1111111111111111_1111011110101111_1001001111001011"; -- -0.03247715273949562
	pesos_i(21385) := b"1111111111111111_1111111111111111_1110101001000110_0000010011000011"; -- -0.0848691010281714
	pesos_i(21386) := b"1111111111111111_1111111111111111_1111110011000101_1110101000011001"; -- -0.012605065198523304
	pesos_i(21387) := b"0000000000000000_0000000000000000_0010110100010000_1011010000010011"; -- 0.17603612379929937
	pesos_i(21388) := b"1111111111111111_1111111111111111_1110101000000110_1010111000110001"; -- -0.08583556476043461
	pesos_i(21389) := b"1111111111111111_1111111111111111_1110111110011110_0100111011011100"; -- -0.06399066099951234
	pesos_i(21390) := b"1111111111111111_1111111111111111_1110101000001010_1001001111110001"; -- -0.0857760941234934
	pesos_i(21391) := b"1111111111111111_1111111111111111_1111100011111110_0111101111000011"; -- -0.02736689074372869
	pesos_i(21392) := b"0000000000000000_0000000000000000_0000100001000100_1010000110101111"; -- 0.03229723468633513
	pesos_i(21393) := b"0000000000000000_0000000000000000_0010010010111001_0000010100001000"; -- 0.14344817592562153
	pesos_i(21394) := b"0000000000000000_0000000000000000_0001001000001000_0111101000100110"; -- 0.07044185100340117
	pesos_i(21395) := b"0000000000000000_0000000000000000_0000110110011110_0001110110010110"; -- 0.053193902094620785
	pesos_i(21396) := b"1111111111111111_1111111111111111_1111101101101010_0001100101100100"; -- -0.01791230498274271
	pesos_i(21397) := b"0000000000000000_0000000000000000_0001010100000000_0101100010001010"; -- 0.08203652727883973
	pesos_i(21398) := b"1111111111111111_1111111111111111_1111000100011111_0110001011010010"; -- -0.05811483733424391
	pesos_i(21399) := b"0000000000000000_0000000000000000_0000100111010000_0011001000001101"; -- 0.0383330614717241
	pesos_i(21400) := b"0000000000000000_0000000000000000_0001010001110011_0100000010000110"; -- 0.07988360657205391
	pesos_i(21401) := b"0000000000000000_0000000000000000_0001000101001111_0000010011011010"; -- 0.06761198358658992
	pesos_i(21402) := b"1111111111111111_1111111111111111_1111001000001100_0111110101000001"; -- -0.05449692870723181
	pesos_i(21403) := b"0000000000000000_0000000000000000_0000011011011111_1111100111110111"; -- 0.02685510907872767
	pesos_i(21404) := b"1111111111111111_1111111111111111_1110100001011010_0111000001101101"; -- -0.09237000791340062
	pesos_i(21405) := b"0000000000000000_0000000000000000_0000010010101011_1010011101110000"; -- 0.018244233064769036
	pesos_i(21406) := b"1111111111111111_1111111111111111_1110100111000101_1000100111010001"; -- -0.08682955415666428
	pesos_i(21407) := b"0000000000000000_0000000000000000_0000000100100110_1000110100110010"; -- 0.004494499915618464
	pesos_i(21408) := b"0000000000000000_0000000000000000_0010010111000111_1111101101111011"; -- 0.14758273853774787
	pesos_i(21409) := b"1111111111111111_1111111111111111_1101111111110010_0111110001011001"; -- -0.1252062112787361
	pesos_i(21410) := b"1111111111111111_1111111111111111_1111001010010111_1001001011101010"; -- -0.05237466600325541
	pesos_i(21411) := b"1111111111111111_1111111111111111_1110011100100001_0110010001101100"; -- -0.09714672431693017
	pesos_i(21412) := b"1111111111111111_1111111111111111_1111100001001101_0011001100111001"; -- -0.030072020190083183
	pesos_i(21413) := b"1111111111111111_1111111111111111_1110111100011010_1101111110110110"; -- -0.06599618734884888
	pesos_i(21414) := b"0000000000000000_0000000000000000_0000000100101000_1000110001011111"; -- 0.00452496830671806
	pesos_i(21415) := b"0000000000000000_0000000000000000_0000100000110010_0100000001001110"; -- 0.03201677237104639
	pesos_i(21416) := b"0000000000000000_0000000000000000_0001111011001000_0111001110110001"; -- 0.12024615364073256
	pesos_i(21417) := b"0000000000000000_0000000000000000_0001010110101010_0101010001110100"; -- 0.08463027791136721
	pesos_i(21418) := b"0000000000000000_0000000000000000_0010000001001011_1111000101111101"; -- 0.12615880293922677
	pesos_i(21419) := b"0000000000000000_0000000000000000_0010000000001100_1001110111111010"; -- 0.12519252171077122
	pesos_i(21420) := b"1111111111111111_1111111111111111_1111000110000001_1111110101000000"; -- -0.056610271364176824
	pesos_i(21421) := b"0000000000000000_0000000000000000_0001011100111001_1010000110110010"; -- 0.09072313879870253
	pesos_i(21422) := b"1111111111111111_1111111111111111_1111010010100100_1110110000100000"; -- -0.0443584844187931
	pesos_i(21423) := b"1111111111111111_1111111111111111_1111001000000010_1111000011111101"; -- -0.05464261843755696
	pesos_i(21424) := b"1111111111111111_1111111111111111_1111100000100110_0110011110011111"; -- -0.030663989829119505
	pesos_i(21425) := b"0000000000000000_0000000000000000_0000110001011111_0100101110000001"; -- 0.04832908539849445
	pesos_i(21426) := b"0000000000000000_0000000000000000_0001111100000001_1110011011110010"; -- 0.12112277424321122
	pesos_i(21427) := b"0000000000000000_0000000000000000_0001000110100011_1101110100100111"; -- 0.06890661431915403
	pesos_i(21428) := b"0000000000000000_0000000000000000_0000101100100000_0100011101000011"; -- 0.04346127873191397
	pesos_i(21429) := b"0000000000000000_0000000000000000_0001111000011001_0000110000011111"; -- 0.11756969212547373
	pesos_i(21430) := b"0000000000000000_0000000000000000_0001000001100011_1010111011010110"; -- 0.0640210410708091
	pesos_i(21431) := b"0000000000000000_0000000000000000_0001111111110010_1100011011111011"; -- 0.12479823713019544
	pesos_i(21432) := b"0000000000000000_0000000000000000_0001111010011101_1010110001011001"; -- 0.11959340264621429
	pesos_i(21433) := b"1111111111111111_1111111111111111_1111000111001001_0001110100101100"; -- -0.05552499461520703
	pesos_i(21434) := b"0000000000000000_0000000000000000_0001010110000001_1110001010111111"; -- 0.08401314891637056
	pesos_i(21435) := b"1111111111111111_1111111111111111_1111101100110111_1101010010000100"; -- -0.01867934972080084
	pesos_i(21436) := b"1111111111111111_1111111111111111_1101100000100010_0011000001100110"; -- -0.15572831638580645
	pesos_i(21437) := b"1111111111111111_1111111111111111_1110110110011100_1110010111111111"; -- -0.07182467012416152
	pesos_i(21438) := b"0000000000000000_0000000000000000_0001011111111011_1101011100011101"; -- 0.0936865278301106
	pesos_i(21439) := b"0000000000000000_0000000000000000_0000001001110011_0010000101001110"; -- 0.009569245850308557
	pesos_i(21440) := b"1111111111111111_1111111111111111_1111111011010001_0001110100101110"; -- -0.004621673892554745
	pesos_i(21441) := b"1111111111111111_1111111111111111_1101111110110001_0110011100111101"; -- -0.12619929084299206
	pesos_i(21442) := b"0000000000000000_0000000000000000_0000000111001000_0000111100001100"; -- 0.006958904734150891
	pesos_i(21443) := b"1111111111111111_1111111111111111_1101110001101010_0010000101100111"; -- -0.13900557740689312
	pesos_i(21444) := b"0000000000000000_0000000000000000_0001101011011011_0000010111011100"; -- 0.10490452403476185
	pesos_i(21445) := b"1111111111111111_1111111111111111_1110011111011100_1001101111110110"; -- -0.0942900203611065
	pesos_i(21446) := b"0000000000000000_0000000000000000_0000001010100001_0011111110011100"; -- 0.0102729565358513
	pesos_i(21447) := b"0000000000000000_0000000000000000_0000000101000010_1101110001100100"; -- 0.004926466361083528
	pesos_i(21448) := b"0000000000000000_0000000000000000_0000101000001110_1000001011001100"; -- 0.0392839192293574
	pesos_i(21449) := b"1111111111111111_1111111111111111_1101110000001111_0010001010110111"; -- -0.14039404909707423
	pesos_i(21450) := b"0000000000000000_0000000000000000_0001001011110000_1100100111000111"; -- 0.073986636286423
	pesos_i(21451) := b"1111111111111111_1111111111111111_1111100010110100_0101100110110111"; -- -0.02849807050100435
	pesos_i(21452) := b"1111111111111111_1111111111111111_1110011111111001_0110011100100101"; -- -0.0938506635410227
	pesos_i(21453) := b"1111111111111111_1111111111111111_1110010000001001_1110110010010100"; -- -0.10922356965773003
	pesos_i(21454) := b"0000000000000000_0000000000000000_0000000111001101_0000100100000110"; -- 0.007034839693477468
	pesos_i(21455) := b"0000000000000000_0000000000000000_0000100010011110_1010111001011101"; -- 0.033671281508774666
	pesos_i(21456) := b"1111111111111111_1111111111111111_1111100000110001_0100110111110101"; -- -0.030497672798594475
	pesos_i(21457) := b"0000000000000000_0000000000000000_0000110110000000_0110000011100101"; -- 0.052740150383476674
	pesos_i(21458) := b"1111111111111111_1111111111111111_1110101100110111_1001010111010000"; -- -0.08118308703165693
	pesos_i(21459) := b"1111111111111111_1111111111111111_1110010001000000_1100010000011010"; -- -0.10838674883986348
	pesos_i(21460) := b"0000000000000000_0000000000000000_0001100001010100_0001000101100101"; -- 0.09503277511108807
	pesos_i(21461) := b"0000000000000000_0000000000000000_0000111010001010_1000110110011100"; -- 0.05680165354945838
	pesos_i(21462) := b"0000000000000000_0000000000000000_0000001001110011_0100010101101110"; -- 0.009571398975412754
	pesos_i(21463) := b"1111111111111111_1111111111111111_1110100011111011_1001100000011100"; -- -0.08991097760973187
	pesos_i(21464) := b"0000000000000000_0000000000000000_0010001100111111_1100111010111101"; -- 0.1376923763088381
	pesos_i(21465) := b"1111111111111111_1111111111111111_1111010001110010_1001000110000011"; -- -0.04512682483514256
	pesos_i(21466) := b"0000000000000000_0000000000000000_0000110111101000_0101101100111110"; -- 0.05432672754864175
	pesos_i(21467) := b"1111111111111111_1111111111111111_1111111011001101_0010111101000001"; -- -0.004681631767159124
	pesos_i(21468) := b"0000000000000000_0000000000000000_0010011001101101_0101011101000110"; -- 0.15010590995042572
	pesos_i(21469) := b"1111111111111111_1111111111111111_1111101000001010_0000111100100101"; -- -0.02328400941690712
	pesos_i(21470) := b"0000000000000000_0000000000000000_0000111111001111_1100011010101000"; -- 0.06176416018132377
	pesos_i(21471) := b"0000000000000000_0000000000000000_0000110100011001_1110111001001101"; -- 0.05117692354412699
	pesos_i(21472) := b"1111111111111111_1111111111111111_1110011111111111_0001100110000001"; -- -0.09376373865943591
	pesos_i(21473) := b"1111111111111111_1111111111111111_1101110101100001_1100100110110010"; -- -0.13522662542768654
	pesos_i(21474) := b"1111111111111111_1111111111111111_1111000011001010_0000011101001111"; -- -0.05941728900598573
	pesos_i(21475) := b"0000000000000000_0000000000000000_0000111110010001_1001100000100011"; -- 0.06081534257744976
	pesos_i(21476) := b"0000000000000000_0000000000000000_0001011101101000_0010010001000110"; -- 0.09143282614694286
	pesos_i(21477) := b"0000000000000000_0000000000000000_0001101000001101_1001100110111101"; -- 0.10177002784049127
	pesos_i(21478) := b"0000000000000000_0000000000000000_0010100010000111_1111100110010100"; -- 0.15832481244900262
	pesos_i(21479) := b"1111111111111111_1111111111111111_1111100111111101_1111111111001111"; -- -0.023468028919085115
	pesos_i(21480) := b"1111111111111111_1111111111111111_1101110101111010_1001110111010010"; -- -0.1348477708777894
	pesos_i(21481) := b"0000000000000000_0000000000000000_0000101011111111_1111011111111110"; -- 0.04296827272675912
	pesos_i(21482) := b"1111111111111111_1111111111111111_1101101100100011_1101001010010000"; -- -0.1439846418873109
	pesos_i(21483) := b"1111111111111111_1111111111111111_1111110000101100_0100100011101001"; -- -0.01494926760457443
	pesos_i(21484) := b"0000000000000000_0000000000000000_0000100101011000_1111011101101010"; -- 0.03651377055364719
	pesos_i(21485) := b"0000000000000000_0000000000000000_0000100100011100_0110010010110111"; -- 0.035589499100582685
	pesos_i(21486) := b"0000000000000000_0000000000000000_0000110100110111_1010011011001110"; -- 0.05163042565884364
	pesos_i(21487) := b"1111111111111111_1111111111111111_1111101101101001_0011010101000001"; -- -0.017925902946602963
	pesos_i(21488) := b"0000000000000000_0000000000000000_0000000101011011_0010110111101101"; -- 0.0052975371391557275
	pesos_i(21489) := b"0000000000000000_0000000000000000_0000111010110011_1111100110111011"; -- 0.057433708271215994
	pesos_i(21490) := b"1111111111111111_1111111111111111_1110101011011000_1111011010110110"; -- -0.08262689653916086
	pesos_i(21491) := b"1111111111111111_1111111111111111_1110011110111100_1110001001010101"; -- -0.09477410731934882
	pesos_i(21492) := b"1111111111111111_1111111111111111_1111101101001101_1110110101110010"; -- -0.018342170310421707
	pesos_i(21493) := b"0000000000000000_0000000000000000_0010011011101011_0011100001110100"; -- 0.15202668030917865
	pesos_i(21494) := b"1111111111111111_1111111111111111_1111111011101011_1011101001011100"; -- -0.004215576730401603
	pesos_i(21495) := b"1111111111111111_1111111111111111_1101110010101001_0100011011011010"; -- -0.13804204157850916
	pesos_i(21496) := b"0000000000000000_0000000000000000_0001001010100101_0001000111001100"; -- 0.07283126101810983
	pesos_i(21497) := b"0000000000000000_0000000000000000_0000011101010110_1110101111001011"; -- 0.02867006032063916
	pesos_i(21498) := b"1111111111111111_1111111111111111_1110000010011001_0111000010100001"; -- -0.1226586920873941
	pesos_i(21499) := b"1111111111111111_1111111111111111_1110010100111100_1101011111001011"; -- -0.10454036044074103
	pesos_i(21500) := b"1111111111111111_1111111111111111_1110001100101111_0011110100010110"; -- -0.11256044600677459
	pesos_i(21501) := b"1111111111111111_1111111111111111_1110010011101110_0111100100000100"; -- -0.10573619507939602
	pesos_i(21502) := b"0000000000000000_0000000000000000_0010011110010100_1101100010101001"; -- 0.15461496474309686
	pesos_i(21503) := b"0000000000000000_0000000000000000_0000010001100011_0001110010000111"; -- 0.01713732056426106
	pesos_i(21504) := b"0000000000000000_0000000000000000_0001111100000100_0001000110000100"; -- 0.12115582928488285
	pesos_i(21505) := b"0000000000000000_0000000000000000_0001111001101000_0001001101111110"; -- 0.11877557580824026
	pesos_i(21506) := b"1111111111111111_1111111111111111_1110000001001010_1011110111000100"; -- -0.12385953877190423
	pesos_i(21507) := b"0000000000000000_0000000000000000_0000111011100000_1111100100011111"; -- 0.05812031752185605
	pesos_i(21508) := b"1111111111111111_1111111111111111_1111011011111000_1001001001011001"; -- -0.03526959740289113
	pesos_i(21509) := b"0000000000000000_0000000000000000_0001000011100001_0100110100001011"; -- 0.06593781972399324
	pesos_i(21510) := b"0000000000000000_0000000000000000_0010001001011001_0010001101100101"; -- 0.1341726419119405
	pesos_i(21511) := b"0000000000000000_0000000000000000_0000000011100100_1100010011101011"; -- 0.0034907410361827685
	pesos_i(21512) := b"1111111111111111_1111111111111111_1111010001010101_0101000111000110"; -- -0.045573128892714455
	pesos_i(21513) := b"1111111111111111_1111111111111111_1101111000101011_1011001110000010"; -- -0.1321456726547726
	pesos_i(21514) := b"1111111111111111_1111111111111111_1110000110001111_1000001101100011"; -- -0.1189039118628846
	pesos_i(21515) := b"0000000000000000_0000000000000000_0000111010100101_0111010110111110"; -- 0.05721221815781634
	pesos_i(21516) := b"1111111111111111_1111111111111111_1110110010100101_1000101001100011"; -- -0.07559905141480976
	pesos_i(21517) := b"0000000000000000_0000000000000000_0000000100000110_1000110101110001"; -- 0.004006233328163806
	pesos_i(21518) := b"1111111111111111_1111111111111111_1111100000111100_1101100001110011"; -- -0.030321571176145066
	pesos_i(21519) := b"1111111111111111_1111111111111111_1101111010101011_1110100011000000"; -- -0.13018937415186996
	pesos_i(21520) := b"0000000000000000_0000000000000000_0000001100000011_1110011111011110"; -- 0.011778346838950063
	pesos_i(21521) := b"0000000000000000_0000000000000000_0001110010010011_1000010110000000"; -- 0.11162599916540521
	pesos_i(21522) := b"0000000000000000_0000000000000000_0001111100000111_0100000010010000"; -- 0.12120440985970644
	pesos_i(21523) := b"1111111111111111_1111111111111111_1101110011001001_0110100100010011"; -- -0.13755172048178213
	pesos_i(21524) := b"1111111111111111_1111111111111111_1111110011101010_0111101110010010"; -- -0.012047077965806334
	pesos_i(21525) := b"0000000000000000_0000000000000000_0001111111010000_0000111010001110"; -- 0.12426844565449478
	pesos_i(21526) := b"0000000000000000_0000000000000000_0000101111011111_0010101110111011"; -- 0.04637406653393867
	pesos_i(21527) := b"0000000000000000_0000000000000000_0001101010011100_1011101000010101"; -- 0.10395396241268702
	pesos_i(21528) := b"0000000000000000_0000000000000000_0000011001100100_1101011100100110"; -- 0.024976202720255646
	pesos_i(21529) := b"0000000000000000_0000000000000000_0000011100111001_1011011001011011"; -- 0.028224370282941655
	pesos_i(21530) := b"0000000000000000_0000000000000000_0000101011101010_1000111100111001"; -- 0.04264159342342365
	pesos_i(21531) := b"1111111111111111_1111111111111111_1110000101001001_0110000110001000"; -- -0.11997404518815098
	pesos_i(21532) := b"1111111111111111_1111111111111111_1110001000110011_1110011101000011"; -- -0.11639551739230689
	pesos_i(21533) := b"1111111111111111_1111111111111111_1111011000011100_0100101110101010"; -- -0.038630743893411534
	pesos_i(21534) := b"0000000000000000_0000000000000000_0010001000110010_0011110011001011"; -- 0.13357906303540856
	pesos_i(21535) := b"1111111111111111_1111111111111111_1111111000010110_1001111010010101"; -- -0.007467354479135766
	pesos_i(21536) := b"1111111111111111_1111111111111111_1110101010110001_0011110011100001"; -- -0.08323306561134083
	pesos_i(21537) := b"0000000000000000_0000000000000000_0001101001001001_1110110111100011"; -- 0.1026905707163028
	pesos_i(21538) := b"1111111111111111_1111111111111111_1110010100111011_0101011110001001"; -- -0.10456326399516007
	pesos_i(21539) := b"1111111111111111_1111111111111111_1111010000001110_0101111000001101"; -- -0.04665577100596983
	pesos_i(21540) := b"1111111111111111_1111111111111111_1111011110001000_0110000110111100"; -- -0.03307522925228617
	pesos_i(21541) := b"0000000000000000_0000000000000000_0001111010101001_1000111111010000"; -- 0.11977480726915185
	pesos_i(21542) := b"0000000000000000_0000000000000000_0001001010011111_1001110000010111"; -- 0.0727479511513561
	pesos_i(21543) := b"0000000000000000_0000000000000000_0000000110000111_1110110001011001"; -- 0.005980273905197965
	pesos_i(21544) := b"1111111111111111_1111111111111111_1111101111100011_0100110100111011"; -- -0.01606290156311659
	pesos_i(21545) := b"0000000000000000_0000000000000000_0010000001101001_1110101001000101"; -- 0.12661613631880983
	pesos_i(21546) := b"1111111111111111_1111111111111111_1110111001110001_0111011001000111"; -- -0.0685812069934216
	pesos_i(21547) := b"0000000000000000_0000000000000000_0000111101011100_0011001101001101"; -- 0.06000061643722481
	pesos_i(21548) := b"1111111111111111_1111111111111111_1111111000011010_1101011011001100"; -- -0.007402968520422625
	pesos_i(21549) := b"0000000000000000_0000000000000000_0001110111001111_0000100001110100"; -- 0.11644032310070078
	pesos_i(21550) := b"0000000000000000_0000000000000000_0001010000100001_1001001111001001"; -- 0.07863734867927209
	pesos_i(21551) := b"1111111111111111_1111111111111111_1110101000101000_0100001111100001"; -- -0.08532310260168234
	pesos_i(21552) := b"1111111111111111_1111111111111111_1110000010001101_0100110011011011"; -- -0.12284392970783393
	pesos_i(21553) := b"0000000000000000_0000000000000000_0001010100100100_1110011100010100"; -- 0.08259433974819941
	pesos_i(21554) := b"1111111111111111_1111111111111111_1111001110100101_0100101000001100"; -- -0.0482591363582614
	pesos_i(21555) := b"0000000000000000_0000000000000000_0000001100001000_0011100111101101"; -- 0.011844273022146098
	pesos_i(21556) := b"1111111111111111_1111111111111111_1110101000111001_0000011110110001"; -- -0.08506729050862484
	pesos_i(21557) := b"1111111111111111_1111111111111111_1101101100111010_1100110001000100"; -- -0.14363406504861287
	pesos_i(21558) := b"0000000000000000_0000000000000000_0001000011011101_0000001111000011"; -- 0.06587241664279045
	pesos_i(21559) := b"1111111111111111_1111111111111111_1111000111011110_1111001011011000"; -- -0.05519182428571353
	pesos_i(21560) := b"0000000000000000_0000000000000000_0010000011110010_1101110000100011"; -- 0.12870574819172106
	pesos_i(21561) := b"0000000000000000_0000000000000000_0001100101111100_1001100101010100"; -- 0.09955747882501925
	pesos_i(21562) := b"1111111111111111_1111111111111111_1110101011011111_1000110111001111"; -- -0.0825263375580449
	pesos_i(21563) := b"0000000000000000_0000000000000000_0000010001001111_0111001011101110"; -- 0.01683729460836759
	pesos_i(21564) := b"1111111111111111_1111111111111111_1111100010101101_1011101110011110"; -- -0.02859904670057464
	pesos_i(21565) := b"0000000000000000_0000000000000000_0001101010001101_0100001001111110"; -- 0.10371795241254943
	pesos_i(21566) := b"0000000000000000_0000000000000000_0001101010001101_0001100010100011"; -- 0.10371545779620207
	pesos_i(21567) := b"0000000000000000_0000000000000000_0000011101111101_0011011110100100"; -- 0.029254415150869406
	pesos_i(21568) := b"1111111111111111_1111111111111111_1111101000011110_1100100000010000"; -- -0.022967811667023517
	pesos_i(21569) := b"0000000000000000_0000000000000000_0000101101000100_1010001001101101"; -- 0.044016028888672835
	pesos_i(21570) := b"0000000000000000_0000000000000000_0010001111101001_0111001011110011"; -- 0.14028089932361051
	pesos_i(21571) := b"0000000000000000_0000000000000000_0000100010110110_0110100011101001"; -- 0.0340333527928831
	pesos_i(21572) := b"1111111111111111_1111111111111111_1110110101100111_0111101110101001"; -- -0.07263972411051897
	pesos_i(21573) := b"0000000000000000_0000000000000000_0000101110010101_0111100110010100"; -- 0.0452495561301081
	pesos_i(21574) := b"0000000000000000_0000000000000000_0001011000011101_0110010100001111"; -- 0.08638602839092012
	pesos_i(21575) := b"0000000000000000_0000000000000000_0000011111101111_0001111000010101"; -- 0.03099239362180064
	pesos_i(21576) := b"0000000000000000_0000000000000000_0010001101101010_1000111000011100"; -- 0.1383446520110435
	pesos_i(21577) := b"1111111111111111_1111111111111111_1111010110010000_0100110100000110"; -- -0.04076689331054882
	pesos_i(21578) := b"0000000000000000_0000000000000000_0001100111101101_0001011111100100"; -- 0.101274007086623
	pesos_i(21579) := b"1111111111111111_1111111111111111_1101110001101010_0010100110000101"; -- -0.1390050934866692
	pesos_i(21580) := b"1111111111111111_1111111111111111_1111100110100010_0010011111000101"; -- -0.024869455649606298
	pesos_i(21581) := b"1111111111111111_1111111111111111_1110111101110110_0001100010100000"; -- -0.06460424516852306
	pesos_i(21582) := b"0000000000000000_0000000000000000_0000010111100010_1100101101000111"; -- 0.022991852680944214
	pesos_i(21583) := b"0000000000000000_0000000000000000_0001110110110000_1011100100010101"; -- 0.1159778285447438
	pesos_i(21584) := b"1111111111111111_1111111111111111_1111010001011001_0000110010101010"; -- -0.04551621292074459
	pesos_i(21585) := b"0000000000000000_0000000000000000_0000010101010100_1111100001110101"; -- 0.020827797398413304
	pesos_i(21586) := b"1111111111111111_1111111111111111_1110110010100001_1011001001001011"; -- -0.07565770794495269
	pesos_i(21587) := b"1111111111111111_1111111111111111_1101101100010101_1010111110101100"; -- -0.14420034459652545
	pesos_i(21588) := b"0000000000000000_0000000000000000_0001010011001000_0011111000101011"; -- 0.08118046329558241
	pesos_i(21589) := b"1111111111111111_1111111111111111_1101110110110001_1011001000000111"; -- -0.13400733315244434
	pesos_i(21590) := b"1111111111111111_1111111111111111_1110001101101100_0100100111110001"; -- -0.11162889354735145
	pesos_i(21591) := b"1111111111111111_1111111111111111_1110011110010001_1010101011000000"; -- -0.09543354813961187
	pesos_i(21592) := b"0000000000000000_0000000000000000_0000101000010100_0011000001111100"; -- 0.0393705657574454
	pesos_i(21593) := b"1111111111111111_1111111111111111_1111101111001110_0000000000001001"; -- -0.016387937244618365
	pesos_i(21594) := b"1111111111111111_1111111111111111_1111000100100101_0111100110111110"; -- -0.05802191847304364
	pesos_i(21595) := b"1111111111111111_1111111111111111_1110111011100101_0100100010100011"; -- -0.06681390782501752
	pesos_i(21596) := b"1111111111111111_1111111111111111_1111010100100100_0110000000110001"; -- -0.042413700043893755
	pesos_i(21597) := b"1111111111111111_1111111111111111_1111001011100111_0010110101110110"; -- -0.05116000996026472
	pesos_i(21598) := b"0000000000000000_0000000000000000_0000101101100100_1111111010011111"; -- 0.044509805438942944
	pesos_i(21599) := b"1111111111111111_1111111111111111_1111101100101010_1000110000101100"; -- -0.018882025944869894
	pesos_i(21600) := b"1111111111111111_1111111111111111_1110110010000000_0101010010111100"; -- -0.07616682439926503
	pesos_i(21601) := b"1111111111111111_1111111111111111_1101100100001101_0001110000101101"; -- -0.15214370644544606
	pesos_i(21602) := b"1111111111111111_1111111111111111_1111010111000101_1110010011100111"; -- -0.0399491250255067
	pesos_i(21603) := b"1111111111111111_1111111111111111_1110110001000000_1100101110110000"; -- -0.07713629670327557
	pesos_i(21604) := b"1111111111111111_1111111111111111_1111110010001101_1111011110010001"; -- -0.013458754660789378
	pesos_i(21605) := b"0000000000000000_0000000000000000_0000100101001010_1000001111101011"; -- 0.03629326324826376
	pesos_i(21606) := b"1111111111111111_1111111111111111_1111011001100000_0101000101100110"; -- -0.03759280453865638
	pesos_i(21607) := b"1111111111111111_1111111111111111_1110011101001100_1010000000011010"; -- -0.09648703926396093
	pesos_i(21608) := b"0000000000000000_0000000000000000_0000001111010110_0101111101110010"; -- 0.014989819938357747
	pesos_i(21609) := b"1111111111111111_1111111111111111_1111000100010000_0001000110101010"; -- -0.05834855643539057
	pesos_i(21610) := b"0000000000000000_0000000000000000_0000010000010010_0111010111011101"; -- 0.015906683331954732
	pesos_i(21611) := b"0000000000000000_0000000000000000_0001111101010010_0000011110001100"; -- 0.12234542059469469
	pesos_i(21612) := b"1111111111111111_1111111111111111_1111001100000011_1100110010011010"; -- -0.05072327839129808
	pesos_i(21613) := b"0000000000000000_0000000000000000_0000100011011001_0110011110110001"; -- 0.03456733770702466
	pesos_i(21614) := b"0000000000000000_0000000000000000_0010011100111110_0000011101111000"; -- 0.15329024011157383
	pesos_i(21615) := b"1111111111111111_1111111111111111_1101100101110101_1101010000100010"; -- -0.15054582747686118
	pesos_i(21616) := b"1111111111111111_1111111111111111_1111100111011110_0010001000100101"; -- -0.023954263766651177
	pesos_i(21617) := b"0000000000000000_0000000000000000_0000011100111010_0101011100011001"; -- 0.028233951297296996
	pesos_i(21618) := b"1111111111111111_1111111111111111_1111110100001011_1101110010110000"; -- -0.011537749319835613
	pesos_i(21619) := b"0000000000000000_0000000000000000_0001100101100110_0000011010000111"; -- 0.09921303542874321
	pesos_i(21620) := b"1111111111111111_1111111111111111_1101110001001001_1001110100010110"; -- -0.13950174537488913
	pesos_i(21621) := b"1111111111111111_1111111111111111_1111000101001100_1110001110100111"; -- -0.05742051278902262
	pesos_i(21622) := b"0000000000000000_0000000000000000_0000010101011000_0001101011100101"; -- 0.020875626520347704
	pesos_i(21623) := b"1111111111111111_1111111111111111_1101111010001101_0111101111000010"; -- -0.130653634225279
	pesos_i(21624) := b"0000000000000000_0000000000000000_0010001111011110_0101101010110001"; -- 0.1401116068309078
	pesos_i(21625) := b"0000000000000000_0000000000000000_0000011101011110_0000110110001101"; -- 0.0287788838549892
	pesos_i(21626) := b"1111111111111111_1111111111111111_1111111011000011_0000101010100111"; -- -0.0048364011780736025
	pesos_i(21627) := b"1111111111111111_1111111111111111_1110011101101100_0101110000100000"; -- -0.09600280976322025
	pesos_i(21628) := b"1111111111111111_1111111111111111_1110001100010011_1000111100111101"; -- -0.11298279529589461
	pesos_i(21629) := b"1111111111111111_1111111111111111_1111101010100001_0010111001011000"; -- -0.020978072604609717
	pesos_i(21630) := b"1111111111111111_1111111111111111_1111000011100000_0101111010110011"; -- -0.059076386703963715
	pesos_i(21631) := b"1111111111111111_1111111111111111_1111111000011100_1101000110100001"; -- -0.0073727590774848
	pesos_i(21632) := b"1111111111111111_1111111111111111_1111100011010101_1000011100011110"; -- -0.027991824211603043
	pesos_i(21633) := b"0000000000000000_0000000000000000_0000100111111000_0010110010100000"; -- 0.03894308952569228
	pesos_i(21634) := b"1111111111111111_1111111111111111_1110101011100010_1001111100100100"; -- -0.08247952823988519
	pesos_i(21635) := b"0000000000000000_0000000000000000_0001011100100101_0000011010000001"; -- 0.09040871283654019
	pesos_i(21636) := b"1111111111111111_1111111111111111_1110011000011000_0011010110110010"; -- -0.1011930885509733
	pesos_i(21637) := b"0000000000000000_0000000000000000_0000011000101000_1100001111111110"; -- 0.024059533698678186
	pesos_i(21638) := b"1111111111111111_1111111111111111_1111011001100100_0111011001100101"; -- -0.03752956417085827
	pesos_i(21639) := b"1111111111111111_1111111111111111_1110110000100100_0110100010100010"; -- -0.07756944705886898
	pesos_i(21640) := b"0000000000000000_0000000000000000_0000111101010110_1001111111000010"; -- 0.05991552820050837
	pesos_i(21641) := b"0000000000000000_0000000000000000_0000100111010010_0110110111001101"; -- 0.038367140240996904
	pesos_i(21642) := b"1111111111111111_1111111111111111_1110011111010001_0010101011011010"; -- -0.09446460889792763
	pesos_i(21643) := b"1111111111111111_1111111111111111_1111110110101111_0000010000011001"; -- -0.009048217662018451
	pesos_i(21644) := b"1111111111111111_1111111111111111_1111101000001000_0110101110011110"; -- -0.02330901530969975
	pesos_i(21645) := b"0000000000000000_0000000000000000_0000110001000101_1001100000010111"; -- 0.04793692163582666
	pesos_i(21646) := b"0000000000000000_0000000000000000_0001011101010010_1100101100110100"; -- 0.09110708266832965
	pesos_i(21647) := b"1111111111111111_1111111111111111_1110001100000011_0001010001101111"; -- -0.11323425558733259
	pesos_i(21648) := b"1111111111111111_1111111111111111_1110101000011100_1101010101111000"; -- -0.0854975302879661
	pesos_i(21649) := b"0000000000000000_0000000000000000_0001110101100011_0010101101110110"; -- 0.11479446062860796
	pesos_i(21650) := b"0000000000000000_0000000000000000_0001100100000101_1011010011010110"; -- 0.0977433225406883
	pesos_i(21651) := b"0000000000000000_0000000000000000_0001110101001101_0011011011100010"; -- 0.11445944799326169
	pesos_i(21652) := b"0000000000000000_0000000000000000_0000111010001101_1010110001011011"; -- 0.056849262475360006
	pesos_i(21653) := b"1111111111111111_1111111111111111_1111111110011001_0011110011101110"; -- -0.0015680235258565668
	pesos_i(21654) := b"1111111111111111_1111111111111111_1111101110000011_0011101101000111"; -- -0.017528815517701784
	pesos_i(21655) := b"0000000000000000_0000000000000000_0000110010001100_1101000111000100"; -- 0.04902373336390263
	pesos_i(21656) := b"1111111111111111_1111111111111111_1110101011111111_0111001100101011"; -- -0.08203964430995533
	pesos_i(21657) := b"1111111111111111_1111111111111111_1110101000101000_0101010111111010"; -- -0.08532202372493747
	pesos_i(21658) := b"1111111111111111_1111111111111111_1111111110010001_0110110010011010"; -- -0.0016872523834103447
	pesos_i(21659) := b"1111111111111111_1111111111111111_1111110101010010_0100011110001010"; -- -0.010463265345153856
	pesos_i(21660) := b"1111111111111111_1111111111111111_1101100001010100_1110111001110000"; -- -0.15495404984607994
	pesos_i(21661) := b"0000000000000000_0000000000000000_0001000010110111_0101101101110011"; -- 0.0652978091550075
	pesos_i(21662) := b"1111111111111111_1111111111111111_1101110001111011_1101101000111011"; -- -0.13873516146346287
	pesos_i(21663) := b"0000000000000000_0000000000000000_0001011010100111_1100111010010011"; -- 0.08849803056246731
	pesos_i(21664) := b"0000000000000000_0000000000000000_0001010011000110_1101111001111111"; -- 0.0811595021237286
	pesos_i(21665) := b"0000000000000000_0000000000000000_0000000101101101_1001001101101100"; -- 0.005578245011016558
	pesos_i(21666) := b"1111111111111111_1111111111111111_1111100011011111_0000000011000101"; -- -0.02784724422925001
	pesos_i(21667) := b"0000000000000000_0000000000000000_0001101000010111_1101101101001110"; -- 0.10192652383968259
	pesos_i(21668) := b"0000000000000000_0000000000000000_0001111010100000_0001001010010010"; -- 0.11963001308159224
	pesos_i(21669) := b"0000000000000000_0000000000000000_0010010100111010_0010110100101001"; -- 0.14541895154824203
	pesos_i(21670) := b"1111111111111111_1111111111111111_1110111000010001_0111110000011011"; -- -0.07004570330536082
	pesos_i(21671) := b"1111111111111111_1111111111111111_1111111000001100_1010110001001001"; -- -0.007619125480488272
	pesos_i(21672) := b"0000000000000000_0000000000000000_0010010100100101_0001110111110100"; -- 0.1450976106420139
	pesos_i(21673) := b"1111111111111111_1111111111111111_1110111010111000_1010000000100001"; -- -0.06749533846536898
	pesos_i(21674) := b"0000000000000000_0000000000000000_0000001100000001_0111010110000110"; -- 0.011741013689631315
	pesos_i(21675) := b"0000000000000000_0000000000000000_0010001011001001_0101111110101011"; -- 0.13588521891512745
	pesos_i(21676) := b"0000000000000000_0000000000000000_0001000111001011_0101101001000010"; -- 0.06950916401917881
	pesos_i(21677) := b"0000000000000000_0000000000000000_0010000010100100_1000010100110110"; -- 0.1275103815122964
	pesos_i(21678) := b"1111111111111111_1111111111111111_1110000110001101_1000100001010111"; -- -0.11893413431847685
	pesos_i(21679) := b"0000000000000000_0000000000000000_0000110111000100_1000011000110110"; -- 0.05377997236276857
	pesos_i(21680) := b"1111111111111111_1111111111111111_1111111011011101_1111011100010000"; -- -0.004425581475636871
	pesos_i(21681) := b"1111111111111111_1111111111111111_1101100101010011_0101100001011110"; -- -0.15107200333726303
	pesos_i(21682) := b"0000000000000000_0000000000000000_0001100100101110_0001000010010101"; -- 0.09835914265885708
	pesos_i(21683) := b"0000000000000000_0000000000000000_0001011011001011_1101111010001011"; -- 0.08904829886845998
	pesos_i(21684) := b"1111111111111111_1111111111111111_1111001010110111_1000110010101110"; -- -0.051886756415372506
	pesos_i(21685) := b"0000000000000000_0000000000000000_0000110000101011_0010100011011011"; -- 0.04753356302383305
	pesos_i(21686) := b"1111111111111111_1111111111111111_1111011110000110_0011100110100010"; -- -0.033108137153427177
	pesos_i(21687) := b"0000000000000000_0000000000000000_0001001111101110_0010011100001110"; -- 0.07785266969170064
	pesos_i(21688) := b"0000000000000000_0000000000000000_0000111010011111_0100110110110101"; -- 0.057118279243980614
	pesos_i(21689) := b"0000000000000000_0000000000000000_0000011000110000_1111011000000011"; -- 0.024184585338479937
	pesos_i(21690) := b"1111111111111111_1111111111111111_1110001001110000_0110111000101010"; -- -0.11547194925665694
	pesos_i(21691) := b"0000000000000000_0000000000000000_0001001000011101_1010010101010110"; -- 0.07076485956546873
	pesos_i(21692) := b"0000000000000000_0000000000000000_0010000011110100_0011100110010111"; -- 0.1287265772441853
	pesos_i(21693) := b"1111111111111111_1111111111111111_1110011101101001_0101101000010001"; -- -0.09604870886615889
	pesos_i(21694) := b"0000000000000000_0000000000000000_0000001101011010_1010010101100010"; -- 0.013101898619535864
	pesos_i(21695) := b"0000000000000000_0000000000000000_0010010110101001_0000000111001101"; -- 0.14711009266714262
	pesos_i(21696) := b"1111111111111111_1111111111111111_1110111110111110_1001111100101110"; -- -0.06349759221523818
	pesos_i(21697) := b"0000000000000000_0000000000000000_0001011111111101_0110010001101001"; -- 0.09371020847705568
	pesos_i(21698) := b"1111111111111111_1111111111111111_1101101010010111_1101000010101100"; -- -0.14612098492887185
	pesos_i(21699) := b"1111111111111111_1111111111111111_1111101110000111_1011100111100011"; -- -0.01746023379641066
	pesos_i(21700) := b"0000000000000000_0000000000000000_0001111000111000_0001001011010001"; -- 0.11804311378178484
	pesos_i(21701) := b"1111111111111111_1111111111111111_1110011101000110_1110111000000101"; -- -0.09657394772708987
	pesos_i(21702) := b"0000000000000000_0000000000000000_0001100100110100_1000101100010011"; -- 0.09845799654505037
	pesos_i(21703) := b"0000000000000000_0000000000000000_0001001011100111_0000100100100101"; -- 0.07383782541146396
	pesos_i(21704) := b"1111111111111111_1111111111111111_1110011101100111_1100110111010000"; -- -0.09607232740460389
	pesos_i(21705) := b"1111111111111111_1111111111111111_1111000101000000_1000110001110001"; -- -0.05760881644395853
	pesos_i(21706) := b"0000000000000000_0000000000000000_0001101101110000_0010100001111000"; -- 0.10718014649609822
	pesos_i(21707) := b"1111111111111111_1111111111111111_1101011100110011_1000101110010110"; -- -0.15936973175990585
	pesos_i(21708) := b"1111111111111111_1111111111111111_1110101111110101_0101000011001010"; -- -0.07828803118198158
	pesos_i(21709) := b"1111111111111111_1111111111111111_1110001110101110_1100101000101100"; -- -0.11061417020462272
	pesos_i(21710) := b"0000000000000000_0000000000000000_0001111111110111_1101011101100001"; -- 0.12487550846273554
	pesos_i(21711) := b"0000000000000000_0000000000000000_0000000000101010_0110011100010100"; -- 0.0006470131691113894
	pesos_i(21712) := b"1111111111111111_1111111111111111_1111101101101001_0110111000111110"; -- -0.01792250617319998
	pesos_i(21713) := b"1111111111111111_1111111111111111_1110010101100010_1100110111101110"; -- -0.10396111440559212
	pesos_i(21714) := b"0000000000000000_0000000000000000_0010001000011000_1101001110010110"; -- 0.13319132247766977
	pesos_i(21715) := b"1111111111111111_1111111111111111_1101110110000111_0110000010011010"; -- -0.13465305559220325
	pesos_i(21716) := b"0000000000000000_0000000000000000_0001011111110000_0000011010001100"; -- 0.0935062495806519
	pesos_i(21717) := b"1111111111111111_1111111111111111_1101111110000001_0101101010010001"; -- -0.12693246807440325
	pesos_i(21718) := b"0000000000000000_0000000000000000_0000101111010000_1111010001110101"; -- 0.04615714886846363
	pesos_i(21719) := b"0000000000000000_0000000000000000_0000011110011011_1100101101110101"; -- 0.02972098919648991
	pesos_i(21720) := b"0000000000000000_0000000000000000_0000100011110001_1101100001000111"; -- 0.034940259327158614
	pesos_i(21721) := b"0000000000000000_0000000000000000_0010010111111011_1100101110000000"; -- 0.14837333564001598
	pesos_i(21722) := b"0000000000000000_0000000000000000_0001100101000000_1000011011011010"; -- 0.09864085026504772
	pesos_i(21723) := b"1111111111111111_1111111111111111_1110100100101001_1000111111110101"; -- -0.08920955906761847
	pesos_i(21724) := b"0000000000000000_0000000000000000_0001000100011101_0111111010110111"; -- 0.06685630765663711
	pesos_i(21725) := b"0000000000000000_0000000000000000_0000111110100000_1100011010111100"; -- 0.06104700173008238
	pesos_i(21726) := b"1111111111111111_1111111111111111_1110011111110000_1110100100100101"; -- -0.09398024403191224
	pesos_i(21727) := b"1111111111111111_1111111111111111_1110001101011100_1011111110000001"; -- -0.11186602681844995
	pesos_i(21728) := b"1111111111111111_1111111111111111_1111101010100100_0011110101101100"; -- -0.02093139746254814
	pesos_i(21729) := b"1111111111111111_1111111111111111_1111000001111000_1001101001010101"; -- -0.06065974649396363
	pesos_i(21730) := b"0000000000000000_0000000000000000_0000011001100011_1011100001001010"; -- 0.02495910452387682
	pesos_i(21731) := b"1111111111111111_1111111111111111_1110001111110101_1011101010101000"; -- -0.10953172116179535
	pesos_i(21732) := b"1111111111111111_1111111111111111_1111110010100011_0010010111011100"; -- -0.013135560878476811
	pesos_i(21733) := b"1111111111111111_1111111111111111_1111111101010111_0011100100010101"; -- -0.0025753330018757348
	pesos_i(21734) := b"1111111111111111_1111111111111111_1110100111110111_1000010001100000"; -- -0.08606693893541953
	pesos_i(21735) := b"1111111111111111_1111111111111111_1110010110111111_1110000111010000"; -- -0.10254086184663026
	pesos_i(21736) := b"1111111111111111_1111111111111111_1111010110010100_1001100011001101"; -- -0.04070134155728791
	pesos_i(21737) := b"1111111111111111_1111111111111111_1110100010111010_1001010101110100"; -- -0.09090295715969325
	pesos_i(21738) := b"1111111111111111_1111111111111111_1111111010010100_0011010101111100"; -- -0.005551011257663171
	pesos_i(21739) := b"1111111111111111_1111111111111111_1111000000001000_0110110011101100"; -- -0.062371437395044964
	pesos_i(21740) := b"1111111111111111_1111111111111111_1110001111000001_1001011000010111"; -- -0.11032735769182543
	pesos_i(21741) := b"1111111111111111_1111111111111111_1110101011100110_1100101100001111"; -- -0.08241587525949064
	pesos_i(21742) := b"0000000000000000_0000000000000000_0000001101011001_1000100100110001"; -- 0.013084959564229158
	pesos_i(21743) := b"0000000000000000_0000000000000000_0010010110011000_0100111010011011"; -- 0.14685527109591404
	pesos_i(21744) := b"1111111111111111_1111111111111111_1111101010001010_0010101011001110"; -- -0.02132923580692484
	pesos_i(21745) := b"1111111111111111_1111111111111111_1110110101110000_0100011101010010"; -- -0.07250551462065638
	pesos_i(21746) := b"0000000000000000_0000000000000000_0001000110101001_0100001001000101"; -- 0.06898893536592499
	pesos_i(21747) := b"1111111111111111_1111111111111111_1111010010101000_1001110001010100"; -- -0.04430220552299568
	pesos_i(21748) := b"1111111111111111_1111111111111111_1110101100101100_0001001110101010"; -- -0.08135869120031576
	pesos_i(21749) := b"0000000000000000_0000000000000000_0010000010011010_1110101011001100"; -- 0.12736384843456708
	pesos_i(21750) := b"1111111111111111_1111111111111111_1110000001110100_0010011010000000"; -- -0.12322768564833621
	pesos_i(21751) := b"1111111111111111_1111111111111111_1110000100110011_0011011110100010"; -- -0.120312235715573
	pesos_i(21752) := b"0000000000000000_0000000000000000_0001010001111001_1010010010100101"; -- 0.07998112714963283
	pesos_i(21753) := b"0000000000000000_0000000000000000_0000110010010100_1001000011100011"; -- 0.04914193666784889
	pesos_i(21754) := b"0000000000000000_0000000000000000_0001011111110000_1010101011111110"; -- 0.09351605121089955
	pesos_i(21755) := b"0000000000000000_0000000000000000_0000011111111000_1111100110010000"; -- 0.031142804694945812
	pesos_i(21756) := b"1111111111111111_1111111111111111_1111000111000110_1111111010010000"; -- -0.055557336643793025
	pesos_i(21757) := b"0000000000000000_0000000000000000_0001011101011101_0111010110100001"; -- 0.09126982855817135
	pesos_i(21758) := b"0000000000000000_0000000000000000_0000010001010101_1011101010100111"; -- 0.016933122395982814
	pesos_i(21759) := b"1111111111111111_1111111111111111_1110011101111101_1010000001011110"; -- -0.09573934270895315
	pesos_i(21760) := b"1111111111111111_1111111111111111_1111000000111010_0000010000100001"; -- -0.061614744173691297
	pesos_i(21761) := b"0000000000000000_0000000000000000_0001011010000100_0110101011101110"; -- 0.08795803357238356
	pesos_i(21762) := b"0000000000000000_0000000000000000_0001001011001100_1101010001111100"; -- 0.07343795797795873
	pesos_i(21763) := b"0000000000000000_0000000000000000_0000110001111111_0011000111101000"; -- 0.04881584091884211
	pesos_i(21764) := b"0000000000000000_0000000000000000_0001000110011101_1101101111110011"; -- 0.06881498976198748
	pesos_i(21765) := b"1111111111111111_1111111111111111_1101101011110100_0001001111101100"; -- -0.14471316805340909
	pesos_i(21766) := b"1111111111111111_1111111111111111_1110010100101011_1001000001101101"; -- -0.10480401350663981
	pesos_i(21767) := b"0000000000000000_0000000000000000_0001000111000001_1011111001011101"; -- 0.06936254289488392
	pesos_i(21768) := b"1111111111111111_1111111111111111_1111111101110101_1101100100101110"; -- -0.0021080268098153353
	pesos_i(21769) := b"0000000000000000_0000000000000000_0000111100010000_0111001100101101"; -- 0.05884475556348969
	pesos_i(21770) := b"0000000000000000_0000000000000000_0001111100000011_1011011100000100"; -- 0.12115043486881778
	pesos_i(21771) := b"0000000000000000_0000000000000000_0000101011011101_1111101001010010"; -- 0.04244961266048944
	pesos_i(21772) := b"0000000000000000_0000000000000000_0001011000001010_1010101000100011"; -- 0.08610022878186903
	pesos_i(21773) := b"0000000000000000_0000000000000000_0000011001111110_0011011101100110"; -- 0.025363409402959405
	pesos_i(21774) := b"0000000000000000_0000000000000000_0001100101101000_1001000101001100"; -- 0.09925182449083603
	pesos_i(21775) := b"0000000000000000_0000000000000000_0010010011010000_1001101111111100"; -- 0.14380812559105585
	pesos_i(21776) := b"1111111111111111_1111111111111111_1110011100111100_0011001010101011"; -- -0.09673770260371047
	pesos_i(21777) := b"0000000000000000_0000000000000000_0000111010011110_1010111101000000"; -- 0.05710883428156887
	pesos_i(21778) := b"0000000000000000_0000000000000000_0010001101110101_1100001100111001"; -- 0.13851566446474736
	pesos_i(21779) := b"0000000000000000_0000000000000000_0001001010100011_1110100001010111"; -- 0.07281353106315178
	pesos_i(21780) := b"0000000000000000_0000000000000000_0000110001111010_1001100100100111"; -- 0.048745700775579874
	pesos_i(21781) := b"1111111111111111_1111111111111111_1110001010011101_0100110011101010"; -- -0.11478728569683425
	pesos_i(21782) := b"0000000000000000_0000000000000000_0000000001110011_1111100100110100"; -- 0.0017696145153766267
	pesos_i(21783) := b"1111111111111111_1111111111111111_1101011101110110_1001010110101101"; -- -0.15834679163438523
	pesos_i(21784) := b"0000000000000000_0000000000000000_0001111001100110_0001101101011110"; -- 0.11874552776137667
	pesos_i(21785) := b"1111111111111111_1111111111111111_1110001011000011_0110011010111111"; -- -0.11420591192828713
	pesos_i(21786) := b"0000000000000000_0000000000000000_0010010010011001_0001001100011101"; -- 0.14296073394883121
	pesos_i(21787) := b"1111111111111111_1111111111111111_1111001001111001_0010111100011111"; -- -0.05283837779318088
	pesos_i(21788) := b"0000000000000000_0000000000000000_0001011010000010_1100100111010010"; -- 0.08793317207227462
	pesos_i(21789) := b"0000000000000000_0000000000000000_0001010001001111_0110001011001101"; -- 0.07933633324784006
	pesos_i(21790) := b"0000000000000000_0000000000000000_0001110000111000_0001101111100111"; -- 0.1102311553580784
	pesos_i(21791) := b"1111111111111111_1111111111111111_1110000010101100_0001111010110011"; -- -0.12237365847902372
	pesos_i(21792) := b"1111111111111111_1111111111111111_1110110101100101_0100000001101100"; -- -0.07267377254008048
	pesos_i(21793) := b"0000000000000000_0000000000000000_0000110100111100_0110011001000100"; -- 0.05170287274600275
	pesos_i(21794) := b"1111111111111111_1111111111111111_1110011001001010_0011100110101011"; -- -0.10042991236183497
	pesos_i(21795) := b"1111111111111111_1111111111111111_1111000111111110_0100100001011010"; -- -0.05471370497565452
	pesos_i(21796) := b"0000000000000000_0000000000000000_0000100110110101_0110101111100101"; -- 0.03792452189868996
	pesos_i(21797) := b"0000000000000000_0000000000000000_0010000101100001_1100001001110110"; -- 0.1303979432920397
	pesos_i(21798) := b"1111111111111111_1111111111111111_1111000111100010_1000101000111000"; -- -0.0551370251397107
	pesos_i(21799) := b"1111111111111111_1111111111111111_1110011111111100_1101101101001111"; -- -0.09379796325246836
	pesos_i(21800) := b"1111111111111111_1111111111111111_1110010001101001_1101110011000101"; -- -0.1077596682477339
	pesos_i(21801) := b"1111111111111111_1111111111111111_1110111110011100_0001000001011111"; -- -0.06402490314976243
	pesos_i(21802) := b"1111111111111111_1111111111111111_1111110110101110_1000010110111000"; -- -0.00905575039350578
	pesos_i(21803) := b"0000000000000000_0000000000000000_0010001010111100_0111110111111011"; -- 0.1356886612767932
	pesos_i(21804) := b"0000000000000000_0000000000000000_0010001010111101_1111100001000011"; -- 0.13571120869732964
	pesos_i(21805) := b"0000000000000000_0000000000000000_0000101010011001_0001000101011110"; -- 0.04139812988382026
	pesos_i(21806) := b"0000000000000000_0000000000000000_0001100100110110_1011111010110000"; -- 0.09849159037086722
	pesos_i(21807) := b"1111111111111111_1111111111111111_1110101010001011_1000101000110101"; -- -0.08380829065432344
	pesos_i(21808) := b"1111111111111111_1111111111111111_1111101001111011_1011101000100001"; -- -0.021549574817774877
	pesos_i(21809) := b"1111111111111111_1111111111111111_1110100111001001_0011010100110000"; -- -0.08677356326479184
	pesos_i(21810) := b"1111111111111111_1111111111111111_1111111000000010_1111011010010111"; -- -0.007767284416397786
	pesos_i(21811) := b"1111111111111111_1111111111111111_1111110010001100_1111000110010000"; -- -0.013474371286543042
	pesos_i(21812) := b"0000000000000000_0000000000000000_0001000101101011_0110100101101110"; -- 0.06804522454245596
	pesos_i(21813) := b"0000000000000000_0000000000000000_0001100001111111_0000101010001000"; -- 0.09568849400450657
	pesos_i(21814) := b"0000000000000000_0000000000000000_0010000001000011_1101111001100011"; -- 0.1260355941880593
	pesos_i(21815) := b"1111111111111111_1111111111111111_1110111011001000_1001000111000110"; -- -0.06725205331772176
	pesos_i(21816) := b"0000000000000000_0000000000000000_0001010110100110_0100001010011100"; -- 0.0845681792184926
	pesos_i(21817) := b"1111111111111111_1111111111111111_1111011110110011_1100010101110001"; -- -0.03241315838341137
	pesos_i(21818) := b"1111111111111111_1111111111111111_1111000001110101_1011001101010100"; -- -0.06070403279797198
	pesos_i(21819) := b"1111111111111111_1111111111111111_1101101101100011_0101010110111100"; -- -0.1430155197994953
	pesos_i(21820) := b"1111111111111111_1111111111111111_1110010000100100_0100010000110011"; -- -0.10882161870717619
	pesos_i(21821) := b"1111111111111111_1111111111111111_1110110100111000_0100001001000101"; -- -0.07336030776033746
	pesos_i(21822) := b"1111111111111111_1111111111111111_1111011010000100_1111110001001000"; -- -0.03703330264761354
	pesos_i(21823) := b"0000000000000000_0000000000000000_0001111110011010_0100010001001010"; -- 0.12344767380058483
	pesos_i(21824) := b"0000000000000000_0000000000000000_0000100111101100_0100111111110001"; -- 0.03876208907042596
	pesos_i(21825) := b"0000000000000000_0000000000000000_0000101001100010_0111110000100000"; -- 0.04056525980552151
	pesos_i(21826) := b"1111111111111111_1111111111111111_1101111000011100_1010100101110111"; -- -0.13237515304796413
	pesos_i(21827) := b"1111111111111111_1111111111111111_1110111001101000_1111011110001100"; -- -0.068710830947657
	pesos_i(21828) := b"0000000000000000_0000000000000000_0000110010100100_0100100001010011"; -- 0.04938175232241887
	pesos_i(21829) := b"1111111111111111_1111111111111111_1111101010110010_0000111100001111"; -- -0.02072053788083013
	pesos_i(21830) := b"1111111111111111_1111111111111111_1110001111111111_1110101011000001"; -- -0.10937626636954853
	pesos_i(21831) := b"0000000000000000_0000000000000000_0000101110000001_1111100000000111"; -- 0.044951917389154515
	pesos_i(21832) := b"0000000000000000_0000000000000000_0001100011111010_1111001011101001"; -- 0.09757917593446468
	pesos_i(21833) := b"0000000000000000_0000000000000000_0001011010001011_0111110000101000"; -- 0.08806587194102822
	pesos_i(21834) := b"1111111111111111_1111111111111111_1110010111100110_1001011001011111"; -- -0.1019502657813782
	pesos_i(21835) := b"1111111111111111_1111111111111111_1101110100011101_0111110111110010"; -- -0.13626873812762538
	pesos_i(21836) := b"0000000000000000_0000000000000000_0001100110111100_1100001101110111"; -- 0.10053655298597927
	pesos_i(21837) := b"1111111111111111_1111111111111111_1111111100111000_1110001100100001"; -- -0.003038219866634337
	pesos_i(21838) := b"1111111111111111_1111111111111111_1110011100010010_1000011110011101"; -- -0.09737350873013478
	pesos_i(21839) := b"1111111111111111_1111111111111111_1111111011001100_0101101100011011"; -- -0.00469427674969822
	pesos_i(21840) := b"1111111111111111_1111111111111111_1111000000001110_0100010110001001"; -- -0.06228223238446458
	pesos_i(21841) := b"1111111111111111_1111111111111111_1110010100010011_1010110010000100"; -- -0.10516855027547804
	pesos_i(21842) := b"0000000000000000_0000000000000000_0000101000100100_1001011100100010"; -- 0.039620824739509654
	pesos_i(21843) := b"1111111111111111_1111111111111111_1101111110000110_1001101010001011"; -- -0.1268523608799359
	pesos_i(21844) := b"1111111111111111_1111111111111111_1101111000011011_0010110101101100"; -- -0.1323978053035814
	pesos_i(21845) := b"0000000000000000_0000000000000000_0010000111011110_0000001000100001"; -- 0.13229382805359688
	pesos_i(21846) := b"0000000000000000_0000000000000000_0001111100110001_1000101101111011"; -- 0.12184974441740641
	pesos_i(21847) := b"0000000000000000_0000000000000000_0001111111001100_1001101011111111"; -- 0.12421578143093906
	pesos_i(21848) := b"1111111111111111_1111111111111111_1101101110010001_0110001100011110"; -- -0.14231281785450697
	pesos_i(21849) := b"1111111111111111_1111111111111111_1101100010001000_0101100100011111"; -- -0.15416949254101195
	pesos_i(21850) := b"0000000000000000_0000000000000000_0010000100001101_1110000100101010"; -- 0.129118034970898
	pesos_i(21851) := b"1111111111111111_1111111111111111_1101011101100010_0101100110001101"; -- -0.15865555096627415
	pesos_i(21852) := b"0000000000000000_0000000000000000_0001001010000101_0011111100111001"; -- 0.07234568734441474
	pesos_i(21853) := b"0000000000000000_0000000000000000_0000000001101000_0001100011010100"; -- 0.0015883938621782628
	pesos_i(21854) := b"0000000000000000_0000000000000000_0000000001011111_1100101100011011"; -- 0.0014616910330470037
	pesos_i(21855) := b"1111111111111111_1111111111111111_1111010101010010_0100000010010000"; -- -0.04171368110143334
	pesos_i(21856) := b"0000000000000000_0000000000000000_0001111101110101_0000000100000110"; -- 0.12287908937240004
	pesos_i(21857) := b"1111111111111111_1111111111111111_1110100111101110_1110111100000101"; -- -0.08619791142555673
	pesos_i(21858) := b"1111111111111111_1111111111111111_1101111101101111_1000011110010001"; -- -0.1272044439202167
	pesos_i(21859) := b"0000000000000000_0000000000000000_0001011101101000_0001011101011010"; -- 0.09143205588660126
	pesos_i(21860) := b"0000000000000000_0000000000000000_0000011101001101_0100111100001001"; -- 0.028523387677546135
	pesos_i(21861) := b"1111111111111111_1111111111111111_1111000011001111_1101100101000100"; -- -0.05932848070487267
	pesos_i(21862) := b"1111111111111111_1111111111111111_1111011111000101_0101000010001110"; -- -0.0321454672185149
	pesos_i(21863) := b"1111111111111111_1111111111111111_1110110100011101_0000111110101010"; -- -0.07377531156975939
	pesos_i(21864) := b"0000000000000000_0000000000000000_0001010100000110_0001011101010111"; -- 0.08212419391427776
	pesos_i(21865) := b"1111111111111111_1111111111111111_1111100011110010_0001111100010110"; -- -0.02755552011081146
	pesos_i(21866) := b"1111111111111111_1111111111111111_1111111111110001_1000101110100011"; -- -0.00022055878619588545
	pesos_i(21867) := b"1111111111111111_1111111111111111_1110011011100011_1101100100111001"; -- -0.09808580750649495
	pesos_i(21868) := b"0000000000000000_0000000000000000_0000101111110110_0000111101111011"; -- 0.046723334861164416
	pesos_i(21869) := b"0000000000000000_0000000000000000_0001001100101100_1010111001101000"; -- 0.07490053218630661
	pesos_i(21870) := b"0000000000000000_0000000000000000_0001000011101000_0000110001111001"; -- 0.06604078248376725
	pesos_i(21871) := b"0000000000000000_0000000000000000_0001111001010100_1000111011010101"; -- 0.11847775171974906
	pesos_i(21872) := b"0000000000000000_0000000000000000_0000001010111101_1000001101001010"; -- 0.010704236516857969
	pesos_i(21873) := b"0000000000000000_0000000000000000_0010010110110101_0101010100111100"; -- 0.14729817115943514
	pesos_i(21874) := b"1111111111111111_1111111111111111_1111110011001010_1001111001111110"; -- -0.01253327779997515
	pesos_i(21875) := b"1111111111111111_1111111111111111_1101101111000010_0010010100001011"; -- -0.14156883705047282
	pesos_i(21876) := b"1111111111111111_1111111111111111_1111000111110111_1111010100001010"; -- -0.05481022373562083
	pesos_i(21877) := b"1111111111111111_1111111111111111_1111010001001000_1011011100011011"; -- -0.04576545325621064
	pesos_i(21878) := b"1111111111111111_1111111111111111_1110101010110001_1011111111010001"; -- -0.08322526113292873
	pesos_i(21879) := b"0000000000000000_0000000000000000_0000101111001011_1011001000010011"; -- 0.04607689814840081
	pesos_i(21880) := b"1111111111111111_1111111111111111_1110010100010100_0011110001001110"; -- -0.10515997975053187
	pesos_i(21881) := b"0000000000000000_0000000000000000_0000011101011011_0001111011001100"; -- 0.028734135355656137
	pesos_i(21882) := b"0000000000000000_0000000000000000_0010010111110110_0010101000110101"; -- 0.1482874277662642
	pesos_i(21883) := b"0000000000000000_0000000000000000_0000001111101110_0010010000011101"; -- 0.015352494359019288
	pesos_i(21884) := b"0000000000000000_0000000000000000_0001111011110000_1010110000100101"; -- 0.12085987008748283
	pesos_i(21885) := b"0000000000000000_0000000000000000_0001101000111000_1001100010000011"; -- 0.10242608262940137
	pesos_i(21886) := b"1111111111111111_1111111111111111_1101101000001010_0101001100101110"; -- -0.14827995430277932
	pesos_i(21887) := b"1111111111111111_1111111111111111_1111101000111100_1010110101001001"; -- -0.022511643985795568
	pesos_i(21888) := b"0000000000000000_0000000000000000_0001001001110000_1001001010110010"; -- 0.07203022800358296
	pesos_i(21889) := b"1111111111111111_1111111111111111_1110111011100100_0010001110001101"; -- -0.06683137721742442
	pesos_i(21890) := b"0000000000000000_0000000000000000_0001110110000011_1010010010011011"; -- 0.11528996265019135
	pesos_i(21891) := b"0000000000000000_0000000000000000_0000101010011101_0001001000010011"; -- 0.04145920713123906
	pesos_i(21892) := b"0000000000000000_0000000000000000_0000111100100101_1011111100111100"; -- 0.059169723747790774
	pesos_i(21893) := b"1111111111111111_1111111111111111_1101101010000010_1100111000011000"; -- -0.14644157327357055
	pesos_i(21894) := b"1111111111111111_1111111111111111_1110000010100110_1111110111111010"; -- -0.12245190290823421
	pesos_i(21895) := b"1111111111111111_1111111111111111_1111100011111001_0111110010111101"; -- -0.027443126655718644
	pesos_i(21896) := b"1111111111111111_1111111111111111_1110000101101011_1111001000010110"; -- -0.11944663004735069
	pesos_i(21897) := b"0000000000000000_0000000000000000_0000101000011111_0110100110101001"; -- 0.039541820343344594
	pesos_i(21898) := b"1111111111111111_1111111111111111_1111111111001111_0011000001000001"; -- -0.0007448045110379174
	pesos_i(21899) := b"1111111111111111_1111111111111111_1111110010100110_1000100100101010"; -- -0.013083865509883916
	pesos_i(21900) := b"0000000000000000_0000000000000000_0001101001110011_0111010110100000"; -- 0.1033242718244394
	pesos_i(21901) := b"1111111111111111_1111111111111111_1110111101111101_1101010111010011"; -- -0.06448615633610356
	pesos_i(21902) := b"0000000000000000_0000000000000000_0001010100101111_1011110001111111"; -- 0.08275964829393091
	pesos_i(21903) := b"0000000000000000_0000000000000000_0010010011110101_0111101001001111"; -- 0.14437069341556047
	pesos_i(21904) := b"0000000000000000_0000000000000000_0001110011110010_0101110000100001"; -- 0.11307311836523175
	pesos_i(21905) := b"1111111111111111_1111111111111111_1110010100011110_0100100101111101"; -- -0.10500660619703543
	pesos_i(21906) := b"0000000000000000_0000000000000000_0000011000111100_0010000110011111"; -- 0.024355031301672242
	pesos_i(21907) := b"0000000000000000_0000000000000000_0000000111010000_0111001111110111"; -- 0.007086990054587898
	pesos_i(21908) := b"0000000000000000_0000000000000000_0010000000011001_1011001010011101"; -- 0.12539211602184186
	pesos_i(21909) := b"1111111111111111_1111111111111111_1110010001100110_0010100011101100"; -- -0.10781616433748105
	pesos_i(21910) := b"0000000000000000_0000000000000000_0001001101000001_1010000001011110"; -- 0.07522012999609735
	pesos_i(21911) := b"0000000000000000_0000000000000000_0001001011101110_1000011001001110"; -- 0.0739520970643413
	pesos_i(21912) := b"1111111111111111_1111111111111111_1110010011111011_1010101101111111"; -- -0.1055348219751541
	pesos_i(21913) := b"0000000000000000_0000000000000000_0000000011011101_0000111010001001"; -- 0.0033730586451017133
	pesos_i(21914) := b"0000000000000000_0000000000000000_0010000000111010_0010010011001100"; -- 0.1258872029261216
	pesos_i(21915) := b"0000000000000000_0000000000000000_0001101111010000_1010110011010011"; -- 0.1086528792766909
	pesos_i(21916) := b"0000000000000000_0000000000000000_0001000101101110_0001011111011001"; -- 0.06808613833212804
	pesos_i(21917) := b"1111111111111111_1111111111111111_1110111111000000_1110111101111011"; -- -0.06346228839705731
	pesos_i(21918) := b"0000000000000000_0000000000000000_0001100010010000_0110000011101111"; -- 0.09595304328168666
	pesos_i(21919) := b"0000000000000000_0000000000000000_0001111110101111_1000000011000100"; -- 0.12377171322547975
	pesos_i(21920) := b"1111111111111111_1111111111111111_1110100001111101_1111000100100100"; -- -0.09182827817851143
	pesos_i(21921) := b"1111111111111111_1111111111111111_1111011000101110_1000010110001000"; -- -0.03835263672261399
	pesos_i(21922) := b"1111111111111111_1111111111111111_1111110011000110_0100100011111011"; -- -0.012599409887510534
	pesos_i(21923) := b"1111111111111111_1111111111111111_1111001100001010_1100011011111110"; -- -0.05061680122320975
	pesos_i(21924) := b"0000000000000000_0000000000000000_0001100011110110_0011010100100100"; -- 0.09750682942650464
	pesos_i(21925) := b"0000000000000000_0000000000000000_0000001101111011_0011110000101001"; -- 0.013599166898603184
	pesos_i(21926) := b"1111111111111111_1111111111111111_1111110110011011_1111101000001110"; -- -0.00933873333284917
	pesos_i(21927) := b"0000000000000000_0000000000000000_0001011111101011_1100100000100000"; -- 0.09344149376178203
	pesos_i(21928) := b"1111111111111111_1111111111111111_1111110111011010_0001000011011101"; -- -0.00839132896638834
	pesos_i(21929) := b"1111111111111111_1111111111111111_1111010010111111_0001100010000110"; -- -0.043959109646618484
	pesos_i(21930) := b"0000000000000000_0000000000000000_0010011001000011_1010000111111000"; -- 0.14946949293415696
	pesos_i(21931) := b"0000000000000000_0000000000000000_0000101111111011_1110011111101010"; -- 0.046812529113930954
	pesos_i(21932) := b"1111111111111111_1111111111111111_1111100111111010_1100001100001000"; -- -0.023517428051059542
	pesos_i(21933) := b"0000000000000000_0000000000000000_0001110101010111_0001101011100011"; -- 0.11461036712959945
	pesos_i(21934) := b"1111111111111111_1111111111111111_1101110001011011_1110000111111101"; -- -0.13922298026344568
	pesos_i(21935) := b"0000000000000000_0000000000000000_0010010010100100_0010001000100001"; -- 0.1431294757059439
	pesos_i(21936) := b"1111111111111111_1111111111111111_1110011110000011_0100001000100100"; -- -0.09565340626086494
	pesos_i(21937) := b"1111111111111111_1111111111111111_1111010010001001_0001000100001011"; -- -0.044783530026901844
	pesos_i(21938) := b"0000000000000000_0000000000000000_0000000001100111_0101100101000000"; -- 0.0015769749373811294
	pesos_i(21939) := b"0000000000000000_0000000000000000_0010000010001101_1000110101011010"; -- 0.12715991455792014
	pesos_i(21940) := b"0000000000000000_0000000000000000_0001100001011000_1001000111110010"; -- 0.09510147240847344
	pesos_i(21941) := b"0000000000000000_0000000000000000_0001111100011100_0000110110101011"; -- 0.12152181088373079
	pesos_i(21942) := b"1111111111111111_1111111111111111_1101110010001011_0100101101100001"; -- -0.13849953538061843
	pesos_i(21943) := b"1111111111111111_1111111111111111_1111101110000010_0100001111110010"; -- -0.017543557579031206
	pesos_i(21944) := b"1111111111111111_1111111111111111_1111000110011101_1010000110001011"; -- -0.056188491511756276
	pesos_i(21945) := b"0000000000000000_0000000000000000_0001100100000001_0101101111100101"; -- 0.09767698617745366
	pesos_i(21946) := b"1111111111111111_1111111111111111_1101110000011010_0110101001110011"; -- -0.14022192670295708
	pesos_i(21947) := b"1111111111111111_1111111111111111_1110110000001100_1000100100101110"; -- -0.07793371809681797
	pesos_i(21948) := b"0000000000000000_0000000000000000_0000011110011001_1110111001110000"; -- 0.0296925566009647
	pesos_i(21949) := b"1111111111111111_1111111111111111_1110110101000010_0000001101111101"; -- -0.07321146203435541
	pesos_i(21950) := b"0000000000000000_0000000000000000_0001110000000110_1000001000011110"; -- 0.10947430841639298
	pesos_i(21951) := b"0000000000000000_0000000000000000_0000000110000000_1101011100011111"; -- 0.005872197162662219
	pesos_i(21952) := b"0000000000000000_0000000000000000_0001011101111001_1101100000111111"; -- 0.09170295280418096
	pesos_i(21953) := b"1111111111111111_1111111111111111_1110010011110110_1010111010000011"; -- -0.10561093629153316
	pesos_i(21954) := b"1111111111111111_1111111111111111_1111100000000101_0010001010101100"; -- -0.031171639559504503
	pesos_i(21955) := b"0000000000000000_0000000000000000_0001110111001110_0110001000110111"; -- 0.11643041468700417
	pesos_i(21956) := b"1111111111111111_1111111111111111_1111100000111001_1000111111011100"; -- -0.030371674237871567
	pesos_i(21957) := b"1111111111111111_1111111111111111_1110100000101110_0110100101100100"; -- -0.09304181391577067
	pesos_i(21958) := b"0000000000000000_0000000000000000_0000100011000010_0010110101000111"; -- 0.034212903880120146
	pesos_i(21959) := b"0000000000000000_0000000000000000_0000111110100100_1000001011000110"; -- 0.06110398619383606
	pesos_i(21960) := b"1111111111111111_1111111111111111_1111001100011011_0000111101010111"; -- -0.05036834826038599
	pesos_i(21961) := b"1111111111111111_1111111111111111_1101101111100000_1011010110100001"; -- -0.1411024553194967
	pesos_i(21962) := b"0000000000000000_0000000000000000_0000110010100010_0100110110101100"; -- 0.04935155350232456
	pesos_i(21963) := b"0000000000000000_0000000000000000_0000011011010111_0110111001001110"; -- 0.026724714338804186
	pesos_i(21964) := b"1111111111111111_1111111111111111_1111111100101101_0110000111111010"; -- -0.003213764573207759
	pesos_i(21965) := b"0000000000000000_0000000000000000_0000100001111101_1011010011111100"; -- 0.03316813615760409
	pesos_i(21966) := b"1111111111111111_1111111111111111_1111010100111001_1001101100000101"; -- -0.042089759067297595
	pesos_i(21967) := b"1111111111111111_1111111111111111_1110000110100011_1001101101001101"; -- -0.11859731083840404
	pesos_i(21968) := b"0000000000000000_0000000000000000_0010000010101000_1010011001011101"; -- 0.12757339260780742
	pesos_i(21969) := b"0000000000000000_0000000000000000_0000010010000111_0001000100111001"; -- 0.01768596303582918
	pesos_i(21970) := b"1111111111111111_1111111111111111_1111000011101010_0011110100101010"; -- -0.058925797756196774
	pesos_i(21971) := b"1111111111111111_1111111111111111_1110010111000101_1010011100100111"; -- -0.10245280560907943
	pesos_i(21972) := b"0000000000000000_0000000000000000_0010010101101100_0101010011010101"; -- 0.14618425562037274
	pesos_i(21973) := b"1111111111111111_1111111111111111_1110101001111100_0000000011000010"; -- -0.08404536508073085
	pesos_i(21974) := b"0000000000000000_0000000000000000_0010010000001011_0001010100111001"; -- 0.1407941115354686
	pesos_i(21975) := b"1111111111111111_1111111111111111_1111100001000001_1111110111110000"; -- -0.030243042927582998
	pesos_i(21976) := b"0000000000000000_0000000000000000_0000101001111011_0101010110001100"; -- 0.040944430115084834
	pesos_i(21977) := b"1111111111111111_1111111111111111_1110101011111000_0101000011011011"; -- -0.08214850083621311
	pesos_i(21978) := b"1111111111111111_1111111111111111_1101111010101001_0010001111111000"; -- -0.130231620833787
	pesos_i(21979) := b"0000000000000000_0000000000000000_0000110111000001_1111110111010011"; -- 0.05374132539384674
	pesos_i(21980) := b"1111111111111111_1111111111111111_1111010111010011_0010010010010110"; -- -0.03974696486392151
	pesos_i(21981) := b"1111111111111111_1111111111111111_1111010010011001_1110100101011100"; -- -0.044526496084939214
	pesos_i(21982) := b"1111111111111111_1111111111111111_1111011011000100_1010011010110100"; -- -0.03606184111042753
	pesos_i(21983) := b"0000000000000000_0000000000000000_0000111000010110_1000110000100000"; -- 0.05503154546262036
	pesos_i(21984) := b"1111111111111111_1111111111111111_1111010110000010_0000100111101000"; -- -0.04098451700250449
	pesos_i(21985) := b"1111111111111111_1111111111111111_1101101101001000_0111111100111111"; -- -0.1434250326303867
	pesos_i(21986) := b"1111111111111111_1111111111111111_1110000001001110_0100000010101111"; -- -0.12380595904407242
	pesos_i(21987) := b"1111111111111111_1111111111111111_1110101010100111_1011111111001110"; -- -0.08337784972372124
	pesos_i(21988) := b"0000000000000000_0000000000000000_0001011000001010_0100100010010101"; -- 0.08609441416714052
	pesos_i(21989) := b"0000000000000000_0000000000000000_0001011110111001_0101000110001100"; -- 0.09267148661515885
	pesos_i(21990) := b"0000000000000000_0000000000000000_0001000110110100_1111111011010011"; -- 0.06916802079962146
	pesos_i(21991) := b"1111111111111111_1111111111111111_1110000000101010_1110010101000110"; -- -0.12434546510322335
	pesos_i(21992) := b"0000000000000000_0000000000000000_0000010101011011_0011000111000101"; -- 0.020922766229975836
	pesos_i(21993) := b"0000000000000000_0000000000000000_0001001111110100_0101100100100110"; -- 0.0779472081821135
	pesos_i(21994) := b"0000000000000000_0000000000000000_0001001011000000_1010010001000001"; -- 0.07325197779006784
	pesos_i(21995) := b"0000000000000000_0000000000000000_0010010010001011_0001111110110100"; -- 0.14274786139239642
	pesos_i(21996) := b"0000000000000000_0000000000000000_0000001101001010_1011100110110010"; -- 0.012858968596719778
	pesos_i(21997) := b"0000000000000000_0000000000000000_0000010111010011_0110100110101001"; -- 0.02275715228522374
	pesos_i(21998) := b"1111111111111111_1111111111111111_1111000110100001_1101010011010001"; -- -0.056124400200913874
	pesos_i(21999) := b"1111111111111111_1111111111111111_1110011111100110_0110000110101001"; -- -0.0941409076215092
	pesos_i(22000) := b"0000000000000000_0000000000000000_0000011000001011_0011100001000101"; -- 0.02360870056565765
	pesos_i(22001) := b"0000000000000000_0000000000000000_0000111011100111_0100111001100111"; -- 0.058216953503923585
	pesos_i(22002) := b"0000000000000000_0000000000000000_0001000110110010_1111110011111111"; -- 0.06913739426893316
	pesos_i(22003) := b"1111111111111111_1111111111111111_1111001100110010_0101100001001010"; -- -0.050013048149726354
	pesos_i(22004) := b"0000000000000000_0000000000000000_0001110100100001_0111111101011001"; -- 0.11379238066456318
	pesos_i(22005) := b"1111111111111111_1111111111111111_1101101011110000_0101001100000100"; -- -0.14477044240654832
	pesos_i(22006) := b"1111111111111111_1111111111111111_1111111000000010_1011000000000000"; -- -0.007771491938573726
	pesos_i(22007) := b"1111111111111111_1111111111111111_1111010111010000_1101000100111010"; -- -0.03978245095631421
	pesos_i(22008) := b"1111111111111111_1111111111111111_1111101110010111_1010101110100100"; -- -0.017216942225582378
	pesos_i(22009) := b"1111111111111111_1111111111111111_1110010100010101_1111100110101101"; -- -0.10513343352966875
	pesos_i(22010) := b"0000000000000000_0000000000000000_0001011111110011_0011001111010011"; -- 0.09355472470578269
	pesos_i(22011) := b"1111111111111111_1111111111111111_1101110110000100_1100001100111110"; -- -0.13469295238830897
	pesos_i(22012) := b"0000000000000000_0000000000000000_0001101110010100_1100001010000101"; -- 0.10773864512698579
	pesos_i(22013) := b"1111111111111111_1111111111111111_1110100011010101_1110010111010000"; -- -0.0904861800244759
	pesos_i(22014) := b"1111111111111111_1111111111111111_1111110001111001_1111011010000011"; -- -0.013763993181585185
	pesos_i(22015) := b"0000000000000000_0000000000000000_0000111110100100_0011111000000111"; -- 0.06109988861581603
	pesos_i(22016) := b"1111111111111111_1111111111111111_1110001110110100_0010101101000111"; -- -0.11053208847846234
	pesos_i(22017) := b"1111111111111111_1111111111111111_1110011101110100_0100101011000110"; -- -0.09588177363992272
	pesos_i(22018) := b"1111111111111111_1111111111111111_1111010111011001_0011001110011001"; -- -0.03965451720445163
	pesos_i(22019) := b"0000000000000000_0000000000000000_0000001101000100_1011100111111010"; -- 0.012767432750921914
	pesos_i(22020) := b"1111111111111111_1111111111111111_1110111010101100_0010001110010100"; -- -0.0676858676315456
	pesos_i(22021) := b"0000000000000000_0000000000000000_0001000100101110_1010111111111000"; -- 0.06711864294554216
	pesos_i(22022) := b"1111111111111111_1111111111111111_1101101110100101_1101001010111000"; -- -0.14200098990278048
	pesos_i(22023) := b"1111111111111111_1111111111111111_1110001110011000_0100001110001100"; -- -0.11095788800428352
	pesos_i(22024) := b"0000000000000000_0000000000000000_0001011101000001_0011100100100010"; -- 0.09083897672040624
	pesos_i(22025) := b"0000000000000000_0000000000000000_0001001111111110_1100111000100101"; -- 0.07810676958967981
	pesos_i(22026) := b"1111111111111111_1111111111111111_1111011010011001_0100110000010000"; -- -0.03672337159828949
	pesos_i(22027) := b"0000000000000000_0000000000000000_0001111100111011_1001110100101111"; -- 0.12200338731724686
	pesos_i(22028) := b"0000000000000000_0000000000000000_0000011101110001_0000101010101100"; -- 0.02906862923397253
	pesos_i(22029) := b"1111111111111111_1111111111111111_1111110110100111_0001100111000111"; -- -0.009168995789722176
	pesos_i(22030) := b"1111111111111111_1111111111111111_1111000110011010_1001000001110000"; -- -0.05623528728554696
	pesos_i(22031) := b"1111111111111111_1111111111111111_1111001101100111_1100011101101011"; -- -0.049197708593289834
	pesos_i(22032) := b"0000000000000000_0000000000000000_0001001011001000_0100000010101101"; -- 0.07336811267876091
	pesos_i(22033) := b"1111111111111111_1111111111111111_1111010100100001_0100011011100110"; -- -0.0424609841537302
	pesos_i(22034) := b"0000000000000000_0000000000000000_0001110000101100_0001100001111001"; -- 0.11004784545597633
	pesos_i(22035) := b"0000000000000000_0000000000000000_0001011101000000_1010000000010010"; -- 0.09082985354120424
	pesos_i(22036) := b"1111111111111111_1111111111111111_1111010100000101_1010100011000100"; -- -0.04288239673296112
	pesos_i(22037) := b"1111111111111111_1111111111111111_1111110110101111_1101010001111111"; -- -0.00903579626358104
	pesos_i(22038) := b"1111111111111111_1111111111111111_1110011010110010_1110000011001110"; -- -0.09883303606523905
	pesos_i(22039) := b"1111111111111111_1111111111111111_1110110000001010_1010000000110000"; -- -0.07796286421506884
	pesos_i(22040) := b"0000000000000000_0000000000000000_0001001111010011_0001100111010111"; -- 0.07743989468560611
	pesos_i(22041) := b"0000000000000000_0000000000000000_0001111111011000_1011001111001110"; -- 0.12440036564834403
	pesos_i(22042) := b"1111111111111111_1111111111111111_1110100010111001_0111100100011100"; -- -0.09091990544321553
	pesos_i(22043) := b"0000000000000000_0000000000000000_0000111101011110_0100001100101111"; -- 0.06003208052773564
	pesos_i(22044) := b"0000000000000000_0000000000000000_0001011101001100_1001010010110100"; -- 0.091012281270739
	pesos_i(22045) := b"1111111111111111_1111111111111111_1111000111011011_1111110001011100"; -- -0.05523703343095682
	pesos_i(22046) := b"1111111111111111_1111111111111111_1101101110000010_0010110010101010"; -- -0.14254494514757712
	pesos_i(22047) := b"1111111111111111_1111111111111111_1110110001101110_0101101100000000"; -- -0.0764411092097278
	pesos_i(22048) := b"0000000000000000_0000000000000000_0010011010101110_0000001010001001"; -- 0.15109268042045626
	pesos_i(22049) := b"0000000000000000_0000000000000000_0001010101001100_1011001011101001"; -- 0.08320158175315119
	pesos_i(22050) := b"1111111111111111_1111111111111111_1110000010000111_1011011000101100"; -- -0.12292920515742123
	pesos_i(22051) := b"1111111111111111_1111111111111111_1111111011001000_0010010011010010"; -- -0.0047585475785533885
	pesos_i(22052) := b"0000000000000000_0000000000000000_0001010010100100_0110011010100110"; -- 0.08063355966244436
	pesos_i(22053) := b"1111111111111111_1111111111111111_1110000101100100_0001011111101110"; -- -0.11956644480084097
	pesos_i(22054) := b"0000000000000000_0000000000000000_0001010010111100_0111001101110000"; -- 0.08100053287350681
	pesos_i(22055) := b"1111111111111111_1111111111111111_1101100110010001_0111000110000100"; -- -0.15012445958341603
	pesos_i(22056) := b"0000000000000000_0000000000000000_0001101001000001_1100110000011101"; -- 0.10256648749320169
	pesos_i(22057) := b"0000000000000000_0000000000000000_0010000101010111_0101111101001011"; -- 0.13023944443763036
	pesos_i(22058) := b"0000000000000000_0000000000000000_0001001011111011_1010010001011010"; -- 0.07415225205510954
	pesos_i(22059) := b"1111111111111111_1111111111111111_1111001100010010_1101110001011100"; -- -0.05049345729895002
	pesos_i(22060) := b"1111111111111111_1111111111111111_1110110111101010_1111101000111101"; -- -0.07063327805727522
	pesos_i(22061) := b"1111111111111111_1111111111111111_1111110100011011_1110100011111110"; -- -0.011292875252788399
	pesos_i(22062) := b"0000000000000000_0000000000000000_0001011011100001_1010010000010111"; -- 0.08938050809382708
	pesos_i(22063) := b"1111111111111111_1111111111111111_1111000111010001_0111001011001001"; -- -0.05539782130391603
	pesos_i(22064) := b"0000000000000000_0000000000000000_0000011111100000_0011011010110001"; -- 0.030764978710071895
	pesos_i(22065) := b"1111111111111111_1111111111111111_1111111111011000_1011011111011000"; -- -0.0005993935809641359
	pesos_i(22066) := b"0000000000000000_0000000000000000_0001100011001011_1010001101010101"; -- 0.09685726945060677
	pesos_i(22067) := b"1111111111111111_1111111111111111_1110000111000011_0101110111110111"; -- -0.1181126854635645
	pesos_i(22068) := b"0000000000000000_0000000000000000_0001100000100111_0100011101101111"; -- 0.09434935054769236
	pesos_i(22069) := b"1111111111111111_1111111111111111_1110010101010000_1111111011111001"; -- -0.10423284939003273
	pesos_i(22070) := b"1111111111111111_1111111111111111_1111110110000111_0101111001011101"; -- -0.00965318905082264
	pesos_i(22071) := b"0000000000000000_0000000000000000_0010010100110100_1010111000110101"; -- 0.14533509056110702
	pesos_i(22072) := b"1111111111111111_1111111111111111_1110101110110101_1010111111001001"; -- -0.07925893150330157
	pesos_i(22073) := b"1111111111111111_1111111111111111_1101101101100110_0001111110000011"; -- -0.14297297529428069
	pesos_i(22074) := b"1111111111111111_1111111111111111_1110111001000101_1011110001001101"; -- -0.0692484199670458
	pesos_i(22075) := b"1111111111111111_1111111111111111_1111110110110110_0010111110010011"; -- -0.008938814773403185
	pesos_i(22076) := b"1111111111111111_1111111111111111_1110011001011101_0100001100001001"; -- -0.10013943697249526
	pesos_i(22077) := b"1111111111111111_1111111111111111_1111110111001011_0100101010111000"; -- -0.008616762192292468
	pesos_i(22078) := b"0000000000000000_0000000000000000_0000101111000110_1111011101111100"; -- 0.04600474154005876
	pesos_i(22079) := b"0000000000000000_0000000000000000_0000010011100111_1000010000011110"; -- 0.01915765497628587
	pesos_i(22080) := b"0000000000000000_0000000000000000_0000101001011110_1011111110111100"; -- 0.04050825444647543
	pesos_i(22081) := b"1111111111111111_1111111111111111_1110111110100010_0110010100100010"; -- -0.06392829809077534
	pesos_i(22082) := b"0000000000000000_0000000000000000_0001011110111111_1111110011001000"; -- 0.09277324560056305
	pesos_i(22083) := b"0000000000000000_0000000000000000_0000101110100101_0111000111111001"; -- 0.04549324349683178
	pesos_i(22084) := b"1111111111111111_1111111111111111_1111011001001011_0000010010110101"; -- -0.037917810180925236
	pesos_i(22085) := b"1111111111111111_1111111111111111_1101101111100111_0100010011110110"; -- -0.1410023593965742
	pesos_i(22086) := b"0000000000000000_0000000000000000_0001001011110100_1001101101001010"; -- 0.07404490043787901
	pesos_i(22087) := b"0000000000000000_0000000000000000_0001100010111010_0110100001111011"; -- 0.09659436232232137
	pesos_i(22088) := b"1111111111111111_1111111111111111_1110011111010111_0011101000011100"; -- -0.09437214672399628
	pesos_i(22089) := b"1111111111111111_1111111111111111_1110001001110100_1100011000000010"; -- -0.1154056783281944
	pesos_i(22090) := b"0000000000000000_0000000000000000_0001110111000110_0011100001111000"; -- 0.11630585604739245
	pesos_i(22091) := b"1111111111111111_1111111111111111_1111101101000000_0000101011010000"; -- -0.018554042953031587
	pesos_i(22092) := b"0000000000000000_0000000000000000_0000100100001011_0000001000010001"; -- 0.03532421977136955
	pesos_i(22093) := b"0000000000000000_0000000000000000_0001100011100010_1011111100010101"; -- 0.09720987562180866
	pesos_i(22094) := b"0000000000000000_0000000000000000_0000000100011010_0001010100111110"; -- 0.004304244652465802
	pesos_i(22095) := b"0000000000000000_0000000000000000_0000100111000000_1100110100100010"; -- 0.03809816431370983
	pesos_i(22096) := b"0000000000000000_0000000000000000_0001001011010111_1110110000101001"; -- 0.07360721590628017
	pesos_i(22097) := b"0000000000000000_0000000000000000_0001001101110100_1011011010110010"; -- 0.07599965898007954
	pesos_i(22098) := b"0000000000000000_0000000000000000_0000111111001111_1011011001010100"; -- 0.06176318700690847
	pesos_i(22099) := b"0000000000000000_0000000000000000_0000100100010011_1110101101110001"; -- 0.03546020041665764
	pesos_i(22100) := b"0000000000000000_0000000000000000_0001101110100010_0110111001001110"; -- 0.1079472485504488
	pesos_i(22101) := b"0000000000000000_0000000000000000_0000110110101010_1101011010111100"; -- 0.05338804341894199
	pesos_i(22102) := b"0000000000000000_0000000000000000_0001111100110011_0001101001010101"; -- 0.121873517742352
	pesos_i(22103) := b"1111111111111111_1111111111111111_1110010010110010_0001010101101101"; -- -0.10665765842526133
	pesos_i(22104) := b"0000000000000000_0000000000000000_0001011001000000_1010011010100000"; -- 0.08692399424033062
	pesos_i(22105) := b"0000000000000000_0000000000000000_0001110100011111_0111100101100101"; -- 0.11376150807285694
	pesos_i(22106) := b"1111111111111111_1111111111111111_1110111010100101_0110101000001011"; -- -0.06778847914488957
	pesos_i(22107) := b"1111111111111111_1111111111111111_1111000000011010_1000100101011000"; -- -0.062095085100055666
	pesos_i(22108) := b"0000000000000000_0000000000000000_0001110011000110_0000110100001000"; -- 0.11239701692076692
	pesos_i(22109) := b"0000000000000000_0000000000000000_0001100010100011_0100101011110011"; -- 0.09624164994765008
	pesos_i(22110) := b"1111111111111111_1111111111111111_1111010011101110_1111000001001011"; -- -0.04322908571412521
	pesos_i(22111) := b"0000000000000000_0000000000000000_0010000101010011_0000110010011011"; -- 0.13017348084721267
	pesos_i(22112) := b"0000000000000000_0000000000000000_0001111101010001_1010010010110101"; -- 0.12233952919567447
	pesos_i(22113) := b"0000000000000000_0000000000000000_0000000010111101_1100010011101100"; -- 0.0028956487067771414
	pesos_i(22114) := b"0000000000000000_0000000000000000_0001000011110100_0000100000111100"; -- 0.06622363532638542
	pesos_i(22115) := b"1111111111111111_1111111111111111_1110001011011011_0101001110110101"; -- -0.1138408357544668
	pesos_i(22116) := b"0000000000000000_0000000000000000_0010001000011100_1110001110000001"; -- 0.133253306354431
	pesos_i(22117) := b"0000000000000000_0000000000000000_0001001011101111_1101011110000000"; -- 0.073972195376497
	pesos_i(22118) := b"0000000000000000_0000000000000000_0001100111110111_0010001101001011"; -- 0.10142727444097008
	pesos_i(22119) := b"1111111111111111_1111111111111111_1110011000010011_0110011010000001"; -- -0.10126647332260189
	pesos_i(22120) := b"0000000000000000_0000000000000000_0000110011111111_0001010001001100"; -- 0.050767200926134896
	pesos_i(22121) := b"1111111111111111_1111111111111111_1101111110000101_1111011001101100"; -- -0.12686214307768817
	pesos_i(22122) := b"0000000000000000_0000000000000000_0001011110010011_1001110101011110"; -- 0.09209617174047811
	pesos_i(22123) := b"0000000000000000_0000000000000000_0010011110111100_0000110100101101"; -- 0.15521318761161151
	pesos_i(22124) := b"1111111111111111_1111111111111111_1110001111000110_0011101110110001"; -- -0.11025645199175951
	pesos_i(22125) := b"0000000000000000_0000000000000000_0000011110000000_1000001001100111"; -- 0.029304647575001123
	pesos_i(22126) := b"1111111111111111_1111111111111111_1111010010011000_0001000100010100"; -- -0.04455464606261672
	pesos_i(22127) := b"1111111111111111_1111111111111111_1101111111011100_1100110011000101"; -- -0.1255371111613292
	pesos_i(22128) := b"0000000000000000_0000000000000000_0001011010111000_0100101000100110"; -- 0.08874953668951
	pesos_i(22129) := b"1111111111111111_1111111111111111_1110010100100011_1011011111111000"; -- -0.10492372704587513
	pesos_i(22130) := b"1111111111111111_1111111111111111_1101100100000111_1001110111001111"; -- -0.15222753227499786
	pesos_i(22131) := b"0000000000000000_0000000000000000_0001000000101111_1100000011110100"; -- 0.06322866387307309
	pesos_i(22132) := b"0000000000000000_0000000000000000_0000000100111000_0011100011101001"; -- 0.0047641343896065716
	pesos_i(22133) := b"0000000000000000_0000000000000000_0000100100111100_1110110100001010"; -- 0.03608590596817322
	pesos_i(22134) := b"1111111111111111_1111111111111111_1111100111011010_0001010001111011"; -- -0.024016113362429214
	pesos_i(22135) := b"0000000000000000_0000000000000000_0010001011111001_0001000001101101"; -- 0.13661291763698294
	pesos_i(22136) := b"1111111111111111_1111111111111111_1111011001000011_0010010100111010"; -- -0.038037942171650456
	pesos_i(22137) := b"0000000000000000_0000000000000000_0001001101000110_0010010111010100"; -- 0.07528911996450584
	pesos_i(22138) := b"0000000000000000_0000000000000000_0001000110000011_1011000100111000"; -- 0.06841571451591565
	pesos_i(22139) := b"0000000000000000_0000000000000000_0000001110010110_0100000010110111"; -- 0.014011425556836299
	pesos_i(22140) := b"0000000000000000_0000000000000000_0000000111101011_0001101000011010"; -- 0.007493621315903774
	pesos_i(22141) := b"0000000000000000_0000000000000000_0000001100111111_0100000101010000"; -- 0.01268394667423944
	pesos_i(22142) := b"0000000000000000_0000000000000000_0001101100000010_0110011100000001"; -- 0.10550540698621212
	pesos_i(22143) := b"1111111111111111_1111111111111111_1101101001001011_0000001001101000"; -- -0.14729294745227722
	pesos_i(22144) := b"1111111111111111_1111111111111111_1110001011010110_0001000100011010"; -- -0.1139210998676781
	pesos_i(22145) := b"1111111111111111_1111111111111111_1110101000010010_0001000101111100"; -- -0.08566179973671058
	pesos_i(22146) := b"0000000000000000_0000000000000000_0001001101101111_1001010010011100"; -- 0.07592133335520054
	pesos_i(22147) := b"0000000000000000_0000000000000000_0000100101011100_0101011000011001"; -- 0.036565190503041516
	pesos_i(22148) := b"1111111111111111_1111111111111111_1110011111111110_1000000100100111"; -- -0.09377281958637645
	pesos_i(22149) := b"0000000000000000_0000000000000000_0001111001100100_0010010000010010"; -- 0.11871552879037416
	pesos_i(22150) := b"1111111111111111_1111111111111111_1111011011011111_1010010100110010"; -- -0.03564994355773084
	pesos_i(22151) := b"0000000000000000_0000000000000000_0000100100001011_0001111010111000"; -- 0.03532592773609075
	pesos_i(22152) := b"0000000000000000_0000000000000000_0000110111001001_0101101110000011"; -- 0.05385372109217732
	pesos_i(22153) := b"0000000000000000_0000000000000000_0010001110000000_1011011100101111"; -- 0.13868279358160296
	pesos_i(22154) := b"0000000000000000_0000000000000000_0010001000011000_1011101011001000"; -- 0.13318984402091222
	pesos_i(22155) := b"1111111111111111_1111111111111111_1111000001011111_1000111110010111"; -- -0.06104185634314038
	pesos_i(22156) := b"1111111111111111_1111111111111111_1110000101011010_1010011110111011"; -- -0.11971046143416873
	pesos_i(22157) := b"1111111111111111_1111111111111111_1111100111011000_0100101001110111"; -- -0.024043413188380627
	pesos_i(22158) := b"0000000000000000_0000000000000000_0001000111100000_0111000001011101"; -- 0.06983091608997435
	pesos_i(22159) := b"1111111111111111_1111111111111111_1101101101100001_0000011011101101"; -- -0.14305073471803093
	pesos_i(22160) := b"0000000000000000_0000000000000000_0001010000100101_0011000111100110"; -- 0.07869254926828638
	pesos_i(22161) := b"1111111111111111_1111111111111111_1111111001011110_1001100110100001"; -- -0.006369016818716011
	pesos_i(22162) := b"0000000000000000_0000000000000000_0000000100010100_1110011001100011"; -- 0.004225157787338866
	pesos_i(22163) := b"0000000000000000_0000000000000000_0000011011110101_0000100000101111"; -- 0.02717639106393989
	pesos_i(22164) := b"0000000000000000_0000000000000000_0000110110111111_1100001000000000"; -- 0.05370724205182985
	pesos_i(22165) := b"1111111111111111_1111111111111111_1110101001010100_0011011111101100"; -- -0.08465242844928858
	pesos_i(22166) := b"0000000000000000_0000000000000000_0001100100101111_1010011001011011"; -- 0.09838332864948
	pesos_i(22167) := b"1111111111111111_1111111111111111_1110100010011011_1110111011101000"; -- -0.0913706476790602
	pesos_i(22168) := b"0000000000000000_0000000000000000_0000000011010111_1010010000100110"; -- 0.003290423621153302
	pesos_i(22169) := b"1111111111111111_1111111111111111_1101111010011101_0000101001010000"; -- -0.1304162554099157
	pesos_i(22170) := b"0000000000000000_0000000000000000_0010010011000010_0000100111000101"; -- 0.14358578733903418
	pesos_i(22171) := b"1111111111111111_1111111111111111_1101110100111000_1000111001010111"; -- -0.13585577370318067
	pesos_i(22172) := b"1111111111111111_1111111111111111_1110100111110010_1110001100110110"; -- -0.08613758031988417
	pesos_i(22173) := b"0000000000000000_0000000000000000_0010110101110001_1010001101101000"; -- 0.1775152329118031
	pesos_i(22174) := b"0000000000000000_0000000000000000_0001111001110101_0001110000000111"; -- 0.11897444892061074
	pesos_i(22175) := b"0000000000000000_0000000000000000_0001000111010001_0000000111111001"; -- 0.06959545454776345
	pesos_i(22176) := b"0000000000000000_0000000000000000_0001101000010110_0010010111110110"; -- 0.10190045607771045
	pesos_i(22177) := b"0000000000000000_0000000000000000_0001001000010011_0100010101011101"; -- 0.07060655137581388
	pesos_i(22178) := b"1111111111111111_1111111111111111_1101110001010110_1011000100110011"; -- -0.13930218235123948
	pesos_i(22179) := b"0000000000000000_0000000000000000_0001011001110001_0100000010111111"; -- 0.08766560230894524
	pesos_i(22180) := b"1111111111111111_1111111111111111_1101101100000111_1110111000011001"; -- -0.14441024667042487
	pesos_i(22181) := b"1111111111111111_1111111111111111_1110100100111100_0111011010001111"; -- -0.0889211560171711
	pesos_i(22182) := b"0000000000000000_0000000000000000_0010100100111101_1010110011110011"; -- 0.16109734461418432
	pesos_i(22183) := b"1111111111111111_1111111111111111_1110110011001011_1000100000101110"; -- -0.07501934891112567
	pesos_i(22184) := b"0000000000000000_0000000000000000_0000000100110001_1101011100010100"; -- 0.004666750351587253
	pesos_i(22185) := b"0000000000000000_0000000000000000_0000011101010010_1101111000110001"; -- 0.028608214253923705
	pesos_i(22186) := b"0000000000000000_0000000000000000_0001010011111111_0001100000001110"; -- 0.08201742509033436
	pesos_i(22187) := b"1111111111111111_1111111111111111_1111011000101110_0010000011111111"; -- -0.03835862898898964
	pesos_i(22188) := b"1111111111111111_1111111111111111_1101111001001000_1001000101001101"; -- -0.1317052064992316
	pesos_i(22189) := b"1111111111111111_1111111111111111_1111000100011101_1000000010110101"; -- -0.05814357352576633
	pesos_i(22190) := b"1111111111111111_1111111111111111_1110101011101011_0110010000110101"; -- -0.0823457118642256
	pesos_i(22191) := b"1111111111111111_1111111111111111_1110001101010110_1101000010010111"; -- -0.11195656116073639
	pesos_i(22192) := b"0000000000000000_0000000000000000_0000111010111101_0011111111001000"; -- 0.05757521269429501
	pesos_i(22193) := b"0000000000000000_0000000000000000_0000001110001101_0001100111010110"; -- 0.013871779296489873
	pesos_i(22194) := b"0000000000000000_0000000000000000_0000011111000100_1010110011101100"; -- 0.030344779586999417
	pesos_i(22195) := b"1111111111111111_1111111111111111_1111101011000101_0111110111010001"; -- -0.02042401941067079
	pesos_i(22196) := b"0000000000000000_0000000000000000_0000100010100110_0000011001001101"; -- 0.03378333464372258
	pesos_i(22197) := b"0000000000000000_0000000000000000_0001100100111101_0001111101000011"; -- 0.09858889949317835
	pesos_i(22198) := b"1111111111111111_1111111111111111_1111010001010011_0100111011010111"; -- -0.04560382139292708
	pesos_i(22199) := b"1111111111111111_1111111111111111_1101111010101111_0000000110010010"; -- -0.13014211826513203
	pesos_i(22200) := b"0000000000000000_0000000000000000_0000011100010000_1110111000010000"; -- 0.027602080177631036
	pesos_i(22201) := b"0000000000000000_0000000000000000_0000110101011011_0101010100001101"; -- 0.05217486911177442
	pesos_i(22202) := b"1111111111111111_1111111111111111_1110101111000111_0111010101010011"; -- -0.07898775802455589
	pesos_i(22203) := b"1111111111111111_1111111111111111_1111010110110100_0001111101011110"; -- -0.040220298315866695
	pesos_i(22204) := b"0000000000000000_0000000000000000_0000001001001001_1000001010011010"; -- 0.008934175974151193
	pesos_i(22205) := b"1111111111111111_1111111111111111_1110110011110100_0100011111010000"; -- -0.07439757511285797
	pesos_i(22206) := b"0000000000000000_0000000000000000_0001000101000100_0110010010100101"; -- 0.06744984657358759
	pesos_i(22207) := b"1111111111111111_1111111111111111_1101100011101111_0000101010111110"; -- -0.1526025091531857
	pesos_i(22208) := b"1111111111111111_1111111111111111_1110110001000011_1000110100011110"; -- -0.07709424991786144
	pesos_i(22209) := b"0000000000000000_0000000000000000_0000111001111100_1111011010101010"; -- 0.056594292188592146
	pesos_i(22210) := b"0000000000000000_0000000000000000_0000000001001101_0011000101001111"; -- 0.0011778656982047316
	pesos_i(22211) := b"1111111111111111_1111111111111111_1110110101010011_0000101100111101"; -- -0.07295160057055369
	pesos_i(22212) := b"1111111111111111_1111111111111111_1111011111010100_1111110111101111"; -- -0.03190625105228827
	pesos_i(22213) := b"1111111111111111_1111111111111111_1111001100110111_0001111010001110"; -- -0.049940195429483115
	pesos_i(22214) := b"0000000000000000_0000000000000000_0001000100101110_0001101100101101"; -- 0.06710977409679825
	pesos_i(22215) := b"1111111111111111_1111111111111111_1101100110000010_0000001111101101"; -- -0.15035987347332788
	pesos_i(22216) := b"1111111111111111_1111111111111111_1101101110000011_1000101011001011"; -- -0.14252407587062957
	pesos_i(22217) := b"1111111111111111_1111111111111111_1110111011011010_0011010011111101"; -- -0.06698292552551156
	pesos_i(22218) := b"0000000000000000_0000000000000000_0000000101111010_0001010011000111"; -- 0.0057690607259991075
	pesos_i(22219) := b"0000000000000000_0000000000000000_0001001101101101_0110010101101000"; -- 0.07588800220498997
	pesos_i(22220) := b"1111111111111111_1111111111111111_1111111101000100_0110001111101101"; -- -0.0028626961927390067
	pesos_i(22221) := b"1111111111111111_1111111111111111_1110011011100100_1001001000111000"; -- -0.098074780671673
	pesos_i(22222) := b"1111111111111111_1111111111111111_1101110011001101_1110010111001110"; -- -0.13748325090421684
	pesos_i(22223) := b"1111111111111111_1111111111111111_1111010000101011_1110010010110100"; -- -0.046205240398877453
	pesos_i(22224) := b"1111111111111111_1111111111111111_1110000001110101_0001010001001100"; -- -0.123213512003916
	pesos_i(22225) := b"1111111111111111_1111111111111111_1110101111111001_1100101001010100"; -- -0.0782197517438255
	pesos_i(22226) := b"0000000000000000_0000000000000000_0010000001101000_1110010000111000"; -- 0.12660051697429348
	pesos_i(22227) := b"1111111111111111_1111111111111111_1111000010101101_0000001000000101"; -- -0.05986010910786475
	pesos_i(22228) := b"1111111111111111_1111111111111111_1111010110101010_0000100101001000"; -- -0.0403742025901688
	pesos_i(22229) := b"1111111111111111_1111111111111111_1111000001011111_0000110011101000"; -- -0.06104964566655841
	pesos_i(22230) := b"1111111111111111_1111111111111111_1111100101110010_1010100001000110"; -- -0.025594218226432312
	pesos_i(22231) := b"0000000000000000_0000000000000000_0001111010101110_0101000001101100"; -- 0.1198473228477899
	pesos_i(22232) := b"0000000000000000_0000000000000000_0010001111110110_0101101100010101"; -- 0.14047784093092963
	pesos_i(22233) := b"0000000000000000_0000000000000000_0010001100011001_1100011001001111"; -- 0.137112039887976
	pesos_i(22234) := b"1111111111111111_1111111111111111_1111110111001000_1010001000101110"; -- -0.008657325592366589
	pesos_i(22235) := b"1111111111111111_1111111111111111_1110100011011010_1011101011001101"; -- -0.0904124498695209
	pesos_i(22236) := b"1111111111111111_1111111111111111_1111011110110001_1000010010100011"; -- -0.03244753861600452
	pesos_i(22237) := b"0000000000000000_0000000000000000_0001111010011010_1100100110110011"; -- 0.11954937561406725
	pesos_i(22238) := b"0000000000000000_0000000000000000_0001011101010000_0000111100011011"; -- 0.09106535344203702
	pesos_i(22239) := b"1111111111111111_1111111111111111_1111001111010100_1001101000110001"; -- -0.04753719610701087
	pesos_i(22240) := b"1111111111111111_1111111111111111_1111110000001000_1001001000101110"; -- -0.015494216634034498
	pesos_i(22241) := b"1111111111111111_1111111111111111_1110101100101011_0011111000000011"; -- -0.08137142584061399
	pesos_i(22242) := b"0000000000000000_0000000000000000_0001110000100111_0110001110001000"; -- 0.10997602538515647
	pesos_i(22243) := b"1111111111111111_1111111111111111_1111011100110101_0110000011101000"; -- -0.034341758213335266
	pesos_i(22244) := b"0000000000000000_0000000000000000_0010100101001100_1100111110011001"; -- 0.16132829165479445
	pesos_i(22245) := b"1111111111111111_1111111111111111_1110100000100000_0101101111111010"; -- -0.09325623644233245
	pesos_i(22246) := b"1111111111111111_1111111111111111_1111000000001100_1101001111110101"; -- -0.06230426099985006
	pesos_i(22247) := b"1111111111111111_1111111111111111_1111001001110000_0011101000011101"; -- -0.052975051845981794
	pesos_i(22248) := b"1111111111111111_1111111111111111_1111010110101100_0111101011101010"; -- -0.04033691210662663
	pesos_i(22249) := b"0000000000000000_0000000000000000_0000100011101111_0100011001110100"; -- 0.0349010499916802
	pesos_i(22250) := b"0000000000000000_0000000000000000_0000101010110111_0110000011010101"; -- 0.04186063013782093
	pesos_i(22251) := b"0000000000000000_0000000000000000_0001001101000011_0001011110011011"; -- 0.0752424957589806
	pesos_i(22252) := b"1111111111111111_1111111111111111_1111011100001001_0001010101101110"; -- -0.03501764354435576
	pesos_i(22253) := b"1111111111111111_1111111111111111_1101111111110001_1000011000100100"; -- -0.1252208863492784
	pesos_i(22254) := b"0000000000000000_0000000000000000_0000110110111101_0110001101100111"; -- 0.0536710859618771
	pesos_i(22255) := b"1111111111111111_1111111111111111_1101111000010111_1110101010100111"; -- -0.13244756137483768
	pesos_i(22256) := b"0000000000000000_0000000000000000_0001000101001110_0010101010010000"; -- 0.06759897235763322
	pesos_i(22257) := b"1111111111111111_1111111111111111_1101101010000111_1111110011001001"; -- -0.14636249621183306
	pesos_i(22258) := b"0000000000000000_0000000000000000_0000011101001101_1110010000010000"; -- 0.02853227029525215
	pesos_i(22259) := b"1111111111111111_1111111111111111_1110110111111101_0110100010011101"; -- -0.0703520408197875
	pesos_i(22260) := b"0000000000000000_0000000000000000_0001000110100001_1011100111110110"; -- 0.0688739992256264
	pesos_i(22261) := b"0000000000000000_0000000000000000_0001111110100011_1111100010010011"; -- 0.12359574869155265
	pesos_i(22262) := b"0000000000000000_0000000000000000_0000111110111010_1101111100111111"; -- 0.06144519119141467
	pesos_i(22263) := b"1111111111111111_1111111111111111_1110101010110001_1001010111111101"; -- -0.08322775430687504
	pesos_i(22264) := b"1111111111111111_1111111111111111_1110000001100110_0110001010001010"; -- -0.12343773011568138
	pesos_i(22265) := b"0000000000000000_0000000000000000_0000111111000110_0010000001101100"; -- 0.06161692268564447
	pesos_i(22266) := b"0000000000000000_0000000000000000_0001010100010111_0011010101101001"; -- 0.08238538574239888
	pesos_i(22267) := b"0000000000000000_0000000000000000_0000100011101101_1111111010011110"; -- 0.03488150948331235
	pesos_i(22268) := b"0000000000000000_0000000000000000_0010000001001110_1111110111100110"; -- 0.1262053191255384
	pesos_i(22269) := b"0000000000000000_0000000000000000_0001100010000100_1010001010000110"; -- 0.09577384730156738
	pesos_i(22270) := b"0000000000000000_0000000000000000_0000001000111011_1011011100111110"; -- 0.008723690714908465
	pesos_i(22271) := b"1111111111111111_1111111111111111_1101011101111001_0110101011000011"; -- -0.15830357304575005
	pesos_i(22272) := b"1111111111111111_1111111111111111_1101110000110010_1111000111000000"; -- -0.13984765107136193
	pesos_i(22273) := b"1111111111111111_1111111111111111_1110100111110111_1011110100111000"; -- -0.08606355081086106
	pesos_i(22274) := b"0000000000000000_0000000000000000_0000101010000011_0111010001100111"; -- 0.04106833939078968
	pesos_i(22275) := b"1111111111111111_1111111111111111_1101110010000000_1001111110101001"; -- -0.1386623584591971
	pesos_i(22276) := b"0000000000000000_0000000000000000_0010000011101111_1000111111001110"; -- 0.12865542206783212
	pesos_i(22277) := b"1111111111111111_1111111111111111_1111000100000110_0000100110100010"; -- -0.05850162320185919
	pesos_i(22278) := b"1111111111111111_1111111111111111_1101101100010000_0011011101000010"; -- -0.14428381570938978
	pesos_i(22279) := b"0000000000000000_0000000000000000_0001001011011111_1010100100111000"; -- 0.07372529626901489
	pesos_i(22280) := b"0000000000000000_0000000000000000_0000100001011010_0011011110100100"; -- 0.0326266074379252
	pesos_i(22281) := b"0000000000000000_0000000000000000_0000111111111000_1000001001001100"; -- 0.06238569587054726
	pesos_i(22282) := b"1111111111111111_1111111111111111_1101110011100101_1010001011111110"; -- -0.13712102218911995
	pesos_i(22283) := b"0000000000000000_0000000000000000_0001111111100011_0011111001001110"; -- 0.12456120884955527
	pesos_i(22284) := b"0000000000000000_0000000000000000_0010001000001011_1010111010100101"; -- 0.132990756221116
	pesos_i(22285) := b"1111111111111111_1111111111111111_1110101001101000_1001110100010011"; -- -0.08434122364209419
	pesos_i(22286) := b"0000000000000000_0000000000000000_0001011110010110_0000100011111010"; -- 0.0921331034648774
	pesos_i(22287) := b"1111111111111111_1111111111111111_1111011110100011_1010100111110111"; -- -0.032658936580440195
	pesos_i(22288) := b"1111111111111111_1111111111111111_1110000011010100_0000100010100100"; -- -0.12176462177075646
	pesos_i(22289) := b"1111111111111111_1111111111111111_1111000010110101_0010001100111101"; -- -0.05973605874221935
	pesos_i(22290) := b"1111111111111111_1111111111111111_1111010100111101_0011000010111010"; -- -0.04203505951372648
	pesos_i(22291) := b"0000000000000000_0000000000000000_0000001001101100_0100100011101100"; -- 0.00946479560214459
	pesos_i(22292) := b"0000000000000000_0000000000000000_0000001000101011_1010010001101110"; -- 0.008478428694765517
	pesos_i(22293) := b"0000000000000000_0000000000000000_0010000110110010_0001000010110000"; -- 0.1316233091851989
	pesos_i(22294) := b"0000000000000000_0000000000000000_0001110010110110_0101110111110110"; -- 0.11215770010140823
	pesos_i(22295) := b"0000000000000000_0000000000000000_0000000000111000_0000000000111111"; -- 0.0008545068625406504
	pesos_i(22296) := b"0000000000000000_0000000000000000_0000111111011100_1010101110001110"; -- 0.061960909158779866
	pesos_i(22297) := b"1111111111111111_1111111111111111_1110001101111111_0100100010001101"; -- -0.1113390594848528
	pesos_i(22298) := b"0000000000000000_0000000000000000_0000010111011111_0010111011010000"; -- 0.02293675026877108
	pesos_i(22299) := b"1111111111111111_1111111111111111_1110011110100101_0010111000000101"; -- -0.09513580680307428
	pesos_i(22300) := b"0000000000000000_0000000000000000_0000101000001011_1100110111001000"; -- 0.03924261208198011
	pesos_i(22301) := b"0000000000000000_0000000000000000_0000010110010000_0111000101100001"; -- 0.02173527343248496
	pesos_i(22302) := b"0000000000000000_0000000000000000_0001010100101100_1001101001010100"; -- 0.08271183548721162
	pesos_i(22303) := b"1111111111111111_1111111111111111_1110000000110100_0100100111000000"; -- -0.12420214719688377
	pesos_i(22304) := b"0000000000000000_0000000000000000_0000101110101001_0110110001001111"; -- 0.04555394095265005
	pesos_i(22305) := b"1111111111111111_1111111111111111_1111011000001100_1001100111110001"; -- -0.038870218913363466
	pesos_i(22306) := b"0000000000000000_0000000000000000_0000101101111001_1010011011111001"; -- 0.04482501574379371
	pesos_i(22307) := b"1111111111111111_1111111111111111_1111000000010011_1011101011000010"; -- -0.062198951332056066
	pesos_i(22308) := b"1111111111111111_1111111111111111_1111010000000111_0100111011111111"; -- -0.04676347995792645
	pesos_i(22309) := b"1111111111111111_1111111111111111_1111001000111100_0110000110000111"; -- -0.0537661596633458
	pesos_i(22310) := b"0000000000000000_0000000000000000_0000110111100110_0111100101000011"; -- 0.05429799920673491
	pesos_i(22311) := b"1111111111111111_1111111111111111_1111010010011001_0110000111011111"; -- -0.044534571736557164
	pesos_i(22312) := b"1111111111111111_1111111111111111_1111111011011110_0100111011111111"; -- -0.004420340271585676
	pesos_i(22313) := b"1111111111111111_1111111111111111_1111111011101110_1100111110010101"; -- -0.004168535375432745
	pesos_i(22314) := b"0000000000000000_0000000000000000_0010011000010011_0011000000111110"; -- 0.14873029255249762
	pesos_i(22315) := b"1111111111111111_1111111111111111_1110001001011100_0000100011111111"; -- -0.11578315513818463
	pesos_i(22316) := b"1111111111111111_1111111111111111_1110010001010000_0101110100010010"; -- -0.10814874935783829
	pesos_i(22317) := b"0000000000000000_0000000000000000_0000001000011100_1011011010010110"; -- 0.008250629136676341
	pesos_i(22318) := b"1111111111111111_1111111111111111_1111011010100011_0110111111101110"; -- -0.0365686458975862
	pesos_i(22319) := b"0000000000000000_0000000000000000_0001011111000111_0000100101101010"; -- 0.09288081023397934
	pesos_i(22320) := b"0000000000000000_0000000000000000_0000101001001010_0100110010100111"; -- 0.04019621924780756
	pesos_i(22321) := b"0000000000000000_0000000000000000_0000011000010110_1011000110011111"; -- 0.023783780285609474
	pesos_i(22322) := b"1111111111111111_1111111111111111_1111111110100101_0100011011000110"; -- -0.001384331290358419
	pesos_i(22323) := b"1111111111111111_1111111111111111_1111010110101011_0000000000000101"; -- -0.04035949582555259
	pesos_i(22324) := b"0000000000000000_0000000000000000_0010001110000111_0011111001100110"; -- 0.1387824058352715
	pesos_i(22325) := b"1111111111111111_1111111111111111_1101111111000000_1001111111001001"; -- -0.12596703862118436
	pesos_i(22326) := b"0000000000000000_0000000000000000_0001111110010100_1011000001110100"; -- 0.12336256812851754
	pesos_i(22327) := b"1111111111111111_1111111111111111_1111100001010111_0010000000001011"; -- -0.0299205754765523
	pesos_i(22328) := b"1111111111111111_1111111111111111_1110001010111011_1111000011111010"; -- -0.11431974310163955
	pesos_i(22329) := b"1111111111111111_1111111111111111_1110111111011101_1011101110010001"; -- -0.06302287768735262
	pesos_i(22330) := b"0000000000000000_0000000000000000_0000101001000000_0110011011001111"; -- 0.04004519046203021
	pesos_i(22331) := b"0000000000000000_0000000000000000_0010010001101010_1010110000100101"; -- 0.14225269217383682
	pesos_i(22332) := b"1111111111111111_1111111111111111_1110010110101010_0001101001111101"; -- -0.10287317709029607
	pesos_i(22333) := b"0000000000000000_0000000000000000_0001111000011100_1010010100011110"; -- 0.1176245879491354
	pesos_i(22334) := b"1111111111111111_1111111111111111_1111001110111111_1101101110001110"; -- -0.047853734829719136
	pesos_i(22335) := b"0000000000000000_0000000000000000_0001100110111010_1110110110100001"; -- 0.10050854863774254
	pesos_i(22336) := b"1111111111111111_1111111111111111_1110000000110110_1000111001010101"; -- -0.12416754173369941
	pesos_i(22337) := b"0000000000000000_0000000000000000_0001100110100101_0111110100110001"; -- 0.10018141221729499
	pesos_i(22338) := b"1111111111111111_1111111111111111_1111001010101110_1101010011011101"; -- -0.052019782974330186
	pesos_i(22339) := b"0000000000000000_0000000000000000_0000110010010000_1100100110101011"; -- 0.049084285965027126
	pesos_i(22340) := b"0000000000000000_0000000000000000_0001010001101101_0110010011111001"; -- 0.07979422647407494
	pesos_i(22341) := b"1111111111111111_1111111111111111_1111000001011000_1110011101111101"; -- -0.061143428879900284
	pesos_i(22342) := b"1111111111111111_1111111111111111_1110000100000110_1010010111001110"; -- -0.12099231445854104
	pesos_i(22343) := b"0000000000000000_0000000000000000_0000110010011011_1001111010101110"; -- 0.04924957029465372
	pesos_i(22344) := b"0000000000000000_0000000000000000_0001100100110101_0000000110010111"; -- 0.09846506063103565
	pesos_i(22345) := b"1111111111111111_1111111111111111_1110100010101110_0011000101001101"; -- -0.09109203213048311
	pesos_i(22346) := b"0000000000000000_0000000000000000_0000011001000010_0110000111011010"; -- 0.024450412416667833
	pesos_i(22347) := b"0000000000000000_0000000000000000_0000111101100010_0101011010100000"; -- 0.06009427460012703
	pesos_i(22348) := b"1111111111111111_1111111111111111_1110110000110100_1010011100001011"; -- -0.07732158645040005
	pesos_i(22349) := b"1111111111111111_1111111111111111_1110011111100001_0101010111011110"; -- -0.09421790448967952
	pesos_i(22350) := b"0000000000000000_0000000000000000_0001000000101110_0101101000010111"; -- 0.06320727405747913
	pesos_i(22351) := b"1111111111111111_1111111111111111_1111010000111110_1011001010111010"; -- -0.045918302191318434
	pesos_i(22352) := b"0000000000000000_0000000000000000_0010010010101010_1001000010101111"; -- 0.14322761795173536
	pesos_i(22353) := b"0000000000000000_0000000000000000_0001100101001101_1100110000110010"; -- 0.09884334783979411
	pesos_i(22354) := b"1111111111111111_1111111111111111_1111101111111011_0010001111000100"; -- -0.01569916205548789
	pesos_i(22355) := b"0000000000000000_0000000000000000_0001100001110110_1110111101111110"; -- 0.09556481192760556
	pesos_i(22356) := b"0000000000000000_0000000000000000_0000100101101101_0001110000111010"; -- 0.03682114037677489
	pesos_i(22357) := b"0000000000000000_0000000000000000_0001011100111001_1101000111111010"; -- 0.09072601646234513
	pesos_i(22358) := b"0000000000000000_0000000000000000_0001100100111010_1010110000000110"; -- 0.0985515130569454
	pesos_i(22359) := b"1111111111111111_1111111111111111_1111111101110101_1110101111011110"; -- -0.0021069128135786544
	pesos_i(22360) := b"1111111111111111_1111111111111111_1111010010100001_1110010101011001"; -- -0.044404664765028
	pesos_i(22361) := b"1111111111111111_1111111111111111_1111000111111100_0100001111001000"; -- -0.05474449512913738
	pesos_i(22362) := b"0000000000000000_0000000000000000_0000110000011001_1000110001100111"; -- 0.04726483834949996
	pesos_i(22363) := b"1111111111111111_1111111111111111_1101110100101111_0100101100011111"; -- -0.13599710924409208
	pesos_i(22364) := b"1111111111111111_1111111111111111_1101111000000001_0100011111011000"; -- -0.13279295910554473
	pesos_i(22365) := b"1111111111111111_1111111111111111_1101100001101110_0011011001010010"; -- -0.15456829538587463
	pesos_i(22366) := b"1111111111111111_1111111111111111_1111110110111100_1111000101010011"; -- -0.0088357137101077
	pesos_i(22367) := b"0000000000000000_0000000000000000_0000010011111100_1000100100110110"; -- 0.019478393320913667
	pesos_i(22368) := b"1111111111111111_1111111111111111_1101110100011001_0110111101110111"; -- -0.13633063655970676
	pesos_i(22369) := b"1111111111111111_1111111111111111_1101110010111011_0101110110011010"; -- -0.13776602746869265
	pesos_i(22370) := b"0000000000000000_0000000000000000_0001100010010101_1101011010001110"; -- 0.09603634800785806
	pesos_i(22371) := b"1111111111111111_1111111111111111_1101110111000010_0100000001010011"; -- -0.13375471079566248
	pesos_i(22372) := b"0000000000000000_0000000000000000_0000100001111101_0011011101000100"; -- 0.033160642665333986
	pesos_i(22373) := b"1111111111111111_1111111111111111_1111111101001110_1111000011100010"; -- -0.0027017066247675982
	pesos_i(22374) := b"1111111111111111_1111111111111111_1111011001110101_0010000101100000"; -- -0.03727523240528877
	pesos_i(22375) := b"0000000000000000_0000000000000000_0000101111001111_0100101101001100"; -- 0.04613180748743894
	pesos_i(22376) := b"1111111111111111_1111111111111111_1110100111000001_0001000101101101"; -- -0.08689776497703762
	pesos_i(22377) := b"1111111111111111_1111111111111111_1111111101011011_1000001001000100"; -- -0.002509935799051491
	pesos_i(22378) := b"0000000000000000_0000000000000000_0010000100001100_1010110100111111"; -- 0.1290996817757231
	pesos_i(22379) := b"0000000000000000_0000000000000000_0010001000001111_1010101011111000"; -- 0.13305157243306803
	pesos_i(22380) := b"1111111111111111_1111111111111111_1111110000010011_0010111110110101"; -- -0.015332239331456774
	pesos_i(22381) := b"0000000000000000_0000000000000000_0000001110110000_0110011110110001"; -- 0.014410477381085751
	pesos_i(22382) := b"1111111111111111_1111111111111111_1111101000011000_1101011001011010"; -- -0.023058512811211088
	pesos_i(22383) := b"0000000000000000_0000000000000000_0000011001000001_0001010100000000"; -- 0.024430572959298413
	pesos_i(22384) := b"0000000000000000_0000000000000000_0010011001110110_1011111011110011"; -- 0.1502494186856177
	pesos_i(22385) := b"0000000000000000_0000000000000000_0000100010011110_0100101100111011"; -- 0.03366537273095097
	pesos_i(22386) := b"0000000000000000_0000000000000000_0000110001110011_1000110110000010"; -- 0.048638195312837425
	pesos_i(22387) := b"1111111111111111_1111111111111111_1111100011000100_1010110101100011"; -- -0.028248942706928973
	pesos_i(22388) := b"0000000000000000_0000000000000000_0000110001100001_1100111001010101"; -- 0.04836740077470611
	pesos_i(22389) := b"1111111111111111_1111111111111111_1111100001101110_1000010100001010"; -- -0.029563603392192033
	pesos_i(22390) := b"0000000000000000_0000000000000000_0001001001111001_1111010000111011"; -- 0.07217337066834913
	pesos_i(22391) := b"0000000000000000_0000000000000000_0010010110111100_0101011110111110"; -- 0.1474051321834029
	pesos_i(22392) := b"1111111111111111_1111111111111111_1111101010101000_0100001011111111"; -- -0.020870030259110186
	pesos_i(22393) := b"0000000000000000_0000000000000000_0001001100011011_1110010010000110"; -- 0.0746443583766361
	pesos_i(22394) := b"0000000000000000_0000000000000000_0001001001001011_0110110111000101"; -- 0.07146345199726507
	pesos_i(22395) := b"0000000000000000_0000000000000000_0000010010100100_1010010011010001"; -- 0.0181372651681359
	pesos_i(22396) := b"1111111111111111_1111111111111111_1111000110111001_0000010110010000"; -- -0.05577054243789786
	pesos_i(22397) := b"1111111111111111_1111111111111111_1111011110010001_0101011011010101"; -- -0.03293854987722661
	pesos_i(22398) := b"1111111111111111_1111111111111111_1110010010110001_0111001010010011"; -- -0.10666736525382334
	pesos_i(22399) := b"0000000000000000_0000000000000000_0000101110010110_0110101111101001"; -- 0.04526400032994228
	pesos_i(22400) := b"0000000000000000_0000000000000000_0000000001000111_0010001000100101"; -- 0.0010854092810173108
	pesos_i(22401) := b"0000000000000000_0000000000000000_0001110001011001_1000001011110011"; -- 0.1107408373182065
	pesos_i(22402) := b"0000000000000000_0000000000000000_0001010100111000_1100011100110111"; -- 0.08289761628155472
	pesos_i(22403) := b"1111111111111111_1111111111111111_1110111110101101_1000010001001010"; -- -0.06375859448059763
	pesos_i(22404) := b"1111111111111111_1111111111111111_1111101111001011_1110001101000010"; -- -0.016420170188376316
	pesos_i(22405) := b"1111111111111111_1111111111111111_1110001010100100_1001000010011111"; -- -0.11467643846037692
	pesos_i(22406) := b"0000000000000000_0000000000000000_0010000101000000_0111001111010100"; -- 0.1298897163456877
	pesos_i(22407) := b"0000000000000000_0000000000000000_0000101100011010_1100110001100110"; -- 0.043377661651609806
	pesos_i(22408) := b"0000000000000000_0000000000000000_0000111010001011_0100100101100011"; -- 0.056812845799536736
	pesos_i(22409) := b"1111111111111111_1111111111111111_1111101101000001_1110110001000011"; -- -0.01852534645263384
	pesos_i(22410) := b"1111111111111111_1111111111111111_1110010110101101_0111100101110101"; -- -0.10282174014015404
	pesos_i(22411) := b"1111111111111111_1111111111111111_1110000011000101_1010101010011101"; -- -0.12198384918952798
	pesos_i(22412) := b"1111111111111111_1111111111111111_1111101101101101_1101000000110110"; -- -0.01785563164870499
	pesos_i(22413) := b"1111111111111111_1111111111111111_1111001010110001_1111000111111100"; -- -0.05197227087234503
	pesos_i(22414) := b"1111111111111111_1111111111111111_1111011010100100_0101001001110111"; -- -0.036555143195625514
	pesos_i(22415) := b"0000000000000000_0000000000000000_0001111111101101_0100110111001001"; -- 0.12471471931061727
	pesos_i(22416) := b"1111111111111111_1111111111111111_1111111101111110_0010000011010011"; -- -0.001981686005861074
	pesos_i(22417) := b"1111111111111111_1111111111111111_1111111111001011_1010000111011000"; -- -0.0007990692730132884
	pesos_i(22418) := b"1111111111111111_1111111111111111_1111001111001111_0011000110010111"; -- -0.04761972484298829
	pesos_i(22419) := b"0000000000000000_0000000000000000_0001001100111111_1001111111001001"; -- 0.07518957770757748
	pesos_i(22420) := b"1111111111111111_1111111111111111_1110011010100000_0100111100011001"; -- -0.09911637911800637
	pesos_i(22421) := b"1111111111111111_1111111111111111_1111101100101100_0100110111001110"; -- -0.018855225700585385
	pesos_i(22422) := b"0000000000000000_0000000000000000_0001001010110011_0100111010001001"; -- 0.07304850425019516
	pesos_i(22423) := b"0000000000000000_0000000000000000_0000100011100011_1011100101010010"; -- 0.03472479109535619
	pesos_i(22424) := b"1111111111111111_1111111111111111_1101111011100011_0101000010100101"; -- -0.12934394801270654
	pesos_i(22425) := b"0000000000000000_0000000000000000_0001101001111001_0000111010000001"; -- 0.10340967786075873
	pesos_i(22426) := b"0000000000000000_0000000000000000_0000101001001111_0000111011110000"; -- 0.040268834645725844
	pesos_i(22427) := b"1111111111111111_1111111111111111_1111101011110101_1011010000101101"; -- -0.01968835725721986
	pesos_i(22428) := b"1111111111111111_1111111111111111_1101101100011010_0010100111010001"; -- -0.14413202910083672
	pesos_i(22429) := b"1111111111111111_1111111111111111_1101101100101101_0100100010101001"; -- -0.14384027355486265
	pesos_i(22430) := b"0000000000000000_0000000000000000_0001111000101000_1100001101111000"; -- 0.11780950237590222
	pesos_i(22431) := b"1111111111111111_1111111111111111_1111001001000100_0000000100110101"; -- -0.05364983036386231
	pesos_i(22432) := b"0000000000000000_0000000000000000_0001110100001101_0100110100101001"; -- 0.11348421344507281
	pesos_i(22433) := b"0000000000000000_0000000000000000_0000011110110100_1011010001010100"; -- 0.030101080379065837
	pesos_i(22434) := b"1111111111111111_1111111111111111_1101110100000001_1000110001000010"; -- -0.1366951311757897
	pesos_i(22435) := b"1111111111111111_1111111111111111_1101101101110010_1000001101000010"; -- -0.14278392454861252
	pesos_i(22436) := b"0000000000000000_0000000000000000_0000110111101111_1100101010101100"; -- 0.05444018085810794
	pesos_i(22437) := b"0000000000000000_0000000000000000_0000110010100101_1000011100111100"; -- 0.04940076081137405
	pesos_i(22438) := b"0000000000000000_0000000000000000_0000100111001011_0001001011010010"; -- 0.03825490588856171
	pesos_i(22439) := b"0000000000000000_0000000000000000_0010010110011111_0100101101111111"; -- 0.14696189738747115
	pesos_i(22440) := b"1111111111111111_1111111111111111_1110001010100001_1110000110011000"; -- -0.1147173884093066
	pesos_i(22441) := b"1111111111111111_1111111111111111_1111100010101011_0000111001011010"; -- -0.02863989168486359
	pesos_i(22442) := b"1111111111111111_1111111111111111_1111000111000011_1011010100101000"; -- -0.05560748847084538
	pesos_i(22443) := b"1111111111111111_1111111111111111_1101110010010110_0111110110101000"; -- -0.13832869196748487
	pesos_i(22444) := b"1111111111111111_1111111111111111_1110100001110111_0100101100011011"; -- -0.09192972736733832
	pesos_i(22445) := b"0000000000000000_0000000000000000_0000111010100100_0001011110000110"; -- 0.057191343568735876
	pesos_i(22446) := b"1111111111111111_1111111111111111_1110000010000101_1010011111111111"; -- -0.12296056779065966
	pesos_i(22447) := b"0000000000000000_0000000000000000_0001111110001001_1110101110000011"; -- 0.12319824164148047
	pesos_i(22448) := b"1111111111111111_1111111111111111_1110100001000010_0111100100000001"; -- -0.09273570747979279
	pesos_i(22449) := b"0000000000000000_0000000000000000_0001011010000100_1000100100101001"; -- 0.08795983544648393
	pesos_i(22450) := b"0000000000000000_0000000000000000_0001101001101101_1000111001110000"; -- 0.10323419799876551
	pesos_i(22451) := b"0000000000000000_0000000000000000_0000110001010100_1101111101011101"; -- 0.04817005170210407
	pesos_i(22452) := b"0000000000000000_0000000000000000_0000100110010000_1010010100101111"; -- 0.03736336131170877
	pesos_i(22453) := b"1111111111111111_1111111111111111_1111111010100100_0111000001110101"; -- -0.005303355606757907
	pesos_i(22454) := b"0000000000000000_0000000000000000_0001011001111101_0100111101000011"; -- 0.08784957297281754
	pesos_i(22455) := b"1111111111111111_1111111111111111_1110011101101001_0110101110000100"; -- -0.09604766867851364
	pesos_i(22456) := b"0000000000000000_0000000000000000_0001111110111101_1110001111111110"; -- 0.1239912506034345
	pesos_i(22457) := b"1111111111111111_1111111111111111_1110110010110111_1001001010000101"; -- -0.07532390846137438
	pesos_i(22458) := b"1111111111111111_1111111111111111_1101111001100010_1110011011001110"; -- -0.13130338175230913
	pesos_i(22459) := b"1111111111111111_1111111111111111_1111110010111010_0111000110011110"; -- -0.012780093149342387
	pesos_i(22460) := b"1111111111111111_1111111111111111_1110011000010011_1001001000111101"; -- -0.1012638665879858
	pesos_i(22461) := b"0000000000000000_0000000000000000_0000011101000010_0111010111010010"; -- 0.028357852637381928
	pesos_i(22462) := b"1111111111111111_1111111111111111_1111100101110101_0100100011110110"; -- -0.025554122940129046
	pesos_i(22463) := b"0000000000000000_0000000000000000_0010011110101000_1110101011111101"; -- 0.15492123301051716
	pesos_i(22464) := b"1111111111111111_1111111111111111_1110100101100011_1000001100100100"; -- -0.08832531322197358
	pesos_i(22465) := b"1111111111111111_1111111111111111_1111100101001110_0010101101100011"; -- -0.026150978451495294
	pesos_i(22466) := b"1111111111111111_1111111111111111_1111100011011011_1010110110111111"; -- -0.02789796923591522
	pesos_i(22467) := b"1111111111111111_1111111111111111_1111101110111100_0011011010010101"; -- -0.016659344413640937
	pesos_i(22468) := b"1111111111111111_1111111111111111_1111100000011100_0111110001111010"; -- -0.030815334622393782
	pesos_i(22469) := b"0000000000000000_0000000000000000_0000000110110110_0101111000010001"; -- 0.006688956377516751
	pesos_i(22470) := b"0000000000000000_0000000000000000_0000010001001011_1110111011001001"; -- 0.016783641814050305
	pesos_i(22471) := b"1111111111111111_1111111111111111_1111000111101100_1110001011011101"; -- -0.05497915366121369
	pesos_i(22472) := b"0000000000000000_0000000000000000_0000110110101011_1011101110100100"; -- 0.053401687168362674
	pesos_i(22473) := b"1111111111111111_1111111111111111_1111111010111011_0000101110011100"; -- -0.004958414539099395
	pesos_i(22474) := b"0000000000000000_0000000000000000_0001001000010101_1110100001001111"; -- 0.07064678128978981
	pesos_i(22475) := b"1111111111111111_1111111111111111_1111000001011111_1110011101010011"; -- -0.06103662699707274
	pesos_i(22476) := b"0000000000000000_0000000000000000_0000000101000010_0010000111010111"; -- 0.004915347027599665
	pesos_i(22477) := b"0000000000000000_0000000000000000_0001000101110011_1100010100110011"; -- 0.0681727648223796
	pesos_i(22478) := b"0000000000000000_0000000000000000_0001001010000110_0100000100001110"; -- 0.07236105537145862
	pesos_i(22479) := b"1111111111111111_1111111111111111_1110101110100011_0110011101110100"; -- -0.07953790100804647
	pesos_i(22480) := b"1111111111111111_1111111111111111_1111001101111101_1011011001101111"; -- -0.048863027472356206
	pesos_i(22481) := b"1111111111111111_1111111111111111_1111011110101011_1011010101110101"; -- -0.032536181377157185
	pesos_i(22482) := b"0000000000000000_0000000000000000_0000101000000011_1001000011010000"; -- 0.039116907964637015
	pesos_i(22483) := b"1111111111111111_1111111111111111_1111011100110110_1000000110111110"; -- -0.034324542127274454
	pesos_i(22484) := b"1111111111111111_1111111111111111_1111100101011001_0110101111111110"; -- -0.02597928103788233
	pesos_i(22485) := b"1111111111111111_1111111111111111_1110111000000001_1111001110101111"; -- -0.07028271658070934
	pesos_i(22486) := b"0000000000000000_0000000000000000_0000011000110111_1010110000000111"; -- 0.024286986953592077
	pesos_i(22487) := b"1111111111111111_1111111111111111_1110010110011001_1110010100101110"; -- -0.10312049502517283
	pesos_i(22488) := b"1111111111111111_1111111111111111_1110101001111011_1101100101000101"; -- -0.08404771858703677
	pesos_i(22489) := b"0000000000000000_0000000000000000_0001011001111110_0111101111001110"; -- 0.08786748675028451
	pesos_i(22490) := b"1111111111111111_1111111111111111_1111110011001001_1111011011110010"; -- -0.012543264274196239
	pesos_i(22491) := b"0000000000000000_0000000000000000_0000111001111011_1011110101001101"; -- 0.056575614367660586
	pesos_i(22492) := b"1111111111111111_1111111111111111_1101101000001010_0110110010111001"; -- -0.14827843174343708
	pesos_i(22493) := b"0000000000000000_0000000000000000_0000110001000001_0000111101000101"; -- 0.0478677313292878
	pesos_i(22494) := b"1111111111111111_1111111111111111_1111001110011000_0000010000111011"; -- -0.04846166198819893
	pesos_i(22495) := b"0000000000000000_0000000000000000_0000000001110111_1010011110100110"; -- 0.0018257885475898908
	pesos_i(22496) := b"1111111111111111_1111111111111111_1110110001111110_0101111111101100"; -- -0.07619667515391473
	pesos_i(22497) := b"1111111111111111_1111111111111111_1111001000000010_0001101001010011"; -- -0.05465541339760686
	pesos_i(22498) := b"0000000000000000_0000000000000000_0001000010111010_1110010010011001"; -- 0.06535176032563123
	pesos_i(22499) := b"1111111111111111_1111111111111111_1110011101111110_1001001001000011"; -- -0.09572492465806177
	pesos_i(22500) := b"0000000000000000_0000000000000000_0000010011111100_1100000110000100"; -- 0.019481749251632517
	pesos_i(22501) := b"0000000000000000_0000000000000000_0001110000101011_1001111101010100"; -- 0.1100406246798563
	pesos_i(22502) := b"0000000000000000_0000000000000000_0000001100100101_1001011010011100"; -- 0.012292302295676771
	pesos_i(22503) := b"0000000000000000_0000000000000000_0010001111011110_1101000111001101"; -- 0.14011870628475442
	pesos_i(22504) := b"1111111111111111_1111111111111111_1110100110010100_0101110001101010"; -- -0.08757994084945647
	pesos_i(22505) := b"1111111111111111_1111111111111111_1111101001000100_1110011100011110"; -- -0.022386126784941115
	pesos_i(22506) := b"0000000000000000_0000000000000000_0001000011110111_0101011101111001"; -- 0.06627413477678451
	pesos_i(22507) := b"0000000000000000_0000000000000000_0000110101010110_1111100111011011"; -- 0.052108398482277815
	pesos_i(22508) := b"0000000000000000_0000000000000000_0001111111110111_1100111010101110"; -- 0.12487498991821683
	pesos_i(22509) := b"1111111111111111_1111111111111111_1110101111010101_0010000101001100"; -- -0.07877914329747104
	pesos_i(22510) := b"1111111111111111_1111111111111111_1111000001110011_1011111101001010"; -- -0.060733837520360934
	pesos_i(22511) := b"1111111111111111_1111111111111111_1110001111010001_1011011000101101"; -- -0.1100813045908727
	pesos_i(22512) := b"0000000000000000_0000000000000000_0001000000011111_0110001111111011"; -- 0.06297898166720015
	pesos_i(22513) := b"0000000000000000_0000000000000000_0001100000100111_1100000000001101"; -- 0.09435653989144505
	pesos_i(22514) := b"1111111111111111_1111111111111111_1110100001010100_0011010010001001"; -- -0.09246513042817675
	pesos_i(22515) := b"1111111111111111_1111111111111111_1110011010110100_0001000010011011"; -- -0.09881492828485289
	pesos_i(22516) := b"0000000000000000_0000000000000000_0001100010001000_1100110101111110"; -- 0.09583744349520985
	pesos_i(22517) := b"1111111111111111_1111111111111111_1111011111000110_1000100111011010"; -- -0.032126793285219474
	pesos_i(22518) := b"1111111111111111_1111111111111111_1110001100010011_0000000101001011"; -- -0.11299125602808463
	pesos_i(22519) := b"1111111111111111_1111111111111111_1110001101111001_0001001110101111"; -- -0.11143376337556925
	pesos_i(22520) := b"0000000000000000_0000000000000000_0001001011010101_1110101100000100"; -- 0.07357663008548557
	pesos_i(22521) := b"0000000000000000_0000000000000000_0001100010111011_1001010011111000"; -- 0.09661227279166722
	pesos_i(22522) := b"1111111111111111_1111111111111111_1111000111110001_1001101001010111"; -- -0.05490718254298739
	pesos_i(22523) := b"1111111111111111_1111111111111111_1111011000101111_0111011111011011"; -- -0.03833819303506929
	pesos_i(22524) := b"0000000000000000_0000000000000000_0001011111110000_0100111110101011"; -- 0.09351060796258513
	pesos_i(22525) := b"0000000000000000_0000000000000000_0000101001000100_1111011111100101"; -- 0.04011487343283416
	pesos_i(22526) := b"0000000000000000_0000000000000000_0001000110110101_0101101000011010"; -- 0.06917346134074866
	pesos_i(22527) := b"1111111111111111_1111111111111111_1111111011110100_1100111111000001"; -- -0.004076972350149624
	pesos_i(22528) := b"0000000000000000_0000000000000000_0001001001111000_0111011001011110"; -- 0.07215060992388134
	pesos_i(22529) := b"1111111111111111_1111111111111111_1101101011000110_0111011011011101"; -- -0.1454091750161278
	pesos_i(22530) := b"1111111111111111_1111111111111111_1101101111111111_0011110111111100"; -- -0.14063656418428477
	pesos_i(22531) := b"0000000000000000_0000000000000000_0001111001100011_0001010111001100"; -- 0.1186994191976061
	pesos_i(22532) := b"1111111111111111_1111111111111111_1111110010110001_1000000001001100"; -- -0.012916547190272574
	pesos_i(22533) := b"1111111111111111_1111111111111111_1111111110001100_1010101001101000"; -- -0.0017598625348073486
	pesos_i(22534) := b"1111111111111111_1111111111111111_1110100111111111_0111101000010011"; -- -0.0859454826074839
	pesos_i(22535) := b"0000000000000000_0000000000000000_0001100100100011_1010010100010101"; -- 0.09820014734921653
	pesos_i(22536) := b"1111111111111111_1111111111111111_1111000000101010_0010110100111011"; -- -0.06185643499320301
	pesos_i(22537) := b"1111111111111111_1111111111111111_1110110011101110_0101100010111111"; -- -0.07448811848481215
	pesos_i(22538) := b"1111111111111111_1111111111111111_1101101011101010_0000000111100010"; -- -0.14486683117793936
	pesos_i(22539) := b"0000000000000000_0000000000000000_0000110000010110_1001010111101010"; -- 0.047219629014732575
	pesos_i(22540) := b"1111111111111111_1111111111111111_1110000011001001_0000010010011100"; -- -0.12193270857497175
	pesos_i(22541) := b"0000000000000000_0000000000000000_0000010001011011_1001011111100101"; -- 0.017022603355989745
	pesos_i(22542) := b"0000000000000000_0000000000000000_0001010110110001_1100010000000101"; -- 0.08474373945342868
	pesos_i(22543) := b"0000000000000000_0000000000000000_0000001100110011_0101111011110101"; -- 0.012502608049872625
	pesos_i(22544) := b"1111111111111111_1111111111111111_1110000111001110_1011001100111110"; -- -0.11793975566987484
	pesos_i(22545) := b"0000000000000000_0000000000000000_0000011100011010_1101011001010000"; -- 0.027753252450288955
	pesos_i(22546) := b"0000000000000000_0000000000000000_0001001001001000_1000001011100000"; -- 0.07141893353147169
	pesos_i(22547) := b"1111111111111111_1111111111111111_1110101101111101_0100110011000011"; -- -0.08011932604697014
	pesos_i(22548) := b"0000000000000000_0000000000000000_0000100110111100_0111111011101000"; -- 0.038032466552779975
	pesos_i(22549) := b"1111111111111111_1111111111111111_1111000101111101_0001100100101111"; -- -0.0566849003363897
	pesos_i(22550) := b"0000000000000000_0000000000000000_0000000100001001_1100001100000001"; -- 0.0040552022913698865
	pesos_i(22551) := b"0000000000000000_0000000000000000_0010010010111000_1100001110110100"; -- 0.14344428209060386
	pesos_i(22552) := b"1111111111111111_1111111111111111_1101100100010010_1001001100011100"; -- -0.15206032342582973
	pesos_i(22553) := b"0000000000000000_0000000000000000_0010010001110000_1111101011101000"; -- 0.14234893950542493
	pesos_i(22554) := b"1111111111111111_1111111111111111_1110110111001011_0010010110100001"; -- -0.0711189729748327
	pesos_i(22555) := b"1111111111111111_1111111111111111_1110111001110000_0000001010110110"; -- -0.06860335406526724
	pesos_i(22556) := b"0000000000000000_0000000000000000_0001101000010000_0101000100100111"; -- 0.10181147757250275
	pesos_i(22557) := b"1111111111111111_1111111111111111_1111100101111010_1001000011111111"; -- -0.025473535296028
	pesos_i(22558) := b"1111111111111111_1111111111111111_1101101010110000_0110100111101001"; -- -0.1457456402764583
	pesos_i(22559) := b"1111111111111111_1111111111111111_1111010000001001_0111011001011101"; -- -0.04673061583212501
	pesos_i(22560) := b"0000000000000000_0000000000000000_0000111100011010_1000000101010110"; -- 0.05899818751843014
	pesos_i(22561) := b"1111111111111111_1111111111111111_1111111101001000_0110000100010011"; -- -0.002801831075074837
	pesos_i(22562) := b"1111111111111111_1111111111111111_1111111001011001_0100101001111100"; -- -0.006450028252724562
	pesos_i(22563) := b"0000000000000000_0000000000000000_0000001110110111_1100000001101111"; -- 0.014522578314117952
	pesos_i(22564) := b"1111111111111111_1111111111111111_1110011011010110_1111010000110010"; -- -0.09828256403595612
	pesos_i(22565) := b"1111111111111111_1111111111111111_1111011010000010_1011101011111011"; -- -0.03706771246072695
	pesos_i(22566) := b"1111111111111111_1111111111111111_1110101111101100_1000101101001111"; -- -0.07842187230227735
	pesos_i(22567) := b"1111111111111111_1111111111111111_1111010100100100_1011000010101101"; -- -0.04240890297078065
	pesos_i(22568) := b"1111111111111111_1111111111111111_1110001011101101_0010100111110001"; -- -0.11356866716189853
	pesos_i(22569) := b"0000000000000000_0000000000000000_0010000100000100_0001101111111111"; -- 0.12896895396276617
	pesos_i(22570) := b"0000000000000000_0000000000000000_0000010111101100_0110101110000001"; -- 0.0231387320297373
	pesos_i(22571) := b"0000000000000000_0000000000000000_0000011010001001_1111000111101001"; -- 0.025542373030931306
	pesos_i(22572) := b"1111111111111111_1111111111111111_1110110111001101_0001000101101011"; -- -0.07108966013988284
	pesos_i(22573) := b"0000000000000000_0000000000000000_0010010001010110_0100000011000111"; -- 0.14194111692664
	pesos_i(22574) := b"0000000000000000_0000000000000000_0000110101111101_1110110000000101"; -- 0.052702666475694056
	pesos_i(22575) := b"0000000000000000_0000000000000000_0010010111010101_0010100011010101"; -- 0.14778380596492235
	pesos_i(22576) := b"0000000000000000_0000000000000000_0001000010101100_1011110101110110"; -- 0.06513580447173718
	pesos_i(22577) := b"0000000000000000_0000000000000000_0001110111111111_1110111100001110"; -- 0.11718648988034606
	pesos_i(22578) := b"1111111111111111_1111111111111111_1110101100110011_0011110101101110"; -- -0.08124939027794385
	pesos_i(22579) := b"0000000000000000_0000000000000000_0001000111100110_0110100111001101"; -- 0.06992207763472748
	pesos_i(22580) := b"0000000000000000_0000000000000000_0010010111011001_1011101010010011"; -- 0.14785352787203251
	pesos_i(22581) := b"1111111111111111_1111111111111111_1110101001111110_0011001110001110"; -- -0.08401181964778329
	pesos_i(22582) := b"1111111111111111_1111111111111111_1110001001100110_0110101111000010"; -- -0.11562468060888816
	pesos_i(22583) := b"0000000000000000_0000000000000000_0010000100110011_1101001101101011"; -- 0.12969704968771192
	pesos_i(22584) := b"0000000000000000_0000000000000000_0001010101101001_0010111101011000"; -- 0.08363624471935538
	pesos_i(22585) := b"0000000000000000_0000000000000000_0000010110010001_1010100010110110"; -- 0.021753830368844033
	pesos_i(22586) := b"0000000000000000_0000000000000000_0000101100001111_0110001010011111"; -- 0.04320351006350073
	pesos_i(22587) := b"0000000000000000_0000000000000000_0000010100111101_0011000000011101"; -- 0.02046490379790501
	pesos_i(22588) := b"1111111111111111_1111111111111111_1101110010001001_1100010000000000"; -- -0.138522863347748
	pesos_i(22589) := b"1111111111111111_1111111111111111_1101111011110101_0101001011101001"; -- -0.1290691547455334
	pesos_i(22590) := b"1111111111111111_1111111111111111_1111110001000010_1110001101000100"; -- -0.014604373827117895
	pesos_i(22591) := b"0000000000000000_0000000000000000_0010011101010110_1001110000001111"; -- 0.153665307595596
	pesos_i(22592) := b"0000000000000000_0000000000000000_0000010110010101_1000011101111000"; -- 0.021812884078585032
	pesos_i(22593) := b"1111111111111111_1111111111111111_1110010011010000_0010101011010110"; -- -0.10619861861529287
	pesos_i(22594) := b"1111111111111111_1111111111111111_1111100011111100_1011000001000110"; -- -0.027394278522564288
	pesos_i(22595) := b"1111111111111111_1111111111111111_1111110011111111_1110100001011000"; -- -0.0117201599897192
	pesos_i(22596) := b"0000000000000000_0000000000000000_0000111000111111_1000110011100010"; -- 0.05565720107003444
	pesos_i(22597) := b"1111111111111111_1111111111111111_1101100101010010_1000100001110101"; -- -0.15108439586372685
	pesos_i(22598) := b"1111111111111111_1111111111111111_1110111010101001_1100010101101110"; -- -0.06772199703095239
	pesos_i(22599) := b"0000000000000000_0000000000000000_0000101101101000_1111110010000000"; -- 0.044570714138887094
	pesos_i(22600) := b"1111111111111111_1111111111111111_1110101111111000_1000100110001010"; -- -0.07823887237448104
	pesos_i(22601) := b"0000000000000000_0000000000000000_0000011011000011_0000010101010001"; -- 0.026413280659400438
	pesos_i(22602) := b"1111111111111111_1111111111111111_1110110110101101_1000111011100011"; -- -0.07157046269859266
	pesos_i(22603) := b"1111111111111111_1111111111111111_1111101001100101_1110101111001000"; -- -0.021882308573889415
	pesos_i(22604) := b"1111111111111111_1111111111111111_1111010010000010_0000011000000001"; -- -0.04489099956184754
	pesos_i(22605) := b"0000000000000000_0000000000000000_0000100100001000_0000001010101101"; -- 0.03527847969828319
	pesos_i(22606) := b"0000000000000000_0000000000000000_0010000100000110_1100111101111110"; -- 0.12901017019477287
	pesos_i(22607) := b"1111111111111111_1111111111111111_1101111100000100_0000001010101100"; -- -0.12884505559245465
	pesos_i(22608) := b"1111111111111111_1111111111111111_1111000011011101_1110100011101100"; -- -0.05911392433659795
	pesos_i(22609) := b"0000000000000000_0000000000000000_0010010010100000_1100100111111001"; -- 0.1430784447287438
	pesos_i(22610) := b"0000000000000000_0000000000000000_0001111011001100_0000100000001111"; -- 0.12030077327180884
	pesos_i(22611) := b"0000000000000000_0000000000000000_0000010000001010_0101101100110010"; -- 0.015783023492661953
	pesos_i(22612) := b"0000000000000000_0000000000000000_0001101000011001_0101101010010111"; -- 0.10194936929928103
	pesos_i(22613) := b"0000000000000000_0000000000000000_0000011010111111_1111110111111111"; -- 0.026367068127551862
	pesos_i(22614) := b"1111111111111111_1111111111111111_1111001110011110_1111110010111011"; -- -0.04835529742315372
	pesos_i(22615) := b"0000000000000000_0000000000000000_0001000110101001_0111011101111010"; -- 0.06899210675269303
	pesos_i(22616) := b"0000000000000000_0000000000000000_0000111100010100_0110011000001001"; -- 0.05890500751962918
	pesos_i(22617) := b"1111111111111111_1111111111111111_1111000100111100_0110110010000100"; -- -0.05767175470443484
	pesos_i(22618) := b"1111111111111111_1111111111111111_1110111110001110_1100010100101110"; -- -0.0642277492413634
	pesos_i(22619) := b"0000000000000000_0000000000000000_0000011111000101_1011011110101010"; -- 0.030360678587980347
	pesos_i(22620) := b"1111111111111111_1111111111111111_1111101010110101_1001011000110101"; -- -0.020666706186031312
	pesos_i(22621) := b"1111111111111111_1111111111111111_1101100111011000_0100000000110100"; -- -0.1490440247533303
	pesos_i(22622) := b"0000000000000000_0000000000000000_0000110001001001_0100010001010011"; -- 0.04799296407046058
	pesos_i(22623) := b"0000000000000000_0000000000000000_0000000100100010_1011110110100000"; -- 0.004436351447113197
	pesos_i(22624) := b"0000000000000000_0000000000000000_0000100111010000_0110100011111110"; -- 0.03833633614623184
	pesos_i(22625) := b"0000000000000000_0000000000000000_0001000010110101_0101110110110011"; -- 0.06526742577852236
	pesos_i(22626) := b"0000000000000000_0000000000000000_0010000000111111_0101001110000111"; -- 0.1259662824359553
	pesos_i(22627) := b"1111111111111111_1111111111111111_1110110011010000_1110011110100011"; -- -0.07493736528180685
	pesos_i(22628) := b"1111111111111111_1111111111111111_1101101110101011_1101111010000110"; -- -0.1419087336907441
	pesos_i(22629) := b"0000000000000000_0000000000000000_0000010100110101_0000010001100001"; -- 0.020340226799670565
	pesos_i(22630) := b"1111111111111111_1111111111111111_1110110001111000_0011100110101101"; -- -0.07629050761035619
	pesos_i(22631) := b"1111111111111111_1111111111111111_1111001000001011_1000000100001101"; -- -0.054511961239709646
	pesos_i(22632) := b"1111111111111111_1111111111111111_1111110001000100_1011100111000101"; -- -0.014576329634149197
	pesos_i(22633) := b"1111111111111111_1111111111111111_1111101111011001_0100011110011011"; -- -0.016215824671766108
	pesos_i(22634) := b"0000000000000000_0000000000000000_0000101100110010_1010101011011000"; -- 0.04374187242419259
	pesos_i(22635) := b"1111111111111111_1111111111111111_1110111010111011_1110000000010001"; -- -0.06744575100406329
	pesos_i(22636) := b"0000000000000000_0000000000000000_0001000111111011_1000111000000100"; -- 0.0702446708153715
	pesos_i(22637) := b"0000000000000000_0000000000000000_0001110010101010_1010100011100000"; -- 0.11197905984701607
	pesos_i(22638) := b"1111111111111111_1111111111111111_1111011110001010_1100111101011000"; -- -0.03303817849354106
	pesos_i(22639) := b"0000000000000000_0000000000000000_0000000001011000_0111010100010100"; -- 0.0013497519412224075
	pesos_i(22640) := b"1111111111111111_1111111111111111_1110000010111010_1101011001010111"; -- -0.12214908959321406
	pesos_i(22641) := b"1111111111111111_1111111111111111_1111000101001011_1111110011001011"; -- -0.05743427329048324
	pesos_i(22642) := b"1111111111111111_1111111111111111_1101110100110011_1101010010011001"; -- -0.1359278799606131
	pesos_i(22643) := b"1111111111111111_1111111111111111_1111100001001010_1010000010010111"; -- -0.03011127776669252
	pesos_i(22644) := b"0000000000000000_0000000000000000_0001001000111010_1100100011111011"; -- 0.07120948922782976
	pesos_i(22645) := b"1111111111111111_1111111111111111_1111011100100001_1011101001010100"; -- -0.034641603863981074
	pesos_i(22646) := b"1111111111111111_1111111111111111_1111000100001100_1110111110000000"; -- -0.058396369150227556
	pesos_i(22647) := b"1111111111111111_1111111111111111_1110100011100101_0101000111101110"; -- -0.09025085395937289
	pesos_i(22648) := b"0000000000000000_0000000000000000_0000111110001001_0110011100100001"; -- 0.060690351119773334
	pesos_i(22649) := b"0000000000000000_0000000000000000_0000011011110010_1000101011110101"; -- 0.027138409368640804
	pesos_i(22650) := b"0000000000000000_0000000000000000_0010010000010100_1111110011011100"; -- 0.1409452472990777
	pesos_i(22651) := b"1111111111111111_1111111111111111_1101011010110110_0101010111110110"; -- -0.16128027683506474
	pesos_i(22652) := b"0000000000000000_0000000000000000_0001011101011111_1001110110101111"; -- 0.0913027336301155
	pesos_i(22653) := b"1111111111111111_1111111111111111_1101100011011010_1100010001111111"; -- -0.15291187197243572
	pesos_i(22654) := b"0000000000000000_0000000000000000_0000010010111111_1010000001000011"; -- 0.018548981055336443
	pesos_i(22655) := b"0000000000000000_0000000000000000_0010010110011011_1001101000001001"; -- 0.1469055434933687
	pesos_i(22656) := b"0000000000000000_0000000000000000_0000000100110111_0100100011110000"; -- 0.004749830708617543
	pesos_i(22657) := b"1111111111111111_1111111111111111_1110111101100001_0001001000010000"; -- -0.0649250708006688
	pesos_i(22658) := b"1111111111111111_1111111111111111_1110100000011011_1111101010111011"; -- -0.09332306801482163
	pesos_i(22659) := b"1111111111111111_1111111111111111_1110101101011010_0111101001001001"; -- -0.08065067014591283
	pesos_i(22660) := b"1111111111111111_1111111111111111_1111100001000010_1111010011110010"; -- -0.03022832010460149
	pesos_i(22661) := b"0000000000000000_0000000000000000_0000000010001000_0011100011101100"; -- 0.0020785880864480134
	pesos_i(22662) := b"1111111111111111_1111111111111111_1110010011001100_0100001100001001"; -- -0.1062582113186228
	pesos_i(22663) := b"0000000000000000_0000000000000000_0000101010101111_0110001110001100"; -- 0.04173872153018336
	pesos_i(22664) := b"0000000000000000_0000000000000000_0000100010100111_0110100001000001"; -- 0.03380443182875822
	pesos_i(22665) := b"1111111111111111_1111111111111111_1110001111001101_1010001110000001"; -- -0.1101434526304257
	pesos_i(22666) := b"1111111111111111_1111111111111111_1101111011011110_1000001110101011"; -- -0.12941720076879815
	pesos_i(22667) := b"1111111111111111_1111111111111111_1110100000111110_0111101011001011"; -- -0.09279663608895418
	pesos_i(22668) := b"0000000000000000_0000000000000000_0001101111100011_0110001101011101"; -- 0.10893841760035086
	pesos_i(22669) := b"1111111111111111_1111111111111111_1111100001101100_0111110010111100"; -- -0.029594616106648555
	pesos_i(22670) := b"1111111111111111_1111111111111111_1111001101011110_0001000110011001"; -- -0.0493458748297102
	pesos_i(22671) := b"0000000000000000_0000000000000000_0010000101101111_0100100101010001"; -- 0.1306043455574169
	pesos_i(22672) := b"0000000000000000_0000000000000000_0001110011110110_1000101010001010"; -- 0.11313691972530775
	pesos_i(22673) := b"0000000000000000_0000000000000000_0010011110000101_1110010110111011"; -- 0.15438686200124815
	pesos_i(22674) := b"0000000000000000_0000000000000000_0010001010000000_0010000000001111"; -- 0.13476753575235625
	pesos_i(22675) := b"0000000000000000_0000000000000000_0001001111111110_1001101111000111"; -- 0.07810376752966837
	pesos_i(22676) := b"1111111111111111_1111111111111111_1110000101101101_0010011100101010"; -- -0.11942820761642244
	pesos_i(22677) := b"0000000000000000_0000000000000000_0001010000101110_0110110010000101"; -- 0.07883337259070766
	pesos_i(22678) := b"1111111111111111_1111111111111111_1101101000001100_0010111000100011"; -- -0.1482516444532841
	pesos_i(22679) := b"1111111111111111_1111111111111111_1101110101010111_1101110000000100"; -- -0.13537812145845274
	pesos_i(22680) := b"0000000000000000_0000000000000000_0000010011110010_0000000110110111"; -- 0.019317729219367717
	pesos_i(22681) := b"0000000000000000_0000000000000000_0001110001001101_1100010100110010"; -- 0.11056168039902078
	pesos_i(22682) := b"0000000000000000_0000000000000000_0001100110001100_0011110011000011"; -- 0.0997961021575118
	pesos_i(22683) := b"0000000000000000_0000000000000000_0000110010110101_1000001001100001"; -- 0.04964461194473461
	pesos_i(22684) := b"0000000000000000_0000000000000000_0001111110010000_1101000110000001"; -- 0.12330350308267313
	pesos_i(22685) := b"1111111111111111_1111111111111111_1110110001111110_0001000001101001"; -- -0.07620141445001563
	pesos_i(22686) := b"0000000000000000_0000000000000000_0000101110101100_0100000110010000"; -- 0.045597169517041125
	pesos_i(22687) := b"1111111111111111_1111111111111111_1101101111000101_1111010101001101"; -- -0.1415106474746566
	pesos_i(22688) := b"1111111111111111_1111111111111111_1111101110101110_0000000010000010"; -- -0.0168761903861225
	pesos_i(22689) := b"0000000000000000_0000000000000000_0010010000010011_1101000101011010"; -- 0.14092739540810892
	pesos_i(22690) := b"0000000000000000_0000000000000000_0001111010100100_1010111110101101"; -- 0.11970041253781896
	pesos_i(22691) := b"1111111111111111_1111111111111111_1111101101010001_1111000001011111"; -- -0.018280960822760522
	pesos_i(22692) := b"0000000000000000_0000000000000000_0010001011010000_1110111011001001"; -- 0.1360005609105877
	pesos_i(22693) := b"0000000000000000_0000000000000000_0010010010010111_0001011111001011"; -- 0.14293049538719282
	pesos_i(22694) := b"1111111111111111_1111111111111111_1111101010010100_1001110000110001"; -- -0.0211698894077039
	pesos_i(22695) := b"1111111111111111_1111111111111111_1111100111011101_1111100101110111"; -- -0.023956688339459572
	pesos_i(22696) := b"1111111111111111_1111111111111111_1110100100000001_1101110011010011"; -- -0.08981532900717644
	pesos_i(22697) := b"1111111111111111_1111111111111111_1111101000110111_0111001000111010"; -- -0.02259145813717396
	pesos_i(22698) := b"0000000000000000_0000000000000000_0000101001011100_0000000000100011"; -- 0.040466316826964735
	pesos_i(22699) := b"0000000000000000_0000000000000000_0001110011010100_0101010010010100"; -- 0.11261490463316087
	pesos_i(22700) := b"1111111111111111_1111111111111111_1111101000101100_0011010011001110"; -- -0.02276296581788124
	pesos_i(22701) := b"0000000000000000_0000000000000000_0001001111011011_0101100111011001"; -- 0.07756578024665188
	pesos_i(22702) := b"1111111111111111_1111111111111111_1110100100001011_1000110101010111"; -- -0.08966747886190397
	pesos_i(22703) := b"0000000000000000_0000000000000000_0000000011100001_1110001010110000"; -- 0.0034467392364443887
	pesos_i(22704) := b"0000000000000000_0000000000000000_0000000100001100_1111111011110101"; -- 0.0041045521663177174
	pesos_i(22705) := b"0000000000000000_0000000000000000_0000010010110011_0110110011000010"; -- 0.01836280571882478
	pesos_i(22706) := b"0000000000000000_0000000000000000_0000111010101000_1100010101100000"; -- 0.05726274098494765
	pesos_i(22707) := b"1111111111111111_1111111111111111_1111000011000001_0000110100100101"; -- -0.05955427034666417
	pesos_i(22708) := b"0000000000000000_0000000000000000_0001111111110110_1101101010110101"; -- 0.12486044807314944
	pesos_i(22709) := b"0000000000000000_0000000000000000_0001111000110011_1110001001011110"; -- 0.11797919086899951
	pesos_i(22710) := b"0000000000000000_0000000000000000_0010000000101101_0111010000001111"; -- 0.12569356321175504
	pesos_i(22711) := b"0000000000000000_0000000000000000_0010000011101100_0110100010001000"; -- 0.12860730482555494
	pesos_i(22712) := b"1111111111111111_1111111111111111_1110100010111111_1110011111011000"; -- -0.0908217523304914
	pesos_i(22713) := b"0000000000000000_0000000000000000_0000000011000000_1100101111111100"; -- 0.0029418458365165247
	pesos_i(22714) := b"1111111111111111_1111111111111111_1111000000000111_1010101111100111"; -- -0.062382942281519124
	pesos_i(22715) := b"1111111111111111_1111111111111111_1101100110000010_0011011000000110"; -- -0.1503568874223883
	pesos_i(22716) := b"0000000000000000_0000000000000000_0001100011010111_1110101010000111"; -- 0.09704461853052807
	pesos_i(22717) := b"1111111111111111_1111111111111111_1101101101011100_0111100000011001"; -- -0.14312028292390283
	pesos_i(22718) := b"1111111111111111_1111111111111111_1111010010110000_1000001101010010"; -- -0.04418162593462825
	pesos_i(22719) := b"1111111111111111_1111111111111111_1110100110100010_0000011010011011"; -- -0.0873714324290336
	pesos_i(22720) := b"0000000000000000_0000000000000000_0010000001011000_0000100111101100"; -- 0.1263433647176787
	pesos_i(22721) := b"0000000000000000_0000000000000000_0000110010000011_1010001000100001"; -- 0.04888356511122683
	pesos_i(22722) := b"0000000000000000_0000000000000000_0001000001111110_0000000001000101"; -- 0.06442262358093523
	pesos_i(22723) := b"0000000000000000_0000000000000000_0000101000001100_1111011101110110"; -- 0.039260355307979396
	pesos_i(22724) := b"0000000000000000_0000000000000000_0000100110101001_0111100110010110"; -- 0.037742232489279604
	pesos_i(22725) := b"0000000000000000_0000000000000000_0000111111100000_1000000011100010"; -- 0.06201940071275159
	pesos_i(22726) := b"1111111111111111_1111111111111111_1101101010100101_0100001111111011"; -- -0.1459157477968787
	pesos_i(22727) := b"1111111111111111_1111111111111111_1111001100000010_0000011111110000"; -- -0.05075025932982173
	pesos_i(22728) := b"1111111111111111_1111111111111111_1111010110110000_1000000001011011"; -- -0.04027555259413454
	pesos_i(22729) := b"0000000000000000_0000000000000000_0000011001111111_0011011100000000"; -- 0.025378644460257702
	pesos_i(22730) := b"1111111111111111_1111111111111111_1110011011101001_1010010101110111"; -- -0.09799733965047817
	pesos_i(22731) := b"1111111111111111_1111111111111111_1111001011100000_1111111110101110"; -- -0.05125429157325895
	pesos_i(22732) := b"1111111111111111_1111111111111111_1111100001101000_1100010100010000"; -- -0.029651339987359828
	pesos_i(22733) := b"0000000000000000_0000000000000000_0000010001100011_1000100011101000"; -- 0.01714378036014404
	pesos_i(22734) := b"0000000000000000_0000000000000000_0000111101011001_1010010101110111"; -- 0.059961644702483205
	pesos_i(22735) := b"0000000000000000_0000000000000000_0001000100111011_0110110011101000"; -- 0.06731300992713267
	pesos_i(22736) := b"1111111111111111_1111111111111111_1110001010010100_1111001001000101"; -- -0.11491475887256286
	pesos_i(22737) := b"1111111111111111_1111111111111111_1111011111011001_0101110011100000"; -- -0.031839556964564884
	pesos_i(22738) := b"1111111111111111_1111111111111111_1110110011110001_0000011100011011"; -- -0.0744472082049411
	pesos_i(22739) := b"0000000000000000_0000000000000000_0000110001101011_1100000110100100"; -- 0.04851923223811985
	pesos_i(22740) := b"1111111111111111_1111111111111111_1111000001001000_1011101010001100"; -- -0.061390248090498235
	pesos_i(22741) := b"0000000000000000_0000000000000000_0001110110100100_0110101110001000"; -- 0.11579010079224163
	pesos_i(22742) := b"1111111111111111_1111111111111111_1111010000001011_0100111100001000"; -- -0.046702442712241214
	pesos_i(22743) := b"1111111111111111_1111111111111111_1110110111000001_1110000000101100"; -- -0.07126044196948364
	pesos_i(22744) := b"0000000000000000_0000000000000000_0000110010110111_1110101010110111"; -- 0.049681348585754494
	pesos_i(22745) := b"1111111111111111_1111111111111111_1110100101011001_1111001001000101"; -- -0.08847127727592312
	pesos_i(22746) := b"0000000000000000_0000000000000000_0001011100000101_1100011110100111"; -- 0.08993194408343122
	pesos_i(22747) := b"0000000000000000_0000000000000000_0010001110110100_0111001110101111"; -- 0.1394722273190169
	pesos_i(22748) := b"1111111111111111_1111111111111111_1101110011001010_1101011010010110"; -- -0.1375299343467065
	pesos_i(22749) := b"1111111111111111_1111111111111111_1110000001111110_0111010000100011"; -- -0.12307047038740879
	pesos_i(22750) := b"1111111111111111_1111111111111111_1111110100101111_1100101001110100"; -- -0.010989519736578171
	pesos_i(22751) := b"1111111111111111_1111111111111111_1110001101010101_1011111110001001"; -- -0.11197283663896264
	pesos_i(22752) := b"0000000000000000_0000000000000000_0001100110100001_0101011110110011"; -- 0.10011814240725032
	pesos_i(22753) := b"0000000000000000_0000000000000000_0000011100001111_0101110111100101"; -- 0.027578228340025046
	pesos_i(22754) := b"0000000000000000_0000000000000000_0010010101010101_0001110101000111"; -- 0.14582999213136408
	pesos_i(22755) := b"0000000000000000_0000000000000000_0010000000111011_0011001110010110"; -- 0.1259033433017217
	pesos_i(22756) := b"0000000000000000_0000000000000000_0000100011000000_1100110001011111"; -- 0.03419186897791301
	pesos_i(22757) := b"1111111111111111_1111111111111111_1110001101110111_1110000011011111"; -- -0.111452050830153
	pesos_i(22758) := b"0000000000000000_0000000000000000_0001100110100101_1110000000010001"; -- 0.10018730552819237
	pesos_i(22759) := b"0000000000000000_0000000000000000_0000100110011011_1000100011001111"; -- 0.03752951672060979
	pesos_i(22760) := b"1111111111111111_1111111111111111_1111101001010100_1011101101110010"; -- -0.022144589081422916
	pesos_i(22761) := b"1111111111111111_1111111111111111_1110110001011001_1111011010011010"; -- -0.07675226919324471
	pesos_i(22762) := b"0000000000000000_0000000000000000_0010000000101111_1000110001110100"; -- 0.12572553467272166
	pesos_i(22763) := b"1111111111111111_1111111111111111_1110001111001100_1101001101101110"; -- -0.11015585483617396
	pesos_i(22764) := b"1111111111111111_1111111111111111_1111100000111010_1011010011000111"; -- -0.030354215032436477
	pesos_i(22765) := b"1111111111111111_1111111111111111_1101111000110011_1001110110111111"; -- -0.1320248992631631
	pesos_i(22766) := b"0000000000000000_0000000000000000_0000000100000100_1110010011011110"; -- 0.00398092671534376
	pesos_i(22767) := b"0000000000000000_0000000000000000_0000010100000100_0100101101011110"; -- 0.01959677741088565
	pesos_i(22768) := b"0000000000000000_0000000000000000_0010001101111010_0011110100111101"; -- 0.13858397224441044
	pesos_i(22769) := b"0000000000000000_0000000000000000_0000110101100111_1011011111101111"; -- 0.052363868562929454
	pesos_i(22770) := b"1111111111111111_1111111111111111_1111111011010010_1010111001100010"; -- -0.004597760373465864
	pesos_i(22771) := b"0000000000000000_0000000000000000_0001110101101000_1110001011011101"; -- 0.11488168609660496
	pesos_i(22772) := b"0000000000000000_0000000000000000_0001000001110001_0100111001010001"; -- 0.06422891129023561
	pesos_i(22773) := b"1111111111111111_1111111111111111_1111101010110011_1111011010011000"; -- -0.020691478656215866
	pesos_i(22774) := b"1111111111111111_1111111111111111_1101111111100111_0111011100001111"; -- -0.12537437323341868
	pesos_i(22775) := b"0000000000000000_0000000000000000_0010000011001111_0001011110000111"; -- 0.12815997172684562
	pesos_i(22776) := b"1111111111111111_1111111111111111_1110010010101011_0111111011101001"; -- -0.10675818269987476
	pesos_i(22777) := b"0000000000000000_0000000000000000_0000101011011111_0101001111111111"; -- 0.04247021643191142
	pesos_i(22778) := b"0000000000000000_0000000000000000_0001101101101010_0011011110111001"; -- 0.10708950297200014
	pesos_i(22779) := b"0000000000000000_0000000000000000_0010010101100111_0000001100100111"; -- 0.14610309314052336
	pesos_i(22780) := b"0000000000000000_0000000000000000_0010010010011001_1011001011100001"; -- 0.14297025676389574
	pesos_i(22781) := b"1111111111111111_1111111111111111_1101111010010001_0000110101010011"; -- -0.13059918141400573
	pesos_i(22782) := b"1111111111111111_1111111111111111_1111001010001101_0110111100001010"; -- -0.0525293923189091
	pesos_i(22783) := b"1111111111111111_1111111111111111_1110110111111001_1110111100001010"; -- -0.07040506362556383
	pesos_i(22784) := b"1111111111111111_1111111111111111_1111001100000111_1101110111001001"; -- -0.050661219046645264
	pesos_i(22785) := b"0000000000000000_0000000000000000_0000011110000111_0010010101101111"; -- 0.029405917844485353
	pesos_i(22786) := b"1111111111111111_1111111111111111_1111000000000000_0100110111010110"; -- -0.06249536050435889
	pesos_i(22787) := b"0000000000000000_0000000000000000_0001000011000101_0111100010101110"; -- 0.0655131745038802
	pesos_i(22788) := b"0000000000000000_0000000000000000_0010001011000010_0000011110110100"; -- 0.1357731642326782
	pesos_i(22789) := b"1111111111111111_1111111111111111_1110011000010001_0001000110010001"; -- -0.1013020536506537
	pesos_i(22790) := b"0000000000000000_0000000000000000_0001000011110101_1110101001010111"; -- 0.06625237102396475
	pesos_i(22791) := b"0000000000000000_0000000000000000_0000101110111100_1111000011100001"; -- 0.04585175986993463
	pesos_i(22792) := b"1111111111111111_1111111111111111_1111111110110001_0010100110101011"; -- -0.001202960828950758
	pesos_i(22793) := b"0000000000000000_0000000000000000_0001001010101001_1101100101111000"; -- 0.07290419753606202
	pesos_i(22794) := b"0000000000000000_0000000000000000_0000110110001111_1100011110010111"; -- 0.052975153417398856
	pesos_i(22795) := b"1111111111111111_1111111111111111_1110011110101100_1000010100100101"; -- -0.09502380229669308
	pesos_i(22796) := b"0000000000000000_0000000000000000_0001111101010000_1010101001110001"; -- 0.12232461230890121
	pesos_i(22797) := b"0000000000000000_0000000000000000_0010010000111010_0100111011101101"; -- 0.141514714043645
	pesos_i(22798) := b"0000000000000000_0000000000000000_0001000000011011_0000110101010000"; -- 0.06291278074411305
	pesos_i(22799) := b"0000000000000000_0000000000000000_0001110101100000_0001011000100110"; -- 0.11474741382673838
	pesos_i(22800) := b"0000000000000000_0000000000000000_0001111011111001_1011100010000101"; -- 0.12099793676881146
	pesos_i(22801) := b"0000000000000000_0000000000000000_0010011001010011_0010011100000001"; -- 0.14970630433869028
	pesos_i(22802) := b"0000000000000000_0000000000000000_0001001011110101_1000100101011100"; -- 0.07405909066347194
	pesos_i(22803) := b"0000000000000000_0000000000000000_0001010001010111_1000001011010010"; -- 0.07946031225215582
	pesos_i(22804) := b"1111111111111111_1111111111111111_1110000001010011_1100001101111110"; -- -0.12372186837722295
	pesos_i(22805) := b"0000000000000000_0000000000000000_0000111010110011_0110010101111111"; -- 0.05742487277654726
	pesos_i(22806) := b"0000000000000000_0000000000000000_0001011010000100_1011100100101100"; -- 0.08796269726857946
	pesos_i(22807) := b"1111111111111111_1111111111111111_1101110001100100_1011011110000110"; -- -0.1390881821616555
	pesos_i(22808) := b"0000000000000000_0000000000000000_0000000011010000_0100110111101100"; -- 0.0031784726371815114
	pesos_i(22809) := b"0000000000000000_0000000000000000_0001100111001110_0011110000001010"; -- 0.10080313905768336
	pesos_i(22810) := b"0000000000000000_0000000000000000_0001000011101011_0111110011101101"; -- 0.06609326154670289
	pesos_i(22811) := b"1111111111111111_1111111111111111_1101011111010111_0111100010000101"; -- -0.15686842688346503
	pesos_i(22812) := b"0000000000000000_0000000000000000_0001111001010010_0001101000001100"; -- 0.11844027310806186
	pesos_i(22813) := b"0000000000000000_0000000000000000_0010101010000110_1011010011111011"; -- 0.16611796491549213
	pesos_i(22814) := b"0000000000000000_0000000000000000_0001100010110011_1100101011100010"; -- 0.09649341597755005
	pesos_i(22815) := b"1111111111111111_1111111111111111_1111001111010011_1100110000011110"; -- -0.04754947913449418
	pesos_i(22816) := b"0000000000000000_0000000000000000_0001101001011101_0101111111011011"; -- 0.10298728085857801
	pesos_i(22817) := b"1111111111111111_1111111111111111_1111111011110011_0001001111000001"; -- -0.004103436795686486
	pesos_i(22818) := b"1111111111111111_1111111111111111_1110001111010101_0110111010100110"; -- -0.1100245328480025
	pesos_i(22819) := b"1111111111111111_1111111111111111_1111010000111000_0000001000000100"; -- -0.04602038768841369
	pesos_i(22820) := b"1111111111111111_1111111111111111_1110111111001001_1100111110011100"; -- -0.06332685897958219
	pesos_i(22821) := b"1111111111111111_1111111111111111_1111110000110000_1001110011111111"; -- -0.014883220331354816
	pesos_i(22822) := b"1111111111111111_1111111111111111_1101110001010001_1011101101101010"; -- -0.13937786735902002
	pesos_i(22823) := b"0000000000000000_0000000000000000_0000100110000101_0100110000110100"; -- 0.037190210953339006
	pesos_i(22824) := b"0000000000000000_0000000000000000_0001110111100100_0111011010100111"; -- 0.11676732622907844
	pesos_i(22825) := b"1111111111111111_1111111111111111_1101110100100110_1101110010100010"; -- -0.13612576537685056
	pesos_i(22826) := b"1111111111111111_1111111111111111_1111101101100001_1000111101110101"; -- -0.01804259685247818
	pesos_i(22827) := b"0000000000000000_0000000000000000_0000011110001100_1101101001010111"; -- 0.029492994472690263
	pesos_i(22828) := b"1111111111111111_1111111111111111_1111000111000101_1100101100010001"; -- -0.055575664762426494
	pesos_i(22829) := b"0000000000000000_0000000000000000_0001001011111000_0100101001011000"; -- 0.07410111082257395
	pesos_i(22830) := b"1111111111111111_1111111111111111_1111100101001111_0110111010001100"; -- -0.02613171647604552
	pesos_i(22831) := b"1111111111111111_1111111111111111_1111111101011010_0010011110001111"; -- -0.002530601177192944
	pesos_i(22832) := b"0000000000000000_0000000000000000_0000011101101011_1000100011101001"; -- 0.028984600917169274
	pesos_i(22833) := b"1111111111111111_1111111111111111_1110111000001000_0111010110001111"; -- -0.07018342276162867
	pesos_i(22834) := b"0000000000000000_0000000000000000_0001101001110000_1001101010001101"; -- 0.1032806962698009
	pesos_i(22835) := b"1111111111111111_1111111111111111_1110110111010001_1100000101110110"; -- -0.07101813191619906
	pesos_i(22836) := b"0000000000000000_0000000000000000_0000100111101000_1101000111110011"; -- 0.03870880303446619
	pesos_i(22837) := b"1111111111111111_1111111111111111_1111001011000110_0111111011101100"; -- -0.05165869466381543
	pesos_i(22838) := b"0000000000000000_0000000000000000_0000011100010100_1101011011000101"; -- 0.027661726972480642
	pesos_i(22839) := b"1111111111111111_1111111111111111_1111011011111011_0110110101000010"; -- -0.03522603178621184
	pesos_i(22840) := b"0000000000000000_0000000000000000_0001100001001100_1001101101000100"; -- 0.09491892261161726
	pesos_i(22841) := b"0000000000000000_0000000000000000_0001000000011011_1100001100101100"; -- 0.06292362056716909
	pesos_i(22842) := b"1111111111111111_1111111111111111_1101111100100011_0011101110111000"; -- -0.1283686329605681
	pesos_i(22843) := b"0000000000000000_0000000000000000_0001110110100000_0011010110011011"; -- 0.11572585144488767
	pesos_i(22844) := b"0000000000000000_0000000000000000_0000111110101110_0110111011010101"; -- 0.06125538542554285
	pesos_i(22845) := b"0000000000000000_0000000000000000_0001111100101100_1010110110101110"; -- 0.12177548884836524
	pesos_i(22846) := b"1111111111111111_1111111111111111_1101101110001100_0011011001001001"; -- -0.1423917839227811
	pesos_i(22847) := b"1111111111111111_1111111111111111_1111111000010011_1101010111011100"; -- -0.007509835957656538
	pesos_i(22848) := b"1111111111111111_1111111111111111_1110010110110101_0000010000001010"; -- -0.10270666838015785
	pesos_i(22849) := b"0000000000000000_0000000000000000_0000000010101001_1010100011100001"; -- 0.002588801214207732
	pesos_i(22850) := b"0000000000000000_0000000000000000_0010010011111111_0110110011100101"; -- 0.14452248190519917
	pesos_i(22851) := b"1111111111111111_1111111111111111_1101110110111100_0010010101101000"; -- -0.13384786807704838
	pesos_i(22852) := b"0000000000000000_0000000000000000_0000111010100101_0010001000111100"; -- 0.057207240620191745
	pesos_i(22853) := b"1111111111111111_1111111111111111_1101111100101010_0000101010001001"; -- -0.1282647529871176
	pesos_i(22854) := b"0000000000000000_0000000000000000_0001011111011110_0100100011011111"; -- 0.09323554467872949
	pesos_i(22855) := b"0000000000000000_0000000000000000_0001111010110000_1111010111100010"; -- 0.11988770252758647
	pesos_i(22856) := b"0000000000000000_0000000000000000_0000110001100001_0101010010010100"; -- 0.04836014375256651
	pesos_i(22857) := b"1111111111111111_1111111111111111_1101111100011111_1011010000101110"; -- -0.12842248793578792
	pesos_i(22858) := b"1111111111111111_1111111111111111_1111011000111011_0001110010101110"; -- -0.038160522001669285
	pesos_i(22859) := b"1111111111111111_1111111111111111_1101100100001100_0010110100010011"; -- -0.15215795786684666
	pesos_i(22860) := b"0000000000000000_0000000000000000_0010000001010011_0001000011101111"; -- 0.12626748882872227
	pesos_i(22861) := b"1111111111111111_1111111111111111_1110011101101010_0101010010001110"; -- -0.09603377860514273
	pesos_i(22862) := b"1111111111111111_1111111111111111_1110110100101101_1110110111001111"; -- -0.0735179299970866
	pesos_i(22863) := b"0000000000000000_0000000000000000_0001101111100111_1110101011010000"; -- 0.10900752613089472
	pesos_i(22864) := b"0000000000000000_0000000000000000_0001111011001111_1010001100111000"; -- 0.12035579793198785
	pesos_i(22865) := b"0000000000000000_0000000000000000_0000111011111100_0101011111110100"; -- 0.0585379573153263
	pesos_i(22866) := b"1111111111111111_1111111111111111_1111111011110010_1000001110110101"; -- -0.004112022686248337
	pesos_i(22867) := b"0000000000000000_0000000000000000_0010000010110010_0001011010100001"; -- 0.12771741334688297
	pesos_i(22868) := b"0000000000000000_0000000000000000_0000110011010111_1110100110101111"; -- 0.05016956825159849
	pesos_i(22869) := b"1111111111111111_1111111111111111_1110111010000101_0111100100110001"; -- -0.06827585738795279
	pesos_i(22870) := b"0000000000000000_0000000000000000_0000000100000110_0110101110101111"; -- 0.004004221221652444
	pesos_i(22871) := b"0000000000000000_0000000000000000_0000011001100000_0000100001011101"; -- 0.024902842210114844
	pesos_i(22872) := b"0000000000000000_0000000000000000_0000011001111101_0100100011001010"; -- 0.02534918715121935
	pesos_i(22873) := b"0000000000000000_0000000000000000_0000110010010011_0011100100101011"; -- 0.0491214494252905
	pesos_i(22874) := b"0000000000000000_0000000000000000_0010100001010010_0011001101011100"; -- 0.15750428204117642
	pesos_i(22875) := b"1111111111111111_1111111111111111_1110110010010111_0100100101000111"; -- -0.07581655525101183
	pesos_i(22876) := b"1111111111111111_1111111111111111_1111100111101111_0011001100101100"; -- -0.023693849221247464
	pesos_i(22877) := b"0000000000000000_0000000000000000_0001101111111000_1110110000001111"; -- 0.10926699991639754
	pesos_i(22878) := b"0000000000000000_0000000000000000_0000111000001110_0010011110010011"; -- 0.054903481745604554
	pesos_i(22879) := b"0000000000000000_0000000000000000_0000100010111011_1001110101011111"; -- 0.03411277354970635
	pesos_i(22880) := b"0000000000000000_0000000000000000_0000100101010001_1110100111010110"; -- 0.0364061497278439
	pesos_i(22881) := b"0000000000000000_0000000000000000_0000011001101100_1101110101101100"; -- 0.025098647016629755
	pesos_i(22882) := b"1111111111111111_1111111111111111_1110011011011000_0100101111011001"; -- -0.098262080575901
	pesos_i(22883) := b"1111111111111111_1111111111111111_1110111000101110_1001001000000010"; -- -0.06960189301804176
	pesos_i(22884) := b"1111111111111111_1111111111111111_1111110010100011_0111011111011011"; -- -0.013130673428380056
	pesos_i(22885) := b"1111111111111111_1111111111111111_1101011111111101_1110110011001000"; -- -0.15628166300492302
	pesos_i(22886) := b"1111111111111111_1111111111111111_1101101101010111_0011100011000001"; -- -0.14320035247835958
	pesos_i(22887) := b"1111111111111111_1111111111111111_1110101011100111_1100100010001100"; -- -0.08240076622782898
	pesos_i(22888) := b"1111111111111111_1111111111111111_1110111000010110_1001000011010110"; -- -0.06996817365875581
	pesos_i(22889) := b"0000000000000000_0000000000000000_0001101010010110_0010011011101111"; -- 0.10385363890739348
	pesos_i(22890) := b"1111111111111111_1111111111111111_1111010101001010_1011101100000111"; -- -0.04182845200227595
	pesos_i(22891) := b"1111111111111111_1111111111111111_1101100111010111_0111000010010011"; -- -0.14905640037532158
	pesos_i(22892) := b"0000000000000000_0000000000000000_0001010001001110_1101111001100000"; -- 0.07932844010042062
	pesos_i(22893) := b"1111111111111111_1111111111111111_1111000100000010_0110110111111110"; -- -0.0585566764073866
	pesos_i(22894) := b"1111111111111111_1111111111111111_1101100111001101_1110000010111011"; -- -0.14920230322893327
	pesos_i(22895) := b"0000000000000000_0000000000000000_0001010000101101_0010001001010010"; -- 0.07881369119832349
	pesos_i(22896) := b"1111111111111111_1111111111111111_1110010000010111_0000100100110100"; -- -0.1090234993199875
	pesos_i(22897) := b"1111111111111111_1111111111111111_1111110000011011_1010001011100000"; -- -0.015203304686854872
	pesos_i(22898) := b"1111111111111111_1111111111111111_1111000111010000_0101011000011101"; -- -0.055414789063082774
	pesos_i(22899) := b"0000000000000000_0000000000000000_0000010101010101_1101111111101010"; -- 0.020841593504515178
	pesos_i(22900) := b"1111111111111111_1111111111111111_1110000111101100_1110111010010111"; -- -0.1174784547862269
	pesos_i(22901) := b"0000000000000000_0000000000000000_0000100101101010_0010100111111001"; -- 0.0367761834374305
	pesos_i(22902) := b"1111111111111111_1111111111111111_1111010011011101_1110100000010001"; -- -0.04348897532839967
	pesos_i(22903) := b"1111111111111111_1111111111111111_1110000110100001_0101101110110010"; -- -0.118631619508095
	pesos_i(22904) := b"1111111111111111_1111111111111111_1111011101111011_1011110000000110"; -- -0.033268211875926844
	pesos_i(22905) := b"0000000000000000_0000000000000000_0001011000010100_1111010000001111"; -- 0.08625722288957491
	pesos_i(22906) := b"0000000000000000_0000000000000000_0001101010011111_0000011101001111"; -- 0.10398908310108843
	pesos_i(22907) := b"1111111111111111_1111111111111111_1111111101010111_0110010110110101"; -- -0.002572673121553485
	pesos_i(22908) := b"0000000000000000_0000000000000000_0001100100010100_0000000001001000"; -- 0.09796144244602299
	pesos_i(22909) := b"0000000000000000_0000000000000000_0000100111100001_1000011001100101"; -- 0.038597488067478467
	pesos_i(22910) := b"0000000000000000_0000000000000000_0000001000011000_1110000000011101"; -- 0.008192069241271544
	pesos_i(22911) := b"1111111111111111_1111111111111111_1101110001000101_0100101110101001"; -- -0.1395676337721112
	pesos_i(22912) := b"1111111111111111_1111111111111111_1110000100101010_0101101011001011"; -- -0.12044746910608196
	pesos_i(22913) := b"1111111111111111_1111111111111111_1101100010110010_1110001011111110"; -- -0.15352040585583923
	pesos_i(22914) := b"0000000000000000_0000000000000000_0000001100100010_1100001110000111"; -- 0.012249203282253412
	pesos_i(22915) := b"1111111111111111_1111111111111111_1111000111100111_0010101000100100"; -- -0.05506645798216931
	pesos_i(22916) := b"1111111111111111_1111111111111111_1101111001101101_1100011011101001"; -- -0.13113743596255065
	pesos_i(22917) := b"0000000000000000_0000000000000000_0000100011101011_1101111010011000"; -- 0.03484908294449474
	pesos_i(22918) := b"0000000000000000_0000000000000000_0001110110000110_1011110100011011"; -- 0.11533719923752811
	pesos_i(22919) := b"1111111111111111_1111111111111111_1111110111110010_0001110011110100"; -- -0.00802439739223114
	pesos_i(22920) := b"0000000000000000_0000000000000000_0010010110010010_1001100000111100"; -- 0.14676810707092713
	pesos_i(22921) := b"0000000000000000_0000000000000000_0001101000001011_1111100100010011"; -- 0.10174519256794967
	pesos_i(22922) := b"1111111111111111_1111111111111111_1111010101101001_1111010001000101"; -- -0.04135201757302252
	pesos_i(22923) := b"1111111111111111_1111111111111111_1101110111010100_0101100001101010"; -- -0.13347861682716847
	pesos_i(22924) := b"1111111111111111_1111111111111111_1110110100101010_0000010000010010"; -- -0.07357763822471862
	pesos_i(22925) := b"1111111111111111_1111111111111111_1110000001010011_1101010000110011"; -- -0.12372087238565053
	pesos_i(22926) := b"1111111111111111_1111111111111111_1111110110000101_0101011101001100"; -- -0.009684127703793637
	pesos_i(22927) := b"1111111111111111_1111111111111111_1111001001111101_1000100111011110"; -- -0.05277193395665538
	pesos_i(22928) := b"1111111111111111_1111111111111111_1101110100001010_0000011101101110"; -- -0.13656571935453876
	pesos_i(22929) := b"1111111111111111_1111111111111111_1101111000100100_0111111110110010"; -- -0.13225557237610075
	pesos_i(22930) := b"0000000000000000_0000000000000000_0000100000110000_0011101001101000"; -- 0.03198590314313787
	pesos_i(22931) := b"1111111111111111_1111111111111111_1111000111010100_1000010000111001"; -- -0.055351005660183694
	pesos_i(22932) := b"0000000000000000_0000000000000000_0001110010010001_1111110101100010"; -- 0.11160262718768726
	pesos_i(22933) := b"1111111111111111_1111111111111111_1110111111001011_0100101111010011"; -- -0.06330419644504659
	pesos_i(22934) := b"0000000000000000_0000000000000000_0000011000110101_0101000110011100"; -- 0.024251080007591214
	pesos_i(22935) := b"1111111111111111_1111111111111111_1101100110011100_0100000111000111"; -- -0.14995945815703668
	pesos_i(22936) := b"1111111111111111_1111111111111111_1111011110110001_1001111100010100"; -- -0.032445962567576175
	pesos_i(22937) := b"0000000000000000_0000000000000000_0000001001111010_1110110001111111"; -- 0.00968816845334391
	pesos_i(22938) := b"0000000000000000_0000000000000000_0001110101101101_1101010100000101"; -- 0.11495715499918635
	pesos_i(22939) := b"0000000000000000_0000000000000000_0000011100100001_0001011101100010"; -- 0.027848683672753644
	pesos_i(22940) := b"0000000000000000_0000000000000000_0010001101000001_0011010100011000"; -- 0.13771373602787843
	pesos_i(22941) := b"0000000000000000_0000000000000000_0000000101101000_1101101000010010"; -- 0.005506162036489732
	pesos_i(22942) := b"1111111111111111_1111111111111111_1111000101010110_0101101111110110"; -- -0.057276012878769156
	pesos_i(22943) := b"0000000000000000_0000000000000000_0000000111110111_1011001101100101"; -- 0.007685863564441776
	pesos_i(22944) := b"0000000000000000_0000000000000000_0010000111001001_0101010110010111"; -- 0.1319783682140893
	pesos_i(22945) := b"1111111111111111_1111111111111111_1101111100110000_1101011011010100"; -- -0.1281610234680878
	pesos_i(22946) := b"0000000000000000_0000000000000000_0000010010010010_1111111110111110"; -- 0.01786802657104602
	pesos_i(22947) := b"0000000000000000_0000000000000000_0010000101101110_1110011010011111"; -- 0.13059846298779923
	pesos_i(22948) := b"0000000000000000_0000000000000000_0001000111001010_0010011111000110"; -- 0.0694908961422351
	pesos_i(22949) := b"1111111111111111_1111111111111111_1111010110010001_1111101110001001"; -- -0.04074123296650979
	pesos_i(22950) := b"1111111111111111_1111111111111111_1101011100101111_1001110101101010"; -- -0.1594297043280771
	pesos_i(22951) := b"1111111111111111_1111111111111111_1110110011010111_1100001110101100"; -- -0.07483269739052997
	pesos_i(22952) := b"1111111111111111_1111111111111111_1110100000010101_0011101001110011"; -- -0.09342608156470579
	pesos_i(22953) := b"1111111111111111_1111111111111111_1110010110010000_1101010100110010"; -- -0.10325877695020087
	pesos_i(22954) := b"1111111111111111_1111111111111111_1110000111100110_0001000001110010"; -- -0.11758324825091493
	pesos_i(22955) := b"0000000000000000_0000000000000000_0001010101010010_0000101001010110"; -- 0.08328308680146869
	pesos_i(22956) := b"1111111111111111_1111111111111111_1110101100011110_0000011101011101"; -- -0.08157304733353322
	pesos_i(22957) := b"1111111111111111_1111111111111111_1101110011100101_1011001001111100"; -- -0.13712009891988697
	pesos_i(22958) := b"0000000000000000_0000000000000000_0000010000111100_0110110011101000"; -- 0.01654701874114522
	pesos_i(22959) := b"1111111111111111_1111111111111111_1101110010101000_0001010000110100"; -- -0.13806031924152692
	pesos_i(22960) := b"1111111111111111_1111111111111111_1110101010000010_0111010110010101"; -- -0.08394684891336789
	pesos_i(22961) := b"1111111111111111_1111111111111111_1111000001111101_1101110100000010"; -- -0.06057947825168262
	pesos_i(22962) := b"1111111111111111_1111111111111111_1111100000110111_0001110110001101"; -- -0.030409005124513833
	pesos_i(22963) := b"1111111111111111_1111111111111111_1101011001101111_1000101100110100"; -- -0.1623604771780962
	pesos_i(22964) := b"0000000000000000_0000000000000000_0010011001001010_0110110011011010"; -- 0.14957313848734582
	pesos_i(22965) := b"1111111111111111_1111111111111111_1111010010111011_0100111010101110"; -- -0.04401691667951099
	pesos_i(22966) := b"1111111111111111_1111111111111111_1110000100001011_1001010011111100"; -- -0.12091702306189131
	pesos_i(22967) := b"0000000000000000_0000000000000000_0001110110000000_0101010011011001"; -- 0.11523943236718569
	pesos_i(22968) := b"0000000000000000_0000000000000000_0000101101000001_0011001000100011"; -- 0.043963559563232106
	pesos_i(22969) := b"1111111111111111_1111111111111111_1111010011000111_1110100100001011"; -- -0.043824610644572215
	pesos_i(22970) := b"1111111111111111_1111111111111111_1110011011111101_0110000100101100"; -- -0.09769623455063801
	pesos_i(22971) := b"1111111111111111_1111111111111111_1111000011001101_0011100110001100"; -- -0.05936851811624403
	pesos_i(22972) := b"1111111111111111_1111111111111111_1110001110011001_1111010100110001"; -- -0.1109320408047817
	pesos_i(22973) := b"1111111111111111_1111111111111111_1111010111101011_0011001101100111"; -- -0.03937987085348649
	pesos_i(22974) := b"1111111111111111_1111111111111111_1110011011100000_1000110011110001"; -- -0.09813613038615195
	pesos_i(22975) := b"0000000000000000_0000000000000000_0001011001011010_0101101010000100"; -- 0.08731618623087331
	pesos_i(22976) := b"0000000000000000_0000000000000000_0001100111000100_0001000100010001"; -- 0.10064798983366913
	pesos_i(22977) := b"0000000000000000_0000000000000000_0000001011011000_0001000001101010"; -- 0.011109376731937516
	pesos_i(22978) := b"1111111111111111_1111111111111111_1110100001110010_1110111111011000"; -- -0.09199620226094465
	pesos_i(22979) := b"1111111111111111_1111111111111111_1110101000101101_1111101000000010"; -- -0.08523595291983464
	pesos_i(22980) := b"1111111111111111_1111111111111111_1111110111000001_1111000011101110"; -- -0.008759443231740967
	pesos_i(22981) := b"0000000000000000_0000000000000000_0001001101110001_0011101001100101"; -- 0.07594647371427923
	pesos_i(22982) := b"1111111111111111_1111111111111111_1111101111001110_1110010010001010"; -- -0.016374317517413795
	pesos_i(22983) := b"0000000000000000_0000000000000000_0000000101011110_1111100011010100"; -- 0.00535540749041025
	pesos_i(22984) := b"1111111111111111_1111111111111111_1111101110001000_1000011100101100"; -- -0.017447997802799462
	pesos_i(22985) := b"0000000000000000_0000000000000000_0010010011000100_1110110010100000"; -- 0.14362982669788968
	pesos_i(22986) := b"1111111111111111_1111111111111111_1111111000110100_1010101000011101"; -- -0.00700890350725869
	pesos_i(22987) := b"1111111111111111_1111111111111111_1111001011110001_1011010011000010"; -- -0.050999357904946425
	pesos_i(22988) := b"0000000000000000_0000000000000000_0000111001000101_0111100111010001"; -- 0.05574761720309377
	pesos_i(22989) := b"0000000000000000_0000000000000000_0000101100110000_0100011101111100"; -- 0.04370543272689922
	pesos_i(22990) := b"0000000000000000_0000000000000000_0000100111000000_1111101111100111"; -- 0.03810095195865837
	pesos_i(22991) := b"0000000000000000_0000000000000000_0001011000011111_1011111010001101"; -- 0.08642188013692861
	pesos_i(22992) := b"1111111111111111_1111111111111111_1110011100100110_1001101010101111"; -- -0.09706719611565237
	pesos_i(22993) := b"1111111111111111_1111111111111111_1110000100100111_0011001010110010"; -- -0.1204956356283591
	pesos_i(22994) := b"0000000000000000_0000000000000000_0000010110111010_0101000111011101"; -- 0.022374264313469016
	pesos_i(22995) := b"0000000000000000_0000000000000000_0001010111101101_0110001101110010"; -- 0.08565351033989364
	pesos_i(22996) := b"1111111111111111_1111111111111111_1110001110010111_1111111001011101"; -- -0.11096201162969882
	pesos_i(22997) := b"1111111111111111_1111111111111111_1110011011000000_0010100111010000"; -- -0.0986303203244037
	pesos_i(22998) := b"0000000000000000_0000000000000000_0010010100001101_0001001001011100"; -- 0.14473070867083673
	pesos_i(22999) := b"1111111111111111_1111111111111111_1101110100110111_1011110100110011"; -- -0.13586823947836152
	pesos_i(23000) := b"0000000000000000_0000000000000000_0000101000111001_1011100011101010"; -- 0.039943272655492655
	pesos_i(23001) := b"0000000000000000_0000000000000000_0000100011100110_0111100111111100"; -- 0.03476679241235121
	pesos_i(23002) := b"1111111111111111_1111111111111111_1111100001001100_0010111111111011"; -- -0.030087472256988917
	pesos_i(23003) := b"1111111111111111_1111111111111111_1111001001011011_1110111101000001"; -- -0.05328468964106879
	pesos_i(23004) := b"1111111111111111_1111111111111111_1111000110111001_1011010000111010"; -- -0.05576013159710361
	pesos_i(23005) := b"0000000000000000_0000000000000000_0001010101010111_1100110000100101"; -- 0.08337093266524728
	pesos_i(23006) := b"1111111111111111_1111111111111111_1111010110010111_1110101101010001"; -- -0.04065064695172844
	pesos_i(23007) := b"0000000000000000_0000000000000000_0001010100100000_1010110011111111"; -- 0.08252984253272386
	pesos_i(23008) := b"1111111111111111_1111111111111111_1111111101101000_0101011000111010"; -- -0.0023141963462789093
	pesos_i(23009) := b"1111111111111111_1111111111111111_1110001101100011_0000000110111011"; -- -0.1117705266966382
	pesos_i(23010) := b"1111111111111111_1111111111111111_1110010010000100_0011101000001010"; -- -0.10735738043692485
	pesos_i(23011) := b"0000000000000000_0000000000000000_0000001011000101_0111011110101001"; -- 0.01082561365528663
	pesos_i(23012) := b"1111111111111111_1111111111111111_1101111110011001_0100001111111000"; -- -0.1265676040879472
	pesos_i(23013) := b"0000000000000000_0000000000000000_0001011010111001_0101110010001101"; -- 0.08876589248891543
	pesos_i(23014) := b"1111111111111111_1111111111111111_1101110111101100_0111010110011111"; -- -0.13311066503472505
	pesos_i(23015) := b"1111111111111111_1111111111111111_1110111011111001_1000000010110011"; -- -0.0665053905518846
	pesos_i(23016) := b"0000000000000000_0000000000000000_0001000011111100_0101100111011000"; -- 0.06635056992393018
	pesos_i(23017) := b"1111111111111111_1111111111111111_1110100010100111_0000001011010000"; -- -0.09120161460435011
	pesos_i(23018) := b"0000000000000000_0000000000000000_0000101001100110_0110111110011000"; -- 0.04062554807292372
	pesos_i(23019) := b"0000000000000000_0000000000000000_0010101000110001_1000001111011001"; -- 0.16481803938916523
	pesos_i(23020) := b"1111111111111111_1111111111111111_1101111100001000_0111111010000111"; -- -0.12877663815741655
	pesos_i(23021) := b"0000000000000000_0000000000000000_0000010010010100_0010110101010010"; -- 0.017886002164450066
	pesos_i(23022) := b"1111111111111111_1111111111111111_1101010010100100_0101010011101111"; -- -0.16936749619433825
	pesos_i(23023) := b"0000000000000000_0000000000000000_0000101011001000_1100101001000011"; -- 0.042126313481944615
	pesos_i(23024) := b"1111111111111111_1111111111111111_1110011110110000_1101111101000100"; -- -0.09495739552265053
	pesos_i(23025) := b"0000000000000000_0000000000000000_0010001001011100_1111101001000000"; -- 0.1342312246220703
	pesos_i(23026) := b"0000000000000000_0000000000000000_0000011101001110_0110011110101000"; -- 0.028540113829210866
	pesos_i(23027) := b"0000000000000000_0000000000000000_0010001000011001_0011110000011100"; -- 0.13319755241837508
	pesos_i(23028) := b"1111111111111111_1111111111111111_1101101111101100_0100011010110101"; -- -0.14092596141207694
	pesos_i(23029) := b"0000000000000000_0000000000000000_0000000011111101_0000100110001001"; -- 0.0038610418900443945
	pesos_i(23030) := b"1111111111111111_1111111111111111_1111101010011100_0000111001111011"; -- -0.02105626582220673
	pesos_i(23031) := b"0000000000000000_0000000000000000_0001010010111101_0111110111101010"; -- 0.08101641618360018
	pesos_i(23032) := b"1111111111111111_1111111111111111_1110011011101101_0100001010001011"; -- -0.09794220077154674
	pesos_i(23033) := b"0000000000000000_0000000000000000_0001001000111001_1100000010010011"; -- 0.07119372933019237
	pesos_i(23034) := b"0000000000000000_0000000000000000_0001110111011011_1010011011011001"; -- 0.11663286972262539
	pesos_i(23035) := b"0000000000000000_0000000000000000_0001010100111111_0100001000001011"; -- 0.08299649027686333
	pesos_i(23036) := b"1111111111111111_1111111111111111_1111100101101010_1100011100001011"; -- -0.025714454381181816
	pesos_i(23037) := b"1111111111111111_1111111111111111_1111110101001010_0101101001000100"; -- -0.010584219262274779
	pesos_i(23038) := b"0000000000000000_0000000000000000_0001111001001011_0110110111000001"; -- 0.11833845105607975
	pesos_i(23039) := b"1111111111111111_1111111111111111_1101110111111101_1000000000010101"; -- -0.13285064208935518
	pesos_i(23040) := b"0000000000000000_0000000000000000_0010000001111000_0111101010101100"; -- 0.1268383665901751
	pesos_i(23041) := b"1111111111111111_1111111111111111_1111011110011101_1001110111110000"; -- -0.03275120633973861
	pesos_i(23042) := b"1111111111111111_1111111111111111_1111110101111000_0001001110001110"; -- -0.009886529850758302
	pesos_i(23043) := b"1111111111111111_1111111111111111_1111111001001111_0001000110101100"; -- -0.0066060024127561935
	pesos_i(23044) := b"1111111111111111_1111111111111111_1110011100011010_1000010101001101"; -- -0.09725157618507276
	pesos_i(23045) := b"0000000000000000_0000000000000000_0001101001111001_0110101100111110"; -- 0.10341520553202145
	pesos_i(23046) := b"1111111111111111_1111111111111111_1111010110000100_0010100000111010"; -- -0.04095219204789897
	pesos_i(23047) := b"1111111111111111_1111111111111111_1111100000111100_0100101101101011"; -- -0.030329977352076945
	pesos_i(23048) := b"0000000000000000_0000000000000000_0000000111101010_0011101001101011"; -- 0.007480288525752416
	pesos_i(23049) := b"0000000000000000_0000000000000000_0001010011011000_1011110111110011"; -- 0.08143222034448991
	pesos_i(23050) := b"1111111111111111_1111111111111111_1111010111111000_1010100010110001"; -- -0.0391745154490509
	pesos_i(23051) := b"0000000000000000_0000000000000000_0000000100000011_1101000110100101"; -- 0.003964522075945829
	pesos_i(23052) := b"0000000000000000_0000000000000000_0010000101010100_1000000010110001"; -- 0.1301956587981242
	pesos_i(23053) := b"0000000000000000_0000000000000000_0010001101110010_0000100101111010"; -- 0.13845881670371565
	pesos_i(23054) := b"0000000000000000_0000000000000000_0001101001001000_1100010110100100"; -- 0.10267291308492944
	pesos_i(23055) := b"1111111111111111_1111111111111111_1111110100100111_1010011000100111"; -- -0.011113753802560883
	pesos_i(23056) := b"0000000000000000_0000000000000000_0001011100110000_1001011111010001"; -- 0.09058522072643084
	pesos_i(23057) := b"0000000000000000_0000000000000000_0001111010000101_1110101000100100"; -- 0.11923087473286732
	pesos_i(23058) := b"1111111111111111_1111111111111111_1111011001110011_0001000100001000"; -- -0.037306724131064756
	pesos_i(23059) := b"1111111111111111_1111111111111111_1110001111110000_0010010010101111"; -- -0.10961695411941189
	pesos_i(23060) := b"1111111111111111_1111111111111111_1111111011001100_1111000011011100"; -- -0.0046853506143401565
	pesos_i(23061) := b"0000000000000000_0000000000000000_0000110111110110_0001011111101001"; -- 0.05453633726663361
	pesos_i(23062) := b"0000000000000000_0000000000000000_0010111110011110_0010101100111010"; -- 0.18600721522626126
	pesos_i(23063) := b"0000000000000000_0000000000000000_0000100011110110_0000101001101001"; -- 0.035004282656843244
	pesos_i(23064) := b"0000000000000000_0000000000000000_0000110101011010_0010101111011110"; -- 0.05215715580308592
	pesos_i(23065) := b"0000000000000000_0000000000000000_0000000001000001_1001011111111010"; -- 0.0010008797677697
	pesos_i(23066) := b"1111111111111111_1111111111111111_1111110001100011_0100101101001101"; -- -0.01410989160890047
	pesos_i(23067) := b"1111111111111111_1111111111111111_1101111111101110_0100000011100000"; -- -0.12527079139540917
	pesos_i(23068) := b"1111111111111111_1111111111111111_1101110000110000_1110011000111010"; -- -0.13987885547685017
	pesos_i(23069) := b"1111111111111111_1111111111111111_1110111011010111_0010111001001011"; -- -0.06702910114235389
	pesos_i(23070) := b"1111111111111111_1111111111111111_1101101111011000_1111001100101010"; -- -0.14122085775002208
	pesos_i(23071) := b"0000000000000000_0000000000000000_0001101011110010_1011101011001110"; -- 0.1052662613219513
	pesos_i(23072) := b"1111111111111111_1111111111111111_1111100000000001_0100101101001101"; -- -0.031230252935718936
	pesos_i(23073) := b"0000000000000000_0000000000000000_0000100110111011_0101100100001001"; -- 0.038014950488074316
	pesos_i(23074) := b"0000000000000000_0000000000000000_0001001110101100_1101000010101001"; -- 0.07685569894729169
	pesos_i(23075) := b"0000000000000000_0000000000000000_0001000011010010_1001011100101111"; -- 0.06571335686198754
	pesos_i(23076) := b"0000000000000000_0000000000000000_0010000110001010_1001000111101101"; -- 0.1310206607044847
	pesos_i(23077) := b"1111111111111111_1111111111111111_1110011010111011_1110010000101010"; -- -0.09869550690063468
	pesos_i(23078) := b"0000000000000000_0000000000000000_0001000010101011_1100010001011111"; -- 0.06512095746267031
	pesos_i(23079) := b"0000000000000000_0000000000000000_0000011010111101_1000001101110111"; -- 0.026329247036835538
	pesos_i(23080) := b"1111111111111111_1111111111111111_1111101010001010_1100001111110101"; -- -0.021320107073407202
	pesos_i(23081) := b"0000000000000000_0000000000000000_0001001000000011_0100000000011111"; -- 0.07036209819453022
	pesos_i(23082) := b"0000000000000000_0000000000000000_0000100100000011_0011001010010000"; -- 0.035205040188485685
	pesos_i(23083) := b"1111111111111111_1111111111111111_1110110011001011_1101000001001001"; -- -0.07501505116270432
	pesos_i(23084) := b"0000000000000000_0000000000000000_0010001011010100_0111100010000001"; -- 0.13605454592103727
	pesos_i(23085) := b"0000000000000000_0000000000000000_0000000010100110_0000010010001001"; -- 0.002533229190037479
	pesos_i(23086) := b"0000000000000000_0000000000000000_0000011111011010_0000011011011110"; -- 0.03067057536519144
	pesos_i(23087) := b"1111111111111111_1111111111111111_1111001001100100_0110011011001000"; -- -0.053155494959441135
	pesos_i(23088) := b"0000000000000000_0000000000000000_0000110000010010_0111011101000110"; -- 0.04715676756449374
	pesos_i(23089) := b"1111111111111111_1111111111111111_1111000100000010_1000001000000111"; -- -0.0585554822261073
	pesos_i(23090) := b"0000000000000000_0000000000000000_0001011001111101_1111000001011110"; -- 0.08785917551935804
	pesos_i(23091) := b"0000000000000000_0000000000000000_0001000010011000_0100011000100100"; -- 0.06482351667611869
	pesos_i(23092) := b"0000000000000000_0000000000000000_0010100001000100_1011001000101000"; -- 0.15729821670023855
	pesos_i(23093) := b"0000000000000000_0000000000000000_0010000111001000_1010001101010001"; -- 0.1319677422234779
	pesos_i(23094) := b"1111111111111111_1111111111111111_1111000000101011_0110101111011000"; -- -0.06183744400444486
	pesos_i(23095) := b"1111111111111111_1111111111111111_1111001001110100_0000110111011111"; -- -0.05291665364137731
	pesos_i(23096) := b"0000000000000000_0000000000000000_0000000101111010_0111001111001101"; -- 0.00577472445792392
	pesos_i(23097) := b"1111111111111111_1111111111111111_1111001111101111_1111110010110011"; -- -0.04711933739780027
	pesos_i(23098) := b"0000000000000000_0000000000000000_0000100001100000_0010110110101100"; -- 0.03271756603747779
	pesos_i(23099) := b"1111111111111111_1111111111111111_1110110011100011_0000011101011000"; -- -0.0746608172710253
	pesos_i(23100) := b"0000000000000000_0000000000000000_0000100110010111_0110110111111000"; -- 0.03746688181426637
	pesos_i(23101) := b"1111111111111111_1111111111111111_1111110010011110_0100110000100111"; -- -0.013209572262890863
	pesos_i(23102) := b"1111111111111111_1111111111111111_1110001111100100_0110001000011001"; -- -0.10979639892644055
	pesos_i(23103) := b"0000000000000000_0000000000000000_0001010111110111_0110111001100001"; -- 0.08580674997059015
	pesos_i(23104) := b"0000000000000000_0000000000000000_0001100001001100_1111111011001101"; -- 0.09492485520751434
	pesos_i(23105) := b"1111111111111111_1111111111111111_1110101001010010_0111101001100100"; -- -0.0846789843539053
	pesos_i(23106) := b"1111111111111111_1111111111111111_1101101001110000_0000100110011111"; -- -0.14672794223099922
	pesos_i(23107) := b"0000000000000000_0000000000000000_0000101011101011_0001010010101110"; -- 0.042649547965148554
	pesos_i(23108) := b"0000000000000000_0000000000000000_0001001000010111_0101100011101001"; -- 0.07066875158101384
	pesos_i(23109) := b"1111111111111111_1111111111111111_1101111101101100_1010100000101101"; -- -0.12724827673718148
	pesos_i(23110) := b"0000000000000000_0000000000000000_0000010110110110_0100011010010100"; -- 0.022312556316340666
	pesos_i(23111) := b"1111111111111111_1111111111111111_1110001001011000_0111100110001000"; -- -0.11583748265421574
	pesos_i(23112) := b"0000000000000000_0000000000000000_0000000011101001_1110110011110100"; -- 0.0035694214740786202
	pesos_i(23113) := b"1111111111111111_1111111111111111_1111001111111101_0010011111011011"; -- -0.046918400896024684
	pesos_i(23114) := b"0000000000000000_0000000000000000_0001101110101011_0011111101101010"; -- 0.1080817828146916
	pesos_i(23115) := b"1111111111111111_1111111111111111_1111001101110101_1101001111011101"; -- -0.048983343692077116
	pesos_i(23116) := b"0000000000000000_0000000000000000_0001011001110111_0010111001110111"; -- 0.08775606535483299
	pesos_i(23117) := b"0000000000000000_0000000000000000_0001101000010011_1000001110110110"; -- 0.10186026767643393
	pesos_i(23118) := b"0000000000000000_0000000000000000_0001011110111000_0100000010111101"; -- 0.09265522599523628
	pesos_i(23119) := b"1111111111111111_1111111111111111_1110001110101011_1111010001001100"; -- -0.11065743586212795
	pesos_i(23120) := b"1111111111111111_1111111111111111_1111010101110010_1000000001010110"; -- -0.04122159853257784
	pesos_i(23121) := b"1111111111111111_1111111111111111_1110011010001000_1110111101001111"; -- -0.09947304072338164
	pesos_i(23122) := b"1111111111111111_1111111111111111_1110011000000001_0000010000001000"; -- -0.10154700088114003
	pesos_i(23123) := b"1111111111111111_1111111111111111_1111101011011101_1001011000100011"; -- -0.020056358746964306
	pesos_i(23124) := b"1111111111111111_1111111111111111_1111111110010010_0000010001111110"; -- -0.0016781990475308922
	pesos_i(23125) := b"1111111111111111_1111111111111111_1101110101111001_1000111000010010"; -- -0.1348639684308042
	pesos_i(23126) := b"1111111111111111_1111111111111111_1111001111101101_0111101000011011"; -- -0.04715763884071192
	pesos_i(23127) := b"0000000000000000_0000000000000000_0000000100110111_1011010000010001"; -- 0.0047562162472441685
	pesos_i(23128) := b"0000000000000000_0000000000000000_0010001101100010_0101110111101111"; -- 0.13821971019853602
	pesos_i(23129) := b"0000000000000000_0000000000000000_0000001111100100_1000011000110101"; -- 0.015205753270058525
	pesos_i(23130) := b"0000000000000000_0000000000000000_0000011011101110_0111110101011011"; -- 0.027076563514323186
	pesos_i(23131) := b"0000000000000000_0000000000000000_0001001010101000_0011110000001101"; -- 0.07287955587913054
	pesos_i(23132) := b"0000000000000000_0000000000000000_0001001111000010_0011010101110010"; -- 0.07718214076858171
	pesos_i(23133) := b"0000000000000000_0000000000000000_0000010000011011_0001011100111000"; -- 0.016038371192832
	pesos_i(23134) := b"0000000000000000_0000000000000000_0000100111001001_1110110100100110"; -- 0.03823740185575191
	pesos_i(23135) := b"1111111111111111_1111111111111111_1111011011001010_0000111111011110"; -- -0.03597927882929777
	pesos_i(23136) := b"1111111111111111_1111111111111111_1111100100101011_1111111111110100"; -- -0.026672366100428096
	pesos_i(23137) := b"0000000000000000_0000000000000000_0000111110100011_1101010100001101"; -- 0.0610936314727768
	pesos_i(23138) := b"0000000000000000_0000000000000000_0000111010100010_1100001000000010"; -- 0.057170987503151624
	pesos_i(23139) := b"1111111111111111_1111111111111111_1110011011010110_0101010100111001"; -- -0.09829203958845247
	pesos_i(23140) := b"0000000000000000_0000000000000000_0001111010010100_0011010100010000"; -- 0.11944896348005815
	pesos_i(23141) := b"0000000000000000_0000000000000000_0000011001010010_0110000001000110"; -- 0.02469445913896768
	pesos_i(23142) := b"0000000000000000_0000000000000000_0000110000110010_1100110000001100"; -- 0.047650101695347544
	pesos_i(23143) := b"0000000000000000_0000000000000000_0000001001010001_0000000000100011"; -- 0.009048470075207453
	pesos_i(23144) := b"1111111111111111_1111111111111111_1101110001001011_0100010110101010"; -- -0.13947643846244606
	pesos_i(23145) := b"0000000000000000_0000000000000000_0001010010010001_0100010011000010"; -- 0.08034162259422035
	pesos_i(23146) := b"1111111111111111_1111111111111111_1111010101000111_1001110111101001"; -- -0.04187596387851098
	pesos_i(23147) := b"1111111111111111_1111111111111111_1111010100110100_0100101010010001"; -- -0.04217084846985673
	pesos_i(23148) := b"0000000000000000_0000000000000000_0001010110110001_1000110001011100"; -- 0.08474042163961558
	pesos_i(23149) := b"1111111111111111_1111111111111111_1101010100010110_0100000110110011"; -- -0.16762914056832195
	pesos_i(23150) := b"0000000000000000_0000000000000000_0010111001000111_0010100011001000"; -- 0.1807733047996619
	pesos_i(23151) := b"1111111111111111_1111111111111111_1110010111100111_0011110100011000"; -- -0.10194032816750712
	pesos_i(23152) := b"0000000000000000_0000000000000000_0010010110111000_0101111011100100"; -- 0.1473445230057912
	pesos_i(23153) := b"1111111111111111_1111111111111111_1111001001110101_0011101101011100"; -- -0.05289868355320439
	pesos_i(23154) := b"0000000000000000_0000000000000000_0000000001111100_0000001010011111"; -- 0.0018922460794179798
	pesos_i(23155) := b"0000000000000000_0000000000000000_0000101000010010_0100111010000001"; -- 0.039341837346450366
	pesos_i(23156) := b"1111111111111111_1111111111111111_1110010101000100_1011010011000101"; -- -0.1044203775346104
	pesos_i(23157) := b"1111111111111111_1111111111111111_1101100110101001_0100111001101000"; -- -0.14976034137459085
	pesos_i(23158) := b"0000000000000000_0000000000000000_0000011010000010_1001000110100001"; -- 0.02542982279314406
	pesos_i(23159) := b"0000000000000000_0000000000000000_0001111011000100_1110011111100000"; -- 0.1201920434091736
	pesos_i(23160) := b"0000000000000000_0000000000000000_0000101011001010_1111011001111001"; -- 0.04215946641860615
	pesos_i(23161) := b"1111111111111111_1111111111111111_1110110010010111_1111001101011001"; -- -0.07580641827592546
	pesos_i(23162) := b"1111111111111111_1111111111111111_1110010010011011_0100101100010011"; -- -0.10700541298493509
	pesos_i(23163) := b"1111111111111111_1111111111111111_1110001001100111_1010001011111011"; -- -0.1156061303471285
	pesos_i(23164) := b"0000000000000000_0000000000000000_0001111001101110_1000001000011001"; -- 0.11887372129386968
	pesos_i(23165) := b"1111111111111111_1111111111111111_1110000000110010_0011000000101110"; -- -0.12423418892208508
	pesos_i(23166) := b"0000000000000000_0000000000000000_0001011000011111_0100111001001111"; -- 0.08641519001540872
	pesos_i(23167) := b"0000000000000000_0000000000000000_0000001000100101_1100010001100111"; -- 0.008388781791209344
	pesos_i(23168) := b"1111111111111111_1111111111111111_1101100110110010_1101100011101101"; -- -0.14961475574979752
	pesos_i(23169) := b"1111111111111111_1111111111111111_1110111100101001_0110001000000001"; -- -0.06577479805441935
	pesos_i(23170) := b"1111111111111111_1111111111111111_1111011010000110_0101111010010000"; -- -0.03701218597286222
	pesos_i(23171) := b"1111111111111111_1111111111111111_1110110110010110_0101111110111011"; -- -0.07192422561322036
	pesos_i(23172) := b"1111111111111111_1111111111111111_1101110001001000_1100101000010100"; -- -0.1395143223789254
	pesos_i(23173) := b"0000000000000000_0000000000000000_0001111000101001_0100010111011001"; -- 0.11781727355968233
	pesos_i(23174) := b"0000000000000000_0000000000000000_0000001011101011_0100111011111101"; -- 0.011403023496222773
	pesos_i(23175) := b"1111111111111111_1111111111111111_1101110101111001_0010101010001110"; -- -0.1348699000449574
	pesos_i(23176) := b"1111111111111111_1111111111111111_1111110010000100_1100100010111100"; -- -0.013598875076935734
	pesos_i(23177) := b"0000000000000000_0000000000000000_0000110111000101_1001101110000010"; -- 0.05379650033144836
	pesos_i(23178) := b"1111111111111111_1111111111111111_1110011001100111_0100111000001101"; -- -0.0999861925421831
	pesos_i(23179) := b"0000000000000000_0000000000000000_0010000000011111_0110101001001010"; -- 0.1254793577246323
	pesos_i(23180) := b"0000000000000000_0000000000000000_0001010010001010_1011100110000110"; -- 0.08024177086260832
	pesos_i(23181) := b"0000000000000000_0000000000000000_0000011001111110_1110011001111011"; -- 0.02537384516281907
	pesos_i(23182) := b"1111111111111111_1111111111111111_1110100001001110_0101110101110011"; -- -0.0925542444148137
	pesos_i(23183) := b"1111111111111111_1111111111111111_1111111011100100_1001100000101101"; -- -0.0043244257625119535
	pesos_i(23184) := b"1111111111111111_1111111111111111_1110001010110111_0111100101001110"; -- -0.11438791123636738
	pesos_i(23185) := b"0000000000000000_0000000000000000_0001011100011110_1000111100010010"; -- 0.09031004137754925
	pesos_i(23186) := b"1111111111111111_1111111111111111_1110101011011001_1110010111111101"; -- -0.08261263429581274
	pesos_i(23187) := b"1111111111111111_1111111111111111_1110001111111111_0001011001001010"; -- -0.10938893018033119
	pesos_i(23188) := b"1111111111111111_1111111111111111_1110000101100111_0001011100111010"; -- -0.1195207102993264
	pesos_i(23189) := b"1111111111111111_1111111111111111_1101101111000110_0001001111011110"; -- -0.14150882551857866
	pesos_i(23190) := b"0000000000000000_0000000000000000_0001011100011011_1011010001010110"; -- 0.09026648606005724
	pesos_i(23191) := b"1111111111111111_1111111111111111_1111101010101101_1011000010100011"; -- -0.02078720112809444
	pesos_i(23192) := b"1111111111111111_1111111111111111_1110101101100110_1100001111110011"; -- -0.08046317408116793
	pesos_i(23193) := b"1111111111111111_1111111111111111_1110110010011001_1011100110011110"; -- -0.07577934165746673
	pesos_i(23194) := b"1111111111111111_1111111111111111_1111000000110000_0000111101001000"; -- -0.06176666739380972
	pesos_i(23195) := b"1111111111111111_1111111111111111_1111001100011111_1100011000010101"; -- -0.05029642087009877
	pesos_i(23196) := b"1111111111111111_1111111111111111_1101110100011000_1010101101110010"; -- -0.13634232006732358
	pesos_i(23197) := b"0000000000000000_0000000000000000_0000111101110001_1011000000101101"; -- 0.06032849409733778
	pesos_i(23198) := b"1111111111111111_1111111111111111_1111100000101001_1110111101010011"; -- -0.030610124733774426
	pesos_i(23199) := b"1111111111111111_1111111111111111_1110101111001110_0000010000011101"; -- -0.07888769426918851
	pesos_i(23200) := b"0000000000000000_0000000000000000_0001011111000110_1110010110111000"; -- 0.09287868245964676
	pesos_i(23201) := b"1111111111111111_1111111111111111_1110111001001100_0011011011100110"; -- -0.06914955974886185
	pesos_i(23202) := b"1111111111111111_1111111111111111_1101110110111101_1101001000001000"; -- -0.13382232009005357
	pesos_i(23203) := b"1111111111111111_1111111111111111_1101111000101000_1100100111111000"; -- -0.13219011005627343
	pesos_i(23204) := b"1111111111111111_1111111111111111_1111100110101111_1111101100011111"; -- -0.02465849387419158
	pesos_i(23205) := b"0000000000000000_0000000000000000_0010000100010011_0001000111001110"; -- 0.12919722813839918
	pesos_i(23206) := b"0000000000000000_0000000000000000_0001110000110111_0000000111001010"; -- 0.11021433993719931
	pesos_i(23207) := b"0000000000000000_0000000000000000_0000010001011000_0101000001000100"; -- 0.016972557543290443
	pesos_i(23208) := b"1111111111111111_1111111111111111_1111111000100100_1101000110001001"; -- -0.007250694386739524
	pesos_i(23209) := b"0000000000000000_0000000000000000_0000110111010011_1100011001111100"; -- 0.054012685023680035
	pesos_i(23210) := b"0000000000000000_0000000000000000_0001001101111110_1010110010010000"; -- 0.07615164304345091
	pesos_i(23211) := b"0000000000000000_0000000000000000_0001101101010101_1001111011011010"; -- 0.10677521535969386
	pesos_i(23212) := b"1111111111111111_1111111111111111_1110100101110100_0111000101111100"; -- -0.08806696633278334
	pesos_i(23213) := b"0000000000000000_0000000000000000_0000100010101101_1001001000010011"; -- 0.0338984772307711
	pesos_i(23214) := b"1111111111111111_1111111111111111_1110011100010011_0110100001011110"; -- -0.09736011232790734
	pesos_i(23215) := b"1111111111111111_1111111111111111_1110101111001011_0110010100011011"; -- -0.07892768946778715
	pesos_i(23216) := b"0000000000000000_0000000000000000_0001001101100010_0000010011100001"; -- 0.0757144021096058
	pesos_i(23217) := b"0000000000000000_0000000000000000_0000011110011110_0001000001110110"; -- 0.029755619737392137
	pesos_i(23218) := b"0000000000000000_0000000000000000_0000100110111010_1111000111111010"; -- 0.03800880757849994
	pesos_i(23219) := b"1111111111111111_1111111111111111_1110101110011010_0000011100000110"; -- -0.0796809778660476
	pesos_i(23220) := b"1111111111111111_1111111111111111_1111110111110010_1110110101001101"; -- -0.00801197876994442
	pesos_i(23221) := b"0000000000000000_0000000000000000_0000000101110000_0001101101110100"; -- 0.005616870773755438
	pesos_i(23222) := b"1111111111111111_1111111111111111_1110100010000011_1100000111011111"; -- -0.09173954299129386
	pesos_i(23223) := b"0000000000000000_0000000000000000_0000111110001111_0010110101100111"; -- 0.06077846305038199
	pesos_i(23224) := b"0000000000000000_0000000000000000_0001011111001100_1110111101110101"; -- 0.09297081581756422
	pesos_i(23225) := b"0000000000000000_0000000000000000_0000011010100001_0011100000111110"; -- 0.025897517230059466
	pesos_i(23226) := b"0000000000000000_0000000000000000_0010000010010100_0110100010110010"; -- 0.12726454109302412
	pesos_i(23227) := b"0000000000000000_0000000000000000_0001110011100101_1010011011111110"; -- 0.1128792162388056
	pesos_i(23228) := b"1111111111111111_1111111111111111_1111101001111001_0000000101100100"; -- -0.0215911035786897
	pesos_i(23229) := b"0000000000000000_0000000000000000_0000111010001111_1010110100101110"; -- 0.056879829142188434
	pesos_i(23230) := b"0000000000000000_0000000000000000_0001011100000000_1011100011111001"; -- 0.08985477511497056
	pesos_i(23231) := b"1111111111111111_1111111111111111_1110100010111011_1110011101011000"; -- -0.09088281726683452
	pesos_i(23232) := b"0000000000000000_0000000000000000_0000101000100011_1100110010101011"; -- 0.03960875688416228
	pesos_i(23233) := b"1111111111111111_1111111111111111_1101110001101000_1001110111001000"; -- -0.1390286814391968
	pesos_i(23234) := b"1111111111111111_1111111111111111_1111011010101101_0011010010001111"; -- -0.036419596818456454
	pesos_i(23235) := b"0000000000000000_0000000000000000_0000010001011000_0111000000111111"; -- 0.016974463821628264
	pesos_i(23236) := b"1111111111111111_1111111111111111_1110111111100101_1111110101010100"; -- -0.06289688775155615
	pesos_i(23237) := b"0000000000000000_0000000000000000_0000100111000011_0001000011001000"; -- 0.038132714000757816
	pesos_i(23238) := b"0000000000000000_0000000000000000_0000000101100111_0111101001000111"; -- 0.005485193503199285
	pesos_i(23239) := b"1111111111111111_1111111111111111_1110010111011001_0111111111001100"; -- -0.10214997539959846
	pesos_i(23240) := b"0000000000000000_0000000000000000_0001010011101110_1110111001110000"; -- 0.08177080374524444
	pesos_i(23241) := b"1111111111111111_1111111111111111_1110010000011111_1100111001110101"; -- -0.10888967171506637
	pesos_i(23242) := b"1111111111111111_1111111111111111_1111001000101000_0010011110010101"; -- -0.054074789183393174
	pesos_i(23243) := b"1111111111111111_1111111111111111_1111110000010111_0110111101001000"; -- -0.015267415016743377
	pesos_i(23244) := b"1111111111111111_1111111111111111_1110100111011101_1111110010010001"; -- -0.08645650358998269
	pesos_i(23245) := b"0000000000000000_0000000000000000_0001011101010111_0100000100110110"; -- 0.0911751514082603
	pesos_i(23246) := b"0000000000000000_0000000000000000_0000110110010101_0010101001001101"; -- 0.053057330886036355
	pesos_i(23247) := b"0000000000000000_0000000000000000_0000111001101110_1111010000001010"; -- 0.05638051255275191
	pesos_i(23248) := b"0000000000000000_0000000000000000_0001111111101010_1010010010001100"; -- 0.12467411447742831
	pesos_i(23249) := b"0000000000000000_0000000000000000_0000100001100011_1101111010000001"; -- 0.03277388230638835
	pesos_i(23250) := b"0000000000000000_0000000000000000_0001011000101010_0001001011100001"; -- 0.08657949436224309
	pesos_i(23251) := b"1111111111111111_1111111111111111_1111100111101101_1111010111010001"; -- -0.023712765120226537
	pesos_i(23252) := b"0000000000000000_0000000000000000_0000110111011001_0011110111000110"; -- 0.05409608909546558
	pesos_i(23253) := b"1111111111111111_1111111111111111_1111111001100111_1000011100110011"; -- -0.006232786324471507
	pesos_i(23254) := b"1111111111111111_1111111111111111_1111001000111101_0111101111100000"; -- -0.05374933042093558
	pesos_i(23255) := b"0000000000000000_0000000000000000_0001100101000101_1010100101001110"; -- 0.09871919770785949
	pesos_i(23256) := b"0000000000000000_0000000000000000_0001111110110101_1010001001111111"; -- 0.12386527627458857
	pesos_i(23257) := b"1111111111111111_1111111111111111_1111110000001110_1001011011011001"; -- -0.015402385743610237
	pesos_i(23258) := b"0000000000000000_0000000000000000_0010010010011100_1110101110100000"; -- 0.143019415324919
	pesos_i(23259) := b"1111111111111111_1111111111111111_1111010100010010_1010000111101010"; -- -0.04268444087161388
	pesos_i(23260) := b"1111111111111111_1111111111111111_1111000100110110_1110111001000110"; -- -0.057755573203108077
	pesos_i(23261) := b"0000000000000000_0000000000000000_0010000001101111_0001110101011101"; -- 0.1266954757517389
	pesos_i(23262) := b"0000000000000000_0000000000000000_0010001111101110_1101010110011010"; -- 0.1403630735472052
	pesos_i(23263) := b"0000000000000000_0000000000000000_0001111011010010_1011100000100011"; -- 0.12040282118513365
	pesos_i(23264) := b"1111111111111111_1111111111111111_1101110011110110_1001000000010110"; -- -0.13686274978015228
	pesos_i(23265) := b"0000000000000000_0000000000000000_0000010110100001_0111111010111001"; -- 0.021995468254070002
	pesos_i(23266) := b"1111111111111111_1111111111111111_1110100001000110_1011101101000101"; -- -0.09267072261603335
	pesos_i(23267) := b"1111111111111111_1111111111111111_1101011111000101_0001001011100111"; -- -0.15714914180696574
	pesos_i(23268) := b"1111111111111111_1111111111111111_1110000111110111_0000100111101101"; -- -0.11732423757802647
	pesos_i(23269) := b"0000000000000000_0000000000000000_0000011001101111_1111101100011100"; -- 0.025146192876944022
	pesos_i(23270) := b"1111111111111111_1111111111111111_1111001000100100_0101100100001111"; -- -0.0541328753349946
	pesos_i(23271) := b"0000000000000000_0000000000000000_0010001101110100_0010100111100000"; -- 0.13849126539649084
	pesos_i(23272) := b"0000000000000000_0000000000000000_0001010000101111_1111100100000010"; -- 0.07885700505170487
	pesos_i(23273) := b"0000000000000000_0000000000000000_0001001110111101_1000010010001110"; -- 0.07711056200490873
	pesos_i(23274) := b"1111111111111111_1111111111111111_1111110101000011_0111101010101111"; -- -0.010689098583140377
	pesos_i(23275) := b"0000000000000000_0000000000000000_0001111011100011_1111010011011111"; -- 0.12066584067648391
	pesos_i(23276) := b"1111111111111111_1111111111111111_1111010010000000_0110000001001101"; -- -0.0449161349491907
	pesos_i(23277) := b"0000000000000000_0000000000000000_0000001001101100_1000100011101011"; -- 0.009468610219388125
	pesos_i(23278) := b"1111111111111111_1111111111111111_1110000100111110_1000011100100101"; -- -0.12013964985732634
	pesos_i(23279) := b"0000000000000000_0000000000000000_0000110100111011_1011100101111001"; -- 0.05169257369818964
	pesos_i(23280) := b"0000000000000000_0000000000000000_0000011000010011_1010100111101000"; -- 0.02373754419479593
	pesos_i(23281) := b"1111111111111111_1111111111111111_1110001101010101_0101010010000111"; -- -0.11197921476003533
	pesos_i(23282) := b"1111111111111111_1111111111111111_1110011111111011_1101100111011101"; -- -0.09381330818518185
	pesos_i(23283) := b"0000000000000000_0000000000000000_0001001100010110_0110001110001100"; -- 0.07456037677618939
	pesos_i(23284) := b"0000000000000000_0000000000000000_0000011011101011_1111111011100101"; -- 0.027038508274359416
	pesos_i(23285) := b"1111111111111111_1111111111111111_1111111100011001_0100110000010010"; -- -0.0035202461526992897
	pesos_i(23286) := b"0000000000000000_0000000000000000_0010001001000001_0011110101001001"; -- 0.13380797416818074
	pesos_i(23287) := b"1111111111111111_1111111111111111_1111110001100111_1011101100011001"; -- -0.014042192856486235
	pesos_i(23288) := b"1111111111111111_1111111111111111_1111011001001100_0110000100001110"; -- -0.03789704709195192
	pesos_i(23289) := b"1111111111111111_1111111111111111_1110001001001101_0110111010101110"; -- -0.11600597611359889
	pesos_i(23290) := b"0000000000000000_0000000000000000_0001000011100000_0111101101100010"; -- 0.06592532293645939
	pesos_i(23291) := b"0000000000000000_0000000000000000_0000100011101000_0111101000111011"; -- 0.03479732463453741
	pesos_i(23292) := b"0000000000000000_0000000000000000_0001100101111111_1000101010101010"; -- 0.09960238118319253
	pesos_i(23293) := b"1111111111111111_1111111111111111_1110010101000010_0101101011001011"; -- -0.10445625817102493
	pesos_i(23294) := b"1111111111111111_1111111111111111_1101100100110101_0011101001010100"; -- -0.15153155745505417
	pesos_i(23295) := b"0000000000000000_0000000000000000_0010000101100110_1010010111011111"; -- 0.13047253314686252
	pesos_i(23296) := b"0000000000000000_0000000000000000_0000001101100001_1100100011010100"; -- 0.013210822815705936
	pesos_i(23297) := b"1111111111111111_1111111111111111_1110000111100011_1010010111000011"; -- -0.11762012462857621
	pesos_i(23298) := b"1111111111111111_1111111111111111_1110001100111111_0110011110110001"; -- -0.1123137658073607
	pesos_i(23299) := b"0000000000000000_0000000000000000_0000111000111100_1110101001011110"; -- 0.05561699679231466
	pesos_i(23300) := b"0000000000000000_0000000000000000_0001010011100110_1101101100010110"; -- 0.08164757993749518
	pesos_i(23301) := b"0000000000000000_0000000000000000_0000111001000010_1100110110000100"; -- 0.05570682972710129
	pesos_i(23302) := b"0000000000000000_0000000000000000_0010000000110100_1000000010010011"; -- 0.12580112073455132
	pesos_i(23303) := b"1111111111111111_1111111111111111_1110011011001001_0000000111010000"; -- -0.09849537547009098
	pesos_i(23304) := b"0000000000000000_0000000000000000_0000010100011100_1101011100111100"; -- 0.01997132497665402
	pesos_i(23305) := b"0000000000000000_0000000000000000_0000010010110000_0111100001010100"; -- 0.018317718901192197
	pesos_i(23306) := b"0000000000000000_0000000000000000_0000000001001110_1101001101101101"; -- 0.0012027876163475254
	pesos_i(23307) := b"0000000000000000_0000000000000000_0010011001010000_1000000101001011"; -- 0.14966590955289058
	pesos_i(23308) := b"0000000000000000_0000000000000000_0001001100100011_1111101100010001"; -- 0.07476777228333834
	pesos_i(23309) := b"0000000000000000_0000000000000000_0001000100101000_1001010111111011"; -- 0.0670255409915509
	pesos_i(23310) := b"1111111111111111_1111111111111111_1110000101101000_1010011111010001"; -- -0.11949683331813711
	pesos_i(23311) := b"1111111111111111_1111111111111111_1101110010111010_1000110100001111"; -- -0.13777845749497503
	pesos_i(23312) := b"0000000000000000_0000000000000000_0000001101001110_1010001000111111"; -- 0.012918606180053013
	pesos_i(23313) := b"0000000000000000_0000000000000000_0000101000011000_0010110101111100"; -- 0.0394314219471075
	pesos_i(23314) := b"0000000000000000_0000000000000000_0001101110101010_0010100101001000"; -- 0.10806520463341565
	pesos_i(23315) := b"1111111111111111_1111111111111111_1111011001000100_0011001011110010"; -- -0.038021865666259445
	pesos_i(23316) := b"1111111111111111_1111111111111111_1110100001110101_0101010101110101"; -- -0.09195962801032478
	pesos_i(23317) := b"0000000000000000_0000000000000000_0001110111101110_0010100100111001"; -- 0.11691529885361228
	pesos_i(23318) := b"0000000000000000_0000000000000000_0000001111011110_0000010111100001"; -- 0.015106551644494166
	pesos_i(23319) := b"0000000000000000_0000000000000000_0000011100110110_1010111000010000"; -- 0.028178099508116613
	pesos_i(23320) := b"0000000000000000_0000000000000000_0001011010011011_0011011010111111"; -- 0.08830587542137298
	pesos_i(23321) := b"1111111111111111_1111111111111111_1111110000000010_0001011111110111"; -- -0.015593054076600617
	pesos_i(23322) := b"1111111111111111_1111111111111111_1110101111000011_0110111000101101"; -- -0.07904921906986832
	pesos_i(23323) := b"0000000000000000_0000000000000000_0000000100110010_0111010101000010"; -- 0.004676178620360205
	pesos_i(23324) := b"1111111111111111_1111111111111111_1110101100010100_1101111100000110"; -- -0.08171278094390552
	pesos_i(23325) := b"1111111111111111_1111111111111111_1101111011100101_0001001000111000"; -- -0.12931715131631663
	pesos_i(23326) := b"0000000000000000_0000000000000000_0000011100001010_1010101011001100"; -- 0.027506518132382717
	pesos_i(23327) := b"0000000000000000_0000000000000000_0001001111011011_0111110101100011"; -- 0.07756789837915534
	pesos_i(23328) := b"1111111111111111_1111111111111111_1101110000000110_0111111110110011"; -- -0.14052583591544637
	pesos_i(23329) := b"1111111111111111_1111111111111111_1111100101100001_1110001110001110"; -- -0.025850084222212702
	pesos_i(23330) := b"0000000000000000_0000000000000000_0010001101111010_0001110111110111"; -- 0.13858210826325248
	pesos_i(23331) := b"0000000000000000_0000000000000000_0000011101010111_1101010000010001"; -- 0.02868390473281434
	pesos_i(23332) := b"1111111111111111_1111111111111111_1110000110100101_0111010100111100"; -- -0.11856906204059953
	pesos_i(23333) := b"0000000000000000_0000000000000000_0000111110010110_0111011101101101"; -- 0.060889686761158204
	pesos_i(23334) := b"0000000000000000_0000000000000000_0001000101001110_0011010100110000"; -- 0.0675996058700705
	pesos_i(23335) := b"0000000000000000_0000000000000000_0000010000011010_1110001100110100"; -- 0.01603527083229296
	pesos_i(23336) := b"1111111111111111_1111111111111111_1110111010100001_0110110110011000"; -- -0.06784930256079608
	pesos_i(23337) := b"0000000000000000_0000000000000000_0010000010001110_0101001111111011"; -- 0.1271717536897905
	pesos_i(23338) := b"0000000000000000_0000000000000000_0001011110001100_0101000101110001"; -- 0.09198483480832723
	pesos_i(23339) := b"1111111111111111_1111111111111111_1110001000000001_0001010101100010"; -- -0.11717096661810476
	pesos_i(23340) := b"0000000000000000_0000000000000000_0000110111001101_1010101010011111"; -- 0.05391947157163687
	pesos_i(23341) := b"1111111111111111_1111111111111111_1101101110000111_0010101111010100"; -- -0.14246870102320705
	pesos_i(23342) := b"1111111111111111_1111111111111111_1110100001111110_0000100001101110"; -- -0.09182689001798351
	pesos_i(23343) := b"1111111111111111_1111111111111111_1111010100111111_1100111111101101"; -- -0.04199505290552081
	pesos_i(23344) := b"1111111111111111_1111111111111111_1110000011001001_1011011000011010"; -- -0.12192212927522339
	pesos_i(23345) := b"1111111111111111_1111111111111111_1110100100010101_0011101000010011"; -- -0.08951985399869244
	pesos_i(23346) := b"1111111111111111_1111111111111111_1111001011100000_1100000100001101"; -- -0.05125802447747113
	pesos_i(23347) := b"1111111111111111_1111111111111111_1111010000101111_0011110011001001"; -- -0.04615421390041107
	pesos_i(23348) := b"0000000000000000_0000000000000000_0000111011010010_1000001110000011"; -- 0.05789968432333339
	pesos_i(23349) := b"1111111111111111_1111111111111111_1111011010100000_1111000111010001"; -- -0.036606680469056185
	pesos_i(23350) := b"0000000000000000_0000000000000000_0001111111011110_0011000011010001"; -- 0.12448411092357042
	pesos_i(23351) := b"1111111111111111_1111111111111111_1110110000101001_1111101101011101"; -- -0.07748440719993897
	pesos_i(23352) := b"0000000000000000_0000000000000000_0001010100001101_1111100001101011"; -- 0.08224442122292933
	pesos_i(23353) := b"0000000000000000_0000000000000000_0001000001100111_1011010110100011"; -- 0.06408248176203503
	pesos_i(23354) := b"1111111111111111_1111111111111111_1111111100000110_1010011111001100"; -- -0.0038046957272397483
	pesos_i(23355) := b"1111111111111111_1111111111111111_1110101010000010_1100011000100101"; -- -0.08394204712236836
	pesos_i(23356) := b"1111111111111111_1111111111111111_1110110111110100_0111110011110101"; -- -0.07048815734833508
	pesos_i(23357) := b"1111111111111111_1111111111111111_1110110100010011_0111111010011001"; -- -0.07392128730472382
	pesos_i(23358) := b"1111111111111111_1111111111111111_1110010011111001_0010011010100010"; -- -0.10557325878069554
	pesos_i(23359) := b"0000000000000000_0000000000000000_0001001110001110_1001000101100000"; -- 0.07639416303484615
	pesos_i(23360) := b"1111111111111111_1111111111111111_1111011101111100_0100011001000010"; -- -0.03325997253451501
	pesos_i(23361) := b"0000000000000000_0000000000000000_0000101110000001_0001000111110110"; -- 0.04493820442716896
	pesos_i(23362) := b"1111111111111111_1111111111111111_1101101011011000_1010100100000011"; -- -0.1451315276131041
	pesos_i(23363) := b"1111111111111111_1111111111111111_1110000011100111_1101000110111010"; -- -0.12146271906293529
	pesos_i(23364) := b"0000000000000000_0000000000000000_0010011100101001_1001001010101111"; -- 0.15297810340519272
	pesos_i(23365) := b"1111111111111111_1111111111111111_1111001101011001_1100110100011011"; -- -0.04941099244954112
	pesos_i(23366) := b"1111111111111111_1111111111111111_1111110101001011_0000101011011010"; -- -0.010573694025534477
	pesos_i(23367) := b"0000000000000000_0000000000000000_0001001111101100_1010110100001110"; -- 0.0778301389739321
	pesos_i(23368) := b"1111111111111111_1111111111111111_1111000011010000_0101101011000010"; -- -0.05932076227296108
	pesos_i(23369) := b"1111111111111111_1111111111111111_1101101100101100_0000100100011011"; -- -0.1438593205826716
	pesos_i(23370) := b"0000000000000000_0000000000000000_0001111011010010_1101101101100000"; -- 0.12040492157618456
	pesos_i(23371) := b"0000000000000000_0000000000000000_0001100001110100_1101001000100011"; -- 0.09553254458514884
	pesos_i(23372) := b"0000000000000000_0000000000000000_0010001101110101_0010000100001110"; -- 0.13850599862636837
	pesos_i(23373) := b"1111111111111111_1111111111111111_1111010111111011_1110010011111010"; -- -0.039125145904635984
	pesos_i(23374) := b"1111111111111111_1111111111111111_1111100100000111_0100100100000111"; -- -0.02723258578790962
	pesos_i(23375) := b"1111111111111111_1111111111111111_1101100000100110_0110100011001101"; -- -0.15566391936955834
	pesos_i(23376) := b"0000000000000000_0000000000000000_0001110001010110_1011100110001101"; -- 0.11069831545276657
	pesos_i(23377) := b"0000000000000000_0000000000000000_0000011011000100_1110110010110010"; -- 0.026442330698931468
	pesos_i(23378) := b"0000000000000000_0000000000000000_0001001011100111_1001111111100010"; -- 0.07384681006911341
	pesos_i(23379) := b"1111111111111111_1111111111111111_1101101111110011_1010011101111000"; -- -0.14081338234784305
	pesos_i(23380) := b"0000000000000000_0000000000000000_0001011111001100_0000111101111011"; -- 0.09295746557841668
	pesos_i(23381) := b"0000000000000000_0000000000000000_0001000100101101_0001011110101001"; -- 0.06709430569919224
	pesos_i(23382) := b"0000000000000000_0000000000000000_0000111000101110_1110011100110011"; -- 0.05540318482565806
	pesos_i(23383) := b"1111111111111111_1111111111111111_1101111010100101_1011111010000001"; -- -0.13028344499291292
	pesos_i(23384) := b"0000000000000000_0000000000000000_0000000000000001_1000101011000111"; -- 2.353048998665878e-05
	pesos_i(23385) := b"1111111111111111_1111111111111111_1111010111101011_1001001011010101"; -- -0.03937418265970408
	pesos_i(23386) := b"1111111111111111_1111111111111111_1111000010110000_0111100100001101"; -- -0.059807237920915614
	pesos_i(23387) := b"1111111111111111_1111111111111111_1111111111001101_1100011001100001"; -- -0.00076637404026504
	pesos_i(23388) := b"1111111111111111_1111111111111111_1111011000001101_1110111100001111"; -- -0.038849886720457145
	pesos_i(23389) := b"0000000000000000_0000000000000000_0001010111000000_1101111011101101"; -- 0.08497422497068495
	pesos_i(23390) := b"0000000000000000_0000000000000000_0000101111010010_0000001101111001"; -- 0.04617330261108434
	pesos_i(23391) := b"0000000000000000_0000000000000000_0001101010001001_1110111000100011"; -- 0.10366714804254588
	pesos_i(23392) := b"1111111111111111_1111111111111111_1110010010011001_0001100001001101"; -- -0.10703895689558358
	pesos_i(23393) := b"1111111111111111_1111111111111111_1110110101110000_0001011010111111"; -- -0.07250840987848668
	pesos_i(23394) := b"0000000000000000_0000000000000000_0000010111011111_1011101010000110"; -- 0.022945077535557315
	pesos_i(23395) := b"0000000000000000_0000000000000000_0000010010110010_1111000011111010"; -- 0.018355427758102068
	pesos_i(23396) := b"0000000000000000_0000000000000000_0001101101001110_1101000100100110"; -- 0.10667140165222716
	pesos_i(23397) := b"0000000000000000_0000000000000000_0000101000010110_1100110011010001"; -- 0.03941040131714901
	pesos_i(23398) := b"0000000000000000_0000000000000000_0001000011110111_1010011001000111"; -- 0.06627883189692302
	pesos_i(23399) := b"1111111111111111_1111111111111111_1111010001100001_1010010000110101"; -- -0.04538510989100395
	pesos_i(23400) := b"1111111111111111_1111111111111111_1111000000111101_1001110000111010"; -- -0.0615599019759946
	pesos_i(23401) := b"0000000000000000_0000000000000000_0001001110110110_1000101101010000"; -- 0.07700415320241868
	pesos_i(23402) := b"1111111111111111_1111111111111111_1110111000011001_0011110011100000"; -- -0.06992740176046162
	pesos_i(23403) := b"0000000000000000_0000000000000000_0010001100101100_1111000110000010"; -- 0.13740453163369248
	pesos_i(23404) := b"1111111111111111_1111111111111111_1110000011011001_1110000011000000"; -- -0.1216754466630026
	pesos_i(23405) := b"0000000000000000_0000000000000000_0010001111100110_0011110100111111"; -- 0.14023192193039993
	pesos_i(23406) := b"0000000000000000_0000000000000000_0000110010110011_0100101000011011"; -- 0.04961074021180171
	pesos_i(23407) := b"1111111111111111_1111111111111111_1101111101100101_0011111011001011"; -- -0.1273613695139392
	pesos_i(23408) := b"1111111111111111_1111111111111111_1110010111000010_1000111000101110"; -- -0.10250007043248842
	pesos_i(23409) := b"1111111111111111_1111111111111111_1111111000111001_0011101100100010"; -- -0.006939224333644241
	pesos_i(23410) := b"1111111111111111_1111111111111111_1110010111111000_0101000110011101"; -- -0.10167970582165203
	pesos_i(23411) := b"1111111111111111_1111111111111111_1111111010011011_1010001110010100"; -- -0.005437637713918741
	pesos_i(23412) := b"1111111111111111_1111111111111111_1101101110110110_0010100100101010"; -- -0.141751696888302
	pesos_i(23413) := b"1111111111111111_1111111111111111_1101101011101110_1111101011010001"; -- -0.14479095832426273
	pesos_i(23414) := b"0000000000000000_0000000000000000_0000011100011110_0101001101001001"; -- 0.02780647777585239
	pesos_i(23415) := b"1111111111111111_1111111111111111_1111000110000011_0010111000000000"; -- -0.0565921067617475
	pesos_i(23416) := b"0000000000000000_0000000000000000_0001010101010100_1001110001011000"; -- 0.08332230698813341
	pesos_i(23417) := b"1111111111111111_1111111111111111_1110111001000000_1101100001101010"; -- -0.06932303828034027
	pesos_i(23418) := b"1111111111111111_1111111111111111_1110101000011111_0111110111100011"; -- -0.08545697402125635
	pesos_i(23419) := b"0000000000000000_0000000000000000_0000101000010101_1011000100100111"; -- 0.039393493562649165
	pesos_i(23420) := b"0000000000000000_0000000000000000_0000000100110111_1000110001011011"; -- 0.004753849284907721
	pesos_i(23421) := b"0000000000000000_0000000000000000_0010010000110001_1001011001111001"; -- 0.14138164943876055
	pesos_i(23422) := b"1111111111111111_1111111111111111_1111010101010010_0101010100010110"; -- -0.04171245779376857
	pesos_i(23423) := b"0000000000000000_0000000000000000_0001001111100100_0000011001010100"; -- 0.07769813099948432
	pesos_i(23424) := b"1111111111111111_1111111111111111_1110111110010000_0111001110011011"; -- -0.06420209376293314
	pesos_i(23425) := b"1111111111111111_1111111111111111_1101110100011000_1010100111100110"; -- -0.13634241239451475
	pesos_i(23426) := b"0000000000000000_0000000000000000_0000001010001101_1110001101111001"; -- 0.009977547666714218
	pesos_i(23427) := b"1111111111111111_1111111111111111_1111010110001000_1111011001000001"; -- -0.040878876758874784
	pesos_i(23428) := b"1111111111111111_1111111111111111_1110111001101011_0100000001101011"; -- -0.06867597001272085
	pesos_i(23429) := b"1111111111111111_1111111111111111_1111111011001001_0100100011110011"; -- -0.00474113527842824
	pesos_i(23430) := b"1111111111111111_1111111111111111_1110010111110000_1010011000101011"; -- -0.1017967361961674
	pesos_i(23431) := b"0000000000000000_0000000000000000_0001110110011000_0100101111111100"; -- 0.11560511493541102
	pesos_i(23432) := b"0000000000000000_0000000000000000_0001001111101010_1010100011111011"; -- 0.07779937868678975
	pesos_i(23433) := b"1111111111111111_1111111111111111_1111010000111001_1110101000100111"; -- -0.04599129244424166
	pesos_i(23434) := b"0000000000000000_0000000000000000_0001001111111010_0100011110111001"; -- 0.07803772233023602
	pesos_i(23435) := b"0000000000000000_0000000000000000_0010000010011010_1001111000001111"; -- 0.12735927456804363
	pesos_i(23436) := b"1111111111111111_1111111111111111_1111111000001010_0100000001010001"; -- -0.007656078502194444
	pesos_i(23437) := b"1111111111111111_1111111111111111_1110011101110100_1010001111100011"; -- -0.09587646212052076
	pesos_i(23438) := b"0000000000000000_0000000000000000_0001100111001010_0111000101100111"; -- 0.10074528470012917
	pesos_i(23439) := b"0000000000000000_0000000000000000_0000000000011111_0001110001010100"; -- 0.0004747109663192182
	pesos_i(23440) := b"0000000000000000_0000000000000000_0001001100111010_0110110110111010"; -- 0.0751103000826475
	pesos_i(23441) := b"1111111111111111_1111111111111111_1110111100101000_1111011101000000"; -- -0.06578116107621049
	pesos_i(23442) := b"0000000000000000_0000000000000000_0001100011010001_0000111001110011"; -- 0.09693994819460162
	pesos_i(23443) := b"1111111111111111_1111111111111111_1110011110111010_1001111010100010"; -- -0.09480866004522273
	pesos_i(23444) := b"1111111111111111_1111111111111111_1110100100011111_1111000110111011"; -- -0.08935631936245234
	pesos_i(23445) := b"0000000000000000_0000000000000000_0010000001110011_1010110100110101"; -- 0.1267650847647263
	pesos_i(23446) := b"0000000000000000_0000000000000000_0010000000010011_0110100100010000"; -- 0.12529617930211542
	pesos_i(23447) := b"0000000000000000_0000000000000000_0001111000111010_1010111100100100"; -- 0.11808294896004487
	pesos_i(23448) := b"1111111111111111_1111111111111111_1101100101111011_0000110101110101"; -- -0.15046611686650105
	pesos_i(23449) := b"0000000000000000_0000000000000000_0010000010110100_1101101011010010"; -- 0.12775962473472444
	pesos_i(23450) := b"0000000000000000_0000000000000000_0001101110111100_0011111000010111"; -- 0.1083411032654653
	pesos_i(23451) := b"1111111111111111_1111111111111111_1110011000010011_0111001001101111"; -- -0.10126576218261794
	pesos_i(23452) := b"1111111111111111_1111111111111111_1110001111101001_1111110111111010"; -- -0.10971081390292974
	pesos_i(23453) := b"0000000000000000_0000000000000000_0001110101000001_0010010011010110"; -- 0.11427526682851946
	pesos_i(23454) := b"1111111111111111_1111111111111111_1111000100001100_0000001111011010"; -- -0.05841041500024171
	pesos_i(23455) := b"0000000000000000_0000000000000000_0001110010010000_0000010010001001"; -- 0.1115725359826879
	pesos_i(23456) := b"1111111111111111_1111111111111111_1111100110000111_0100000100101111"; -- -0.025279928294340236
	pesos_i(23457) := b"0000000000000000_0000000000000000_0010100010111001_0111011011001010"; -- 0.15907995638775627
	pesos_i(23458) := b"1111111111111111_1111111111111111_1111101010000100_1010110101001110"; -- -0.02141301011284647
	pesos_i(23459) := b"0000000000000000_0000000000000000_0000111001000000_1110011000111001"; -- 0.05567778490577866
	pesos_i(23460) := b"1111111111111111_1111111111111111_1111010011101010_0101000010100111"; -- -0.043299636133981655
	pesos_i(23461) := b"1111111111111111_1111111111111111_1110000001011101_1000011101010100"; -- -0.12357286632502085
	pesos_i(23462) := b"1111111111111111_1111111111111111_1110010101100110_1110000110111001"; -- -0.10389889939318868
	pesos_i(23463) := b"1111111111111111_1111111111111111_1101111011111111_0011011101110100"; -- -0.1289182035190288
	pesos_i(23464) := b"0000000000000000_0000000000000000_0010001011000001_0000101101010000"; -- 0.13575812051567201
	pesos_i(23465) := b"0000000000000000_0000000000000000_0001010111001000_1000001100001000"; -- 0.08509081789534848
	pesos_i(23466) := b"1111111111111111_1111111111111111_1111001011101000_0011011000100001"; -- -0.05114423456070852
	pesos_i(23467) := b"0000000000000000_0000000000000000_0001000101010000_0110100100101001"; -- 0.06763322118241304
	pesos_i(23468) := b"0000000000000000_0000000000000000_0001010010111001_0011101010110001"; -- 0.08095137426029515
	pesos_i(23469) := b"0000000000000000_0000000000000000_0001001101010011_1001100011010100"; -- 0.0754943387986166
	pesos_i(23470) := b"1111111111111111_1111111111111111_1111110001111111_1101100100110110"; -- -0.013674186913529321
	pesos_i(23471) := b"1111111111111111_1111111111111111_1110111101010110_1000011010101110"; -- -0.06508596659781181
	pesos_i(23472) := b"0000000000000000_0000000000000000_0001101000010101_1001001111110011"; -- 0.10189175299215052
	pesos_i(23473) := b"0000000000000000_0000000000000000_0000110011110110_0010101000111011"; -- 0.05063117923673894
	pesos_i(23474) := b"1111111111111111_1111111111111111_1110000001011001_0100100000000011"; -- -0.1236376754681333
	pesos_i(23475) := b"1111111111111111_1111111111111111_1111111100010010_1000111110000110"; -- -0.0036230372417623826
	pesos_i(23476) := b"0000000000000000_0000000000000000_0001010101001001_0000101101100100"; -- 0.08314582064464543
	pesos_i(23477) := b"1111111111111111_1111111111111111_1111100011001001_1101001011000001"; -- -0.028170421561236614
	pesos_i(23478) := b"1111111111111111_1111111111111111_1110110000011111_0101111001000010"; -- -0.07764635942535045
	pesos_i(23479) := b"0000000000000000_0000000000000000_0001110111100110_0000111001110011"; -- 0.11679163272751325
	pesos_i(23480) := b"1111111111111111_1111111111111111_1110110101011000_0101011101111111"; -- -0.07287076145891466
	pesos_i(23481) := b"1111111111111111_1111111111111111_1110011000011011_1011111111011110"; -- -0.10113907652298136
	pesos_i(23482) := b"1111111111111111_1111111111111111_1111101011110011_0110011010011111"; -- -0.01972349761979366
	pesos_i(23483) := b"1111111111111111_1111111111111111_1110010011101001_1100110111110111"; -- -0.10580742566622706
	pesos_i(23484) := b"1111111111111111_1111111111111111_1111000011100010_0001101000000111"; -- -0.059049962304867615
	pesos_i(23485) := b"1111111111111111_1111111111111111_1111100001011011_1100110110001010"; -- -0.02984919909323854
	pesos_i(23486) := b"1111111111111111_1111111111111111_1101101111100111_1111011101000011"; -- -0.14099173171448753
	pesos_i(23487) := b"0000000000000000_0000000000000000_0000110010100101_1110110001000010"; -- 0.049406782150954516
	pesos_i(23488) := b"1111111111111111_1111111111111111_1111000011110010_1111010101100010"; -- -0.05879274718067633
	pesos_i(23489) := b"1111111111111111_1111111111111111_1111110110010100_1100101101100000"; -- -0.009448327089972204
	pesos_i(23490) := b"1111111111111111_1111111111111111_1110011000101101_0111001010100001"; -- -0.10086902217964695
	pesos_i(23491) := b"1111111111111111_1111111111111111_1110001111100111_0101011010110010"; -- -0.10975130236212866
	pesos_i(23492) := b"1111111111111111_1111111111111111_1110000001011011_0111101111000110"; -- -0.12360407273025971
	pesos_i(23493) := b"1111111111111111_1111111111111111_1101111101111011_0110011001000110"; -- -0.1270233228807648
	pesos_i(23494) := b"0000000000000000_0000000000000000_0001000111110011_0011001010100111"; -- 0.07011715487781786
	pesos_i(23495) := b"1111111111111111_1111111111111111_1110011100100011_1111110100001010"; -- -0.0971071100215069
	pesos_i(23496) := b"0000000000000000_0000000000000000_0010001100011101_0000100011101100"; -- 0.137161786737593
	pesos_i(23497) := b"0000000000000000_0000000000000000_0001110000100100_1011000000101101"; -- 0.10993481718594278
	pesos_i(23498) := b"1111111111111111_1111111111111111_1110100011000110_1101001000000001"; -- -0.09071624253338056
	pesos_i(23499) := b"0000000000000000_0000000000000000_0010011000001101_1001111110001011"; -- 0.14864537385003485
	pesos_i(23500) := b"0000000000000000_0000000000000000_0001001100110110_1000100011001011"; -- 0.0750508780542554
	pesos_i(23501) := b"0000000000000000_0000000000000000_0001011101110111_0110111101110010"; -- 0.0916661884911515
	pesos_i(23502) := b"1111111111111111_1111111111111111_1110010010000001_1010101011100100"; -- -0.10739643022878058
	pesos_i(23503) := b"0000000000000000_0000000000000000_0000100010010000_0000101101010011"; -- 0.033447940504786486
	pesos_i(23504) := b"0000000000000000_0000000000000000_0001011000111001_0001000110001111"; -- 0.08680829752677853
	pesos_i(23505) := b"0000000000000000_0000000000000000_0000011110100111_1111100111110010"; -- 0.02990686576163289
	pesos_i(23506) := b"1111111111111111_1111111111111111_1110110101111110_0010100101101100"; -- -0.07229367353830633
	pesos_i(23507) := b"1111111111111111_1111111111111111_1110101010011110_1111101110000101"; -- -0.08351161955958537
	pesos_i(23508) := b"1111111111111111_1111111111111111_1111101111000010_0100001110111100"; -- -0.016567007692284804
	pesos_i(23509) := b"1111111111111111_1111111111111111_1110111100011110_0100110111001110"; -- -0.0659438489009587
	pesos_i(23510) := b"0000000000000000_0000000000000000_0001101110100101_1100011010010101"; -- 0.10799828664887152
	pesos_i(23511) := b"1111111111111111_1111111111111111_1111001000110011_1001111000111000"; -- -0.05389987112425091
	pesos_i(23512) := b"0000000000000000_0000000000000000_0001010100100001_0011000100101010"; -- 0.08253772054384607
	pesos_i(23513) := b"1111111111111111_1111111111111111_1110000100001111_0001001010000011"; -- -0.12086376473736725
	pesos_i(23514) := b"0000000000000000_0000000000000000_0001011001110001_0101010010100110"; -- 0.08766678870650442
	pesos_i(23515) := b"0000000000000000_0000000000000000_0001011011000100_0110110100000111"; -- 0.08893472126213235
	pesos_i(23516) := b"1111111111111111_1111111111111111_1111010011001011_1001110010011010"; -- -0.0437681317054251
	pesos_i(23517) := b"0000000000000000_0000000000000000_0001001101000011_0001011001010001"; -- 0.0752424190395831
	pesos_i(23518) := b"1111111111111111_1111111111111111_1110110010110010_1001110010111110"; -- -0.07539959296403931
	pesos_i(23519) := b"0000000000000000_0000000000000000_0000001001011000_0100101011110111"; -- 0.00915974175096481
	pesos_i(23520) := b"0000000000000000_0000000000000000_0001000011000100_1110011001101010"; -- 0.06550445645598078
	pesos_i(23521) := b"1111111111111111_1111111111111111_1101110100100000_0001001111111011"; -- -0.13622927776785937
	pesos_i(23522) := b"1111111111111111_1111111111111111_1111010000010001_1001110001100110"; -- -0.04660627848529777
	pesos_i(23523) := b"0000000000000000_0000000000000000_0000111100000100_0100000110100111"; -- 0.05865869828400152
	pesos_i(23524) := b"1111111111111111_1111111111111111_1110110001010000_1111101101110110"; -- -0.07688930868067577
	pesos_i(23525) := b"0000000000000000_0000000000000000_0000110000111001_1111100010011011"; -- 0.04775956891541664
	pesos_i(23526) := b"1111111111111111_1111111111111111_1110100010011011_0000111101100110"; -- -0.09138396985693104
	pesos_i(23527) := b"0000000000000000_0000000000000000_0000111110010000_0001111001110100"; -- 0.06079283085292595
	pesos_i(23528) := b"1111111111111111_1111111111111111_1111110110011111_0010111111110110"; -- -0.009289743836835476
	pesos_i(23529) := b"0000000000000000_0000000000000000_0001011001010011_1001100100100100"; -- 0.08721310732999214
	pesos_i(23530) := b"0000000000000000_0000000000000000_0000111101101100_0101111101110001"; -- 0.060247387989279685
	pesos_i(23531) := b"1111111111111111_1111111111111111_1111000010111010_1111010011110101"; -- -0.05964726474523335
	pesos_i(23532) := b"1111111111111111_1111111111111111_1111000000000111_1110111111100011"; -- -0.062378890021834
	pesos_i(23533) := b"1111111111111111_1111111111111111_1101101000011101_1000011111111100"; -- -0.1479868897239426
	pesos_i(23534) := b"1111111111111111_1111111111111111_1111110001010001_1101010101011101"; -- -0.014376320649087882
	pesos_i(23535) := b"0000000000000000_0000000000000000_0000101011001000_1010111100000011"; -- 0.04212468922223486
	pesos_i(23536) := b"1111111111111111_1111111111111111_1101101100000100_0111011001000001"; -- -0.14446316636214138
	pesos_i(23537) := b"1111111111111111_1111111111111111_1111010011000111_1000110101011101"; -- -0.043830075144846554
	pesos_i(23538) := b"0000000000000000_0000000000000000_0001100101101111_1011001011110100"; -- 0.09936064209368412
	pesos_i(23539) := b"0000000000000000_0000000000000000_0001001101010011_0110010010000000"; -- 0.07549121972842916
	pesos_i(23540) := b"1111111111111111_1111111111111111_1110011000001000_1111111010101101"; -- -0.10142524982830613
	pesos_i(23541) := b"1111111111111111_1111111111111111_1111101011101011_0110001101000000"; -- -0.01984576871443826
	pesos_i(23542) := b"0000000000000000_0000000000000000_0001000000110110_1100011110111101"; -- 0.06333588001601922
	pesos_i(23543) := b"0000000000000000_0000000000000000_0010001111100110_1110100100010111"; -- 0.14024216468635559
	pesos_i(23544) := b"1111111111111111_1111111111111111_1111010000100110_0001110010110001"; -- -0.04629345585254796
	pesos_i(23545) := b"0000000000000000_0000000000000000_0000010110101011_1110000011010001"; -- 0.02215390309427682
	pesos_i(23546) := b"0000000000000000_0000000000000000_0010001101000011_1101001110100001"; -- 0.13775370294497652
	pesos_i(23547) := b"1111111111111111_1111111111111111_1111100000111101_0101100000100010"; -- -0.030313960782919935
	pesos_i(23548) := b"1111111111111111_1111111111111111_1101111111110101_1110001110111101"; -- -0.12515427235655066
	pesos_i(23549) := b"1111111111111111_1111111111111111_1101110101110101_0000010011110000"; -- -0.13493317731739576
	pesos_i(23550) := b"0000000000000000_0000000000000000_0000000110000100_1110111000000101"; -- 0.0059345972630502715
	pesos_i(23551) := b"1111111111111111_1111111111111111_1110001111000100_1110001100011110"; -- -0.11027699020299234
	pesos_i(23552) := b"0000000000000000_0000000000000000_0000110100000001_1001010000011110"; -- 0.05080533733615937
	pesos_i(23553) := b"0000000000000000_0000000000000000_0000011101111001_1001101010011010"; -- 0.029199278331614616
	pesos_i(23554) := b"0000000000000000_0000000000000000_0000100011110100_1000011101000001"; -- 0.03498120617939705
	pesos_i(23555) := b"1111111111111111_1111111111111111_1110100010100111_1010111111100111"; -- -0.0911912976667574
	pesos_i(23556) := b"0000000000000000_0000000000000000_0010000010011100_0100100001011110"; -- 0.12738468444469742
	pesos_i(23557) := b"1111111111111111_1111111111111111_1111001011101001_0100001000111101"; -- -0.05112825412254592
	pesos_i(23558) := b"0000000000000000_0000000000000000_0001000101001100_0001100001111100"; -- 0.06756737731739464
	pesos_i(23559) := b"0000000000000000_0000000000000000_0000110010111010_0010110111001100"; -- 0.049715864559879315
	pesos_i(23560) := b"1111111111111111_1111111111111111_1111010110001100_0100001001100000"; -- -0.04082856323484454
	pesos_i(23561) := b"1111111111111111_1111111111111111_1111001101010010_0001101111001101"; -- -0.04952837226819669
	pesos_i(23562) := b"0000000000000000_0000000000000000_0001111001000110_1000001100100111"; -- 0.11826343250245272
	pesos_i(23563) := b"0000000000000000_0000000000000000_0000110000110000_1101000011001011"; -- 0.047619866916009196
	pesos_i(23564) := b"0000000000000000_0000000000000000_0001110000111110_1001001110101000"; -- 0.11032984580677647
	pesos_i(23565) := b"0000000000000000_0000000000000000_0001011010000011_0110110000011011"; -- 0.0879428449904578
	pesos_i(23566) := b"1111111111111111_1111111111111111_1111000001000001_0010100110111111"; -- -0.061505690560182374
	pesos_i(23567) := b"0000000000000000_0000000000000000_0000110111010111_1011011011101001"; -- 0.054072792014093346
	pesos_i(23568) := b"1111111111111111_1111111111111111_1111101001010000_0101011010001100"; -- -0.022211638173873633
	pesos_i(23569) := b"0000000000000000_0000000000000000_0001110001101110_1110111000001011"; -- 0.11106765516539277
	pesos_i(23570) := b"0000000000000000_0000000000000000_0000101100111011_1010000010111000"; -- 0.04387859806413029
	pesos_i(23571) := b"0000000000000000_0000000000000000_0001001000011100_0011110101011010"; -- 0.07074340294164116
	pesos_i(23572) := b"1111111111111111_1111111111111111_1111111011110010_0011100101000101"; -- -0.004116459477060526
	pesos_i(23573) := b"0000000000000000_0000000000000000_0000100101100100_1010100111110000"; -- 0.036692258077736045
	pesos_i(23574) := b"1111111111111111_1111111111111111_1101011010011000_1111100110000001"; -- -0.16172829242119918
	pesos_i(23575) := b"0000000000000000_0000000000000000_0010000011001011_1010110100010110"; -- 0.1281078509052721
	pesos_i(23576) := b"1111111111111111_1111111111111111_1111100010111011_1001101000000010"; -- -0.028387426919706457
	pesos_i(23577) := b"0000000000000000_0000000000000000_0001011000101010_1101101001100001"; -- 0.08659138547682435
	pesos_i(23578) := b"0000000000000000_0000000000000000_0001010011101111_0101100000000100"; -- 0.08177709682082746
	pesos_i(23579) := b"1111111111111111_1111111111111111_1110001000100000_0111110010000010"; -- -0.11669179748054322
	pesos_i(23580) := b"1111111111111111_1111111111111111_1111001010010100_0010100000110111"; -- -0.05242680215105069
	pesos_i(23581) := b"0000000000000000_0000000000000000_0001100100011101_1010011010100011"; -- 0.09810868708930501
	pesos_i(23582) := b"0000000000000000_0000000000000000_0001001010001111_0001011011011110"; -- 0.07249586977564013
	pesos_i(23583) := b"1111111111111111_1111111111111111_1110000101101000_0001000001000010"; -- -0.11950586681778672
	pesos_i(23584) := b"1111111111111111_1111111111111111_1101111000001011_1101000110110100"; -- -0.13263215415073512
	pesos_i(23585) := b"1111111111111111_1111111111111111_1111001111111110_0011101001011000"; -- -0.04690203994863325
	pesos_i(23586) := b"0000000000000000_0000000000000000_0001001100000100_0100110101100110"; -- 0.07428439844935264
	pesos_i(23587) := b"1111111111111111_1111111111111111_1111111101010010_0111101101001010"; -- -0.0026476807927682984
	pesos_i(23588) := b"0000000000000000_0000000000000000_0000101010000110_0001010110100111"; -- 0.04110846830323426
	pesos_i(23589) := b"0000000000000000_0000000000000000_0001000101111110_0011011011100010"; -- 0.068332128625674
	pesos_i(23590) := b"1111111111111111_1111111111111111_1101101011110010_1111100001011000"; -- -0.14473007064341228
	pesos_i(23591) := b"0000000000000000_0000000000000000_0000011001100001_0010111000011111"; -- 0.024920351658339134
	pesos_i(23592) := b"0000000000000000_0000000000000000_0001100111111011_0110111001000100"; -- 0.10149277851140516
	pesos_i(23593) := b"0000000000000000_0000000000000000_0001100011001011_0010011001111111"; -- 0.09684982871312789
	pesos_i(23594) := b"1111111111111111_1111111111111111_1110110101000010_0000110011111111"; -- -0.073210895319105
	pesos_i(23595) := b"1111111111111111_1111111111111111_1101110100110000_1011010101101010"; -- -0.13597551493198803
	pesos_i(23596) := b"1111111111111111_1111111111111111_1110101001011100_1010000100101111"; -- -0.08452408409893211
	pesos_i(23597) := b"1111111111111111_1111111111111111_1111101011111101_0101101111000000"; -- -0.01957155768489253
	pesos_i(23598) := b"1111111111111111_1111111111111111_1101101011010110_1000010011110110"; -- -0.14516419414383003
	pesos_i(23599) := b"1111111111111111_1111111111111111_1110001101010110_0001101011011000"; -- -0.11196739416987316
	pesos_i(23600) := b"1111111111111111_1111111111111111_1101111111000001_0100110000000000"; -- -0.12595677367570993
	pesos_i(23601) := b"0000000000000000_0000000000000000_0001110000101011_0010111001001010"; -- 0.11003388691584375
	pesos_i(23602) := b"1111111111111111_1111111111111111_1101101011110011_1001010010011000"; -- -0.14472075746999882
	pesos_i(23603) := b"0000000000000000_0000000000000000_0000011101110100_1010011100110010"; -- 0.029123735195354203
	pesos_i(23604) := b"1111111111111111_1111111111111111_1111101000010010_0111011010001100"; -- -0.02315577594509199
	pesos_i(23605) := b"1111111111111111_1111111111111111_1110101000000011_1011000001011111"; -- -0.08588121099020775
	pesos_i(23606) := b"1111111111111111_1111111111111111_1110110101110111_0000101101101000"; -- -0.07240227429122587
	pesos_i(23607) := b"1111111111111111_1111111111111111_1110011010010010_1100110110101111"; -- -0.0993224569976125
	pesos_i(23608) := b"1111111111111111_1111111111111111_1101101100011010_1010001001110100"; -- -0.14412483861136083
	pesos_i(23609) := b"1111111111111111_1111111111111111_1110110011001000_0010000101111111"; -- -0.0750712456560679
	pesos_i(23610) := b"0000000000000000_0000000000000000_0010010001001010_0011111010011000"; -- 0.1417578812742393
	pesos_i(23611) := b"1111111111111111_1111111111111111_1110001111011111_0000110010110010"; -- -0.10987778322590465
	pesos_i(23612) := b"0000000000000000_0000000000000000_0000000101110101_1000000010000011"; -- 0.005699188163839006
	pesos_i(23613) := b"0000000000000000_0000000000000000_0001101101100100_1010110110111010"; -- 0.10700498371547833
	pesos_i(23614) := b"0000000000000000_0000000000000000_0000110000011010_1000010101101101"; -- 0.04727968132130196
	pesos_i(23615) := b"1111111111111111_1111111111111111_1111101010101101_1000100010110110"; -- -0.020789580897074965
	pesos_i(23616) := b"1111111111111111_1111111111111111_1101111000100011_1000010100010100"; -- -0.13227051023461975
	pesos_i(23617) := b"1111111111111111_1111111111111111_1111111000110001_0011001010100000"; -- -0.007061801740669042
	pesos_i(23618) := b"1111111111111111_1111111111111111_1110110101010000_0000010111001011"; -- -0.07299770164195987
	pesos_i(23619) := b"1111111111111111_1111111111111111_1111110111100010_1101101010000010"; -- -0.008257239597257373
	pesos_i(23620) := b"0000000000000000_0000000000000000_0000011101011010_1100010100010100"; -- 0.02872878775962841
	pesos_i(23621) := b"1111111111111111_1111111111111111_1111010111110000_0100111000010001"; -- -0.03930198741913641
	pesos_i(23622) := b"1111111111111111_1111111111111111_1111000001110000_0111000001111011"; -- -0.06078431135669825
	pesos_i(23623) := b"0000000000000000_0000000000000000_0001111110100001_0100001101011000"; -- 0.12355442904354018
	pesos_i(23624) := b"0000000000000000_0000000000000000_0000010100001001_1000001000001010"; -- 0.01967632995124326
	pesos_i(23625) := b"1111111111111111_1111111111111111_1110011000000110_0011100011001011"; -- -0.10146756223984255
	pesos_i(23626) := b"0000000000000000_0000000000000000_0000011100101011_1010000011001110"; -- 0.028009462685648825
	pesos_i(23627) := b"0000000000000000_0000000000000000_0001011111101110_0010100000010000"; -- 0.09347772968559362
	pesos_i(23628) := b"1111111111111111_1111111111111111_1111001010000100_1100011111110011"; -- -0.052661421980359925
	pesos_i(23629) := b"1111111111111111_1111111111111111_1111100111110110_0101111110010101"; -- -0.02358439072755268
	pesos_i(23630) := b"0000000000000000_0000000000000000_0000100111100110_0010100011100000"; -- 0.038668207862732576
	pesos_i(23631) := b"0000000000000000_0000000000000000_0000011010110010_0001110011110001"; -- 0.026155289473383334
	pesos_i(23632) := b"1111111111111111_1111111111111111_1111101101110001_0011001101011111"; -- -0.017803944797761824
	pesos_i(23633) := b"0000000000000000_0000000000000000_0010011000000001_1001001101011110"; -- 0.1484615425603015
	pesos_i(23634) := b"1111111111111111_1111111111111111_1110001001001111_0110001110010001"; -- -0.11597612096199546
	pesos_i(23635) := b"0000000000000000_0000000000000000_0001000100010001_1110010101000101"; -- 0.06667931487687247
	pesos_i(23636) := b"0000000000000000_0000000000000000_0000111000100011_1100000000001101"; -- 0.05523300471348246
	pesos_i(23637) := b"1111111111111111_1111111111111111_1110110100010010_0000010111101101"; -- -0.07394373857915205
	pesos_i(23638) := b"1111111111111111_1111111111111111_1110010011011000_1110100111010000"; -- -0.10606516522465956
	pesos_i(23639) := b"0000000000000000_0000000000000000_0000011000111000_1010000110111100"; -- 0.024301632225550915
	pesos_i(23640) := b"0000000000000000_0000000000000000_0010010100001111_1010101010111011"; -- 0.14477030815717737
	pesos_i(23641) := b"0000000000000000_0000000000000000_0001111111100111_1010011111110001"; -- 0.12462854026182407
	pesos_i(23642) := b"1111111111111111_1111111111111111_1111101010101010_0010000001110111"; -- -0.020841570821096896
	pesos_i(23643) := b"1111111111111111_1111111111111111_1101111010001110_0101000101111101"; -- -0.13064089490021602
	pesos_i(23644) := b"1111111111111111_1111111111111111_1110011110000000_1011011010001100"; -- -0.09569224446008652
	pesos_i(23645) := b"1111111111111111_1111111111111111_1101111010111110_1000001000011101"; -- -0.12990557468444294
	pesos_i(23646) := b"1111111111111111_1111111111111111_1110001000001010_0001100101100010"; -- -0.11703339921639966
	pesos_i(23647) := b"1111111111111111_1111111111111111_1110100100100001_0000100100111101"; -- -0.08933965920932148
	pesos_i(23648) := b"1111111111111111_1111111111111111_1101111010010110_1001110101011101"; -- -0.13051430203993644
	pesos_i(23649) := b"0000000000000000_0000000000000000_0010000011101000_1000011001111011"; -- 0.12854805478805856
	pesos_i(23650) := b"1111111111111111_1111111111111111_1110000010001110_0101001110101010"; -- -0.1228282652877232
	pesos_i(23651) := b"1111111111111111_1111111111111111_1111100100010001_1001001010111110"; -- -0.027075604012354614
	pesos_i(23652) := b"0000000000000000_0000000000000000_0000001010011001_0100101111111010"; -- 0.010151623341079835
	pesos_i(23653) := b"1111111111111111_1111111111111111_1110100100000111_0101000011110001"; -- -0.08973211405229664
	pesos_i(23654) := b"0000000000000000_0000000000000000_0001101110010011_1010110010110001"; -- 0.10772208512804238
	pesos_i(23655) := b"0000000000000000_0000000000000000_0001100010111010_1111011011010011"; -- 0.09660284662568641
	pesos_i(23656) := b"1111111111111111_1111111111111111_1101101100001100_0011010111010000"; -- -0.14434493707412477
	pesos_i(23657) := b"0000000000000000_0000000000000000_0001010101101011_0011000100000101"; -- 0.08366686223718503
	pesos_i(23658) := b"1111111111111111_1111111111111111_1101100000101011_1000101101111011"; -- -0.15558555840236346
	pesos_i(23659) := b"0000000000000000_0000000000000000_0000110011011001_1100000110111000"; -- 0.05019770368717758
	pesos_i(23660) := b"0000000000000000_0000000000000000_0010000101011001_1011001011000110"; -- 0.1302749379959354
	pesos_i(23661) := b"0000000000000000_0000000000000000_0001111000011110_0011110010111011"; -- 0.11764888351991866
	pesos_i(23662) := b"1111111111111111_1111111111111111_1111101101000111_0111001101110110"; -- -0.01844099405317512
	pesos_i(23663) := b"0000000000000000_0000000000000000_0000101101010110_1111111010011010"; -- 0.04429618132387249
	pesos_i(23664) := b"1111111111111111_1111111111111111_1110101011010111_0010101010110010"; -- -0.082654315604873
	pesos_i(23665) := b"1111111111111111_1111111111111111_1111001010111111_1000010110010111"; -- -0.05176510880377144
	pesos_i(23666) := b"1111111111111111_1111111111111111_1111000001110101_1111110010011010"; -- -0.06069966537436744
	pesos_i(23667) := b"1111111111111111_1111111111111111_1110110010000101_0100100010101010"; -- -0.076091249933024
	pesos_i(23668) := b"0000000000000000_0000000000000000_0010001101010100_1111001011000100"; -- 0.13801495828028837
	pesos_i(23669) := b"0000000000000000_0000000000000000_0010001011010001_1000001011011000"; -- 0.13600938579950078
	pesos_i(23670) := b"0000000000000000_0000000000000000_0010001010011100_0101101010010010"; -- 0.13519826953273453
	pesos_i(23671) := b"1111111111111111_1111111111111111_1101111101101110_0111100101010111"; -- -0.1272205507528845
	pesos_i(23672) := b"1111111111111111_1111111111111111_1101100101101111_1100000000010010"; -- -0.15063857622235727
	pesos_i(23673) := b"1111111111111111_1111111111111111_1110010011101100_0110110110101000"; -- -0.10576738970055674
	pesos_i(23674) := b"0000000000000000_0000000000000000_0000110001010001_0000010010001101"; -- 0.048111233053806934
	pesos_i(23675) := b"1111111111111111_1111111111111111_1110101010110010_0011010001001111"; -- -0.08321831773334616
	pesos_i(23676) := b"1111111111111111_1111111111111111_1111011010000110_1001100010100100"; -- -0.037008724168499416
	pesos_i(23677) := b"0000000000000000_0000000000000000_0000110011110010_0100010001101011"; -- 0.050571705097767844
	pesos_i(23678) := b"1111111111111111_1111111111111111_1110010111010100_0110101110101110"; -- -0.10222746851788189
	pesos_i(23679) := b"0000000000000000_0000000000000000_0010010000101010_0111100110000110"; -- 0.14127311245261234
	pesos_i(23680) := b"0000000000000000_0000000000000000_0000110100101111_0010111010000101"; -- 0.051501185893868505
	pesos_i(23681) := b"1111111111111111_1111111111111111_1111101100011010_0100110110111110"; -- -0.019129887723154066
	pesos_i(23682) := b"0000000000000000_0000000000000000_0001011001101010_0010111011000100"; -- 0.08755771911575987
	pesos_i(23683) := b"1111111111111111_1111111111111111_1110010100110010_1100110111111011"; -- -0.10469353305167975
	pesos_i(23684) := b"0000000000000000_0000000000000000_0000111111001010_1100111001100011"; -- 0.061688326944025436
	pesos_i(23685) := b"0000000000000000_0000000000000000_0001100001000010_1000000110111110"; -- 0.0947648133178812
	pesos_i(23686) := b"0000000000000000_0000000000000000_0010011100100001_0101111010000110"; -- 0.15285292411315066
	pesos_i(23687) := b"0000000000000000_0000000000000000_0001110001000001_1001101010001100"; -- 0.11037603311274999
	pesos_i(23688) := b"0000000000000000_0000000000000000_0001001000001101_0111110001111011"; -- 0.07051828386618293
	pesos_i(23689) := b"0000000000000000_0000000000000000_0000001001010001_1011101010011000"; -- 0.009059583730073525
	pesos_i(23690) := b"0000000000000000_0000000000000000_0001101000001010_1000100101010011"; -- 0.10172327301740469
	pesos_i(23691) := b"0000000000000000_0000000000000000_0010011100010000_1111111010001100"; -- 0.1526030628574247
	pesos_i(23692) := b"1111111111111111_1111111111111111_1111100101110000_1001101111000101"; -- -0.02562548095012838
	pesos_i(23693) := b"0000000000000000_0000000000000000_0001000001010110_1010101101001100"; -- 0.06382246603196043
	pesos_i(23694) := b"0000000000000000_0000000000000000_0000101010011110_0000010100001111"; -- 0.04147369023740308
	pesos_i(23695) := b"0000000000000000_0000000000000000_0000101001100110_1110000010110111"; -- 0.04063229046455154
	pesos_i(23696) := b"1111111111111111_1111111111111111_1111100010011100_1101110100101011"; -- -0.028856446331079293
	pesos_i(23697) := b"1111111111111111_1111111111111111_1110110010011010_0001001110110111"; -- -0.07577397129064159
	pesos_i(23698) := b"1111111111111111_1111111111111111_1111111110100010_0001000111110101"; -- -0.0014332559168799507
	pesos_i(23699) := b"1111111111111111_1111111111111111_1110100111011010_1010111010000100"; -- -0.08650693211452636
	pesos_i(23700) := b"1111111111111111_1111111111111111_1110000100110001_1101111011110100"; -- -0.12033278038886625
	pesos_i(23701) := b"1111111111111111_1111111111111111_1110000100010010_0110101011001001"; -- -0.12081272694139356
	pesos_i(23702) := b"0000000000000000_0000000000000000_0001001111001001_1101000100110001"; -- 0.07729823537757072
	pesos_i(23703) := b"1111111111111111_1111111111111111_1111100011001010_1111110110100111"; -- -0.02815260568925706
	pesos_i(23704) := b"1111111111111111_1111111111111111_1110101100110011_0001101000001111"; -- -0.08125149847229352
	pesos_i(23705) := b"1111111111111111_1111111111111111_1110111101010001_0010010111111110"; -- -0.06516802361212978
	pesos_i(23706) := b"1111111111111111_1111111111111111_1101110001100110_0010011100111011"; -- -0.13906626515107062
	pesos_i(23707) := b"0000000000000000_0000000000000000_0010000011001100_1001100111001111"; -- 0.12812196076823507
	pesos_i(23708) := b"1111111111111111_1111111111111111_1110001100001001_0111001010111001"; -- -0.11313708283306359
	pesos_i(23709) := b"0000000000000000_0000000000000000_0000110010000000_0011000100110001"; -- 0.048831056960094085
	pesos_i(23710) := b"1111111111111111_1111111111111111_1111110010001110_0011110101101011"; -- -0.01345459121147959
	pesos_i(23711) := b"1111111111111111_1111111111111111_1111001001100000_1001011110000000"; -- -0.0532136262365728
	pesos_i(23712) := b"1111111111111111_1111111111111111_1101100100110100_1101111010111000"; -- -0.15153701799081606
	pesos_i(23713) := b"0000000000000000_0000000000000000_0010010001010001_0001111000101001"; -- 0.14186275953149546
	pesos_i(23714) := b"1111111111111111_1111111111111111_1110110011000111_0101001100001001"; -- -0.07508355160277147
	pesos_i(23715) := b"0000000000000000_0000000000000000_0001111001111000_1010100100111101"; -- 0.11902864208002228
	pesos_i(23716) := b"0000000000000000_0000000000000000_0001000110000100_1010000001011101"; -- 0.06842996862729833
	pesos_i(23717) := b"1111111111111111_1111111111111111_1101001100011110_0001011110100101"; -- -0.1753220770239819
	pesos_i(23718) := b"0000000000000000_0000000000000000_0010010011100100_0001010111100110"; -- 0.14410530909705205
	pesos_i(23719) := b"0000000000000000_0000000000000000_0000000110100111_0100101001010110"; -- 0.006458898460694394
	pesos_i(23720) := b"1111111111111111_1111111111111111_1110110111101101_1101100101110100"; -- -0.07058945580920388
	pesos_i(23721) := b"0000000000000000_0000000000000000_0001010110111010_0101001001001011"; -- 0.08487428969846686
	pesos_i(23722) := b"0000000000000000_0000000000000000_0001100000101011_1010011101010011"; -- 0.09441610124948553
	pesos_i(23723) := b"0000000000000000_0000000000000000_0000110001100111_1110000000001010"; -- 0.048460009134917895
	pesos_i(23724) := b"1111111111111111_1111111111111111_1110111110101101_1100011011011101"; -- -0.06375462626647231
	pesos_i(23725) := b"0000000000000000_0000000000000000_0000111100101101_0011101100011000"; -- 0.059283917654940975
	pesos_i(23726) := b"0000000000000000_0000000000000000_0000100011110101_1010111011110110"; -- 0.034998831709794155
	pesos_i(23727) := b"1111111111111111_1111111111111111_1111110110101100_1111001110100011"; -- -0.009079716487455028
	pesos_i(23728) := b"0000000000000000_0000000000000000_0001101100001111_1110110010100110"; -- 0.10571173719302976
	pesos_i(23729) := b"1111111111111111_1111111111111111_1111111111000100_1001011010100010"; -- -0.0009065490265777311
	pesos_i(23730) := b"0000000000000000_0000000000000000_0000111001010111_0111000000000011"; -- 0.056021691073534205
	pesos_i(23731) := b"1111111111111111_1111111111111111_1101111100101010_0101011110111110"; -- -0.1282601510145457
	pesos_i(23732) := b"0000000000000000_0000000000000000_0001000101110010_1101010110100000"; -- 0.06815848498449983
	pesos_i(23733) := b"1111111111111111_1111111111111111_1110011001001111_0000000001101000"; -- -0.10035703154065909
	pesos_i(23734) := b"1111111111111111_1111111111111111_1111101100111010_1101110011111101"; -- -0.018633068418818878
	pesos_i(23735) := b"0000000000000000_0000000000000000_0001001001111001_1010110001101001"; -- 0.07216908989195513
	pesos_i(23736) := b"1111111111111111_1111111111111111_1101111110010110_0101100110000110"; -- -0.12661209552244357
	pesos_i(23737) := b"1111111111111111_1111111111111111_1111011110100000_1001101000111001"; -- -0.032705651315523304
	pesos_i(23738) := b"1111111111111111_1111111111111111_1101101010110100_0010110001001111"; -- -0.14568827702685191
	pesos_i(23739) := b"0000000000000000_0000000000000000_0000101001010110_1110111100000010"; -- 0.040389001837743195
	pesos_i(23740) := b"1111111111111111_1111111111111111_1111001010010011_1001100000110000"; -- -0.05243538692541619
	pesos_i(23741) := b"0000000000000000_0000000000000000_0010001010111001_1100110001101111"; -- 0.13564756123646482
	pesos_i(23742) := b"0000000000000000_0000000000000000_0010100110101101_1111101010000101"; -- 0.1628109527135378
	pesos_i(23743) := b"1111111111111111_1111111111111111_1101011000011111_1110001111111011"; -- -0.16357588873616058
	pesos_i(23744) := b"0000000000000000_0000000000000000_0001110011111011_1011111011001101"; -- 0.11321632871391615
	pesos_i(23745) := b"0000000000000000_0000000000000000_0001110101001101_0110011100100011"; -- 0.11446232421206033
	pesos_i(23746) := b"0000000000000000_0000000000000000_0001100000101110_0011100000110100"; -- 0.09445525423734245
	pesos_i(23747) := b"0000000000000000_0000000000000000_0001001100110100_0011111011011000"; -- 0.07501595273605473
	pesos_i(23748) := b"1111111111111111_1111111111111111_1111101010111101_0110101100101011"; -- -0.020547201150987966
	pesos_i(23749) := b"1111111111111111_1111111111111111_1101100000110011_1111011000111100"; -- -0.15545712499036574
	pesos_i(23750) := b"1111111111111111_1111111111111111_1111110110011000_0111110101100100"; -- -0.009391940206273193
	pesos_i(23751) := b"1111111111111111_1111111111111111_1110001101101110_1110100010010010"; -- -0.111588920909915
	pesos_i(23752) := b"0000000000000000_0000000000000000_0010010010101100_1110111011011011"; -- 0.1432637487219354
	pesos_i(23753) := b"0000000000000000_0000000000000000_0000010101010100_0101101010110111"; -- 0.020818395323646845
	pesos_i(23754) := b"1111111111111111_1111111111111111_1111011011101110_1001010100101011"; -- -0.03542201714383692
	pesos_i(23755) := b"0000000000000000_0000000000000000_0010000101001101_1000010111111110"; -- 0.1300891633044523
	pesos_i(23756) := b"1111111111111111_1111111111111111_1111011000101011_1010010101001001"; -- -0.03839652040039214
	pesos_i(23757) := b"0000000000000000_0000000000000000_0000100001111101_0111101110010000"; -- 0.03316471342919088
	pesos_i(23758) := b"0000000000000000_0000000000000000_0001110100000101_0111101010000100"; -- 0.11336484650690853
	pesos_i(23759) := b"0000000000000000_0000000000000000_0001001001101101_1110001011111101"; -- 0.07198923759700733
	pesos_i(23760) := b"1111111111111111_1111111111111111_1111011101101110_0111101010010101"; -- -0.03347047663714975
	pesos_i(23761) := b"1111111111111111_1111111111111111_1110100000100000_0001001110001101"; -- -0.09326055343299613
	pesos_i(23762) := b"0000000000000000_0000000000000000_0000110010110100_1101101000111101"; -- 0.049634590078915734
	pesos_i(23763) := b"1111111111111111_1111111111111111_1111100110011101_1101001101111001"; -- -0.02493551535747133
	pesos_i(23764) := b"1111111111111111_1111111111111111_1111000011101011_1011001000110100"; -- -0.05890356293471611
	pesos_i(23765) := b"1111111111111111_1111111111111111_1111010000100111_1111011110011000"; -- -0.04626514945945316
	pesos_i(23766) := b"0000000000000000_0000000000000000_0001001100101011_0100101011000100"; -- 0.07487933425789266
	pesos_i(23767) := b"1111111111111111_1111111111111111_1101100110000000_1011001110011110"; -- -0.15037991899523834
	pesos_i(23768) := b"0000000000000000_0000000000000000_0010011100101001_1011011101111010"; -- 0.152980296481341
	pesos_i(23769) := b"0000000000000000_0000000000000000_0001000000000011_1011011101010110"; -- 0.06255670395912113
	pesos_i(23770) := b"0000000000000000_0000000000000000_0010001000000111_1111110100011001"; -- 0.1329343972345355
	pesos_i(23771) := b"1111111111111111_1111111111111111_1111001111110101_0001100110111101"; -- -0.04704131261974475
	pesos_i(23772) := b"1111111111111111_1111111111111111_1101100010101101_1100110100011110"; -- -0.15359800357694456
	pesos_i(23773) := b"1111111111111111_1111111111111111_1101011010001000_0111110001100011"; -- -0.16197989059486106
	pesos_i(23774) := b"0000000000000000_0000000000000000_0001100100011100_1010111001010110"; -- 0.09809388725263304
	pesos_i(23775) := b"1111111111111111_1111111111111111_1111011010000000_0011011011100001"; -- -0.03710610386923358
	pesos_i(23776) := b"0000000000000000_0000000000000000_0000110101010010_1111110011010000"; -- 0.05204753946030723
	pesos_i(23777) := b"0000000000000000_0000000000000000_0000000010001001_1100110110100100"; -- 0.002102711226205941
	pesos_i(23778) := b"1111111111111111_1111111111111111_1110011011100000_0011111000110111"; -- -0.09814082304831412
	pesos_i(23779) := b"1111111111111111_1111111111111111_1110001000111011_0111000110011000"; -- -0.11628046066714284
	pesos_i(23780) := b"0000000000000000_0000000000000000_0001001001000011_1111111000001100"; -- 0.07134998113503999
	pesos_i(23781) := b"1111111111111111_1111111111111111_1110001000000100_0010001110011000"; -- -0.11712434320701477
	pesos_i(23782) := b"1111111111111111_1111111111111111_1101111101010100_0100011000001100"; -- -0.12762033658910193
	pesos_i(23783) := b"1111111111111111_1111111111111111_1110011110111111_1001100001010000"; -- -0.09473274267732823
	pesos_i(23784) := b"1111111111111111_1111111111111111_1101111111100101_0110000101001010"; -- -0.1254061884314252
	pesos_i(23785) := b"1111111111111111_1111111111111111_1111101101110011_1110101011011010"; -- -0.01776249093306181
	pesos_i(23786) := b"1111111111111111_1111111111111111_1110000000101110_1111110010011010"; -- -0.12428303942162494
	pesos_i(23787) := b"0000000000000000_0000000000000000_0010001100011001_0101011010001111"; -- 0.13710537907311304
	pesos_i(23788) := b"0000000000000000_0000000000000000_0001001011011100_0110011100001111"; -- 0.07367557639269251
	pesos_i(23789) := b"0000000000000000_0000000000000000_0010000100011111_1111001111011110"; -- 0.12939380812027543
	pesos_i(23790) := b"0000000000000000_0000000000000000_0001011101001011_0011001111111011"; -- 0.0909912574623453
	pesos_i(23791) := b"0000000000000000_0000000000000000_0000001010100101_1111011101100110"; -- 0.010344946305489492
	pesos_i(23792) := b"0000000000000000_0000000000000000_0000111100101010_0100001011010111"; -- 0.059238603158900824
	pesos_i(23793) := b"1111111111111111_1111111111111111_1110010101011101_0101010111011001"; -- -0.10404456560749861
	pesos_i(23794) := b"0000000000000000_0000000000000000_0001101001010100_1101100111111110"; -- 0.10285723157189618
	pesos_i(23795) := b"1111111111111111_1111111111111111_1110010100000101_1101110000000101"; -- -0.10537934193377096
	pesos_i(23796) := b"1111111111111111_1111111111111111_1101101110100010_0111110111110001"; -- -0.14205181950812437
	pesos_i(23797) := b"1111111111111111_1111111111111111_1111001010011100_0111101111100100"; -- -0.052299744381705815
	pesos_i(23798) := b"1111111111111111_1111111111111111_1101101110001000_1011010101011100"; -- -0.1424452447109224
	pesos_i(23799) := b"1111111111111111_1111111111111111_1111001011001101_1101111111111111"; -- -0.051546097150094804
	pesos_i(23800) := b"1111111111111111_1111111111111111_1111000010100111_1111010110111000"; -- -0.05993713619432598
	pesos_i(23801) := b"0000000000000000_0000000000000000_0010001101010111_0110100001110001"; -- 0.1380524898498349
	pesos_i(23802) := b"1111111111111111_1111111111111111_1110011111001111_0101011100011011"; -- -0.09449248887019615
	pesos_i(23803) := b"0000000000000000_0000000000000000_0001111110101000_1000100111001001"; -- 0.12366543911043675
	pesos_i(23804) := b"1111111111111111_1111111111111111_1110011001011011_0010010000100001"; -- -0.100171796782957
	pesos_i(23805) := b"1111111111111111_1111111111111111_1110010101000001_0101000001100000"; -- -0.1044721378917686
	pesos_i(23806) := b"1111111111111111_1111111111111111_1111001000011111_0100100100000011"; -- -0.054210125774514784
	pesos_i(23807) := b"0000000000000000_0000000000000000_0001110111110110_1100010000110111"; -- 0.11704660753607882
	pesos_i(23808) := b"0000000000000000_0000000000000000_0000101101011110_1011101110000001"; -- 0.04441425237265906
	pesos_i(23809) := b"1111111111111111_1111111111111111_1111111001001100_0111000101001110"; -- -0.006646078542847842
	pesos_i(23810) := b"0000000000000000_0000000000000000_0001100100111100_1010000111001101"; -- 0.09858142144987778
	pesos_i(23811) := b"0000000000000000_0000000000000000_0000001001101011_1000101001110111"; -- 0.009453443464046064
	pesos_i(23812) := b"0000000000000000_0000000000000000_0010001111001111_0010011101001100"; -- 0.13987966153072795
	pesos_i(23813) := b"1111111111111111_1111111111111111_1111001110011010_1110100111111000"; -- -0.04841745084646635
	pesos_i(23814) := b"0000000000000000_0000000000000000_0001100110001110_0000111001010010"; -- 0.09982385160127326
	pesos_i(23815) := b"0000000000000000_0000000000000000_0000011010010011_0101001010011001"; -- 0.02568546522774054
	pesos_i(23816) := b"0000000000000000_0000000000000000_0000010101001001_1100111011001111"; -- 0.020657468439012026
	pesos_i(23817) := b"0000000000000000_0000000000000000_0010001111001011_0001110000100110"; -- 0.13981796202519955
	pesos_i(23818) := b"0000000000000000_0000000000000000_0010001101001001_0101101001001101"; -- 0.13783802393302877
	pesos_i(23819) := b"1111111111111111_1111111111111111_1110001100101101_0011010011010010"; -- -0.11259145606750082
	pesos_i(23820) := b"1111111111111111_1111111111111111_1111000101100001_0110110000100011"; -- -0.05710720204219876
	pesos_i(23821) := b"0000000000000000_0000000000000000_0010001101110011_1010001100111101"; -- 0.13848324048033855
	pesos_i(23822) := b"1111111111111111_1111111111111111_1110101100100000_0011011110010100"; -- -0.08153965612682708
	pesos_i(23823) := b"1111111111111111_1111111111111111_1111101001011010_1101001111111100"; -- -0.022051573747778812
	pesos_i(23824) := b"1111111111111111_1111111111111111_1110001000011110_0010111101111001"; -- -0.11672690664102113
	pesos_i(23825) := b"0000000000000000_0000000000000000_0001001000100111_1001000111001110"; -- 0.07091628335049689
	pesos_i(23826) := b"1111111111111111_1111111111111111_1111000101100101_1110101100101000"; -- -0.057038595845693235
	pesos_i(23827) := b"0000000000000000_0000000000000000_0001101001010000_0010011001110011"; -- 0.10278549478218689
	pesos_i(23828) := b"1111111111111111_1111111111111111_1111010001101100_1111101011101001"; -- -0.045212095321087456
	pesos_i(23829) := b"0000000000000000_0000000000000000_0000001111000000_1110011100101111"; -- 0.014662217185044008
	pesos_i(23830) := b"1111111111111111_1111111111111111_1101101010011101_1011001011000100"; -- -0.1460312148019686
	pesos_i(23831) := b"0000000000000000_0000000000000000_0010000010101011_0001100100000111"; -- 0.12761074463048247
	pesos_i(23832) := b"1111111111111111_1111111111111111_1111101001101000_1001010011011000"; -- -0.021841714195013864
	pesos_i(23833) := b"1111111111111111_1111111111111111_1111100110010110_0101100000001101"; -- -0.025049683403567335
	pesos_i(23834) := b"1111111111111111_1111111111111111_1111010010010011_1000100110001001"; -- -0.04462376030459436
	pesos_i(23835) := b"0000000000000000_0000000000000000_0001101100001100_0010100001001010"; -- 0.1056542567812504
	pesos_i(23836) := b"0000000000000000_0000000000000000_0001001001100010_1011000001100011"; -- 0.0718183747309701
	pesos_i(23837) := b"1111111111111111_1111111111111111_1110010111000001_1001110000110010"; -- -0.10251449384324277
	pesos_i(23838) := b"1111111111111111_1111111111111111_1110001111110100_0000001100110001"; -- -0.10955791519794025
	pesos_i(23839) := b"1111111111111111_1111111111111111_1111100010100001_1011100110010100"; -- -0.02878227366996085
	pesos_i(23840) := b"1111111111111111_1111111111111111_1111000101000101_1101001100000011"; -- -0.0575283163366814
	pesos_i(23841) := b"0000000000000000_0000000000000000_0000010101111001_0010001100001100"; -- 0.021379652483914147
	pesos_i(23842) := b"1111111111111111_1111111111111111_1111010010110110_0000101101100000"; -- -0.044097222313653664
	pesos_i(23843) := b"0000000000000000_0000000000000000_0000000111111100_1101111110011100"; -- 0.007764793023439129
	pesos_i(23844) := b"1111111111111111_1111111111111111_1111000011010110_1100111101011110"; -- -0.059222259102680884
	pesos_i(23845) := b"1111111111111111_1111111111111111_1110111011101011_0111100010001011"; -- -0.06671949963016269
	pesos_i(23846) := b"0000000000000000_0000000000000000_0001010000111110_1111010101001001"; -- 0.07908566496651641
	pesos_i(23847) := b"1111111111111111_1111111111111111_1101111001011111_1010001011101011"; -- -0.13135320434258307
	pesos_i(23848) := b"1111111111111111_1111111111111111_1101111110111100_1000010010000010"; -- -0.1260296996102522
	pesos_i(23849) := b"1111111111111111_1111111111111111_1110011111101100_1101100001000001"; -- -0.0940422860443451
	pesos_i(23850) := b"0000000000000000_0000000000000000_0010010010110110_1111101101100011"; -- 0.14341708353235122
	pesos_i(23851) := b"1111111111111111_1111111111111111_1111100101110110_0101110101100110"; -- -0.02553764589927097
	pesos_i(23852) := b"0000000000000000_0000000000000000_0010010011010010_1100010101010011"; -- 0.14384110715645232
	pesos_i(23853) := b"1111111111111111_1111111111111111_1111000101000010_0101000110110011"; -- -0.057581800222393044
	pesos_i(23854) := b"1111111111111111_1111111111111111_1111101000101000_0110010111000111"; -- -0.022821081953058604
	pesos_i(23855) := b"0000000000000000_0000000000000000_0000011000100111_1010110010110010"; -- 0.024042886249073997
	pesos_i(23856) := b"1111111111111111_1111111111111111_1110011111100010_1111101111111100"; -- -0.09419274429993502
	pesos_i(23857) := b"1111111111111111_1111111111111111_1110101111110110_1011001111011101"; -- -0.07826686727412384
	pesos_i(23858) := b"1111111111111111_1111111111111111_1110000100101001_0110101011001010"; -- -0.1204617744890403
	pesos_i(23859) := b"1111111111111111_1111111111111111_1101110110011101_0111011000100011"; -- -0.13431607868337503
	pesos_i(23860) := b"1111111111111111_1111111111111111_1111100100100110_0111011001110010"; -- -0.02675685614838792
	pesos_i(23861) := b"1111111111111111_1111111111111111_1111001011110011_1011111110011000"; -- -0.05096819447873778
	pesos_i(23862) := b"0000000000000000_0000000000000000_0000010001111110_0101101100101001"; -- 0.017553041104083723
	pesos_i(23863) := b"1111111111111111_1111111111111111_1111000011111001_0001110001001011"; -- -0.05869887522317661
	pesos_i(23864) := b"1111111111111111_1111111111111111_1110001011100010_1010010011011001"; -- -0.11372918807530828
	pesos_i(23865) := b"0000000000000000_0000000000000000_0000101000110001_1110010100000110"; -- 0.039823831566632696
	pesos_i(23866) := b"1111111111111111_1111111111111111_1111010000000111_1011011101111110"; -- -0.046757251461118914
	pesos_i(23867) := b"1111111111111111_1111111111111111_1111000000011110_1010111111100100"; -- -0.062031752446510206
	pesos_i(23868) := b"1111111111111111_1111111111111111_1110001110110110_0000001100111100"; -- -0.11050395750641688
	pesos_i(23869) := b"1111111111111111_1111111111111111_1110011111100011_0110101100111111"; -- -0.09418611249549218
	pesos_i(23870) := b"0000000000000000_0000000000000000_0000001000011110_1011101101010111"; -- 0.00828143000267983
	pesos_i(23871) := b"1111111111111111_1111111111111111_1110010110110000_1011110101011111"; -- -0.1027719156539336
	pesos_i(23872) := b"0000000000000000_0000000000000000_0000010001100111_1111100010100000"; -- 0.017211474438473123
	pesos_i(23873) := b"1111111111111111_1111111111111111_1110001000001001_0111010001011100"; -- -0.1170432353454189
	pesos_i(23874) := b"1111111111111111_1111111111111111_1101111111111100_0001000010110101"; -- -0.12506003940223517
	pesos_i(23875) := b"0000000000000000_0000000000000000_0010010000110010_1111100000101100"; -- 0.14140273168069115
	pesos_i(23876) := b"1111111111111111_1111111111111111_1111001010011111_1010110010110111"; -- -0.0522510579730063
	pesos_i(23877) := b"0000000000000000_0000000000000000_0000011100010011_1100100100100110"; -- 0.027645656438800553
	pesos_i(23878) := b"0000000000000000_0000000000000000_0000010101000111_0001001001000100"; -- 0.020615712652874565
	pesos_i(23879) := b"0000000000000000_0000000000000000_0010011000110011_1100101110111010"; -- 0.14922784119989593
	pesos_i(23880) := b"0000000000000000_0000000000000000_0001010001100011_1110010010110011"; -- 0.07964925171418558
	pesos_i(23881) := b"1111111111111111_1111111111111111_1110101000100110_0001100001101111"; -- -0.08535620958726559
	pesos_i(23882) := b"0000000000000000_0000000000000000_0000111111111100_1100110000101000"; -- 0.06245113348875401
	pesos_i(23883) := b"1111111111111111_1111111111111111_1110111011000000_0101000101100010"; -- -0.06737796169951978
	pesos_i(23884) := b"1111111111111111_1111111111111111_1110000000010011_1001011110000001"; -- -0.12470105266235725
	pesos_i(23885) := b"1111111111111111_1111111111111111_1111001101101110_1001010011101000"; -- -0.04909390760752144
	pesos_i(23886) := b"0000000000000000_0000000000000000_0000011100010110_0010010011010000"; -- 0.027681637476155763
	pesos_i(23887) := b"0000000000000000_0000000000000000_0000011101100111_1011100110001000"; -- 0.028926463726263386
	pesos_i(23888) := b"0000000000000000_0000000000000000_0010001101010100_0010101000010101"; -- 0.13800299659788054
	pesos_i(23889) := b"1111111111111111_1111111111111111_1111000000001010_0011110100011100"; -- -0.062343769672178556
	pesos_i(23890) := b"1111111111111111_1111111111111111_1110010111101100_1101000000000100"; -- -0.10185527719207572
	pesos_i(23891) := b"0000000000000000_0000000000000000_0001111110011010_1101110001111101"; -- 0.1234567456719041
	pesos_i(23892) := b"0000000000000000_0000000000000000_0000101001001010_0011110111010101"; -- 0.040195335777791406
	pesos_i(23893) := b"1111111111111111_1111111111111111_1110000001001110_0110111101100111"; -- -0.12380317441443894
	pesos_i(23894) := b"0000000000000000_0000000000000000_0000111011110110_1001110100011101"; -- 0.05845052679431937
	pesos_i(23895) := b"0000000000000000_0000000000000000_0000100000100101_0001100011100101"; -- 0.03181605896709774
	pesos_i(23896) := b"1111111111111111_1111111111111111_1110101100011101_0100001001100000"; -- -0.08158478896952709
	pesos_i(23897) := b"1111111111111111_1111111111111111_1111010011100100_0100001010101101"; -- -0.043392021978453175
	pesos_i(23898) := b"0000000000000000_0000000000000000_0001100100001100_0011110011001100"; -- 0.09784297923632083
	pesos_i(23899) := b"1111111111111111_1111111111111111_1110110010011110_0101111110111001"; -- -0.07570840588751007
	pesos_i(23900) := b"0000000000000000_0000000000000000_0001000011111101_0000011010011011"; -- 0.0663608673385131
	pesos_i(23901) := b"1111111111111111_1111111111111111_1101011001111110_1001111100000100"; -- -0.1621304145841233
	pesos_i(23902) := b"0000000000000000_0000000000000000_0000001100010010_1000011101110001"; -- 0.012001481076341455
	pesos_i(23903) := b"1111111111111111_1111111111111111_1110100001000110_0001001111110010"; -- -0.092680695919286
	pesos_i(23904) := b"0000000000000000_0000000000000000_0010000011001010_0011000101101100"; -- 0.12808522118989174
	pesos_i(23905) := b"1111111111111111_1111111111111111_1111001010000111_1100111000101100"; -- -0.052615274747567276
	pesos_i(23906) := b"1111111111111111_1111111111111111_1101111011101110_1011101010010101"; -- -0.12916978712082378
	pesos_i(23907) := b"1111111111111111_1111111111111111_1111101110010111_1000001101011100"; -- -0.017219343235184474
	pesos_i(23908) := b"0000000000000000_0000000000000000_0001101000111111_1001101010001001"; -- 0.10253301470636969
	pesos_i(23909) := b"0000000000000000_0000000000000000_0001110100110001_1011111011001111"; -- 0.11404030381755281
	pesos_i(23910) := b"0000000000000000_0000000000000000_0001010000111010_0101111011001010"; -- 0.079015659560823
	pesos_i(23911) := b"1111111111111111_1111111111111111_1111001111111111_1001000110010011"; -- -0.04688158179280355
	pesos_i(23912) := b"1111111111111111_1111111111111111_1111010000111100_1101101001101100"; -- -0.045946453601600164
	pesos_i(23913) := b"1111111111111111_1111111111111111_1111111011101001_1000010010111011"; -- -0.004249290735310446
	pesos_i(23914) := b"0000000000000000_0000000000000000_0010010000101100_0000100111100010"; -- 0.14129697583277054
	pesos_i(23915) := b"1111111111111111_1111111111111111_1101111110100001_0100111111100110"; -- -0.12644482269400836
	pesos_i(23916) := b"0000000000000000_0000000000000000_0010001001001110_0011111101100010"; -- 0.1340064634238035
	pesos_i(23917) := b"1111111111111111_1111111111111111_1111000101101000_1011010101000010"; -- -0.05699603213641455
	pesos_i(23918) := b"0000000000000000_0000000000000000_0000001110000101_1010001010110100"; -- 0.013757866919838246
	pesos_i(23919) := b"1111111111111111_1111111111111111_1111100111010111_1010000000110110"; -- -0.02405356099560813
	pesos_i(23920) := b"1111111111111111_1111111111111111_1110001110011111_0111001100110110"; -- -0.11084823532961936
	pesos_i(23921) := b"0000000000000000_0000000000000000_0000101101011011_0000111011101101"; -- 0.04435818953116063
	pesos_i(23922) := b"0000000000000000_0000000000000000_0001001001111110_0000110101001110"; -- 0.07223590040173945
	pesos_i(23923) := b"0000000000000000_0000000000000000_0001110110000010_1011010100111000"; -- 0.11527569404293009
	pesos_i(23924) := b"1111111111111111_1111111111111111_1110101111010101_1011000000101010"; -- -0.07877062783581731
	pesos_i(23925) := b"1111111111111111_1111111111111111_1111110010001011_1100110001011101"; -- -0.013491847382803098
	pesos_i(23926) := b"0000000000000000_0000000000000000_0000011101101010_0111110110000110"; -- 0.028968663339115144
	pesos_i(23927) := b"1111111111111111_1111111111111111_1111110010001101_1101101011010001"; -- -0.013460468345847448
	pesos_i(23928) := b"0000000000000000_0000000000000000_0001111010000101_0100011001011101"; -- 0.11922111299909291
	pesos_i(23929) := b"1111111111111111_1111111111111111_1110111111010001_0101111111010101"; -- -0.0632114510842286
	pesos_i(23930) := b"0000000000000000_0000000000000000_0001011111000101_0000011111100100"; -- 0.09285020181212712
	pesos_i(23931) := b"1111111111111111_1111111111111111_1111111011000000_1110110101100110"; -- -0.0048686625563027245
	pesos_i(23932) := b"0000000000000000_0000000000000000_0000000100110011_1011100100101111"; -- 0.004695486048319379
	pesos_i(23933) := b"0000000000000000_0000000000000000_0001010000101101_1010110101100110"; -- 0.07882198094344774
	pesos_i(23934) := b"1111111111111111_1111111111111111_1111111100100111_1111110011100100"; -- -0.0032960836815740004
	pesos_i(23935) := b"1111111111111111_1111111111111111_1111100011101101_1010001010010110"; -- -0.0276239760580709
	pesos_i(23936) := b"0000000000000000_0000000000000000_0000001101111001_1101000101101011"; -- 0.013577545870677221
	pesos_i(23937) := b"1111111111111111_1111111111111111_1110100001110110_1000010100111010"; -- -0.09194152203528841
	pesos_i(23938) := b"1111111111111111_1111111111111111_1110010111100101_1001000011010001"; -- -0.10196585560175703
	pesos_i(23939) := b"0000000000000000_0000000000000000_0000011000000101_1111110111110010"; -- 0.02352893023318408
	pesos_i(23940) := b"1111111111111111_1111111111111111_1101011001000001_0110101000010011"; -- -0.163064356197197
	pesos_i(23941) := b"1111111111111111_1111111111111111_1101111110001110_0100001011011000"; -- -0.12673551771871291
	pesos_i(23942) := b"0000000000000000_0000000000000000_0000110100011010_0000000001001011"; -- 0.0511779958724692
	pesos_i(23943) := b"0000000000000000_0000000000000000_0001010000101101_0000000101100010"; -- 0.07881172802341285
	pesos_i(23944) := b"0000000000000000_0000000000000000_0000110101101001_0010010110011000"; -- 0.052385663566768825
	pesos_i(23945) := b"0000000000000000_0000000000000000_0001011000101101_1010010110000110"; -- 0.08663401151689334
	pesos_i(23946) := b"1111111111111111_1111111111111111_1110000111001100_1101010110101100"; -- -0.1179682212275484
	pesos_i(23947) := b"0000000000000000_0000000000000000_0001101000010000_0101110110011110"; -- 0.10181222052981567
	pesos_i(23948) := b"0000000000000000_0000000000000000_0010001011100001_0101100011101111"; -- 0.13625102836591182
	pesos_i(23949) := b"0000000000000000_0000000000000000_0000110001100100_1100011000101110"; -- 0.04841269144862023
	pesos_i(23950) := b"1111111111111111_1111111111111111_1111101111101110_1001010001111100"; -- -0.01589080791030183
	pesos_i(23951) := b"0000000000000000_0000000000000000_0001011111111011_0001110010111101"; -- 0.09367541908229811
	pesos_i(23952) := b"1111111111111111_1111111111111111_1110000110010000_0101110111101111"; -- -0.118890885452834
	pesos_i(23953) := b"0000000000000000_0000000000000000_0001000000110101_0100010010100111"; -- 0.06331280780920844
	pesos_i(23954) := b"0000000000000000_0000000000000000_0000110010111101_0010001010000010"; -- 0.04976096793855339
	pesos_i(23955) := b"1111111111111111_1111111111111111_1110111001111000_0101100101101110"; -- -0.0684761149694806
	pesos_i(23956) := b"0000000000000000_0000000000000000_0001011010101110_1001110101111100"; -- 0.0886019161368662
	pesos_i(23957) := b"1111111111111111_1111111111111111_1110010010100111_1010101110000011"; -- -0.10681655937886342
	pesos_i(23958) := b"1111111111111111_1111111111111111_1110001011100111_0100011101101110"; -- -0.11365846220678126
	pesos_i(23959) := b"0000000000000000_0000000000000000_0000011011010110_0100111010011001"; -- 0.02670756564767775
	pesos_i(23960) := b"0000000000000000_0000000000000000_0001010111011111_0001111001100011"; -- 0.08543577110232473
	pesos_i(23961) := b"1111111111111111_1111111111111111_1110011100010000_0110011011111010"; -- -0.09740597160284983
	pesos_i(23962) := b"0000000000000000_0000000000000000_0000010001000011_1111001101001110"; -- 0.016661840990980677
	pesos_i(23963) := b"0000000000000000_0000000000000000_0000010110010110_1011100100000100"; -- 0.021831096216568445
	pesos_i(23964) := b"0000000000000000_0000000000000000_0001010110100110_1001101111000100"; -- 0.08457349327986287
	pesos_i(23965) := b"1111111111111111_1111111111111111_1101110100110010_0101101101110010"; -- -0.13595036006072628
	pesos_i(23966) := b"1111111111111111_1111111111111111_1110000000000010_1100011111101111"; -- -0.12495756553658167
	pesos_i(23967) := b"0000000000000000_0000000000000000_0000000100101100_1101111110001010"; -- 0.004590960664715752
	pesos_i(23968) := b"1111111111111111_1111111111111111_1111011001000110_0000011001001011"; -- -0.03799400971360525
	pesos_i(23969) := b"1111111111111111_1111111111111111_1101110001001110_1111001011001111"; -- -0.1394203418456478
	pesos_i(23970) := b"1111111111111111_1111111111111111_1110111011110111_1011001010110100"; -- -0.06653292747441834
	pesos_i(23971) := b"0000000000000000_0000000000000000_0001001100000011_0100000111000000"; -- 0.07426844532459494
	pesos_i(23972) := b"0000000000000000_0000000000000000_0010011000010001_1011101001001011"; -- 0.14870800333230014
	pesos_i(23973) := b"0000000000000000_0000000000000000_0001111011001110_0001000110100101"; -- 0.12033186231763959
	pesos_i(23974) := b"0000000000000000_0000000000000000_0000010000111010_0111100110100110"; -- 0.0165172605560511
	pesos_i(23975) := b"0000000000000000_0000000000000000_0000110110111001_0100101111101101"; -- 0.05360865159744435
	pesos_i(23976) := b"1111111111111111_1111111111111111_1111110110110011_0001111100000110"; -- -0.008985577621729413
	pesos_i(23977) := b"0000000000000000_0000000000000000_0001110000100100_0010111000011101"; -- 0.1099270650761245
	pesos_i(23978) := b"0000000000000000_0000000000000000_0001101000001010_0001001000000000"; -- 0.10171616087065381
	pesos_i(23979) := b"1111111111111111_1111111111111111_1110100011000100_1111100100111101"; -- -0.09074442169021484
	pesos_i(23980) := b"0000000000000000_0000000000000000_0001110110000110_0000100000110101"; -- 0.11532641687778619
	pesos_i(23981) := b"0000000000000000_0000000000000000_0000010001101000_1001000000111111"; -- 0.017220511901861968
	pesos_i(23982) := b"1111111111111111_1111111111111111_1110010000101101_0010110000011010"; -- -0.10868572579302008
	pesos_i(23983) := b"0000000000000000_0000000000000000_0000100100011000_1101101101000100"; -- 0.035535530302164664
	pesos_i(23984) := b"1111111111111111_1111111111111111_1111100011110010_1000101100100000"; -- -0.0275490804433543
	pesos_i(23985) := b"0000000000000000_0000000000000000_0001111111000000_1010000010001011"; -- 0.12403300656980136
	pesos_i(23986) := b"0000000000000000_0000000000000000_0001010001111100_1101100011001110"; -- 0.0800300124353784
	pesos_i(23987) := b"0000000000000000_0000000000000000_0001111011000011_1000011000011110"; -- 0.12017095779704338
	pesos_i(23988) := b"1111111111111111_1111111111111111_1110001100011000_0111110111010011"; -- -0.11290753939637634
	pesos_i(23989) := b"1111111111111111_1111111111111111_1110100101111011_0011101011011011"; -- -0.08796341092543226
	pesos_i(23990) := b"1111111111111111_1111111111111111_1110110101010100_1011010100100110"; -- -0.07292621444701725
	pesos_i(23991) := b"0000000000000000_0000000000000000_0000000101101010_1011110100110101"; -- 0.005534959325227636
	pesos_i(23992) := b"1111111111111111_1111111111111111_1111101000010110_0101111100011110"; -- -0.023096137172013923
	pesos_i(23993) := b"1111111111111111_1111111111111111_1111100110100011_0110111101111111"; -- -0.02484992175262548
	pesos_i(23994) := b"1111111111111111_1111111111111111_1110001100011110_1110110101011111"; -- -0.11280933784495985
	pesos_i(23995) := b"0000000000000000_0000000000000000_0001010101011111_1011001000001101"; -- 0.08349144768816842
	pesos_i(23996) := b"1111111111111111_1111111111111111_1110110000100011_0110010001111101"; -- -0.07758495288213506
	pesos_i(23997) := b"0000000000000000_0000000000000000_0000001111011011_1000101001101110"; -- 0.01506867592683963
	pesos_i(23998) := b"1111111111111111_1111111111111111_1110100011100110_0011100010101011"; -- -0.09023710086273473
	pesos_i(23999) := b"0000000000000000_0000000000000000_0001111000001001_0000110001101000"; -- 0.1173255686657665
	pesos_i(24000) := b"0000000000000000_0000000000000000_0000100000100011_0100000101011010"; -- 0.03178795287357623
	pesos_i(24001) := b"1111111111111111_1111111111111111_1101011101111010_0111101100111000"; -- -0.15828733325824607
	pesos_i(24002) := b"1111111111111111_1111111111111111_1111110111111011_1111101000100100"; -- -0.007873884289867862
	pesos_i(24003) := b"0000000000000000_0000000000000000_0010001011000110_0101101101001111"; -- 0.13583918269218342
	pesos_i(24004) := b"0000000000000000_0000000000000000_0000010101000110_1100010100101111"; -- 0.020611118351690137
	pesos_i(24005) := b"0000000000000000_0000000000000000_0010001011101100_1011101111010010"; -- 0.13642476920520627
	pesos_i(24006) := b"1111111111111111_1111111111111111_1111001001100010_1111110001101010"; -- -0.05317709354766295
	pesos_i(24007) := b"1111111111111111_1111111111111111_1110000001100010_1011101000100000"; -- -0.12349354480043424
	pesos_i(24008) := b"1111111111111111_1111111111111111_1110000100101101_1100100010110010"; -- -0.12039514216866262
	pesos_i(24009) := b"1111111111111111_1111111111111111_1111000010000011_1110011111111001"; -- -0.06048727203413936
	pesos_i(24010) := b"0000000000000000_0000000000000000_0010000011010001_1011101001100100"; -- 0.12820019667084495
	pesos_i(24011) := b"0000000000000000_0000000000000000_0001000110001011_1000000010011110"; -- 0.06853488794362436
	pesos_i(24012) := b"1111111111111111_1111111111111111_1110100101101011_0011011100010100"; -- -0.08820777654319223
	pesos_i(24013) := b"0000000000000000_0000000000000000_0001111001011000_1100100100010011"; -- 0.11854225844419068
	pesos_i(24014) := b"1111111111111111_1111111111111111_1110101011010011_0001000010000110"; -- -0.08271691058374114
	pesos_i(24015) := b"0000000000000000_0000000000000000_0001110101001011_0000110011010000"; -- 0.11442642293826148
	pesos_i(24016) := b"0000000000000000_0000000000000000_0001110001101011_1000110010000011"; -- 0.11101606550988798
	pesos_i(24017) := b"1111111111111111_1111111111111111_1110010001001111_1100100010001011"; -- -0.10815760246505025
	pesos_i(24018) := b"1111111111111111_1111111111111111_1110110011001000_1111000000111000"; -- -0.07505892398971688
	pesos_i(24019) := b"0000000000000000_0000000000000000_0010001011110001_0101000100000010"; -- 0.13649469659004076
	pesos_i(24020) := b"0000000000000000_0000000000000000_0001101110111010_1001000111000011"; -- 0.10831557280685959
	pesos_i(24021) := b"0000000000000000_0000000000000000_0001000000011110_1011010010001001"; -- 0.06296852437338248
	pesos_i(24022) := b"1111111111111111_1111111111111111_1111011001111111_0111000111111100"; -- -0.03711783968252327
	pesos_i(24023) := b"0000000000000000_0000000000000000_0001000010011011_0000100011111100"; -- 0.06486564785759757
	pesos_i(24024) := b"0000000000000000_0000000000000000_0010011100011101_0100111010100001"; -- 0.15279094164338478
	pesos_i(24025) := b"0000000000000000_0000000000000000_0000001111110110_1011101010001100"; -- 0.015483531239479894
	pesos_i(24026) := b"1111111111111111_1111111111111111_1111001010001100_1110010101100110"; -- -0.052537596304999476
	pesos_i(24027) := b"1111111111111111_1111111111111111_1110011100100010_0100111010100000"; -- -0.09713276471643946
	pesos_i(24028) := b"1111111111111111_1111111111111111_1111011110001010_0010111111101001"; -- -0.033047681497701216
	pesos_i(24029) := b"0000000000000000_0000000000000000_0000000100001011_0011000000100001"; -- 0.004076965401938182
	pesos_i(24030) := b"0000000000000000_0000000000000000_0001010000011100_0110010100010000"; -- 0.07855826985769422
	pesos_i(24031) := b"0000000000000000_0000000000000000_0010011100001101_1101101110101011"; -- 0.1525552075926762
	pesos_i(24032) := b"1111111111111111_1111111111111111_1111000010001100_0100100011110000"; -- -0.06035942221720024
	pesos_i(24033) := b"0000000000000000_0000000000000000_0000100100101011_0100111111100010"; -- 0.03581713935542312
	pesos_i(24034) := b"1111111111111111_1111111111111111_1111000001101110_0010000010100100"; -- -0.06081958757987303
	pesos_i(24035) := b"1111111111111111_1111111111111111_1111101100011110_1001001100101010"; -- -0.019064714669899396
	pesos_i(24036) := b"1111111111111111_1111111111111111_1111001001000110_0001110010100111"; -- -0.053617676975999194
	pesos_i(24037) := b"0000000000000000_0000000000000000_0001000001010101_1111100110101100"; -- 0.06381187878682995
	pesos_i(24038) := b"1111111111111111_1111111111111111_1110000111001011_0101010111101111"; -- -0.11799109375667408
	pesos_i(24039) := b"1111111111111111_1111111111111111_1110011001110100_0111101000010110"; -- -0.09978520367468534
	pesos_i(24040) := b"1111111111111111_1111111111111111_1101110110000000_0010010010001011"; -- -0.13476344690382758
	pesos_i(24041) := b"1111111111111111_1111111111111111_1111011000010001_1010011010010111"; -- -0.03879317110811957
	pesos_i(24042) := b"1111111111111111_1111111111111111_1101110010000001_1011001011000100"; -- -0.13864596102264615
	pesos_i(24043) := b"0000000000000000_0000000000000000_0001000101101001_1101100101100111"; -- 0.06802138104197343
	pesos_i(24044) := b"1111111111111111_1111111111111111_1101110010010111_1001010110011110"; -- -0.13831200504576582
	pesos_i(24045) := b"1111111111111111_1111111111111111_1110110111111100_1011100000101011"; -- -0.0703625578852738
	pesos_i(24046) := b"0000000000000000_0000000000000000_0010000101100110_1011110011011110"; -- 0.13047390376596119
	pesos_i(24047) := b"1111111111111111_1111111111111111_1111010110101100_1000001001010001"; -- -0.04033647084620282
	pesos_i(24048) := b"0000000000000000_0000000000000000_0000010111111110_1000100101101100"; -- 0.02341517330877848
	pesos_i(24049) := b"0000000000000000_0000000000000000_0001101000110110_1010110000010001"; -- 0.10239673065360179
	pesos_i(24050) := b"1111111111111111_1111111111111111_1111011010111000_0011110110000101"; -- -0.03625121606770473
	pesos_i(24051) := b"1111111111111111_1111111111111111_1111100010000010_1110110101000001"; -- -0.029252216079715423
	pesos_i(24052) := b"1111111111111111_1111111111111111_1101011010101000_1000110101000001"; -- -0.16149060410110896
	pesos_i(24053) := b"0000000000000000_0000000000000000_0010011100100101_1111110011111000"; -- 0.1529234034105872
	pesos_i(24054) := b"1111111111111111_1111111111111111_1110101010000011_1001101101001110"; -- -0.08392934179394222
	pesos_i(24055) := b"1111111111111111_1111111111111111_1111111011101101_1101110011011110"; -- -0.00418300235488173
	pesos_i(24056) := b"0000000000000000_0000000000000000_0001011001110000_0010111011010011"; -- 0.08764927535631244
	pesos_i(24057) := b"1111111111111111_1111111111111111_1110000101101011_0010110110110110"; -- -0.11945833506217206
	pesos_i(24058) := b"1111111111111111_1111111111111111_1110011010001101_0011011111001000"; -- -0.09940768594156517
	pesos_i(24059) := b"0000000000000000_0000000000000000_0001011100011000_1100011101101011"; -- 0.09022184713735056
	pesos_i(24060) := b"1111111111111111_1111111111111111_1111001110000000_1101110010001100"; -- -0.048814979311780256
	pesos_i(24061) := b"1111111111111111_1111111111111111_1111111110011010_0101001110011101"; -- -0.0015514127612291006
	pesos_i(24062) := b"0000000000000000_0000000000000000_0000101100001000_0010010110110111"; -- 0.04309306825650723
	pesos_i(24063) := b"0000000000000000_0000000000000000_0000111000000000_0110111001100001"; -- 0.05469407911697223
	pesos_i(24064) := b"0000000000000000_0000000000000000_0000000101000101_1111100010111001"; -- 0.004973931454604308
	pesos_i(24065) := b"0000000000000000_0000000000000000_0001100100111100_0111110011110111"; -- 0.0985792258043283
	pesos_i(24066) := b"0000000000000000_0000000000000000_0000111011100101_1001010101101110"; -- 0.05819066932469185
	pesos_i(24067) := b"0000000000000000_0000000000000000_0000111100111100_0001011110010110"; -- 0.05951068324518466
	pesos_i(24068) := b"1111111111111111_1111111111111111_1111010000001111_1100000011011111"; -- -0.04663462225322207
	pesos_i(24069) := b"1111111111111111_1111111111111111_1111111101101110_1110110101000100"; -- -0.002213641165496446
	pesos_i(24070) := b"1111111111111111_1111111111111111_1101101000110001_0010000101011100"; -- -0.1476878308660532
	pesos_i(24071) := b"1111111111111111_1111111111111111_1111100010110100_0100111000110100"; -- -0.028498756800818776
	pesos_i(24072) := b"0000000000000000_0000000000000000_0000111000000110_0001000000100011"; -- 0.05478001444862716
	pesos_i(24073) := b"0000000000000000_0000000000000000_0001000100110001_1110001011001001"; -- 0.06716744807770376
	pesos_i(24074) := b"1111111111111111_1111111111111111_1111110010101100_1011100111101111"; -- -0.012989405886085383
	pesos_i(24075) := b"1111111111111111_1111111111111111_1111010100011010_1110001110010011"; -- -0.04255845707779777
	pesos_i(24076) := b"1111111111111111_1111111111111111_1101101001001100_1001101111001100"; -- -0.14726854577296516
	pesos_i(24077) := b"1111111111111111_1111111111111111_1111100101111110_1110000010101000"; -- -0.025407752005880364
	pesos_i(24078) := b"0000000000000000_0000000000000000_0001011101100111_1111111100010110"; -- 0.09143060948321688
	pesos_i(24079) := b"0000000000000000_0000000000000000_0010000011111000_1000001011010011"; -- 0.1287919773041377
	pesos_i(24080) := b"1111111111111111_1111111111111111_1111001110101100_1111111000001101"; -- -0.04814159570711133
	pesos_i(24081) := b"1111111111111111_1111111111111111_1111100001001011_1111100101100000"; -- -0.03009072696040028
	pesos_i(24082) := b"0000000000000000_0000000000000000_0001010101000101_1110110111011101"; -- 0.0830982841745231
	pesos_i(24083) := b"0000000000000000_0000000000000000_0001000000101000_0101011100101110"; -- 0.06311554781063608
	pesos_i(24084) := b"0000000000000000_0000000000000000_0000110011001000_1100101010100011"; -- 0.04993883583774576
	pesos_i(24085) := b"1111111111111111_1111111111111111_1111111100010000_1011010110011110"; -- -0.0036512840515364447
	pesos_i(24086) := b"0000000000000000_0000000000000000_0001100110010100_1100010001011011"; -- 0.09992625457378859
	pesos_i(24087) := b"1111111111111111_1111111111111111_1110001111000010_0011010101000101"; -- -0.11031786972966771
	pesos_i(24088) := b"1111111111111111_1111111111111111_1110111001100110_0010000010000010"; -- -0.06875416584675237
	pesos_i(24089) := b"0000000000000000_0000000000000000_0000110100000011_1100011100000110"; -- 0.050838889204517755
	pesos_i(24090) := b"1111111111111111_1111111111111111_1110010001000011_0111000110001111"; -- -0.1083458924755298
	pesos_i(24091) := b"0000000000000000_0000000000000000_0000110111110100_0000011100010101"; -- 0.054504816747931194
	pesos_i(24092) := b"1111111111111111_1111111111111111_1101100000110010_0100110001011001"; -- -0.1554825097764574
	pesos_i(24093) := b"0000000000000000_0000000000000000_0000000100001011_0001011011010110"; -- 0.004075457768529181
	pesos_i(24094) := b"0000000000000000_0000000000000000_0001100110100011_0111100100110110"; -- 0.10015065746012819
	pesos_i(24095) := b"1111111111111111_1111111111111111_1101110110010000_0111000011101001"; -- -0.13451475452010853
	pesos_i(24096) := b"0000000000000000_0000000000000000_0000011100111010_1001010110000001"; -- 0.028237670784403215
	pesos_i(24097) := b"0000000000000000_0000000000000000_0001101111011110_1110000000110001"; -- 0.10886956409458737
	pesos_i(24098) := b"0000000000000000_0000000000000000_0001100000100100_1000101101010001"; -- 0.09430762040279478
	pesos_i(24099) := b"1111111111111111_1111111111111111_1110101011011000_0101100101100101"; -- -0.08263627329842549
	pesos_i(24100) := b"1111111111111111_1111111111111111_1111111100101011_1001011100001101"; -- -0.003241118654855204
	pesos_i(24101) := b"1111111111111111_1111111111111111_1111101000001111_1010100111001000"; -- -0.023198498478460214
	pesos_i(24102) := b"0000000000000000_0000000000000000_0000111010010001_0010100000000010"; -- 0.056902409040551064
	pesos_i(24103) := b"1111111111111111_1111111111111111_1110000111100010_0111001101100011"; -- -0.11763838618593357
	pesos_i(24104) := b"0000000000000000_0000000000000000_0000111101101110_0100010011011100"; -- 0.06027632113371841
	pesos_i(24105) := b"1111111111111111_1111111111111111_1111101010000001_1010010110100010"; -- -0.021459243644563523
	pesos_i(24106) := b"0000000000000000_0000000000000000_0001100110111100_0001010110011110"; -- 0.10052619087912977
	pesos_i(24107) := b"0000000000000000_0000000000000000_0000011110011100_0010100110101011"; -- 0.029726604608682986
	pesos_i(24108) := b"0000000000000000_0000000000000000_0000010110010111_0101110000101010"; -- 0.021840820608712667
	pesos_i(24109) := b"1111111111111111_1111111111111111_1110101000010111_0001001001100000"; -- -0.08558545265252197
	pesos_i(24110) := b"0000000000000000_0000000000000000_0000011010111111_1010011010011010"; -- 0.026361858929889445
	pesos_i(24111) := b"1111111111111111_1111111111111111_1110100000110100_1100110001010101"; -- -0.09294436392043284
	pesos_i(24112) := b"1111111111111111_1111111111111111_1111011011111110_1110110010000101"; -- -0.03517266997239702
	pesos_i(24113) := b"1111111111111111_1111111111111111_1111000001100110_1100100001111011"; -- -0.06093165386193952
	pesos_i(24114) := b"0000000000000000_0000000000000000_0001111000001011_1110101001100000"; -- 0.1173693164193919
	pesos_i(24115) := b"1111111111111111_1111111111111111_1110101000001010_1011010111101000"; -- -0.08577406967739512
	pesos_i(24116) := b"0000000000000000_0000000000000000_0000100100111010_0101110111110110"; -- 0.036046860291177325
	pesos_i(24117) := b"0000000000000000_0000000000000000_0001011001000010_0010001101101000"; -- 0.08694669045458558
	pesos_i(24118) := b"1111111111111111_1111111111111111_1111100011010100_0110101111101110"; -- -0.028008703560965385
	pesos_i(24119) := b"0000000000000000_0000000000000000_0001000011011110_0111010001011001"; -- 0.0658943860911918
	pesos_i(24120) := b"0000000000000000_0000000000000000_0000100111001110_1100101101011111"; -- 0.038311682348539634
	pesos_i(24121) := b"1111111111111111_1111111111111111_1111101111111111_1110101010111100"; -- -0.01562626753701338
	pesos_i(24122) := b"1111111111111111_1111111111111111_1111111111000001_1101100000011111"; -- -0.0009484218096657942
	pesos_i(24123) := b"0000000000000000_0000000000000000_0001100111011011_1011010000111100"; -- 0.10100866750952832
	pesos_i(24124) := b"0000000000000000_0000000000000000_0000110110010011_1111010000000101"; -- 0.053038836583362094
	pesos_i(24125) := b"1111111111111111_1111111111111111_1110101000100010_1111011011010011"; -- -0.0854039892011051
	pesos_i(24126) := b"1111111111111111_1111111111111111_1110111000010001_0110001011100110"; -- -0.07004720584142683
	pesos_i(24127) := b"1111111111111111_1111111111111111_1101101100011001_1111101011111001"; -- -0.1441348210389896
	pesos_i(24128) := b"1111111111111111_1111111111111111_1111001011100111_0101101001110011"; -- -0.05115732855937181
	pesos_i(24129) := b"0000000000000000_0000000000000000_0000011000110011_1000000110101111"; -- 0.024223428054566412
	pesos_i(24130) := b"0000000000000000_0000000000000000_0000011011101011_0011100010001011"; -- 0.02702668554624742
	pesos_i(24131) := b"1111111111111111_1111111111111111_1110000000011111_1111111010001100"; -- -0.12451180541694248
	pesos_i(24132) := b"0000000000000000_0000000000000000_0001110111100110_1110011111011100"; -- 0.11680459140097887
	pesos_i(24133) := b"1111111111111111_1111111111111111_1110100011101011_1000110001110011"; -- -0.09015581308866691
	pesos_i(24134) := b"0000000000000000_0000000000000000_0001110100010000_1000111000111001"; -- 0.11353386776730309
	pesos_i(24135) := b"1111111111111111_1111111111111111_1110110001101100_1111000111111100"; -- -0.0764626274138561
	pesos_i(24136) := b"1111111111111111_1111111111111111_1111010000011101_0001000001000110"; -- -0.046431525091471956
	pesos_i(24137) := b"0000000000000000_0000000000000000_0001011011111110_1100000011011100"; -- 0.08982472770938259
	pesos_i(24138) := b"1111111111111111_1111111111111111_1111100010000001_1110111110110010"; -- -0.029267329333205413
	pesos_i(24139) := b"0000000000000000_0000000000000000_0000101001001101_0011010011100100"; -- 0.040240579390189456
	pesos_i(24140) := b"1111111111111111_1111111111111111_1101111011001001_1000010010011101"; -- -0.12973757908136263
	pesos_i(24141) := b"1111111111111111_1111111111111111_1110100111011111_1000110100001100"; -- -0.08643263303191724
	pesos_i(24142) := b"1111111111111111_1111111111111111_1111111111000101_0001000000011010"; -- -0.0008993088976503996
	pesos_i(24143) := b"1111111111111111_1111111111111111_1101111010100000_1110101101001011"; -- -0.13035706914094491
	pesos_i(24144) := b"0000000000000000_0000000000000000_0000100111101110_1011001101100011"; -- 0.038798534075637756
	pesos_i(24145) := b"1111111111111111_1111111111111111_1111111100010001_0101101010011000"; -- -0.0036414508239669277
	pesos_i(24146) := b"1111111111111111_1111111111111111_1111011101100011_0011101000111100"; -- -0.03364215890930612
	pesos_i(24147) := b"0000000000000000_0000000000000000_0001011110011001_0111100001110110"; -- 0.09218552471039491
	pesos_i(24148) := b"1111111111111111_1111111111111111_1110001101010000_1100001000001101"; -- -0.11204898062687213
	pesos_i(24149) := b"1111111111111111_1111111111111111_1110011001111101_1100100011000011"; -- -0.0996431850424691
	pesos_i(24150) := b"0000000000000000_0000000000000000_0000001100110011_1101111010010100"; -- 0.012510214896155043
	pesos_i(24151) := b"1111111111111111_1111111111111111_1101110111000001_0100101010110100"; -- -0.13376935105437252
	pesos_i(24152) := b"0000000000000000_0000000000000000_0000110110100100_1101001001010100"; -- 0.05329622798940907
	pesos_i(24153) := b"0000000000000000_0000000000000000_0000010101011011_1001101100010001"; -- 0.020929042481530397
	pesos_i(24154) := b"1111111111111111_1111111111111111_1110100001000111_1000100011001010"; -- -0.09265847266759024
	pesos_i(24155) := b"0000000000000000_0000000000000000_0000011100100101_0011101011100100"; -- 0.027911835430072585
	pesos_i(24156) := b"0000000000000000_0000000000000000_0001111010100100_0001001100111111"; -- 0.11969108851965027
	pesos_i(24157) := b"0000000000000000_0000000000000000_0000010100111011_0111100000101001"; -- 0.02043868071893761
	pesos_i(24158) := b"0000000000000000_0000000000000000_0000011110001011_0100011000001001"; -- 0.02946889600883555
	pesos_i(24159) := b"1111111111111111_1111111111111111_1110111011000111_1000101001100110"; -- -0.06726775178222891
	pesos_i(24160) := b"0000000000000000_0000000000000000_0000110110110011_1010100011100100"; -- 0.05352264001617931
	pesos_i(24161) := b"0000000000000000_0000000000000000_0001101101101111_0101111010000011"; -- 0.10716810893743636
	pesos_i(24162) := b"1111111111111111_1111111111111111_1110011101001010_0111010011110001"; -- -0.09652012940971207
	pesos_i(24163) := b"0000000000000000_0000000000000000_0000100100011110_1110100101111011"; -- 0.03562793017450008
	pesos_i(24164) := b"1111111111111111_1111111111111111_1110100101000111_1111100101111111"; -- -0.088745504747113
	pesos_i(24165) := b"1111111111111111_1111111111111111_1111111010000000_0001100000110111"; -- -0.005857931653229576
	pesos_i(24166) := b"1111111111111111_1111111111111111_1101111100010010_0110011001100000"; -- -0.1286254897848217
	pesos_i(24167) := b"0000000000000000_0000000000000000_0001001100110001_1000110000100110"; -- 0.07497478410568133
	pesos_i(24168) := b"1111111111111111_1111111111111111_1110000001001000_0100010110110110"; -- -0.12389721220608137
	pesos_i(24169) := b"0000000000000000_0000000000000000_0001000100011110_0110000001111100"; -- 0.06686976465683589
	pesos_i(24170) := b"0000000000000000_0000000000000000_0001111000101011_0001000111110000"; -- 0.11784469712991626
	pesos_i(24171) := b"1111111111111111_1111111111111111_1101111111110011_0100100010100011"; -- -0.1251940347984338
	pesos_i(24172) := b"0000000000000000_0000000000000000_0000010100001111_1000101111110001"; -- 0.019768473055667837
	pesos_i(24173) := b"1111111111111111_1111111111111111_1110111110111101_0000010111000101"; -- -0.0635219949024008
	pesos_i(24174) := b"0000000000000000_0000000000000000_0000000001111110_0001100011100000"; -- 0.0019240900974023386
	pesos_i(24175) := b"0000000000000000_0000000000000000_0001000100111101_1101101011001110"; -- 0.06735007791898012
	pesos_i(24176) := b"1111111111111111_1111111111111111_1101110110011000_0100110010001011"; -- -0.1343948516327225
	pesos_i(24177) := b"1111111111111111_1111111111111111_1110011100000001_0010011011100000"; -- -0.0976386741553048
	pesos_i(24178) := b"1111111111111111_1111111111111111_1111011110011000_0111010111110011"; -- -0.032829883723118854
	pesos_i(24179) := b"1111111111111111_1111111111111111_1111011100011010_1000010100100101"; -- -0.03475158544982884
	pesos_i(24180) := b"1111111111111111_1111111111111111_1110000111011111_1010010101011101"; -- -0.11768118366032213
	pesos_i(24181) := b"1111111111111111_1111111111111111_1111001110011000_0010101011000011"; -- -0.04845936535474596
	pesos_i(24182) := b"0000000000000000_0000000000000000_0001100100010001_1001011111000011"; -- 0.09792469511193592
	pesos_i(24183) := b"0000000000000000_0000000000000000_0001001000111000_1100001010011000"; -- 0.07117859078221883
	pesos_i(24184) := b"0000000000000000_0000000000000000_0000110011000111_0110111000011001"; -- 0.04991806137368623
	pesos_i(24185) := b"0000000000000000_0000000000000000_0000001100010010_1011110111000111"; -- 0.012004719786729854
	pesos_i(24186) := b"0000000000000000_0000000000000000_0010000010101001_1100011101001111"; -- 0.1275906151122136
	pesos_i(24187) := b"0000000000000000_0000000000000000_0001110100011111_0101101011010100"; -- 0.11375968625677119
	pesos_i(24188) := b"0000000000000000_0000000000000000_0000010110100100_0111111011001101"; -- 0.02204124921468109
	pesos_i(24189) := b"1111111111111111_1111111111111111_1111010001100011_0011001100011001"; -- -0.045361334298463785
	pesos_i(24190) := b"0000000000000000_0000000000000000_0010010111010100_1010000100010100"; -- 0.14777571423304592
	pesos_i(24191) := b"0000000000000000_0000000000000000_0000100001010100_0110100111101010"; -- 0.032538051263326866
	pesos_i(24192) := b"0000000000000000_0000000000000000_0000101110011111_1011000011100011"; -- 0.045405440771991615
	pesos_i(24193) := b"1111111111111111_1111111111111111_1110001011010100_1110001001000101"; -- -0.113939150006195
	pesos_i(24194) := b"0000000000000000_0000000000000000_0010010101110001_0111011111010110"; -- 0.14626263585846155
	pesos_i(24195) := b"1111111111111111_1111111111111111_1111010000011100_0111110111010111"; -- -0.04644025334759021
	pesos_i(24196) := b"1111111111111111_1111111111111111_1110100000111100_0000000011000101"; -- -0.09283442675516757
	pesos_i(24197) := b"0000000000000000_0000000000000000_0000110111010011_1010011001001001"; -- 0.05401076577310942
	pesos_i(24198) := b"0000000000000000_0000000000000000_0001111000011100_0001001110110100"; -- 0.11761592050508707
	pesos_i(24199) := b"1111111111111111_1111111111111111_1101111011101110_0011001100110000"; -- -0.1291778571754605
	pesos_i(24200) := b"1111111111111111_1111111111111111_1101100110001110_1110001010001100"; -- -0.15016349875679302
	pesos_i(24201) := b"1111111111111111_1111111111111111_1111000000001000_1000110101111111"; -- -0.06236949588830389
	pesos_i(24202) := b"1111111111111111_1111111111111111_1110111111110000_1110011001000111"; -- -0.062730415088305
	pesos_i(24203) := b"0000000000000000_0000000000000000_0001110011001100_1010111001111101"; -- 0.1124981932169311
	pesos_i(24204) := b"0000000000000000_0000000000000000_0000110110011010_0011100101011000"; -- 0.053134521509450944
	pesos_i(24205) := b"0000000000000000_0000000000000000_0010000001110001_1010101001110101"; -- 0.1267344032242436
	pesos_i(24206) := b"0000000000000000_0000000000000000_0000011001100110_1000100010010011"; -- 0.025002036840277346
	pesos_i(24207) := b"1111111111111111_1111111111111111_1110100011110101_0111101011010010"; -- -0.09000427612626612
	pesos_i(24208) := b"1111111111111111_1111111111111111_1111001111101111_1101100000111011"; -- -0.047121511073010935
	pesos_i(24209) := b"0000000000000000_0000000000000000_0001111000000101_1000110001111100"; -- 0.1172721675770559
	pesos_i(24210) := b"1111111111111111_1111111111111111_1110111111010011_0001010011101010"; -- -0.06318539888878047
	pesos_i(24211) := b"0000000000000000_0000000000000000_0001100000100100_1010101010000100"; -- 0.09430947995874979
	pesos_i(24212) := b"1111111111111111_1111111111111111_1101111110100001_1001110111101001"; -- -0.1264401727966381
	pesos_i(24213) := b"0000000000000000_0000000000000000_0000111000010100_0110001000111100"; -- 0.05499853100890757
	pesos_i(24214) := b"0000000000000000_0000000000000000_0000110011111111_1000000110011011"; -- 0.05077371620525835
	pesos_i(24215) := b"0000000000000000_0000000000000000_0001101010001001_1100000100010011"; -- 0.10366446221107745
	pesos_i(24216) := b"0000000000000000_0000000000000000_0001001100100011_1100010110001101"; -- 0.07476458261854746
	pesos_i(24217) := b"1111111111111111_1111111111111111_1110110001110111_0100110111001000"; -- -0.07630456787586175
	pesos_i(24218) := b"0000000000000000_0000000000000000_0000111111110010_1100001101010001"; -- 0.062298018807618746
	pesos_i(24219) := b"0000000000000000_0000000000000000_0010001001010101_1110011110011010"; -- 0.13412330168457343
	pesos_i(24220) := b"0000000000000000_0000000000000000_0001100110001001_0000100111000000"; -- 0.09974728527132849
	pesos_i(24221) := b"0000000000000000_0000000000000000_0000100010000001_0000101001100110"; -- 0.03321900366424064
	pesos_i(24222) := b"1111111111111111_1111111111111111_1110000111010011_0110101000110011"; -- -0.11786781559871101
	pesos_i(24223) := b"0000000000000000_0000000000000000_0001001110101000_1011110001010010"; -- 0.07679345133774738
	pesos_i(24224) := b"0000000000000000_0000000000000000_0010001011000011_1110100100111011"; -- 0.13580186546933307
	pesos_i(24225) := b"1111111111111111_1111111111111111_1111001110111101_0001100001010111"; -- -0.04789588811162128
	pesos_i(24226) := b"1111111111111111_1111111111111111_1111000011110111_0011111011000000"; -- -0.058727338869754786
	pesos_i(24227) := b"0000000000000000_0000000000000000_0000001010100011_0000011111011111"; -- 0.010300151823166927
	pesos_i(24228) := b"0000000000000000_0000000000000000_0001000000001110_0011111001001010"; -- 0.0627173358268162
	pesos_i(24229) := b"0000000000000000_0000000000000000_0001011100101000_0100101100111001"; -- 0.09045858516814942
	pesos_i(24230) := b"0000000000000000_0000000000000000_0000001110111001_0010001110100111"; -- 0.014543750982652339
	pesos_i(24231) := b"1111111111111111_1111111111111111_1101101011010110_0000100000101101"; -- -0.14517163182850792
	pesos_i(24232) := b"1111111111111111_1111111111111111_1111010010110100_1111100110000000"; -- -0.044113546628302205
	pesos_i(24233) := b"0000000000000000_0000000000000000_0000111101101111_0000111111010011"; -- 0.06028841888312552
	pesos_i(24234) := b"0000000000000000_0000000000000000_0001011010110011_1000010101000011"; -- 0.08867676623348385
	pesos_i(24235) := b"0000000000000000_0000000000000000_0001010001001000_1110000001010101"; -- 0.07923700415739784
	pesos_i(24236) := b"1111111111111111_1111111111111111_1110110001000110_1100010001110001"; -- -0.07704517601475627
	pesos_i(24237) := b"1111111111111111_1111111111111111_1110110111110101_1101111101100010"; -- -0.07046703204239453
	pesos_i(24238) := b"0000000000000000_0000000000000000_0000000101110110_0010101011010110"; -- 0.005709340233411561
	pesos_i(24239) := b"1111111111111111_1111111111111111_1110111101100001_1101000110000010"; -- -0.0649136597139232
	pesos_i(24240) := b"1111111111111111_1111111111111111_1110110010101101_1000110011010010"; -- -0.07547683604505895
	pesos_i(24241) := b"0000000000000000_0000000000000000_0001001000011000_1100101110110000"; -- 0.07069085161839504
	pesos_i(24242) := b"0000000000000000_0000000000000000_0010010011001001_1010001111110100"; -- 0.14370178904268166
	pesos_i(24243) := b"1111111111111111_1111111111111111_1110110111100001_1000110000011010"; -- -0.07077717167772303
	pesos_i(24244) := b"0000000000000000_0000000000000000_0000001010101110_0110101001100011"; -- 0.010473870529590002
	pesos_i(24245) := b"1111111111111111_1111111111111111_1110110111001100_1111001001100111"; -- -0.07109150868285637
	pesos_i(24246) := b"1111111111111111_1111111111111111_1111111111011000_0101010001101101"; -- -0.0006053194274183717
	pesos_i(24247) := b"1111111111111111_1111111111111111_1101110011110110_0101110111000010"; -- -0.13686574959633002
	pesos_i(24248) := b"1111111111111111_1111111111111111_1101101110100100_1010110010011000"; -- -0.14201852121300487
	pesos_i(24249) := b"1111111111111111_1111111111111111_1101110010101010_1010111001010011"; -- -0.13802061540995503
	pesos_i(24250) := b"0000000000000000_0000000000000000_0000100100011110_0101110011011000"; -- 0.03561954763960594
	pesos_i(24251) := b"0000000000000000_0000000000000000_0001011111011100_0100110001000010"; -- 0.09320522896862637
	pesos_i(24252) := b"1111111111111111_1111111111111111_1110001100111101_0011100111010110"; -- -0.11234701660856584
	pesos_i(24253) := b"0000000000000000_0000000000000000_0010010010010000_0001000001111100"; -- 0.142823248237008
	pesos_i(24254) := b"1111111111111111_1111111111111111_1110010110111010_0100000001101000"; -- -0.10262677629922745
	pesos_i(24255) := b"1111111111111111_1111111111111111_1110010100011101_1010011111001000"; -- -0.10501624459711369
	pesos_i(24256) := b"1111111111111111_1111111111111111_1110001111010000_1110110010101110"; -- -0.1100933147145003
	pesos_i(24257) := b"0000000000000000_0000000000000000_0000100100101011_1011011011101011"; -- 0.03582328059267119
	pesos_i(24258) := b"1111111111111111_1111111111111111_1111000110011101_0111001100111010"; -- -0.05619125216019678
	pesos_i(24259) := b"0000000000000000_0000000000000000_0000001011111010_1100000110100011"; -- 0.011638738911839547
	pesos_i(24260) := b"1111111111111111_1111111111111111_1111000011110010_0101000100100100"; -- -0.05880253674437482
	pesos_i(24261) := b"0000000000000000_0000000000000000_0001110011111111_0011100101010111"; -- 0.11326940904017559
	pesos_i(24262) := b"1111111111111111_1111111111111111_1111101001100111_0000101111010111"; -- -0.021865139097142768
	pesos_i(24263) := b"1111111111111111_1111111111111111_1110011011001111_0110010010000100"; -- -0.09839793942193079
	pesos_i(24264) := b"1111111111111111_1111111111111111_1101111000001000_1111010001100010"; -- -0.13267586342491883
	pesos_i(24265) := b"0000000000000000_0000000000000000_0010000010001010_1001111101110100"; -- 0.12711521712408327
	pesos_i(24266) := b"1111111111111111_1111111111111111_1110111110011011_1101010110111100"; -- -0.06402839812014592
	pesos_i(24267) := b"1111111111111111_1111111111111111_1110010001010100_0110110000001000"; -- -0.10808682259984885
	pesos_i(24268) := b"0000000000000000_0000000000000000_0000010010000110_0101001000000100"; -- 0.017674566200858614
	pesos_i(24269) := b"1111111111111111_1111111111111111_1111000001010001_1101001001111000"; -- -0.06125149307150034
	pesos_i(24270) := b"0000000000000000_0000000000000000_0000101010100001_0000010011101010"; -- 0.04151945784539477
	pesos_i(24271) := b"1111111111111111_1111111111111111_1110000110000100_0101100010100110"; -- -0.11907430587757306
	pesos_i(24272) := b"1111111111111111_1111111111111111_1110100011011101_0001101101001010"; -- -0.09037618097927885
	pesos_i(24273) := b"0000000000000000_0000000000000000_0010010000000011_1101001111000110"; -- 0.14068339895253917
	pesos_i(24274) := b"1111111111111111_1111111111111111_1111000011000101_0011100011001110"; -- -0.0594906326503969
	pesos_i(24275) := b"0000000000000000_0000000000000000_0001111000101100_1011001101110100"; -- 0.11786958307433335
	pesos_i(24276) := b"0000000000000000_0000000000000000_0000000001011101_1101010111001001"; -- 0.0014318099558568826
	pesos_i(24277) := b"0000000000000000_0000000000000000_0000101101100000_1000100100010110"; -- 0.04444176481937407
	pesos_i(24278) := b"1111111111111111_1111111111111111_1110110011111111_0010001010111000"; -- -0.0742319393799607
	pesos_i(24279) := b"0000000000000000_0000000000000000_0001111110000010_1100101010011101"; -- 0.12308946926519519
	pesos_i(24280) := b"0000000000000000_0000000000000000_0010000001000110_0001010010111111"; -- 0.12606935189064708
	pesos_i(24281) := b"0000000000000000_0000000000000000_0001001000100110_0110010101001100"; -- 0.07089837167182854
	pesos_i(24282) := b"0000000000000000_0000000000000000_0000111000010110_1111001110111000"; -- 0.05503772016256484
	pesos_i(24283) := b"0000000000000000_0000000000000000_0010010110110010_1100111101110001"; -- 0.14725967903724277
	pesos_i(24284) := b"0000000000000000_0000000000000000_0000110111101110_1010111111101010"; -- 0.05442332697827044
	pesos_i(24285) := b"1111111111111111_1111111111111111_1101111111010111_0101010001100111"; -- -0.12562057956175943
	pesos_i(24286) := b"0000000000000000_0000000000000000_0000101001010010_0100000110000111"; -- 0.040317626463072714
	pesos_i(24287) := b"0000000000000000_0000000000000000_0000110010000000_1011010010010010"; -- 0.04883888779567387
	pesos_i(24288) := b"0000000000000000_0000000000000000_0000000010101001_1011000010101111"; -- 0.002589266542243265
	pesos_i(24289) := b"0000000000000000_0000000000000000_0010000001010110_0010001001110001"; -- 0.12631430870849014
	pesos_i(24290) := b"1111111111111111_1111111111111111_1111010101011101_1001010010100110"; -- -0.04154082247690584
	pesos_i(24291) := b"0000000000000000_0000000000000000_0000010111011100_1010001100101000"; -- 0.02289790849033322
	pesos_i(24292) := b"1111111111111111_1111111111111111_1110000111010101_0000010010011001"; -- -0.11784335395639255
	pesos_i(24293) := b"0000000000000000_0000000000000000_0001001000111111_0100000000101101"; -- 0.07127762887766029
	pesos_i(24294) := b"0000000000000000_0000000000000000_0000001000000100_0111101011011001"; -- 0.007880857495761756
	pesos_i(24295) := b"1111111111111111_1111111111111111_1111110101001011_0111101000101110"; -- -0.010567058252668689
	pesos_i(24296) := b"0000000000000000_0000000000000000_0001101101101111_0100011100011010"; -- 0.1071667134747145
	pesos_i(24297) := b"0000000000000000_0000000000000000_0010000011000010_0001100101000011"; -- 0.12796171082357388
	pesos_i(24298) := b"1111111111111111_1111111111111111_1111111000110101_0101011011111110"; -- -0.006998598936898316
	pesos_i(24299) := b"1111111111111111_1111111111111111_1110110010001100_0110010001000000"; -- -0.07598279407490167
	pesos_i(24300) := b"0000000000000000_0000000000000000_0001000010110100_0111010000000010"; -- 0.06525349660657072
	pesos_i(24301) := b"0000000000000000_0000000000000000_0010000111100111_1001001100110010"; -- 0.13243980379552303
	pesos_i(24302) := b"1111111111111111_1111111111111111_1111000110010011_0110110111101110"; -- -0.056344155643894896
	pesos_i(24303) := b"1111111111111111_1111111111111111_1111001111110100_0101011110000000"; -- -0.047052890158099804
	pesos_i(24304) := b"0000000000000000_0000000000000000_0001110101001110_0011111011101111"; -- 0.11447518675815944
	pesos_i(24305) := b"0000000000000000_0000000000000000_0001000001110100_0010011000111111"; -- 0.06427229909507388
	pesos_i(24306) := b"0000000000000000_0000000000000000_0010100000010111_0011100000111101"; -- 0.15660430411120535
	pesos_i(24307) := b"0000000000000000_0000000000000000_0001111110000101_1001010010111010"; -- 0.12313203375733531
	pesos_i(24308) := b"1111111111111111_1111111111111111_1111100010111101_0101011110001000"; -- -0.028360871608473556
	pesos_i(24309) := b"1111111111111111_1111111111111111_1111100010110110_0101110111011110"; -- -0.02846730546649259
	pesos_i(24310) := b"0000000000000000_0000000000000000_0001010010110101_0110001101111011"; -- 0.08089277026391267
	pesos_i(24311) := b"0000000000000000_0000000000000000_0000011001010110_1010111010101000"; -- 0.024760166085749533
	pesos_i(24312) := b"1111111111111111_1111111111111111_1110101011010000_1011100100111100"; -- -0.08275263099682542
	pesos_i(24313) := b"0000000000000000_0000000000000000_0000000111001010_0011010111001101"; -- 0.006991732079334703
	pesos_i(24314) := b"1111111111111111_1111111111111111_1110100101000111_1010001100010000"; -- -0.08875065673776919
	pesos_i(24315) := b"0000000000000000_0000000000000000_0001010010110101_1010111000100001"; -- 0.08089721969632316
	pesos_i(24316) := b"0000000000000000_0000000000000000_0001000001100100_1011100010111011"; -- 0.06403688964637246
	pesos_i(24317) := b"0000000000000000_0000000000000000_0001101100101101_0111101100001100"; -- 0.10616272959922449
	pesos_i(24318) := b"0000000000000000_0000000000000000_0001101111101101_1110110100100100"; -- 0.10909921777081237
	pesos_i(24319) := b"0000000000000000_0000000000000000_0010000110010011_1100111100001011"; -- 0.13116163278738086
	pesos_i(24320) := b"0000000000000000_0000000000000000_0001110010000001_1001101010111110"; -- 0.11135260704525432
	pesos_i(24321) := b"0000000000000000_0000000000000000_0000111001101111_1101011000000001"; -- 0.056393981262575395
	pesos_i(24322) := b"0000000000000000_0000000000000000_0000010000101001_1110001011001101"; -- 0.016264128664243968
	pesos_i(24323) := b"1111111111111111_1111111111111111_1111100010110010_1000111011100111"; -- -0.028525417818176108
	pesos_i(24324) := b"1111111111111111_1111111111111111_1111010111100111_0000001000100110"; -- -0.039443841668494045
	pesos_i(24325) := b"0000000000000000_0000000000000000_0000011011001001_0011100111000010"; -- 0.02650795911997388
	pesos_i(24326) := b"1111111111111111_1111111111111111_1101011001000001_0010011111011111"; -- -0.16306830217009505
	pesos_i(24327) := b"1111111111111111_1111111111111111_1110111110100111_1001001010111011"; -- -0.06384928638867168
	pesos_i(24328) := b"0000000000000000_0000000000000000_0001100100101111_1010110110010000"; -- 0.09838375812023485
	pesos_i(24329) := b"0000000000000000_0000000000000000_0000010110011001_1100010111000100"; -- 0.02187763240334698
	pesos_i(24330) := b"1111111111111111_1111111111111111_1110100010100000_0101100011100110"; -- -0.09130329508788838
	pesos_i(24331) := b"0000000000000000_0000000000000000_0000000011101001_0110111111101100"; -- 0.003561968917057875
	pesos_i(24332) := b"1111111111111111_1111111111111111_1111110000111110_0000011011001101"; -- -0.014678549755305838
	pesos_i(24333) := b"1111111111111111_1111111111111111_1101101000101010_1110010110111010"; -- -0.14778293814187907
	pesos_i(24334) := b"1111111111111111_1111111111111111_1111101101001110_1100010101001110"; -- -0.018329304079111826
	pesos_i(24335) := b"1111111111111111_1111111111111111_1101101011001100_0110001100001101"; -- -0.14531880325665497
	pesos_i(24336) := b"0000000000000000_0000000000000000_0001101100010000_1101011010101000"; -- 0.10572568503792694
	pesos_i(24337) := b"0000000000000000_0000000000000000_0000111111000111_0111110010111101"; -- 0.06163768393887548
	pesos_i(24338) := b"1111111111111111_1111111111111111_1111101111111111_0001110101000010"; -- -0.01563851492491697
	pesos_i(24339) := b"1111111111111111_1111111111111111_1110111111011101_1010100011010110"; -- -0.06302399419315788
	pesos_i(24340) := b"0000000000000000_0000000000000000_0000100110011101_0010111100010001"; -- 0.03755468531315011
	pesos_i(24341) := b"1111111111111111_1111111111111111_1111001101110011_0101101011000100"; -- -0.0490210792852992
	pesos_i(24342) := b"1111111111111111_1111111111111111_1111100011111001_1101100111011100"; -- -0.02743757608649314
	pesos_i(24343) := b"1111111111111111_1111111111111111_1111010000101101_0011001110000000"; -- -0.046185284828939105
	pesos_i(24344) := b"0000000000000000_0000000000000000_0000000110000101_0011100000010001"; -- 0.005939010729595395
	pesos_i(24345) := b"1111111111111111_1111111111111111_1110000101101111_0111101100100001"; -- -0.11939268544529798
	pesos_i(24346) := b"1111111111111111_1111111111111111_1111001000001100_0001101101011010"; -- -0.05450276421640967
	pesos_i(24347) := b"1111111111111111_1111111111111111_1111100010110001_0100011110001010"; -- -0.028544930293624808
	pesos_i(24348) := b"1111111111111111_1111111111111111_1111000000110011_1011110101000000"; -- -0.06171052158507492
	pesos_i(24349) := b"0000000000000000_0000000000000000_0000100111111010_1011110101100101"; -- 0.03898223611808233
	pesos_i(24350) := b"0000000000000000_0000000000000000_0001001111101001_0110000100110001"; -- 0.07777984079775851
	pesos_i(24351) := b"1111111111111111_1111111111111111_1111111001101101_1100010111101000"; -- -0.006137495929841363
	pesos_i(24352) := b"0000000000000000_0000000000000000_0010000001100100_1010011010101011"; -- 0.1265358130336208
	pesos_i(24353) := b"0000000000000000_0000000000000000_0001001011101001_0111111001001111"; -- 0.07387532632895218
	pesos_i(24354) := b"1111111111111111_1111111111111111_1110100000000011_1011001111010101"; -- -0.09369350469426538
	pesos_i(24355) := b"0000000000000000_0000000000000000_0010100101001100_1000101001010001"; -- 0.1613241622623325
	pesos_i(24356) := b"1111111111111111_1111111111111111_1111111101110110_1100110101101000"; -- -0.0020934696877633694
	pesos_i(24357) := b"1111111111111111_1111111111111111_1111101100001101_0000011100011110"; -- -0.019332461589749307
	pesos_i(24358) := b"1111111111111111_1111111111111111_1111010000001000_0001011000000110"; -- -0.04675161704212192
	pesos_i(24359) := b"0000000000000000_0000000000000000_0001000101001110_1010001111011110"; -- 0.06760620280870383
	pesos_i(24360) := b"1111111111111111_1111111111111111_1110100111100101_1010101100000001"; -- -0.08633929477149002
	pesos_i(24361) := b"0000000000000000_0000000000000000_0010010100000110_0000101010101111"; -- 0.14462343959952598
	pesos_i(24362) := b"1111111111111111_1111111111111111_1110100000111111_0000101111001010"; -- -0.09278799363912542
	pesos_i(24363) := b"0000000000000000_0000000000000000_0010011100111011_1000101000110011"; -- 0.1532522558149611
	pesos_i(24364) := b"0000000000000000_0000000000000000_0000101000101001_0110010001101011"; -- 0.039694095778114835
	pesos_i(24365) := b"1111111111111111_1111111111111111_1110000110011101_1001111100101101"; -- -0.11868863246142325
	pesos_i(24366) := b"0000000000000000_0000000000000000_0010000100100001_0100011100100001"; -- 0.12941402954259743
	pesos_i(24367) := b"1111111111111111_1111111111111111_1110111111110010_0100110111000110"; -- -0.06270898732981361
	pesos_i(24368) := b"0000000000000000_0000000000000000_0000001111011011_1001111011011110"; -- 0.015069894086339682
	pesos_i(24369) := b"0000000000000000_0000000000000000_0000011000100010_0010011000111101"; -- 0.023958578076706694
	pesos_i(24370) := b"0000000000000000_0000000000000000_0000111100111111_1111100001001111"; -- 0.059569854143824714
	pesos_i(24371) := b"1111111111111111_1111111111111111_1110101101100011_0010011000011010"; -- -0.0805183588658222
	pesos_i(24372) := b"1111111111111111_1111111111111111_1111010100111010_0010101010101010"; -- -0.042081197297524596
	pesos_i(24373) := b"0000000000000000_0000000000000000_0000101000000001_1010010000101101"; -- 0.03908754446611295
	pesos_i(24374) := b"1111111111111111_1111111111111111_1110101100011101_0101010000111000"; -- -0.08158372537290344
	pesos_i(24375) := b"0000000000000000_0000000000000000_0001011010111000_0110010111110111"; -- 0.08875119482094593
	pesos_i(24376) := b"1111111111111111_1111111111111111_1111111010011001_1001111010101011"; -- -0.005468447924841856
	pesos_i(24377) := b"0000000000000000_0000000000000000_0000010101000111_0110011101001010"; -- 0.020620780434436357
	pesos_i(24378) := b"0000000000000000_0000000000000000_0001001100001100_0111010111101110"; -- 0.07440888462776221
	pesos_i(24379) := b"0000000000000000_0000000000000000_0010000010000010_0110011100001011"; -- 0.1269897843208342
	pesos_i(24380) := b"0000000000000000_0000000000000000_0000001001011001_1011101101011010"; -- 0.009181699190415176
	pesos_i(24381) := b"1111111111111111_1111111111111111_1110101000010111_1101010011010001"; -- -0.08557386307258522
	pesos_i(24382) := b"1111111111111111_1111111111111111_1111001101110001_0010100001100111"; -- -0.04905459871589756
	pesos_i(24383) := b"0000000000000000_0000000000000000_0001011010000000_1111111100000101"; -- 0.08790582544784199
	pesos_i(24384) := b"0000000000000000_0000000000000000_0010000110111010_0010001000001110"; -- 0.13174641469767115
	pesos_i(24385) := b"0000000000000000_0000000000000000_0000001000111100_0111000111011100"; -- 0.008734813862164544
	pesos_i(24386) := b"0000000000000000_0000000000000000_0000011001100011_1110011111100011"; -- 0.024961941697370895
	pesos_i(24387) := b"0000000000000000_0000000000000000_0000101100111101_0100111101001000"; -- 0.043904261748061155
	pesos_i(24388) := b"0000000000000000_0000000000000000_0001110001110111_1110111010011101"; -- 0.11120501832204144
	pesos_i(24389) := b"1111111111111111_1111111111111111_1111001011111011_1100101010011010"; -- -0.05084546796106639
	pesos_i(24390) := b"1111111111111111_1111111111111111_1111010000010100_0001010001110000"; -- -0.04656860602342968
	pesos_i(24391) := b"1111111111111111_1111111111111111_1110011001001111_1110011110010111"; -- -0.10034325181052575
	pesos_i(24392) := b"0000000000000000_0000000000000000_0010001011111110_0101000111100011"; -- 0.1366931132189467
	pesos_i(24393) := b"0000000000000000_0000000000000000_0000001000100010_1000101000110101"; -- 0.008339536544412666
	pesos_i(24394) := b"1111111111111111_1111111111111111_1110100001111011_1001111100101100"; -- -0.0918636815414158
	pesos_i(24395) := b"0000000000000000_0000000000000000_0000100010010000_0011101111011011"; -- 0.03345083321735889
	pesos_i(24396) := b"1111111111111111_1111111111111111_1110000010011001_0001000001110100"; -- -0.1226644246755013
	pesos_i(24397) := b"0000000000000000_0000000000000000_0010000111001000_0011110010010000"; -- 0.13196161753799585
	pesos_i(24398) := b"1111111111111111_1111111111111111_1110011010001000_0110101010110110"; -- -0.09948094425607248
	pesos_i(24399) := b"0000000000000000_0000000000000000_0000110100000000_1001011100101101"; -- 0.050790260884354156
	pesos_i(24400) := b"1111111111111111_1111111111111111_1111100010111100_1100011011001010"; -- -0.028369498831841852
	pesos_i(24401) := b"1111111111111111_1111111111111111_1111101000011011_1011000110011110"; -- -0.02301492578090713
	pesos_i(24402) := b"1111111111111111_1111111111111111_1110101111100111_1111111011101001"; -- -0.07849127599438412
	pesos_i(24403) := b"1111111111111111_1111111111111111_1110000110001110_1000111010101010"; -- -0.11891849845618177
	pesos_i(24404) := b"0000000000000000_0000000000000000_0001001111111101_1111000101110110"; -- 0.07809361594070724
	pesos_i(24405) := b"0000000000000000_0000000000000000_0010000000101000_0111011011101011"; -- 0.12561743961877672
	pesos_i(24406) := b"1111111111111111_1111111111111111_1110110101000111_1110100111111010"; -- -0.07312142991866227
	pesos_i(24407) := b"1111111111111111_1111111111111111_1111100101010001_0101100010001100"; -- -0.026102510383793336
	pesos_i(24408) := b"1111111111111111_1111111111111111_1111010000111000_0111101011000010"; -- -0.04601319096496002
	pesos_i(24409) := b"0000000000000000_0000000000000000_0000100011001010_0100110101010111"; -- 0.03433688530271595
	pesos_i(24410) := b"1111111111111111_1111111111111111_1110000011010010_0000001110101010"; -- -0.12179543580614766
	pesos_i(24411) := b"1111111111111111_1111111111111111_1101101100100001_0000010111101011"; -- -0.14402735724915133
	pesos_i(24412) := b"1111111111111111_1111111111111111_1110011011000111_0001111100101101"; -- -0.09852414276957963
	pesos_i(24413) := b"1111111111111111_1111111111111111_1101110001010010_1010010110110100"; -- -0.13936390255370412
	pesos_i(24414) := b"1111111111111111_1111111111111111_1111001100101001_0100011001010000"; -- -0.05015144875548591
	pesos_i(24415) := b"1111111111111111_1111111111111111_1110000010100011_1110000101100101"; -- -0.12249938274952536
	pesos_i(24416) := b"0000000000000000_0000000000000000_0000000100010000_1000011101001001"; -- 0.004158454213527555
	pesos_i(24417) := b"0000000000000000_0000000000000000_0000110100110010_0111011111000101"; -- 0.05155132823151441
	pesos_i(24418) := b"1111111111111111_1111111111111111_1101110100001010_0010000001010111"; -- -0.13656423451744662
	pesos_i(24419) := b"0000000000000000_0000000000000000_0001100000010011_1111011000011001"; -- 0.09405458553178968
	pesos_i(24420) := b"0000000000000000_0000000000000000_0001010101001000_0111001101011010"; -- 0.08313675822493433
	pesos_i(24421) := b"0000000000000000_0000000000000000_0010001010001000_0011010100111010"; -- 0.13489086778189344
	pesos_i(24422) := b"0000000000000000_0000000000000000_0000010001000000_0110000111011100"; -- 0.016607395472233586
	pesos_i(24423) := b"1111111111111111_1111111111111111_1111100010110110_0101101101010001"; -- -0.028467457475883348
	pesos_i(24424) := b"1111111111111111_1111111111111111_1110010101000000_1000011010011000"; -- -0.10448416503312508
	pesos_i(24425) := b"1111111111111111_1111111111111111_1111100000101011_1010010001111101"; -- -0.030584067870012575
	pesos_i(24426) := b"0000000000000000_0000000000000000_0001101111000101_0111000010100011"; -- 0.1084814452304653
	pesos_i(24427) := b"1111111111111111_1111111111111111_1101011110100011_1001111011011001"; -- -0.15765959938848942
	pesos_i(24428) := b"0000000000000000_0000000000000000_0000011001000101_1010010001011011"; -- 0.024500152766273948
	pesos_i(24429) := b"0000000000000000_0000000000000000_0001010101010010_0100110101111001"; -- 0.08328708848461158
	pesos_i(24430) := b"1111111111111111_1111111111111111_1101111010110010_0011000010110111"; -- -0.13009353185645664
	pesos_i(24431) := b"0000000000000000_0000000000000000_0010000111101111_0001110100111100"; -- 0.13255484298870518
	pesos_i(24432) := b"0000000000000000_0000000000000000_0001111010010000_0111101110011111"; -- 0.11939213390126469
	pesos_i(24433) := b"1111111111111111_1111111111111111_1111001000111010_0001010010011001"; -- -0.05380126252186566
	pesos_i(24434) := b"0000000000000000_0000000000000000_0000011010010110_0010111111011100"; -- 0.025729170982923842
	pesos_i(24435) := b"0000000000000000_0000000000000000_0001101100111010_1110010101000001"; -- 0.10636742447557744
	pesos_i(24436) := b"0000000000000000_0000000000000000_0001101100100011_0010001111000110"; -- 0.10600493990795412
	pesos_i(24437) := b"0000000000000000_0000000000000000_0010000000011100_0100110111010100"; -- 0.1254318849951959
	pesos_i(24438) := b"1111111111111111_1111111111111111_1101111010010011_0100011101100011"; -- -0.13056520308052977
	pesos_i(24439) := b"0000000000000000_0000000000000000_0001010010010000_0101011001001010"; -- 0.0803274087559142
	pesos_i(24440) := b"0000000000000000_0000000000000000_0001100101101110_1001100110111100"; -- 0.09934388018956199
	pesos_i(24441) := b"1111111111111111_1111111111111111_1110001101100010_0111110110010011"; -- -0.11177840378660403
	pesos_i(24442) := b"1111111111111111_1111111111111111_1101101000011010_0000001111100101"; -- -0.14804053944464463
	pesos_i(24443) := b"0000000000000000_0000000000000000_0000100010011111_1000111000100001"; -- 0.03368461901690349
	pesos_i(24444) := b"0000000000000000_0000000000000000_0000101010111000_1101000100110001"; -- 0.041882585973217715
	pesos_i(24445) := b"0000000000000000_0000000000000000_0010011000010010_1011000001110010"; -- 0.14872267523941157
	pesos_i(24446) := b"0000000000000000_0000000000000000_0000100000001010_0111100000011111"; -- 0.03140974755114222
	pesos_i(24447) := b"1111111111111111_1111111111111111_1101101111010101_0100010110000111"; -- -0.14127698385696763
	pesos_i(24448) := b"1111111111111111_1111111111111111_1111010000111100_1010110111101010"; -- -0.04594910661721836
	pesos_i(24449) := b"1111111111111111_1111111111111111_1101100010110101_1010100011001101"; -- -0.15347809780368657
	pesos_i(24450) := b"1111111111111111_1111111111111111_1110111110100010_0001110010101011"; -- -0.06393261734657961
	pesos_i(24451) := b"1111111111111111_1111111111111111_1110011001100101_1111100100010101"; -- -0.10000651590922872
	pesos_i(24452) := b"0000000000000000_0000000000000000_0000000100000101_0010010110010110"; -- 0.003984784267023384
	pesos_i(24453) := b"0000000000000000_0000000000000000_0000001100010111_0101000100101101"; -- 0.01207454065989335
	pesos_i(24454) := b"0000000000000000_0000000000000000_0001011100101001_0101101111100100"; -- 0.09047483742120609
	pesos_i(24455) := b"1111111111111111_1111111111111111_1111100110110101_0101000011110010"; -- -0.02457708441668096
	pesos_i(24456) := b"1111111111111111_1111111111111111_1101110001101000_1101100111010100"; -- -0.1390251023597862
	pesos_i(24457) := b"0000000000000000_0000000000000000_0000001000100111_1010001001111000"; -- 0.008417276777498607
	pesos_i(24458) := b"0000000000000000_0000000000000000_0001101110010101_0110000101100001"; -- 0.10774811371579784
	pesos_i(24459) := b"1111111111111111_1111111111111111_1110001000110101_1111111000101010"; -- -0.11636363474063964
	pesos_i(24460) := b"0000000000000000_0000000000000000_0000001110110101_0000001101010011"; -- 0.014480788920740836
	pesos_i(24461) := b"1111111111111111_1111111111111111_1110111100101100_0001110101100101"; -- -0.06573311128732694
	pesos_i(24462) := b"0000000000000000_0000000000000000_0000000010001011_0111110011111011"; -- 0.0021284210937073827
	pesos_i(24463) := b"1111111111111111_1111111111111111_1111000101001000_0011011101101001"; -- -0.057491814416935454
	pesos_i(24464) := b"0000000000000000_0000000000000000_0001001111110100_0000011101000001"; -- 0.07794232693492234
	pesos_i(24465) := b"0000000000000000_0000000000000000_0000001010110011_1010000101011010"; -- 0.010553440659041255
	pesos_i(24466) := b"1111111111111111_1111111111111111_1111001110100101_0110101001001011"; -- -0.04825721432711362
	pesos_i(24467) := b"1111111111111111_1111111111111111_1111100010011000_1101000001100101"; -- -0.028918242711732958
	pesos_i(24468) := b"0000000000000000_0000000000000000_0010000101001000_0010000011111100"; -- 0.13000684894274328
	pesos_i(24469) := b"0000000000000000_0000000000000000_0001111001010000_0100011101110111"; -- 0.11841246280286048
	pesos_i(24470) := b"1111111111111111_1111111111111111_1111110011011010_1110101010110011"; -- -0.012284594733756064
	pesos_i(24471) := b"1111111111111111_1111111111111111_1110011011011100_1010110111000110"; -- -0.09819520862253044
	pesos_i(24472) := b"0000000000000000_0000000000000000_0001000111111011_1111010001101001"; -- 0.07025077392643059
	pesos_i(24473) := b"0000000000000000_0000000000000000_0010011000010011_1110000111010010"; -- 0.14874087685459303
	pesos_i(24474) := b"0000000000000000_0000000000000000_0000001110001010_0101110011100111"; -- 0.01383000031086654
	pesos_i(24475) := b"1111111111111111_1111111111111111_1111001001111111_1010010111111100"; -- -0.05273974024565521
	pesos_i(24476) := b"1111111111111111_1111111111111111_1110111001110110_1001001000000000"; -- -0.06850326060613385
	pesos_i(24477) := b"0000000000000000_0000000000000000_0010010011111101_0100110111110110"; -- 0.1444901203678001
	pesos_i(24478) := b"1111111111111111_1111111111111111_1111101110011111_1000001100110110"; -- -0.01709728180961796
	pesos_i(24479) := b"0000000000000000_0000000000000000_0010011001111111_1001010000011111"; -- 0.15038419486512317
	pesos_i(24480) := b"1111111111111111_1111111111111111_1101101000001110_0001101011011001"; -- -0.1482222767264559
	pesos_i(24481) := b"0000000000000000_0000000000000000_0001010001010100_0110110110011111"; -- 0.07941327219877718
	pesos_i(24482) := b"1111111111111111_1111111111111111_1111101101010001_0001110001011001"; -- -0.018293598539228777
	pesos_i(24483) := b"1111111111111111_1111111111111111_1110100111111011_1111110010111000"; -- -0.08599873081999626
	pesos_i(24484) := b"0000000000000000_0000000000000000_0000101111101110_1110101100000111"; -- 0.04661435044348331
	pesos_i(24485) := b"0000000000000000_0000000000000000_0001110110100100_1010110101001101"; -- 0.11579402097251795
	pesos_i(24486) := b"0000000000000000_0000000000000000_0001101011101100_1100001100000100"; -- 0.1051751980328097
	pesos_i(24487) := b"0000000000000000_0000000000000000_0010010101100110_0111000000110101"; -- 0.14609433452357562
	pesos_i(24488) := b"0000000000000000_0000000000000000_0001100100010100_0010100111000010"; -- 0.09796391477845988
	pesos_i(24489) := b"0000000000000000_0000000000000000_0010001011111010_1100111000101101"; -- 0.1366394862788026
	pesos_i(24490) := b"0000000000000000_0000000000000000_0001000010110010_0010100111000011"; -- 0.06521855375424214
	pesos_i(24491) := b"1111111111111111_1111111111111111_1101111101000011_0001000011101101"; -- -0.12788290220651555
	pesos_i(24492) := b"1111111111111111_1111111111111111_1111101110011010_1011010011111011"; -- -0.017170609134961632
	pesos_i(24493) := b"1111111111111111_1111111111111111_1110101010110101_0001111000011010"; -- -0.08317386495424456
	pesos_i(24494) := b"0000000000000000_0000000000000000_0001011000010011_1000000010101101"; -- 0.08623508668211328
	pesos_i(24495) := b"1111111111111111_1111111111111111_1111110011011101_0111010011100110"; -- -0.012245840015830982
	pesos_i(24496) := b"0000000000000000_0000000000000000_0000011001010110_1111011111100101"; -- 0.024764531458336844
	pesos_i(24497) := b"0000000000000000_0000000000000000_0001011110101101_1101101001101011"; -- 0.0924965391906029
	pesos_i(24498) := b"1111111111111111_1111111111111111_1111110100011101_0011001100111110"; -- -0.011273190775034152
	pesos_i(24499) := b"1111111111111111_1111111111111111_1111011000111001_1010110100111010"; -- -0.038182423802053625
	pesos_i(24500) := b"1111111111111111_1111111111111111_1111011010111010_1011011000011111"; -- -0.03621350995857328
	pesos_i(24501) := b"1111111111111111_1111111111111111_1110010100100101_1100111001010110"; -- -0.10489187627712018
	pesos_i(24502) := b"1111111111111111_1111111111111111_1110110000101101_1000010100010101"; -- -0.0774304221629492
	pesos_i(24503) := b"1111111111111111_1111111111111111_1110111100111111_0111010100000001"; -- -0.06543797229470492
	pesos_i(24504) := b"0000000000000000_0000000000000000_0000010001100000_1010100001101110"; -- 0.017099882980966995
	pesos_i(24505) := b"0000000000000000_0000000000000000_0001011000011010_0001010100011001"; -- 0.08633548611650779
	pesos_i(24506) := b"0000000000000000_0000000000000000_0000110110110010_0111001000000010"; -- 0.053504109846012025
	pesos_i(24507) := b"0000000000000000_0000000000000000_0000011000010110_0101100111111100"; -- 0.023778556888322682
	pesos_i(24508) := b"0000000000000000_0000000000000000_0000000011001011_1011111110100110"; -- 0.0031089572143118433
	pesos_i(24509) := b"1111111111111111_1111111111111111_1110110011011000_1101001111111110"; -- -0.0748164658919484
	pesos_i(24510) := b"0000000000000000_0000000000000000_0001000100111110_0010110101101001"; -- 0.06735500147315422
	pesos_i(24511) := b"1111111111111111_1111111111111111_1101110100111100_1111110001101011"; -- -0.13578817726557246
	pesos_i(24512) := b"1111111111111111_1111111111111111_1101111111010010_1000100001100110"; -- -0.12569377428639397
	pesos_i(24513) := b"1111111111111111_1111111111111111_1111100111101000_1000111010001001"; -- -0.023795215241406095
	pesos_i(24514) := b"0000000000000000_0000000000000000_0001111000101100_0010111000010101"; -- 0.11786163343598441
	pesos_i(24515) := b"1111111111111111_1111111111111111_1110000001001110_0000111011001111"; -- -0.12380893174259433
	pesos_i(24516) := b"1111111111111111_1111111111111111_1111100111111000_1101110001001010"; -- -0.023546439999962355
	pesos_i(24517) := b"1111111111111111_1111111111111111_1110100110111110_0110111110100101"; -- -0.08693792546495006
	pesos_i(24518) := b"1111111111111111_1111111111111111_1101110110111011_1101011011000001"; -- -0.13385255601415194
	pesos_i(24519) := b"0000000000000000_0000000000000000_0010010101001111_0001011111010011"; -- 0.14573811428669198
	pesos_i(24520) := b"0000000000000000_0000000000000000_0001101001101110_1000110001011111"; -- 0.10324933362218858
	pesos_i(24521) := b"0000000000000000_0000000000000000_0001110100111001_1000111011101111"; -- 0.11415952050878835
	pesos_i(24522) := b"0000000000000000_0000000000000000_0000001101101000_0000111011100111"; -- 0.013306552259560143
	pesos_i(24523) := b"0000000000000000_0000000000000000_0000011101010001_0000010001101010"; -- 0.028579974974156555
	pesos_i(24524) := b"0000000000000000_0000000000000000_0000111011110011_0011101001001101"; -- 0.05839886082463034
	pesos_i(24525) := b"1111111111111111_1111111111111111_1111100000101110_0011110110010011"; -- -0.030544425650231462
	pesos_i(24526) := b"0000000000000000_0000000000000000_0010010001100011_1011101100001010"; -- 0.14214676839999682
	pesos_i(24527) := b"0000000000000000_0000000000000000_0001110101000011_1101110010110110"; -- 0.11431674435726118
	pesos_i(24528) := b"1111111111111111_1111111111111111_1110100111110010_0001001011011101"; -- -0.0861499987506342
	pesos_i(24529) := b"0000000000000000_0000000000000000_0001011111010001_0010100001000101"; -- 0.09303523722615756
	pesos_i(24530) := b"0000000000000000_0000000000000000_0010011100001101_1000011000010001"; -- 0.1525501052933527
	pesos_i(24531) := b"1111111111111111_1111111111111111_1110000010111010_0110101001011010"; -- -0.12215552628044496
	pesos_i(24532) := b"1111111111111111_1111111111111111_1110010011111011_1101010110110001"; -- -0.1055323069614956
	pesos_i(24533) := b"0000000000000000_0000000000000000_0010001010010110_1111001110010110"; -- 0.13511583719136463
	pesos_i(24534) := b"1111111111111111_1111111111111111_1111100111000010_1100110100010110"; -- -0.02437132083272972
	pesos_i(24535) := b"1111111111111111_1111111111111111_1101111100000000_0100011000000100"; -- -0.1289020766549362
	pesos_i(24536) := b"1111111111111111_1111111111111111_1101111101000000_0110011000100011"; -- -0.12792359961606098
	pesos_i(24537) := b"0000000000000000_0000000000000000_0000100110010110_1000000111100111"; -- 0.037452811043386644
	pesos_i(24538) := b"0000000000000000_0000000000000000_0001000101101011_1000101010110001"; -- 0.06804720717912097
	pesos_i(24539) := b"1111111111111111_1111111111111111_1110011111110100_0110001110110011"; -- -0.0939271630425237
	pesos_i(24540) := b"1111111111111111_1111111111111111_1101110100111010_1110000001100110"; -- -0.1358203649800642
	pesos_i(24541) := b"1111111111111111_1111111111111111_1110000000100010_0000001100111011"; -- -0.12448100855288889
	pesos_i(24542) := b"0000000000000000_0000000000000000_0001000100001011_0000101011000111"; -- 0.06657473897793008
	pesos_i(24543) := b"0000000000000000_0000000000000000_0010010001100000_1000001101110101"; -- 0.14209767918550836
	pesos_i(24544) := b"1111111111111111_1111111111111111_1111101101010011_1011001110010011"; -- -0.018254067145531568
	pesos_i(24545) := b"0000000000000000_0000000000000000_0001111000000101_0011000100000101"; -- 0.11726671579814035
	pesos_i(24546) := b"0000000000000000_0000000000000000_0010011001000100_0001011110010111"; -- 0.1494765036136166
	pesos_i(24547) := b"1111111111111111_1111111111111111_1111011101001011_1000111000000101"; -- -0.03400337578636846
	pesos_i(24548) := b"0000000000000000_0000000000000000_0001110011111010_0001001100101100"; -- 0.11319084010780571
	pesos_i(24549) := b"0000000000000000_0000000000000000_0000110101111011_0111110101001111"; -- 0.052665549982785526
	pesos_i(24550) := b"1111111111111111_1111111111111111_1101110000101011_0101000100001000"; -- -0.1399640421795697
	pesos_i(24551) := b"1111111111111111_1111111111111111_1110001011011011_1111011011000101"; -- -0.1138311166417909
	pesos_i(24552) := b"1111111111111111_1111111111111111_1111101011101011_0011100101100111"; -- -0.019848263028992407
	pesos_i(24553) := b"1111111111111111_1111111111111111_1110110110111100_1110011001000101"; -- -0.07133637259073355
	pesos_i(24554) := b"0000000000000000_0000000000000000_0001001001111000_1000011000111110"; -- 0.0721515562031939
	pesos_i(24555) := b"1111111111111111_1111111111111111_1110011100101001_0101110010100011"; -- -0.09702511809440599
	pesos_i(24556) := b"0000000000000000_0000000000000000_0000011011110010_0100010001110011"; -- 0.02713420675169172
	pesos_i(24557) := b"0000000000000000_0000000000000000_0000111111000111_1100011011110001"; -- 0.06164210696920044
	pesos_i(24558) := b"1111111111111111_1111111111111111_1110010001000110_0110010111000110"; -- -0.10830081868285125
	pesos_i(24559) := b"1111111111111111_1111111111111111_1110100101101010_0100000110000111"; -- -0.08822241255216397
	pesos_i(24560) := b"1111111111111111_1111111111111111_1101110010111001_0001111001000001"; -- -0.13780032081111723
	pesos_i(24561) := b"1111111111111111_1111111111111111_1101100100000001_1110100010101110"; -- -0.15231462237684013
	pesos_i(24562) := b"1111111111111111_1111111111111111_1101101011100000_0101110101110001"; -- -0.14501396169858852
	pesos_i(24563) := b"1111111111111111_1111111111111111_1101101011001100_1110000010011110"; -- -0.14531131885393134
	pesos_i(24564) := b"1111111111111111_1111111111111111_1110000101001011_1111011010010001"; -- -0.1199346442154787
	pesos_i(24565) := b"1111111111111111_1111111111111111_1111001100110011_1111111100110100"; -- -0.04998784051881629
	pesos_i(24566) := b"1111111111111111_1111111111111111_1111110000100001_1001101001001001"; -- -0.0151122638313641
	pesos_i(24567) := b"1111111111111111_1111111111111111_1111111001111100_1101100110010100"; -- -0.005907441566459403
	pesos_i(24568) := b"1111111111111111_1111111111111111_1111001111110000_1001011100001000"; -- -0.04711013849348865
	pesos_i(24569) := b"0000000000000000_0000000000000000_0001000110111011_0111101100000111"; -- 0.06926697659574486
	pesos_i(24570) := b"1111111111111111_1111111111111111_1111011001111001_1100111001100110"; -- -0.03720388417297736
	pesos_i(24571) := b"1111111111111111_1111111111111111_1111100000000111_1000010111010001"; -- -0.031135212344953297
	pesos_i(24572) := b"1111111111111111_1111111111111111_1110000010001100_1101110010100101"; -- -0.12285061805324611
	pesos_i(24573) := b"1111111111111111_1111111111111111_1101101111010110_1001001011000010"; -- -0.1412571215827844
	pesos_i(24574) := b"1111111111111111_1111111111111111_1111000110101001_0010111100011110"; -- -0.05601220629607694
	pesos_i(24575) := b"1111111111111111_1111111111111111_1101110000010101_0100101010010111"; -- -0.14030011954696586
	pesos_i(24576) := b"1111111111111111_1111111111111111_1101011100101111_1100010010010100"; -- -0.15942736995182782
	pesos_i(24577) := b"0000000000000000_0000000000000000_0000000101110000_1100110011101101"; -- 0.0056274488698367315
	pesos_i(24578) := b"0000000000000000_0000000000000000_0010100001001010_1100110111110101"; -- 0.1573914264802679
	pesos_i(24579) := b"1111111111111111_1111111111111111_1101000100010000_0000100110001101"; -- -0.1833490402083972
	pesos_i(24580) := b"0000000000000000_0000000000000000_0010111110000110_0000111001111101"; -- 0.1856392912401388
	pesos_i(24581) := b"0000000000000000_0000000000000000_0011000100101110_0110111100010010"; -- 0.1921147745963534
	pesos_i(24582) := b"1111111111111111_1111111111111111_1101100111110100_0001011000100010"; -- -0.14861928625047044
	pesos_i(24583) := b"0000000000000000_0000000000000000_0001001111001000_1101100011001001"; -- 0.07728342919962337
	pesos_i(24584) := b"1111111111111111_1111111111111111_1111110110111101_1010110100010011"; -- -0.008824522741994134
	pesos_i(24585) := b"0000000000000000_0000000000000000_0010111010111110_0111110010101000"; -- 0.18259410000132803
	pesos_i(24586) := b"1111111111111111_1111111111111111_1110011110101010_0100011110101110"; -- -0.09505798330885533
	pesos_i(24587) := b"1111111111111111_1111111111111111_1110101000111101_1111001111011101"; -- -0.08499217842505527
	pesos_i(24588) := b"0000000000000000_0000000000000000_0000100100101000_1001001001001000"; -- 0.035775320567056
	pesos_i(24589) := b"1111111111111111_1111111111111111_1110011001110000_0101000100101001"; -- -0.0998486781956041
	pesos_i(24590) := b"1111111111111111_1111111111111111_1101110001101101_0001101010000111"; -- -0.13896021078075252
	pesos_i(24591) := b"0000000000000000_0000000000000000_0001001100111011_0001001011111101"; -- 0.07512015023346466
	pesos_i(24592) := b"1111111111111111_1111111111111111_1111111000001101_1011111101110000"; -- -0.007602725268268705
	pesos_i(24593) := b"1111111111111111_1111111111111111_1110000111000000_0001001100111111"; -- -0.11816291524180658
	pesos_i(24594) := b"0000000000000000_0000000000000000_0000001001101111_1101100010000010"; -- 0.009519130433049899
	pesos_i(24595) := b"0000000000000000_0000000000000000_0010110010001111_0010000100011100"; -- 0.17405898030199277
	pesos_i(24596) := b"1111111111111111_1111111111111111_1100110101000101_1010001110101010"; -- -0.1981561383449027
	pesos_i(24597) := b"1111111111111111_1111111111111111_1101101010011011_0000000001010100"; -- -0.14607236810648513
	pesos_i(24598) := b"0000000000000000_0000000000000000_0010001011100101_1111101010001010"; -- 0.13632169598459176
	pesos_i(24599) := b"1111111111111111_1111111111111111_1110111111100110_0111100111010001"; -- -0.06288946778233653
	pesos_i(24600) := b"0000000000000000_0000000000000000_0001010101011000_0000101111101001"; -- 0.08337473324015493
	pesos_i(24601) := b"1111111111111111_1111111111111111_1101010100100111_0000110100100100"; -- -0.16737287407838897
	pesos_i(24602) := b"1111111111111111_1111111111111111_1111010011110011_1010001110001101"; -- -0.04315736583832078
	pesos_i(24603) := b"1111111111111111_1111111111111111_1111101010001010_1011001011111101"; -- -0.021321118633727078
	pesos_i(24604) := b"0000000000000000_0000000000000000_0010101111001100_1001100111111110"; -- 0.17109072173093062
	pesos_i(24605) := b"0000000000000000_0000000000000000_0001011100000110_0111100100010100"; -- 0.08994251955940827
	pesos_i(24606) := b"1111111111111111_1111111111111111_1111000110110011_1101001111011110"; -- -0.055849798466512106
	pesos_i(24607) := b"1111111111111111_1111111111111111_1101010100001001_1011110101111001"; -- -0.16782012752452782
	pesos_i(24608) := b"1111111111111111_1111111111111111_1101000001010010_0001000001100011"; -- -0.18624780259118595
	pesos_i(24609) := b"0000000000000000_0000000000000000_0010010101100000_0110001010000111"; -- 0.1460019663480673
	pesos_i(24610) := b"1111111111111111_1111111111111111_1110101001110100_0000011010110110"; -- -0.08416708049366842
	pesos_i(24611) := b"1111111111111111_1111111111111111_1111001010101010_0100101100011100"; -- -0.052089028933709515
	pesos_i(24612) := b"0000000000000000_0000000000000000_0001101000011101_1001100010010110"; -- 0.10201409979911985
	pesos_i(24613) := b"0000000000000000_0000000000000000_0000000000000100_1000010011101000"; -- 6.895687154225869e-05
	pesos_i(24614) := b"0000000000000000_0000000000000000_0000100111000001_1001000001100010"; -- 0.03810980207993676
	pesos_i(24615) := b"1111111111111111_1111111111111111_1111111110000011_0011110001110001"; -- -0.0019037459906975172
	pesos_i(24616) := b"0000000000000000_0000000000000000_0000010011101000_0101100011010111"; -- 0.01917033422686707
	pesos_i(24617) := b"1111111111111111_1111111111111111_1110111110100101_1011011001111001"; -- -0.0638776735440116
	pesos_i(24618) := b"1111111111111111_1111111111111111_1101101110110100_1010101110111011"; -- -0.1417744319859773
	pesos_i(24619) := b"1111111111111111_1111111111111111_1101011111101101_1001001100100011"; -- -0.1565311469113713
	pesos_i(24620) := b"0000000000000000_0000000000000000_0000101100100100_1110001010101001"; -- 0.04353157640951885
	pesos_i(24621) := b"0000000000000000_0000000000000000_0010110000100100_1000100100010010"; -- 0.17243248649867518
	pesos_i(24622) := b"1111111111111111_1111111111111111_1111100110000011_0100111110110010"; -- -0.025340098372337548
	pesos_i(24623) := b"1111111111111111_1111111111111111_1101000000000111_0010101001101011"; -- -0.18739066008645117
	pesos_i(24624) := b"1111111111111111_1111111111111111_1101011100011000_1101011100010011"; -- -0.15977721964584599
	pesos_i(24625) := b"0000000000000000_0000000000000000_0010101010110011_1000011001111110"; -- 0.16680183966514656
	pesos_i(24626) := b"1111111111111111_1111111111111111_1101011110111111_0010001100000010"; -- -0.15723973467620012
	pesos_i(24627) := b"0000000000000000_0000000000000000_0010101001010110_1010011001010101"; -- 0.1653846699237718
	pesos_i(24628) := b"0000000000000000_0000000000000000_0000100101001011_1010010001111011"; -- 0.03631046287263488
	pesos_i(24629) := b"0000000000000000_0000000000000000_0010001111101111_1101110100001000"; -- 0.14037877512608363
	pesos_i(24630) := b"1111111111111111_1111111111111111_1110100011011000_0110101111110100"; -- -0.09044766697615167
	pesos_i(24631) := b"0000000000000000_0000000000000000_0010000001011101_1111001101100111"; -- 0.12643357531408653
	pesos_i(24632) := b"1111111111111111_1111111111111111_1110110110010110_0001101100100001"; -- -0.0719283145174913
	pesos_i(24633) := b"1111111111111111_1111111111111111_1110011101001011_0111111001001100"; -- -0.09650431291233813
	pesos_i(24634) := b"0000000000000000_0000000000000000_0001000001001010_1010100101001110"; -- 0.06363924167499077
	pesos_i(24635) := b"1111111111111111_1111111111111111_1111011001000110_0011010011001111"; -- -0.03799123708458622
	pesos_i(24636) := b"1111111111111111_1111111111111111_1111011011001001_1111101111001011"; -- -0.03598047529343832
	pesos_i(24637) := b"1111111111111111_1111111111111111_1111010001111000_0011111101111011"; -- -0.04504016158026466
	pesos_i(24638) := b"1111111111111111_1111111111111111_1110101111010000_0010110110000100"; -- -0.07885470884489099
	pesos_i(24639) := b"0000000000000000_0000000000000000_0001111110110001_1010100001110011"; -- 0.12380459593497663
	pesos_i(24640) := b"1111111111111111_1111111111111111_1101001110101111_0000001000010000"; -- -0.17311083891186888
	pesos_i(24641) := b"1111111111111111_1111111111111111_1111111000100100_0110101101110011"; -- -0.007256779013958645
	pesos_i(24642) := b"1111111111111111_1111111111111111_1111010011001111_1111000000110111"; -- -0.04370211280328939
	pesos_i(24643) := b"1111111111111111_1111111111111111_1111101001111010_1000110101101110"; -- -0.021567497787249146
	pesos_i(24644) := b"0000000000000000_0000000000000000_0001001000101101_1011101110110100"; -- 0.07101033351578748
	pesos_i(24645) := b"1111111111111111_1111111111111111_1111010111101111_1010011111100001"; -- -0.03931189308033227
	pesos_i(24646) := b"0000000000000000_0000000000000000_0010111010011111_0100011110110110"; -- 0.18211792178144556
	pesos_i(24647) := b"0000000000000000_0000000000000000_0001110011100111_0000111110101111"; -- 0.11290071513142848
	pesos_i(24648) := b"1111111111111111_1111111111111111_1111000110011000_0111001011111010"; -- -0.05626756097811602
	pesos_i(24649) := b"0000000000000000_0000000000000000_0010101101010100_0001000010010001"; -- 0.16925147578202576
	pesos_i(24650) := b"1111111111111111_1111111111111111_1110000010000000_1111101110101101"; -- -0.12303187402346605
	pesos_i(24651) := b"1111111111111111_1111111111111111_1110111001100100_1011010101101100"; -- -0.06877580759888491
	pesos_i(24652) := b"0000000000000000_0000000000000000_0010111001111100_1101011101110010"; -- 0.18159243127936975
	pesos_i(24653) := b"0000000000000000_0000000000000000_0001001011101000_1001010000000001"; -- 0.07386136067181044
	pesos_i(24654) := b"1111111111111111_1111111111111111_1101010111111100_0011010000011101"; -- -0.16412042887037348
	pesos_i(24655) := b"0000000000000000_0000000000000000_0010010001010011_1000000100100111"; -- 0.14189917754637432
	pesos_i(24656) := b"0000000000000000_0000000000000000_0001101010100110_0111101111111001"; -- 0.10410284842482022
	pesos_i(24657) := b"0000000000000000_0000000000000000_0000011110110101_1010000001101101"; -- 0.030115152987123934
	pesos_i(24658) := b"1111111111111111_1111111111111111_1110110001100010_1010010111010110"; -- -0.07661975408228283
	pesos_i(24659) := b"1111111111111111_1111111111111111_1111100010001001_0101110010100000"; -- -0.02915402507760619
	pesos_i(24660) := b"1111111111111111_1111111111111111_1101111010101111_1111100011111001"; -- -0.13012737190743728
	pesos_i(24661) := b"1111111111111111_1111111111111111_1100111011000101_0101110100000001"; -- -0.1923009751483687
	pesos_i(24662) := b"1111111111111111_1111111111111111_1101001000001111_0111110100010101"; -- -0.17945116263183616
	pesos_i(24663) := b"1111111111111111_1111111111111111_1111011110010100_1001111110111011"; -- -0.032888428455567914
	pesos_i(24664) := b"0000000000000000_0000000000000000_0010101000101000_0101000011011110"; -- 0.16467767171156075
	pesos_i(24665) := b"1111111111111111_1111111111111111_1111110101110000_1110010101011100"; -- -0.009996094732607838
	pesos_i(24666) := b"0000000000000000_0000000000000000_0010000000100000_0001001101101110"; -- 0.1254894392825438
	pesos_i(24667) := b"0000000000000000_0000000000000000_0010101010111110_1101100100001010"; -- 0.16697460652821214
	pesos_i(24668) := b"0000000000000000_0000000000000000_0000110101000101_1101101111111110"; -- 0.051847219059176164
	pesos_i(24669) := b"0000000000000000_0000000000000000_0010000011001011_1011010111111111"; -- 0.12810838196342128
	pesos_i(24670) := b"0000000000000000_0000000000000000_0010101111011000_0001001010000010"; -- 0.17126575147455517
	pesos_i(24671) := b"0000000000000000_0000000000000000_0010010110111010_1011110010111100"; -- 0.1473806341674289
	pesos_i(24672) := b"1111111111111111_1111111111111111_1101000110101001_0000000011110001"; -- -0.18101495842643925
	pesos_i(24673) := b"0000000000000000_0000000000000000_0010111000000111_1100011001010100"; -- 0.17980613290314534
	pesos_i(24674) := b"0000000000000000_0000000000000000_0001010010111011_1110111010111111"; -- 0.08099262396931993
	pesos_i(24675) := b"0000000000000000_0000000000000000_0000111010000000_1101001110101011"; -- 0.056653241443652476
	pesos_i(24676) := b"0000000000000000_0000000000000000_0010111010100111_1010111010101010"; -- 0.1822461285005513
	pesos_i(24677) := b"0000000000000000_0000000000000000_0001100100011010_0010001110110101"; -- 0.09805510693261005
	pesos_i(24678) := b"1111111111111111_1111111111111111_1110000001111110_0010000111000011"; -- -0.12307538027643156
	pesos_i(24679) := b"1111111111111111_1111111111111111_1111101110010001_0110001001001101"; -- -0.017312866324150078
	pesos_i(24680) := b"0000000000000000_0000000000000000_0001100010111011_0011110011110001"; -- 0.09660702597043783
	pesos_i(24681) := b"1111111111111111_1111111111111111_1111001101000100_1101111101110011"; -- -0.04973033376468772
	pesos_i(24682) := b"0000000000000000_0000000000000000_0001001100011101_0001010101000101"; -- 0.07466252272317507
	pesos_i(24683) := b"1111111111111111_1111111111111111_1111010011100010_1100110001101011"; -- -0.04341432942715479
	pesos_i(24684) := b"1111111111111111_1111111111111111_1110000010001100_0000000110010100"; -- -0.12286367536266922
	pesos_i(24685) := b"0000000000000000_0000000000000000_0010011011001000_0100101010010101"; -- 0.15149370331854195
	pesos_i(24686) := b"0000000000000000_0000000000000000_0001101010010000_1010001010010101"; -- 0.10376945637297728
	pesos_i(24687) := b"1111111111111111_1111111111111111_1111010001101011_0000111011100001"; -- -0.045241422732514316
	pesos_i(24688) := b"1111111111111111_1111111111111111_1100110001000111_0001001110001110"; -- -0.20204046050888405
	pesos_i(24689) := b"1111111111111111_1111111111111111_1101110011001110_1011010010011001"; -- -0.1374709249031162
	pesos_i(24690) := b"0000000000000000_0000000000000000_0010011000011001_1111101001101000"; -- 0.14883389520092768
	pesos_i(24691) := b"1111111111111111_1111111111111111_1110100100101111_0101111110010000"; -- -0.08912089083992382
	pesos_i(24692) := b"1111111111111111_1111111111111111_1110001101001010_1111011101111101"; -- -0.11213734809093089
	pesos_i(24693) := b"0000000000000000_0000000000000000_0010111101101001_0101000010101011"; -- 0.1852007310731957
	pesos_i(24694) := b"0000000000000000_0000000000000000_0010100111001010_0000000111101111"; -- 0.16323864062791202
	pesos_i(24695) := b"1111111111111111_1111111111111111_1110111011001111_0000011101011111"; -- -0.0671534912558152
	pesos_i(24696) := b"1111111111111111_1111111111111111_1110010010011111_0010100011010110"; -- -0.10694641858081619
	pesos_i(24697) := b"0000000000000000_0000000000000000_0000001011111010_1100010111101010"; -- 0.011638993898018743
	pesos_i(24698) := b"1111111111111111_1111111111111111_1110110111100000_1001100001011111"; -- -0.07079169920499895
	pesos_i(24699) := b"0000000000000000_0000000000000000_0000101000100111_1011110001101010"; -- 0.039668823026454865
	pesos_i(24700) := b"1111111111111111_1111111111111111_1111011010010000_1110111010011001"; -- -0.03685101280326643
	pesos_i(24701) := b"0000000000000000_0000000000000000_0010101111111100_0010110001010111"; -- 0.17181660759818163
	pesos_i(24702) := b"0000000000000000_0000000000000000_0000111000011000_1011100111000000"; -- 0.05506478240846768
	pesos_i(24703) := b"0000000000000000_0000000000000000_0001100101011001_1101100111110111"; -- 0.09902727395857175
	pesos_i(24704) := b"1111111111111111_1111111111111111_1101111011010101_0100000011011011"; -- -0.12955851218162523
	pesos_i(24705) := b"1111111111111111_1111111111111111_1111101000000100_1001011111001111"; -- -0.023367416306100352
	pesos_i(24706) := b"0000000000000000_0000000000000000_0001000011100000_1101010001111111"; -- 0.0659306344007607
	pesos_i(24707) := b"0000000000000000_0000000000000000_0000011111110100_0000100011111001"; -- 0.031067429389672097
	pesos_i(24708) := b"1111111111111111_1111111111111111_1100110101101010_1000001000100101"; -- -0.19759356104488557
	pesos_i(24709) := b"0000000000000000_0000000000000000_0001100101001111_0011000110000010"; -- 0.09886464529565857
	pesos_i(24710) := b"0000000000000000_0000000000000000_0001110111000011_1110011110101111"; -- 0.11627052338668928
	pesos_i(24711) := b"0000000000000000_0000000000000000_0000011011011100_1111101011010110"; -- 0.026809384606740257
	pesos_i(24712) := b"1111111111111111_1111111111111111_1110110100110110_1110110001001001"; -- -0.07338069162336987
	pesos_i(24713) := b"0000000000000000_0000000000000000_0000100000001111_1000100011001111"; -- 0.0314870363155251
	pesos_i(24714) := b"0000000000000000_0000000000000000_0001100011000001_1000011111111110"; -- 0.09670305208844387
	pesos_i(24715) := b"0000000000000000_0000000000000000_0010011011010001_1101110101011000"; -- 0.15163977994505728
	pesos_i(24716) := b"0000000000000000_0000000000000000_0001110110010000_1011011101101011"; -- 0.11548944818134034
	pesos_i(24717) := b"1111111111111111_1111111111111111_1110001001100100_1101110100101110"; -- -0.11564843782109609
	pesos_i(24718) := b"1111111111111111_1111111111111111_1110011000100001_0111110101000011"; -- -0.10105149382143022
	pesos_i(24719) := b"1111111111111111_1111111111111111_1101001110110101_1110110010100101"; -- -0.17300530396602296
	pesos_i(24720) := b"1111111111111111_1111111111111111_1111111011010001_0000000001110100"; -- -0.004623385980898866
	pesos_i(24721) := b"0000000000000000_0000000000000000_0010100000001111_1011101000101011"; -- 0.15648997827537375
	pesos_i(24722) := b"0000000000000000_0000000000000000_0000001011100110_0110101100010001"; -- 0.01132840305346924
	pesos_i(24723) := b"0000000000000000_0000000000000000_0010011111101101_0101011011001001"; -- 0.15596525577287396
	pesos_i(24724) := b"1111111111111111_1111111111111111_1101101011111110_1100000001000111"; -- -0.14455030688744508
	pesos_i(24725) := b"0000000000000000_0000000000000000_0010011101111010_1011000100110111"; -- 0.15421588503918426
	pesos_i(24726) := b"1111111111111111_1111111111111111_1101001100100100_1110011000001111"; -- -0.1752182209966382
	pesos_i(24727) := b"0000000000000000_0000000000000000_0010000010111011_0100010001111100"; -- 0.1278574754770879
	pesos_i(24728) := b"1111111111111111_1111111111111111_1111100011001011_0001000000011001"; -- -0.02815150641168281
	pesos_i(24729) := b"0000000000000000_0000000000000000_0010011100000110_1010100011010101"; -- 0.15244536601251038
	pesos_i(24730) := b"1111111111111111_1111111111111111_1110000011011111_1100111000000101"; -- -0.12158501027667555
	pesos_i(24731) := b"1111111111111111_1111111111111111_1111100100000011_0010010011001101"; -- -0.027295780202935684
	pesos_i(24732) := b"0000000000000000_0000000000000000_0001111111001101_1100110100001001"; -- 0.12423402289361994
	pesos_i(24733) := b"0000000000000000_0000000000000000_0001000011000100_0100011000110101"; -- 0.06549490725412413
	pesos_i(24734) := b"0000000000000000_0000000000000000_0001101101110111_0110100100100110"; -- 0.10729081333237403
	pesos_i(24735) := b"1111111111111111_1111111111111111_1110010000101110_1000001001011101"; -- -0.1086653253976541
	pesos_i(24736) := b"0000000000000000_0000000000000000_0001110010100001_0010100011000000"; -- 0.11183409404133192
	pesos_i(24737) := b"1111111111111111_1111111111111111_1111010100100110_0010101001111110"; -- -0.04238638333963363
	pesos_i(24738) := b"0000000000000000_0000000000000000_0001011001100001_0111110001100111"; -- 0.08742501759230678
	pesos_i(24739) := b"1111111111111111_1111111111111111_1101001001010110_1111011011001111"; -- -0.17836053308679345
	pesos_i(24740) := b"1111111111111111_1111111111111111_1110111111111000_1000010000101010"; -- -0.06261419277218035
	pesos_i(24741) := b"1111111111111111_1111111111111111_1101110100010001_1011000100000000"; -- -0.13644880053108716
	pesos_i(24742) := b"0000000000000000_0000000000000000_0000101000111010_1011110100011101"; -- 0.03995878173757149
	pesos_i(24743) := b"1111111111111111_1111111111111111_1110010110101111_0010001100110000"; -- -0.10279636459947225
	pesos_i(24744) := b"1111111111111111_1111111111111111_1111010010101110_0110011111010001"; -- -0.04421378281033652
	pesos_i(24745) := b"0000000000000000_0000000000000000_0000000000111110_1100101001101100"; -- 0.0009581101832645058
	pesos_i(24746) := b"1111111111111111_1111111111111111_1111010111000111_1001110100001011"; -- -0.039922890374038275
	pesos_i(24747) := b"1111111111111111_1111111111111111_1110101001101010_0000101101010010"; -- -0.08431939358325509
	pesos_i(24748) := b"1111111111111111_1111111111111111_1110100110100111_0110001110101011"; -- -0.08728959152762053
	pesos_i(24749) := b"1111111111111111_1111111111111111_1110010001101011_1010010011010101"; -- -0.10773248477813357
	pesos_i(24750) := b"0000000000000000_0000000000000000_0000000111001011_1101001100000001"; -- 0.007016361009073265
	pesos_i(24751) := b"0000000000000000_0000000000000000_0010111011011100_0001001010100011"; -- 0.18304554439663687
	pesos_i(24752) := b"1111111111111111_1111111111111111_1101110001011010_0011011100000011"; -- -0.13924843011215549
	pesos_i(24753) := b"1111111111111111_1111111111111111_1111010110100110_0010101111101100"; -- -0.040433172962951326
	pesos_i(24754) := b"0000000000000000_0000000000000000_0010010000010111_0011110010101000"; -- 0.14097956765816338
	pesos_i(24755) := b"0000000000000000_0000000000000000_0001111100010110_0011000000001001"; -- 0.12143230646262583
	pesos_i(24756) := b"1111111111111111_1111111111111111_1101011011101001_0001111010111110"; -- -0.16050536971762985
	pesos_i(24757) := b"0000000000000000_0000000000000000_0011000001010011_0100111110111001"; -- 0.18877123138818425
	pesos_i(24758) := b"1111111111111111_1111111111111111_1110001110001001_1010001101011010"; -- -0.1111810593860698
	pesos_i(24759) := b"0000000000000000_0000000000000000_0011001000001010_1111000101001011"; -- 0.195479470180645
	pesos_i(24760) := b"1111111111111111_1111111111111111_1110000010111111_0101000100001011"; -- -0.12208074074688155
	pesos_i(24761) := b"1111111111111111_1111111111111111_1110010000101000_1101010001111011"; -- -0.10875198357734223
	pesos_i(24762) := b"0000000000000000_0000000000000000_0001010001111010_0100101000100010"; -- 0.07999099097708068
	pesos_i(24763) := b"1111111111111111_1111111111111111_1110011000111010_0010000011111000"; -- -0.10067552508168812
	pesos_i(24764) := b"0000000000000000_0000000000000000_0010100010110010_0111110111001100"; -- 0.15897356243264002
	pesos_i(24765) := b"1111111111111111_1111111111111111_1110110101101010_0000101110000000"; -- -0.07260063284689638
	pesos_i(24766) := b"0000000000000000_0000000000000000_0011001100110011_1000100000101000"; -- 0.2000050638923753
	pesos_i(24767) := b"0000000000000000_0000000000000000_0010011010100000_1000101100011110"; -- 0.1508871982636528
	pesos_i(24768) := b"0000000000000000_0000000000000000_0010011011011000_1001101001101101"; -- 0.1517426030377624
	pesos_i(24769) := b"1111111111111111_1111111111111111_1101011110001000_0001101110110001"; -- -0.15807940413480193
	pesos_i(24770) := b"0000000000000000_0000000000000000_0000101111010001_1010011110110111"; -- 0.04616783340626886
	pesos_i(24771) := b"1111111111111111_1111111111111111_1100111100000001_1010000010000100"; -- -0.19138142376891545
	pesos_i(24772) := b"1111111111111111_1111111111111111_1111111110110000_1111111010111110"; -- -0.0012055192006755876
	pesos_i(24773) := b"1111111111111111_1111111111111111_1110010010100001_0011111001000001"; -- -0.10691462439920832
	pesos_i(24774) := b"1111111111111111_1111111111111111_1111000001011100_0011001000011001"; -- -0.06109320524248864
	pesos_i(24775) := b"1111111111111111_1111111111111111_1110010011110011_0111101010000111"; -- -0.105659810952172
	pesos_i(24776) := b"1111111111111111_1111111111111111_1110100011110011_0111010101111111"; -- -0.090035111026197
	pesos_i(24777) := b"1111111111111111_1111111111111111_1101000110000110_0000011111110110"; -- -0.18154859767828566
	pesos_i(24778) := b"0000000000000000_0000000000000000_0001100011011101_1011010001000010"; -- 0.09713293648838613
	pesos_i(24779) := b"1111111111111111_1111111111111111_1111001010011100_0111100011010000"; -- -0.05229992782818941
	pesos_i(24780) := b"1111111111111111_1111111111111111_1110100110010110_1011000000010110"; -- -0.08754443617949183
	pesos_i(24781) := b"0000000000000000_0000000000000000_0001001001101110_0000100000011010"; -- 0.07199144970743264
	pesos_i(24782) := b"0000000000000000_0000000000000000_0000101110001111_0111110000100101"; -- 0.04515815639510397
	pesos_i(24783) := b"1111111111111111_1111111111111111_1111001000111010_1011011001101001"; -- -0.05379161771068734
	pesos_i(24784) := b"1111111111111111_1111111111111111_1101011101011001_1110101010010011"; -- -0.15878423612534376
	pesos_i(24785) := b"0000000000000000_0000000000000000_0011000011001111_1101000010010011"; -- 0.1906710012939798
	pesos_i(24786) := b"1111111111111111_1111111111111111_1110110000110101_0110111111110111"; -- -0.0773096104571284
	pesos_i(24787) := b"1111111111111111_1111111111111111_1101010110010010_1111001001101011"; -- -0.16572651745687153
	pesos_i(24788) := b"1111111111111111_1111111111111111_1110101101011010_1111111101110110"; -- -0.08064273221539343
	pesos_i(24789) := b"1111111111111111_1111111111111111_1101100111000011_0011010001110001"; -- -0.14936516030546762
	pesos_i(24790) := b"1111111111111111_1111111111111111_1110001100010110_1011001110100101"; -- -0.1129348490328763
	pesos_i(24791) := b"0000000000000000_0000000000000000_0010001011101100_0011001101101111"; -- 0.13641663990172634
	pesos_i(24792) := b"0000000000000000_0000000000000000_0000000101000011_0110010010111111"; -- 0.004934593846798386
	pesos_i(24793) := b"0000000000000000_0000000000000000_0001101100010110_1001001011110000"; -- 0.10581320147162236
	pesos_i(24794) := b"1111111111111111_1111111111111111_1111110101100010_1111111011111001"; -- -0.01020819113248489
	pesos_i(24795) := b"0000000000000000_0000000000000000_0001000000001111_0100000011100110"; -- 0.06273275001052568
	pesos_i(24796) := b"0000000000000000_0000000000000000_0010101110011101_1001011111011111"; -- 0.1703734320722508
	pesos_i(24797) := b"0000000000000000_0000000000000000_0001111001000101_1101001001010110"; -- 0.11825289338566086
	pesos_i(24798) := b"1111111111111111_1111111111111111_1101111011001001_0010111110110111"; -- -0.12974263936212585
	pesos_i(24799) := b"0000000000000000_0000000000000000_0000000000110111_0000110101010100"; -- 0.0008400278054419936
	pesos_i(24800) := b"0000000000000000_0000000000000000_0000010010000001_1101001010100110"; -- 0.01760593945889634
	pesos_i(24801) := b"0000000000000000_0000000000000000_0000101101011000_0000110011111011"; -- 0.04431229722417098
	pesos_i(24802) := b"0000000000000000_0000000000000000_0001001001000101_1010010100100001"; -- 0.0713751988283605
	pesos_i(24803) := b"1111111111111111_1111111111111111_1111010000000111_0000111111111001"; -- -0.046767236443272985
	pesos_i(24804) := b"1111111111111111_1111111111111111_1101000100001011_1011001110001000"; -- -0.1834152024961556
	pesos_i(24805) := b"0000000000000000_0000000000000000_0000100111001100_0011011011001111"; -- 0.03827230989695185
	pesos_i(24806) := b"1111111111111111_1111111111111111_1111011001110100_0100011110111000"; -- -0.037288205597253626
	pesos_i(24807) := b"0000000000000000_0000000000000000_0010000000010011_0011011110111010"; -- 0.12529323844526846
	pesos_i(24808) := b"1111111111111111_1111111111111111_1101101011101100_1110110110110010"; -- -0.1448222579804493
	pesos_i(24809) := b"1111111111111111_1111111111111111_1110001001000110_1010010111000011"; -- -0.11610950455351979
	pesos_i(24810) := b"0000000000000000_0000000000000000_0010011101101110_0101101110100111"; -- 0.15402767968431966
	pesos_i(24811) := b"1111111111111111_1111111111111111_1111010000001110_0010010101010011"; -- -0.04665915231442874
	pesos_i(24812) := b"1111111111111111_1111111111111111_1101000111100001_1011001101111111"; -- -0.1801498236742947
	pesos_i(24813) := b"1111111111111111_1111111111111111_1101111101000100_0101010101111101"; -- -0.1278635569337768
	pesos_i(24814) := b"1111111111111111_1111111111111111_1111010100111010_0110100111011010"; -- -0.04207743089062973
	pesos_i(24815) := b"0000000000000000_0000000000000000_0011010011100010_1001111001100011"; -- 0.20658292684329957
	pesos_i(24816) := b"1111111111111111_1111111111111111_1111010100110100_1010010001100011"; -- -0.042165494705851916
	pesos_i(24817) := b"0000000000000000_0000000000000000_0001000100001111_0001001010100110"; -- 0.06663624331830056
	pesos_i(24818) := b"1111111111111111_1111111111111111_1100101010000011_1111100010101100"; -- -0.2089237765598539
	pesos_i(24819) := b"0000000000000000_0000000000000000_0011000100001000_1010001010100111"; -- 0.19153801526369257
	pesos_i(24820) := b"0000000000000000_0000000000000000_0010000101110000_1010001110101000"; -- 0.13062498905879577
	pesos_i(24821) := b"0000000000000000_0000000000000000_0000111100101001_1110010000111110"; -- 0.059232964712108066
	pesos_i(24822) := b"0000000000000000_0000000000000000_0010100111100001_0111111000101011"; -- 0.163596997745214
	pesos_i(24823) := b"0000000000000000_0000000000000000_0001111111100000_1100000011111110"; -- 0.12452322201352989
	pesos_i(24824) := b"0000000000000000_0000000000000000_0000011100010010_1100111111001110"; -- 0.027630794413243148
	pesos_i(24825) := b"0000000000000000_0000000000000000_0001100000001001_0100110100000000"; -- 0.09389191857328062
	pesos_i(24826) := b"1111111111111111_1111111111111111_1101101011011011_1000000010000111"; -- -0.14508816444274408
	pesos_i(24827) := b"0000000000000000_0000000000000000_0001010101111010_0100011100101001"; -- 0.08389706379211677
	pesos_i(24828) := b"1111111111111111_1111111111111111_1101101111011001_1100111010101001"; -- -0.1412077748272578
	pesos_i(24829) := b"0000000000000000_0000000000000000_0000111101010001_1011111111100001"; -- 0.05984114888130568
	pesos_i(24830) := b"0000000000000000_0000000000000000_0010010011010010_0111101101110100"; -- 0.14383670418378902
	pesos_i(24831) := b"1111111111111111_1111111111111111_1101000111001011_1011001100111110"; -- -0.18048553211474602
	pesos_i(24832) := b"1111111111111111_1111111111111111_1100101100110000_0011111110010110"; -- -0.20629503811925085
	pesos_i(24833) := b"0000000000000000_0000000000000000_0011001001100110_1010100010011101"; -- 0.19687894661883454
	pesos_i(24834) := b"1111111111111111_1111111111111111_1101101101111110_1110011000010100"; -- -0.14259492888723038
	pesos_i(24835) := b"1111111111111111_1111111111111111_1110100000011001_1001100011111001"; -- -0.09335941233092954
	pesos_i(24836) := b"1111111111111111_1111111111111111_1100101110100011_0111110111100001"; -- -0.20453656445306584
	pesos_i(24837) := b"0000000000000000_0000000000000000_0000001110010011_0111110001011110"; -- 0.013969204939404659
	pesos_i(24838) := b"1111111111111111_1111111111111111_1101111000000000_0010010001000001"; -- -0.13281033904896308
	pesos_i(24839) := b"0000000000000000_0000000000000000_0001101000111111_0110111111001110"; -- 0.1025304677011064
	pesos_i(24840) := b"1111111111111111_1111111111111111_1101001010010000_1001010101101111"; -- -0.17748132741386385
	pesos_i(24841) := b"0000000000000000_0000000000000000_0001001101100001_0001100100000110"; -- 0.07570034400478705
	pesos_i(24842) := b"1111111111111111_1111111111111111_1101001101110111_1010111100111000"; -- -0.1739550103470283
	pesos_i(24843) := b"0000000000000000_0000000000000000_0000101001111111_1010011101100110"; -- 0.041010344037917895
	pesos_i(24844) := b"0000000000000000_0000000000000000_0000110001111101_0101011111000101"; -- 0.048787580100600636
	pesos_i(24845) := b"1111111111111111_1111111111111111_1111010111100100_1101001010100111"; -- -0.03947719018235006
	pesos_i(24846) := b"0000000000000000_0000000000000000_0010110101000011_1111110110111111"; -- 0.17681871327018647
	pesos_i(24847) := b"0000000000000000_0000000000000000_0000001100000101_1001011100010110"; -- 0.011804049341692364
	pesos_i(24848) := b"1111111111111111_1111111111111111_1101100001001000_0011110100000111"; -- -0.15514772959631665
	pesos_i(24849) := b"1111111111111111_1111111111111111_1111001110100000_0010010100011100"; -- -0.04833763193178867
	pesos_i(24850) := b"1111111111111111_1111111111111111_1110110010100001_1101111110000011"; -- -0.07565501254085868
	pesos_i(24851) := b"0000000000000000_0000000000000000_0010101010010111_0101111010101101"; -- 0.16637222025944395
	pesos_i(24852) := b"0000000000000000_0000000000000000_0001011000101110_0100001110001010"; -- 0.08664342984156138
	pesos_i(24853) := b"1111111111111111_1111111111111111_1101100011011010_1101111000111110"; -- -0.1529103373885751
	pesos_i(24854) := b"1111111111111111_1111111111111111_1111111001101011_1100000011001111"; -- -0.006168317224244917
	pesos_i(24855) := b"0000000000000000_0000000000000000_0010011001001101_0101011111001000"; -- 0.149617658813014
	pesos_i(24856) := b"0000000000000000_0000000000000000_0010110101100000_1011000110101101"; -- 0.17725668405060863
	pesos_i(24857) := b"1111111111111111_1111111111111111_1110101001011011_1100100111000000"; -- -0.08453692493455217
	pesos_i(24858) := b"1111111111111111_1111111111111111_1110100011111100_0111011000011000"; -- -0.08989774624711055
	pesos_i(24859) := b"0000000000000000_0000000000000000_0011001111100100_0001111000010000"; -- 0.20269954582387126
	pesos_i(24860) := b"0000000000000000_0000000000000000_0010010011110001_0010010111001111"; -- 0.14430462163624233
	pesos_i(24861) := b"0000000000000000_0000000000000000_0011001010111010_0100100011101011"; -- 0.19815498105902077
	pesos_i(24862) := b"1111111111111111_1111111111111111_1111000001010001_1111111111101110"; -- -0.0612487834060512
	pesos_i(24863) := b"1111111111111111_1111111111111111_1111110011001100_0000011000010000"; -- -0.012511845776254076
	pesos_i(24864) := b"1111111111111111_1111111111111111_1110001011100101_0111101000000100"; -- -0.1136859646855034
	pesos_i(24865) := b"0000000000000000_0000000000000000_0000011100111001_1101000111111000"; -- 0.028226016051021645
	pesos_i(24866) := b"1111111111111111_1111111111111111_1100111010100011_0100001001111001"; -- -0.19282135538336276
	pesos_i(24867) := b"0000000000000000_0000000000000000_0000101111110110_0001000101110100"; -- 0.04672345243203657
	pesos_i(24868) := b"1111111111111111_1111111111111111_1101101110110101_1110111011101101"; -- -0.14175516797786597
	pesos_i(24869) := b"0000000000000000_0000000000000000_0011010100001011_0011100011111010"; -- 0.2072024927391009
	pesos_i(24870) := b"0000000000000000_0000000000000000_0001101100101101_1100001100011000"; -- 0.10616702389973068
	pesos_i(24871) := b"1111111111111111_1111111111111111_1100110110001010_0100000100100111"; -- -0.19710915365032694
	pesos_i(24872) := b"1111111111111111_1111111111111111_1111100010010000_0110100100011010"; -- -0.029046469876833698
	pesos_i(24873) := b"1111111111111111_1111111111111111_1101100001010111_1011101011011011"; -- -0.15491134781823174
	pesos_i(24874) := b"1111111111111111_1111111111111111_1101101110100010_1110010110111010"; -- -0.14204563349213228
	pesos_i(24875) := b"1111111111111111_1111111111111111_1101000000010000_1010101111010100"; -- -0.18724561755233327
	pesos_i(24876) := b"0000000000000000_0000000000000000_0010011011010001_1111001110100111"; -- 0.15164110973488953
	pesos_i(24877) := b"0000000000000000_0000000000000000_0000100011100011_0111011111000011"; -- 0.0347208834079444
	pesos_i(24878) := b"0000000000000000_0000000000000000_0001000101011100_0000010111100111"; -- 0.06781041039178987
	pesos_i(24879) := b"0000000000000000_0000000000000000_0000011011101001_0001101101110101"; -- 0.026994434424654597
	pesos_i(24880) := b"1111111111111111_1111111111111111_1110001010001110_1011000000001100"; -- -0.11501025871673433
	pesos_i(24881) := b"1111111111111111_1111111111111111_1111111011000011_1100111011010010"; -- -0.004824708723306592
	pesos_i(24882) := b"1111111111111111_1111111111111111_1110101110110001_1011010001011110"; -- -0.07931969350657353
	pesos_i(24883) := b"1111111111111111_1111111111111111_1111100100010010_0100100100010000"; -- -0.027064737013848865
	pesos_i(24884) := b"0000000000000000_0000000000000000_0001000010010101_1011001010011010"; -- 0.06478420498059242
	pesos_i(24885) := b"0000000000000000_0000000000000000_0001110101110001_0101111111001111"; -- 0.11501120388743993
	pesos_i(24886) := b"0000000000000000_0000000000000000_0000010110110011_1110110111011010"; -- 0.02227675035651339
	pesos_i(24887) := b"0000000000000000_0000000000000000_0010001110111100_0111011111011100"; -- 0.1395945465713414
	pesos_i(24888) := b"1111111111111111_1111111111111111_1111101011101000_0100000000001001"; -- -0.01989364408619878
	pesos_i(24889) := b"1111111111111111_1111111111111111_1100110001101111_1101010010010010"; -- -0.20141860412014395
	pesos_i(24890) := b"0000000000000000_0000000000000000_0000011101010000_0100110100000110"; -- 0.028569044007904474
	pesos_i(24891) := b"1111111111111111_1111111111111111_1111101100001010_0011010011101001"; -- -0.019375508342416376
	pesos_i(24892) := b"1111111111111111_1111111111111111_1110110111011010_0011101010011101"; -- -0.0708888404359153
	pesos_i(24893) := b"1111111111111111_1111111111111111_1101001100111001_1011011101000111"; -- -0.1749005748779839
	pesos_i(24894) := b"0000000000000000_0000000000000000_0011000110100111_0010110110010101"; -- 0.19395718456115782
	pesos_i(24895) := b"0000000000000000_0000000000000000_0000011111011101_1010001011101100"; -- 0.03072565328582453
	pesos_i(24896) := b"0000000000000000_0000000000000000_0010111011100100_0111001011111000"; -- 0.18317335667952903
	pesos_i(24897) := b"1111111111111111_1111111111111111_1110000111000010_0010101011101010"; -- -0.1181309871029654
	pesos_i(24898) := b"0000000000000000_0000000000000000_0010000010110000_1101110110100110"; -- 0.1276987581201976
	pesos_i(24899) := b"1111111111111111_1111111111111111_1111000011110010_0001001101101111"; -- -0.058806214809936
	pesos_i(24900) := b"1111111111111111_1111111111111111_1110101011011111_1111100101000100"; -- -0.08251993265134379
	pesos_i(24901) := b"1111111111111111_1111111111111111_1111111011110010_0101001111011010"; -- -0.004114874991807601
	pesos_i(24902) := b"0000000000000000_0000000000000000_0011000101010001_1010011101001001"; -- 0.19265218299117884
	pesos_i(24903) := b"1111111111111111_1111111111111111_1111101111110001_1010011011110111"; -- -0.0158439299767446
	pesos_i(24904) := b"1111111111111111_1111111111111111_1100111010111100_1010000000011001"; -- -0.19243430518503388
	pesos_i(24905) := b"0000000000000000_0000000000000000_0000100001111111_1100111011100000"; -- 0.03320019698741933
	pesos_i(24906) := b"1111111111111111_1111111111111111_1101000011100010_1100010001101011"; -- -0.18403980615653723
	pesos_i(24907) := b"1111111111111111_1111111111111111_1110100011100001_1101100010001011"; -- -0.0903038654444497
	pesos_i(24908) := b"0000000000000000_0000000000000000_0000000001110100_1100001101001001"; -- 0.001781659523730801
	pesos_i(24909) := b"0000000000000000_0000000000000000_0010000000011100_1100000001001111"; -- 0.1254387086635709
	pesos_i(24910) := b"0000000000000000_0000000000000000_0010000001101000_1001110100100110"; -- 0.12659628083798175
	pesos_i(24911) := b"1111111111111111_1111111111111111_1101110001110101_1110000000001110"; -- -0.13882636705461532
	pesos_i(24912) := b"1111111111111111_1111111111111111_1110000001101000_1100110110111111"; -- -0.12340082261143459
	pesos_i(24913) := b"0000000000000000_0000000000000000_0010111011011100_1011101111000000"; -- 0.18305562431534644
	pesos_i(24914) := b"1111111111111111_1111111111111111_1111011010000111_0100011100010011"; -- -0.036998327185153515
	pesos_i(24915) := b"1111111111111111_1111111111111111_1101010000101111_1000010111011010"; -- -0.17114985867774243
	pesos_i(24916) := b"1111111111111111_1111111111111111_1100111010110111_0100010011011111"; -- -0.19251603662405534
	pesos_i(24917) := b"0000000000000000_0000000000000000_0001111110100010_0000000101110110"; -- 0.12356576079581073
	pesos_i(24918) := b"0000000000000000_0000000000000000_0010100000110001_0010010011101000"; -- 0.15699988043518992
	pesos_i(24919) := b"1111111111111111_1111111111111111_1111010100000001_0010001100111110"; -- -0.04295139069206534
	pesos_i(24920) := b"0000000000000000_0000000000000000_0000001011010011_1101101101000000"; -- 0.01104517276418386
	pesos_i(24921) := b"0000000000000000_0000000000000000_0010000000001100_1001101100111110"; -- 0.12519235857858288
	pesos_i(24922) := b"1111111111111111_1111111111111111_1101100111011001_0101010110010001"; -- -0.14902749257478212
	pesos_i(24923) := b"0000000000000000_0000000000000000_0001101111000000_1111010011011000"; -- 0.10841303135999077
	pesos_i(24924) := b"1111111111111111_1111111111111111_1110101010101001_1011011000010010"; -- -0.08334791248209843
	pesos_i(24925) := b"1111111111111111_1111111111111111_1100111110110001_0110011010001011"; -- -0.188699332303437
	pesos_i(24926) := b"0000000000000000_0000000000000000_0010000011000111_0010110100100100"; -- 0.12803918957635302
	pesos_i(24927) := b"1111111111111111_1111111111111111_1110111110010010_0101001100100101"; -- -0.06417351103705121
	pesos_i(24928) := b"1111111111111111_1111111111111111_1101000010000100_1100000010100100"; -- -0.18547435752588945
	pesos_i(24929) := b"0000000000000000_0000000000000000_0011001010111110_1000100101010110"; -- 0.19821985577597276
	pesos_i(24930) := b"1111111111111111_1111111111111111_1111001011101110_0000011101111110"; -- -0.05105546166059873
	pesos_i(24931) := b"0000000000000000_0000000000000000_0010111001110001_1010101100011111"; -- 0.18142194287125082
	pesos_i(24932) := b"1111111111111111_1111111111111111_1101010100100111_1010011010001010"; -- -0.16736373075403818
	pesos_i(24933) := b"0000000000000000_0000000000000000_0000010110001000_1001001101001111"; -- 0.02161522568512167
	pesos_i(24934) := b"1111111111111111_1111111111111111_1101000001011011_1010011111011010"; -- -0.18610144542500276
	pesos_i(24935) := b"1111111111111111_1111111111111111_1111101101110001_1001111111111100"; -- -0.017797471036142033
	pesos_i(24936) := b"1111111111111111_1111111111111111_1110110001011000_1001111011011011"; -- -0.07677275800338504
	pesos_i(24937) := b"1111111111111111_1111111111111111_1110011100111000_1010001100001110"; -- -0.0967920389385385
	pesos_i(24938) := b"1111111111111111_1111111111111111_1110010010011110_1011111010010110"; -- -0.1069527515954586
	pesos_i(24939) := b"0000000000000000_0000000000000000_0010100011101000_0110011000111000"; -- 0.15979613176067967
	pesos_i(24940) := b"0000000000000000_0000000000000000_0010100100000100_0100100010001101"; -- 0.16022160952725706
	pesos_i(24941) := b"1111111111111111_1111111111111111_1111110100111110_1100100111100010"; -- -0.010760671885797272
	pesos_i(24942) := b"1111111111111111_1111111111111111_1101000111001001_0000110100000101"; -- -0.18052595744834313
	pesos_i(24943) := b"0000000000000000_0000000000000000_0000000000110010_0101000011001011"; -- 0.0007677551387041697
	pesos_i(24944) := b"1111111111111111_1111111111111111_1110000010001110_0101111010011010"; -- -0.12282761322868871
	pesos_i(24945) := b"1111111111111111_1111111111111111_1101000111101101_1101011111011111"; -- -0.17996455010109372
	pesos_i(24946) := b"1111111111111111_1111111111111111_1111010010010111_1100111000110111"; -- -0.04455863138926859
	pesos_i(24947) := b"0000000000000000_0000000000000000_0000111100001101_0010010001101010"; -- 0.05879428473680362
	pesos_i(24948) := b"0000000000000000_0000000000000000_0010011100000010_0100011101010001"; -- 0.15237851832849497
	pesos_i(24949) := b"1111111111111111_1111111111111111_1110111011100001_1011111101101100"; -- -0.0668678627523189
	pesos_i(24950) := b"0000000000000000_0000000000000000_0000010111100010_1011011000100011"; -- 0.022990592432318747
	pesos_i(24951) := b"0000000000000000_0000000000000000_0000110111101000_1011101101001111"; -- 0.05433245349307815
	pesos_i(24952) := b"0000000000000000_0000000000000000_0001000110110100_0000001100111001"; -- 0.06915302422987833
	pesos_i(24953) := b"1111111111111111_1111111111111111_1111000101010011_1111111111110110"; -- -0.057312014076708426
	pesos_i(24954) := b"1111111111111111_1111111111111111_1100110111011010_1111011101111011"; -- -0.19587758289489257
	pesos_i(24955) := b"0000000000000000_0000000000000000_0001101001111011_1010000011010110"; -- 0.10344891769985665
	pesos_i(24956) := b"0000000000000000_0000000000000000_0010110001100001_1010010101000000"; -- 0.17336495216689013
	pesos_i(24957) := b"0000000000000000_0000000000000000_0010000001010110_0110010010001011"; -- 0.12631824873445172
	pesos_i(24958) := b"0000000000000000_0000000000000000_0000010000001110_1110000011100000"; -- 0.01585202665151633
	pesos_i(24959) := b"0000000000000000_0000000000000000_0000100100011111_1001000111101100"; -- 0.035637969974171055
	pesos_i(24960) := b"1111111111111111_1111111111111111_1111010001010000_0011010000111100"; -- -0.04565118352645403
	pesos_i(24961) := b"1111111111111111_1111111111111111_1101010000111010_0100010000111100"; -- -0.17098592310989819
	pesos_i(24962) := b"0000000000000000_0000000000000000_0001110011010001_1110001001110000"; -- 0.11257758353270789
	pesos_i(24963) := b"1111111111111111_1111111111111111_1101010010000110_1101000011010011"; -- -0.16981787532518194
	pesos_i(24964) := b"1111111111111111_1111111111111111_1110101011110001_1100011101100100"; -- -0.08224824724235887
	pesos_i(24965) := b"0000000000000000_0000000000000000_0011010010110011_1001110000100100"; -- 0.2058656299011747
	pesos_i(24966) := b"0000000000000000_0000000000000000_0001010101000110_0101101111111001"; -- 0.08310484722918442
	pesos_i(24967) := b"1111111111111111_1111111111111111_1110000000100110_0111011110010010"; -- -0.1244130390640372
	pesos_i(24968) := b"0000000000000000_0000000000000000_0011000110010010_0111110110110110"; -- 0.19364152624414768
	pesos_i(24969) := b"1111111111111111_1111111111111111_1100110101000100_1111001001001001"; -- -0.19816671112236242
	pesos_i(24970) := b"1111111111111111_1111111111111111_1101110111000010_0100111101110110"; -- -0.1337538087731816
	pesos_i(24971) := b"1111111111111111_1111111111111111_1110000110110001_1001110111001010"; -- -0.11838353934548561
	pesos_i(24972) := b"1111111111111111_1111111111111111_1110101110110011_0101100111110001"; -- -0.07929456593656073
	pesos_i(24973) := b"0000000000000000_0000000000000000_0010110100001010_1011000101100010"; -- 0.17594441077658218
	pesos_i(24974) := b"0000000000000000_0000000000000000_0001001110110001_0101001110101110"; -- 0.07692454332285134
	pesos_i(24975) := b"1111111111111111_1111111111111111_1110100111000000_0110110100111100"; -- -0.08690755156789168
	pesos_i(24976) := b"0000000000000000_0000000000000000_0001100101001100_0001110011001010"; -- 0.09881763388531654
	pesos_i(24977) := b"1111111111111111_1111111111111111_1101111100101000_1111100011000100"; -- -0.12828107088789778
	pesos_i(24978) := b"0000000000000000_0000000000000000_0010000011101011_0000010101010001"; -- 0.12858613236617802
	pesos_i(24979) := b"0000000000000000_0000000000000000_0010010010111100_0010001100100100"; -- 0.14349574699345866
	pesos_i(24980) := b"0000000000000000_0000000000000000_0000000000101101_0100001100110110"; -- 0.0006906516955802831
	pesos_i(24981) := b"0000000000000000_0000000000000000_0000111100110011_0110000100000000"; -- 0.05937772988878626
	pesos_i(24982) := b"1111111111111111_1111111111111111_1101001010001101_1101000111010010"; -- -0.17752350438574785
	pesos_i(24983) := b"0000000000000000_0000000000000000_0010101111101010_0110111101111010"; -- 0.17154595121289182
	pesos_i(24984) := b"0000000000000000_0000000000000000_0000001110000011_0001100010101011"; -- 0.013719121738176137
	pesos_i(24985) := b"1111111111111111_1111111111111111_1110100001111010_1000100101100001"; -- -0.09188023923767717
	pesos_i(24986) := b"0000000000000000_0000000000000000_0001001100001101_1001110100000010"; -- 0.07442647267430125
	pesos_i(24987) := b"0000000000000000_0000000000000000_0001000101011101_0111101010110010"; -- 0.06783263067040946
	pesos_i(24988) := b"1111111111111111_1111111111111111_1110000010011110_1001000001100111"; -- -0.12258050421331883
	pesos_i(24989) := b"0000000000000000_0000000000000000_0001010011100011_0101101100101011"; -- 0.08159417912226198
	pesos_i(24990) := b"1111111111111111_1111111111111111_1101111110001011_0011101101101110"; -- -0.12678173601267487
	pesos_i(24991) := b"1111111111111111_1111111111111111_1101100001101011_1001011001011110"; -- -0.15460834688061556
	pesos_i(24992) := b"0000000000000000_0000000000000000_0001001011101000_1011101000010111"; -- 0.07386363076905476
	pesos_i(24993) := b"1111111111111111_1111111111111111_1111010011000010_1101110110001101"; -- -0.043901589356670975
	pesos_i(24994) := b"1111111111111111_1111111111111111_1111110010011010_1110101100110101"; -- -0.01326112696198924
	pesos_i(24995) := b"0000000000000000_0000000000000000_0000111100101111_0001001000011110"; -- 0.0593119929493521
	pesos_i(24996) := b"1111111111111111_1111111111111111_1111111110010000_1000100011010101"; -- -0.0017008286168583406
	pesos_i(24997) := b"0000000000000000_0000000000000000_0001110010110001_0111111111110111"; -- 0.11208343295228627
	pesos_i(24998) := b"1111111111111111_1111111111111111_1111001001001001_0011000100110110"; -- -0.05357067521190499
	pesos_i(24999) := b"1111111111111111_1111111111111111_1101000111101000_1101001011101111"; -- -0.18004113831605606
	pesos_i(25000) := b"1111111111111111_1111111111111111_1111000100100100_0101000000010111"; -- -0.058039659760426486
	pesos_i(25001) := b"0000000000000000_0000000000000000_0001110100100100_0000001101101101"; -- 0.11383077069724738
	pesos_i(25002) := b"1111111111111111_1111111111111111_1110000000000011_0110110100001101"; -- -0.12494772367461887
	pesos_i(25003) := b"0000000000000000_0000000000000000_0010000100101001_0001000011111010"; -- 0.1295328721176876
	pesos_i(25004) := b"0000000000000000_0000000000000000_0000110101100001_1000010011000100"; -- 0.05226926600814513
	pesos_i(25005) := b"0000000000000000_0000000000000000_0010001100101011_1000011011110010"; -- 0.1373829214074253
	pesos_i(25006) := b"1111111111111111_1111111111111111_1111111001001010_0111110011100010"; -- -0.006675905957398736
	pesos_i(25007) := b"0000000000000000_0000000000000000_0000000000101011_0000000110110010"; -- 0.0006562290553946712
	pesos_i(25008) := b"0000000000000000_0000000000000000_0010010000101011_1110011111101101"; -- 0.1412949518232783
	pesos_i(25009) := b"0000000000000000_0000000000000000_0001001101011101_1101000110101010"; -- 0.07565031426400556
	pesos_i(25010) := b"0000000000000000_0000000000000000_0010111000000011_0010100010011110"; -- 0.17973569743564435
	pesos_i(25011) := b"1111111111111111_1111111111111111_1101111101000001_0000111100111010"; -- -0.12791352120957708
	pesos_i(25012) := b"1111111111111111_1111111111111111_1101010111101100_0011000111010000"; -- -0.1643647067181294
	pesos_i(25013) := b"1111111111111111_1111111111111111_1110111101111100_1110110111011111"; -- -0.06449998188744219
	pesos_i(25014) := b"0000000000000000_0000000000000000_0000010001101001_0101101011100101"; -- 0.01723259053269093
	pesos_i(25015) := b"1111111111111111_1111111111111111_1110101111000111_0001000010110100"; -- -0.0789937554539874
	pesos_i(25016) := b"0000000000000000_0000000000000000_0000110101010011_0011010011101010"; -- 0.05205088333463675
	pesos_i(25017) := b"0000000000000000_0000000000000000_0001000101101000_0110010111101001"; -- 0.06799923840568332
	pesos_i(25018) := b"0000000000000000_0000000000000000_0001101111110101_1010110001001110"; -- 0.10921742341331853
	pesos_i(25019) := b"0000000000000000_0000000000000000_0000011010110101_0111001100110010"; -- 0.026206207072978844
	pesos_i(25020) := b"1111111111111111_1111111111111111_1101111001101011_1011011011110000"; -- -0.13116890570913597
	pesos_i(25021) := b"0000000000000000_0000000000000000_0000101001011110_0101010000111011"; -- 0.04050184671464011
	pesos_i(25022) := b"0000000000000000_0000000000000000_0010101001001110_0100100100111011"; -- 0.16525705041506314
	pesos_i(25023) := b"0000000000000000_0000000000000000_0001100010101110_1011001100110011"; -- 0.09641571033319059
	pesos_i(25024) := b"0000000000000000_0000000000000000_0010100001110000_0010100011101010"; -- 0.15796142314574482
	pesos_i(25025) := b"0000000000000000_0000000000000000_0000110110010100_1000001001001110"; -- 0.05304731763096368
	pesos_i(25026) := b"0000000000000000_0000000000000000_0001101000010111_0101101111111111"; -- 0.10191893557979194
	pesos_i(25027) := b"0000000000000000_0000000000000000_0001101110001010_0101011010100101"; -- 0.10757962724379143
	pesos_i(25028) := b"1111111111111111_1111111111111111_1110100110111100_1000101101001010"; -- -0.08696679530012406
	pesos_i(25029) := b"0000000000000000_0000000000000000_0010011111000010_0100110011110110"; -- 0.15530854232558794
	pesos_i(25030) := b"0000000000000000_0000000000000000_0000011000010000_1111000000111111"; -- 0.023695960468297906
	pesos_i(25031) := b"0000000000000000_0000000000000000_0000010001001110_1100111111010010"; -- 0.016827572542510893
	pesos_i(25032) := b"1111111111111111_1111111111111111_1111001110101100_1100010111010111"; -- -0.04814494600770879
	pesos_i(25033) := b"0000000000000000_0000000000000000_0001000111111011_0110101001000110"; -- 0.07024254051212586
	pesos_i(25034) := b"1111111111111111_1111111111111111_1110101110011100_1000011110000100"; -- -0.07964280151399002
	pesos_i(25035) := b"0000000000000000_0000000000000000_0010001111010011_0111001010101000"; -- 0.13994518852555768
	pesos_i(25036) := b"1111111111111111_1111111111111111_1101111101010001_0111111011011110"; -- -0.1276627261948646
	pesos_i(25037) := b"1111111111111111_1111111111111111_1100110011011001_1101100101110100"; -- -0.19980088156424225
	pesos_i(25038) := b"1111111111111111_1111111111111111_1111010110101100_0010010010111001"; -- -0.0403420494276248
	pesos_i(25039) := b"1111111111111111_1111111111111111_1111110000011111_1100111001001100"; -- -0.015139681360365469
	pesos_i(25040) := b"0000000000000000_0000000000000000_0010010101000011_1000100001110011"; -- 0.14556172193645905
	pesos_i(25041) := b"1111111111111111_1111111111111111_1111100011010101_0000111001110110"; -- -0.0279990159341516
	pesos_i(25042) := b"0000000000000000_0000000000000000_0001010001101101_1101011001010011"; -- 0.07980098272970784
	pesos_i(25043) := b"1111111111111111_1111111111111111_1110101100010000_1010101100001111"; -- -0.08177691358816451
	pesos_i(25044) := b"1111111111111111_1111111111111111_1101011001010011_0010110011110110"; -- -0.16279334055527056
	pesos_i(25045) := b"1111111111111111_1111111111111111_1110000101110110_0111110001101101"; -- -0.11928579660890161
	pesos_i(25046) := b"0000000000000000_0000000000000000_0000001101101001_0100011110010000"; -- 0.013325188391951664
	pesos_i(25047) := b"0000000000000000_0000000000000000_0000111110001110_1011010001001000"; -- 0.060771243580078994
	pesos_i(25048) := b"1111111111111111_1111111111111111_1100111000010111_0111011010100110"; -- -0.19495447593523071
	pesos_i(25049) := b"1111111111111111_1111111111111111_1110101110100011_0111010110010110"; -- -0.07953705862994405
	pesos_i(25050) := b"1111111111111111_1111111111111111_1111001001111101_1001001010111001"; -- -0.052771405950488216
	pesos_i(25051) := b"1111111111111111_1111111111111111_1111011011010101_1000000101001111"; -- -0.0358046706257406
	pesos_i(25052) := b"0000000000000000_0000000000000000_0000111001101010_0111010011100010"; -- 0.056311898356549955
	pesos_i(25053) := b"0000000000000000_0000000000000000_0010111100110101_0001101001010111"; -- 0.18440403586515022
	pesos_i(25054) := b"0000000000000000_0000000000000000_0011001011010101_0000111101111000"; -- 0.19856354418682806
	pesos_i(25055) := b"0000000000000000_0000000000000000_0010001111001111_1011111010100101"; -- 0.13988868273042723
	pesos_i(25056) := b"1111111111111111_1111111111111111_1101010110001110_1101000000110011"; -- -0.16578959229827658
	pesos_i(25057) := b"0000000000000000_0000000000000000_0010101110111000_1011101000111100"; -- 0.17078746770496467
	pesos_i(25058) := b"1111111111111111_1111111111111111_1111000100011110_1101010101101000"; -- -0.05812326621644787
	pesos_i(25059) := b"0000000000000000_0000000000000000_0001001111000011_0011110001001011"; -- 0.07719780766982956
	pesos_i(25060) := b"0000000000000000_0000000000000000_0010011101000010_1011011100110000"; -- 0.15336174889443285
	pesos_i(25061) := b"1111111111111111_1111111111111111_1110000100100000_0000000010111010"; -- -0.12060542540193055
	pesos_i(25062) := b"1111111111111111_1111111111111111_1111001000001001_1111000000001111"; -- -0.05453586235314947
	pesos_i(25063) := b"0000000000000000_0000000000000000_0001100001110100_1101011000011000"; -- 0.09553278047964052
	pesos_i(25064) := b"0000000000000000_0000000000000000_0010011101001100_0011100001110110"; -- 0.15350678323596637
	pesos_i(25065) := b"1111111111111111_1111111111111111_1110110000110011_1011000001111101"; -- -0.07733628221968755
	pesos_i(25066) := b"1111111111111111_1111111111111111_1110111110100010_1110011001010111"; -- -0.06392059686149175
	pesos_i(25067) := b"1111111111111111_1111111111111111_1111010000100010_1000000010001101"; -- -0.04634853906416526
	pesos_i(25068) := b"1111111111111111_1111111111111111_1101011011100011_0101000001101101"; -- -0.1605939610572809
	pesos_i(25069) := b"1111111111111111_1111111111111111_1110110000111010_0001100100101100"; -- -0.07723848981146232
	pesos_i(25070) := b"1111111111111111_1111111111111111_1110101101011000_1011001101011000"; -- -0.0806777867718971
	pesos_i(25071) := b"0000000000000000_0000000000000000_0001100111011010_0110000001000001"; -- 0.10098840323374955
	pesos_i(25072) := b"1111111111111111_1111111111111111_1110001011101001_0010010101110011"; -- -0.11362997002118462
	pesos_i(25073) := b"1111111111111111_1111111111111111_1101000001101001_0100111101111110"; -- -0.18589308895230153
	pesos_i(25074) := b"1111111111111111_1111111111111111_1110000010101110_0001101011111001"; -- -0.12234336302147528
	pesos_i(25075) := b"0000000000000000_0000000000000000_0010110111010010_1000011110110101"; -- 0.17899368446857603
	pesos_i(25076) := b"0000000000000000_0000000000000000_0010000001111101_1101110100111010"; -- 0.12692053486887064
	pesos_i(25077) := b"1111111111111111_1111111111111111_1101101110010100_0000010010111000"; -- -0.14227266797455185
	pesos_i(25078) := b"0000000000000000_0000000000000000_0000110111010011_0001111010111110"; -- 0.05400268688423093
	pesos_i(25079) := b"1111111111111111_1111111111111111_1110011110110111_1110001101101010"; -- -0.09485033661157144
	pesos_i(25080) := b"0000000000000000_0000000000000000_0000110101100110_1111111010101000"; -- 0.05235282527369462
	pesos_i(25081) := b"0000000000000000_0000000000000000_0001100001100011_1001101100110000"; -- 0.09526986999364567
	pesos_i(25082) := b"1111111111111111_1111111111111111_1111100100000111_1001000010110010"; -- -0.02722831385866477
	pesos_i(25083) := b"1111111111111111_1111111111111111_1110011000100000_1010111100001111"; -- -0.10106378443256349
	pesos_i(25084) := b"1111111111111111_1111111111111111_1111011000010100_0111011011000001"; -- -0.03875024595548937
	pesos_i(25085) := b"0000000000000000_0000000000000000_0001001000000110_1010010100011100"; -- 0.07041389409854326
	pesos_i(25086) := b"1111111111111111_1111111111111111_1110010110101101_1101000001011111"; -- -0.10281655950939064
	pesos_i(25087) := b"0000000000000000_0000000000000000_0001101001010100_1010011111110011"; -- 0.10285424884319117
	pesos_i(25088) := b"0000000000000000_0000000000000000_0010000010101111_0011011011010111"; -- 0.1276735569084528
	pesos_i(25089) := b"0000000000000000_0000000000000000_0001101110011011_0100000010111000"; -- 0.10783771989262583
	pesos_i(25090) := b"1111111111111111_1111111111111111_1101110010011011_0110010010100000"; -- -0.1382538898848836
	pesos_i(25091) := b"1111111111111111_1111111111111111_1101100011110100_1001101101011011"; -- -0.1525175955950344
	pesos_i(25092) := b"0000000000000000_0000000000000000_0010010001101110_0011011111111111"; -- 0.14230680431836273
	pesos_i(25093) := b"1111111111111111_1111111111111111_1111010011100100_0011101101010011"; -- -0.04339246016883003
	pesos_i(25094) := b"0000000000000000_0000000000000000_0010011001000110_1001111110110110"; -- 0.14951513466277777
	pesos_i(25095) := b"0000000000000000_0000000000000000_0000010001111100_0111101100110100"; -- 0.017524433345832705
	pesos_i(25096) := b"0000000000000000_0000000000000000_0001110010110110_1100011010111001"; -- 0.11216394448106277
	pesos_i(25097) := b"0000000000000000_0000000000000000_0001101011011110_0001001100111001"; -- 0.10495109694429011
	pesos_i(25098) := b"0000000000000000_0000000000000000_0001101000000010_0110101100110010"; -- 0.1015994069321509
	pesos_i(25099) := b"0000000000000000_0000000000000000_0010110110010011_1100011000100111"; -- 0.17803610287641908
	pesos_i(25100) := b"1111111111111111_1111111111111111_1100111111111001_1010100011101100"; -- -0.1875967429185711
	pesos_i(25101) := b"1111111111111111_1111111111111111_1101010000010101_0000000001100000"; -- -0.17155454315391094
	pesos_i(25102) := b"0000000000000000_0000000000000000_0010001110010101_0100000011010010"; -- 0.1389961731185376
	pesos_i(25103) := b"0000000000000000_0000000000000000_0001100100111110_0110001111001110"; -- 0.09860824381451433
	pesos_i(25104) := b"1111111111111111_1111111111111111_1110111010100100_0010110101100000"; -- -0.0678073539514897
	pesos_i(25105) := b"0000000000000000_0000000000000000_0010011111101011_1100011101010101"; -- 0.15594144644098967
	pesos_i(25106) := b"0000000000000000_0000000000000000_0001000011000010_1100101101000010"; -- 0.06547232017631137
	pesos_i(25107) := b"1111111111111111_1111111111111111_1111000111110111_0100111001001001"; -- -0.054820162940602185
	pesos_i(25108) := b"1111111111111111_1111111111111111_1101010010100000_1111001110110110"; -- -0.16941906737125148
	pesos_i(25109) := b"0000000000000000_0000000000000000_0001000010100111_0110001100100010"; -- 0.06505412652794838
	pesos_i(25110) := b"1111111111111111_1111111111111111_1100110110111010_1000100100101001"; -- -0.19637243993900802
	pesos_i(25111) := b"1111111111111111_1111111111111111_1110110111010000_1100110001011010"; -- -0.07103274162406895
	pesos_i(25112) := b"0000000000000000_0000000000000000_0010000110000100_0101010110000001"; -- 0.13092550667400465
	pesos_i(25113) := b"0000000000000000_0000000000000000_0000010101101111_0111111011110101"; -- 0.02123254280318103
	pesos_i(25114) := b"0000000000000000_0000000000000000_0010111000111100_0110001100001011"; -- 0.1806089307590458
	pesos_i(25115) := b"0000000000000000_0000000000000000_0011001110001000_1101100101111010"; -- 0.2013069079081718
	pesos_i(25116) := b"1111111111111111_1111111111111111_1101000110010111_0100011011000001"; -- -0.18128545548716873
	pesos_i(25117) := b"1111111111111111_1111111111111111_1110000001010111_0011110011111000"; -- -0.12366885122045604
	pesos_i(25118) := b"1111111111111111_1111111111111111_1111001000000100_0011010011101001"; -- -0.054623311167099814
	pesos_i(25119) := b"0000000000000000_0000000000000000_0001001010100111_0010110011000100"; -- 0.07286338605357279
	pesos_i(25120) := b"0000000000000000_0000000000000000_0001010101111110_1000101100000010"; -- 0.08396214294202564
	pesos_i(25121) := b"1111111111111111_1111111111111111_1100111000110010_1111011001110100"; -- -0.1945348708263753
	pesos_i(25122) := b"1111111111111111_1111111111111111_1101001101101111_1000001100101010"; -- -0.17407970650548305
	pesos_i(25123) := b"1111111111111111_1111111111111111_1110000101011100_0001111101010011"; -- -0.11968807429461817
	pesos_i(25124) := b"1111111111111111_1111111111111111_1110101001100101_1000111000111010"; -- -0.08438788491918835
	pesos_i(25125) := b"0000000000000000_0000000000000000_0001101011000100_0010111101110110"; -- 0.10455605146644148
	pesos_i(25126) := b"0000000000000000_0000000000000000_0010000100101010_1100101010010101"; -- 0.12955919400058707
	pesos_i(25127) := b"1111111111111111_1111111111111111_1110010101101101_1011110100111110"; -- -0.10379426217048228
	pesos_i(25128) := b"0000000000000000_0000000000000000_0010110110011011_1110000111001111"; -- 0.17815982156664864
	pesos_i(25129) := b"0000000000000000_0000000000000000_0010110010110111_1010111010110011"; -- 0.17467777120116376
	pesos_i(25130) := b"0000000000000000_0000000000000000_0011000001100110_0101011001111111"; -- 0.18906155216491077
	pesos_i(25131) := b"1111111111111111_1111111111111111_1101111111101001_0110101011111101"; -- -0.1253445751298716
	pesos_i(25132) := b"0000000000000000_0000000000000000_0001011101010101_0000100111110010"; -- 0.09114133984255687
	pesos_i(25133) := b"1111111111111111_1111111111111111_1101000110111110_0001110001000000"; -- -0.1806928962574781
	pesos_i(25134) := b"0000000000000000_0000000000000000_0000110110110100_1010100000000111"; -- 0.05353784722332287
	pesos_i(25135) := b"1111111111111111_1111111111111111_1110110000011101_0101001001110000"; -- -0.07767758139179451
	pesos_i(25136) := b"1111111111111111_1111111111111111_1110100111110001_0100010110010010"; -- -0.08616223512139592
	pesos_i(25137) := b"0000000000000000_0000000000000000_0000100000001000_0110111110011010"; -- 0.03137872234792003
	pesos_i(25138) := b"0000000000000000_0000000000000000_0001110000001101_0110100000010110"; -- 0.1095795683525419
	pesos_i(25139) := b"0000000000000000_0000000000000000_0010100000001011_1110101011001000"; -- 0.15643184075210825
	pesos_i(25140) := b"1111111111111111_1111111111111111_1110110110001100_1101100100011101"; -- -0.07206957863613958
	pesos_i(25141) := b"0000000000000000_0000000000000000_0010010110111001_0101101010111100"; -- 0.14735953407925706
	pesos_i(25142) := b"0000000000000000_0000000000000000_0010100011010111_1010010100100000"; -- 0.15954048192339626
	pesos_i(25143) := b"1111111111111111_1111111111111111_1101101011011101_0101000001110011"; -- -0.1450605125683482
	pesos_i(25144) := b"1111111111111111_1111111111111111_1111100000111010_0010011000101001"; -- -0.03036271572105303
	pesos_i(25145) := b"1111111111111111_1111111111111111_1110100000111000_0011011011101001"; -- -0.09289223492607475
	pesos_i(25146) := b"1111111111111111_1111111111111111_1111111001011011_0111101001000010"; -- -0.006416663165654373
	pesos_i(25147) := b"0000000000000000_0000000000000000_0010001110010010_1111010111001100"; -- 0.13896118374839414
	pesos_i(25148) := b"1111111111111111_1111111111111111_1111110011100011_1010000000110000"; -- -0.012151706891794792
	pesos_i(25149) := b"0000000000000000_0000000000000000_0001000000000101_0101001111110101"; -- 0.06258129825696401
	pesos_i(25150) := b"1111111111111111_1111111111111111_1111101111111101_1001101100001101"; -- -0.015661534547177367
	pesos_i(25151) := b"0000000000000000_0000000000000000_0000011110100100_0010110101010001"; -- 0.029848892536104826
	pesos_i(25152) := b"0000000000000000_0000000000000000_0001000001111001_1111001000000000"; -- 0.06436073769010404
	pesos_i(25153) := b"0000000000000000_0000000000000000_0010010101011100_1100000111100010"; -- 0.14594661488105684
	pesos_i(25154) := b"1111111111111111_1111111111111111_1110010111001001_0101111010111011"; -- -0.1023960870506543
	pesos_i(25155) := b"0000000000000000_0000000000000000_0011000000011111_0100000000101011"; -- 0.18797684711089405
	pesos_i(25156) := b"0000000000000000_0000000000000000_0001000010000000_1010011110111001"; -- 0.0644631219623493
	pesos_i(25157) := b"1111111111111111_1111111111111111_1111000011111111_1000110110000110"; -- -0.058600573427716886
	pesos_i(25158) := b"1111111111111111_1111111111111111_1111101001110101_0100011001011101"; -- -0.021648027786968123
	pesos_i(25159) := b"1111111111111111_1111111111111111_1111101010010011_1000110000100110"; -- -0.021186104564597744
	pesos_i(25160) := b"1111111111111111_1111111111111111_1111110001100110_1110100111011011"; -- -0.014054664576907223
	pesos_i(25161) := b"0000000000000000_0000000000000000_0001010111110001_0100010001110001"; -- 0.08571269750890327
	pesos_i(25162) := b"1111111111111111_1111111111111111_1110100100100111_0010001100101000"; -- -0.08924656174420909
	pesos_i(25163) := b"1111111111111111_1111111111111111_1101100010111111_0101110101011011"; -- -0.15333000687537693
	pesos_i(25164) := b"0000000000000000_0000000000000000_0010100010011101_1110010001100110"; -- 0.15865924352061916
	pesos_i(25165) := b"0000000000000000_0000000000000000_0001100001110011_1100010001001100"; -- 0.09551646097536483
	pesos_i(25166) := b"1111111111111111_1111111111111111_1101001111111100_0000011010110101"; -- -0.1719356352904637
	pesos_i(25167) := b"1111111111111111_1111111111111111_1100110110101000_1101010101010000"; -- -0.19664255896800711
	pesos_i(25168) := b"0000000000000000_0000000000000000_0000011001001111_0001010110001101"; -- 0.024644228893298523
	pesos_i(25169) := b"0000000000000000_0000000000000000_0000111111010010_1011100000101010"; -- 0.061809072653294723
	pesos_i(25170) := b"0000000000000000_0000000000000000_0010001110101000_1000011001110101"; -- 0.13929024077260274
	pesos_i(25171) := b"1111111111111111_1111111111111111_1110101101011011_0110010001010000"; -- -0.08063672108578566
	pesos_i(25172) := b"1111111111111111_1111111111111111_1110111000101111_0101010001000101"; -- -0.06959031411600557
	pesos_i(25173) := b"1111111111111111_1111111111111111_1110000000010111_0000100010110000"; -- -0.12464853007766902
	pesos_i(25174) := b"0000000000000000_0000000000000000_0001000111000001_0011110110101101"; -- 0.06935487238221245
	pesos_i(25175) := b"1111111111111111_1111111111111111_1101001010000100_1101101111111110"; -- -0.17766022739179071
	pesos_i(25176) := b"0000000000000000_0000000000000000_0000101111110100_1100010000000010"; -- 0.046703577523022746
	pesos_i(25177) := b"1111111111111111_1111111111111111_1101001101010110_1100100000101110"; -- -0.17445706249596132
	pesos_i(25178) := b"1111111111111111_1111111111111111_1111011000110100_0001011011100001"; -- -0.03826767919775034
	pesos_i(25179) := b"1111111111111111_1111111111111111_1111011111101011_0100001111001101"; -- -0.03156639333875257
	pesos_i(25180) := b"1111111111111111_1111111111111111_1101100110100011_0101101111111010"; -- -0.14985108517368068
	pesos_i(25181) := b"0000000000000000_0000000000000000_0010011110011001_0011010100110000"; -- 0.15468151502358027
	pesos_i(25182) := b"1111111111111111_1111111111111111_1101010100011101_0101010001101110"; -- -0.16752121266146144
	pesos_i(25183) := b"1111111111111111_1111111111111111_1111110111100010_1000011101001100"; -- -0.008262199259266073
	pesos_i(25184) := b"1111111111111111_1111111111111111_1110111101000011_0010111010111010"; -- -0.0653811260585291
	pesos_i(25185) := b"0000000000000000_0000000000000000_0001001011111111_1101010011111100"; -- 0.07421618610451784
	pesos_i(25186) := b"1111111111111111_1111111111111111_1111000110000100_0001000100011101"; -- -0.05657856988826015
	pesos_i(25187) := b"1111111111111111_1111111111111111_1101111101110111_0011010000100100"; -- -0.12708734624156004
	pesos_i(25188) := b"1111111111111111_1111111111111111_1101101110101100_1101000011100001"; -- -0.14189428821072247
	pesos_i(25189) := b"0000000000000000_0000000000000000_0010100100111110_0111010100111010"; -- 0.16110928211510547
	pesos_i(25190) := b"0000000000000000_0000000000000000_0001011011000111_0101010111010000"; -- 0.08897911395020666
	pesos_i(25191) := b"0000000000000000_0000000000000000_0001001000101011_0110110111001110"; -- 0.07097517288098676
	pesos_i(25192) := b"1111111111111111_1111111111111111_1101100000001001_0100000110100111"; -- -0.15610875770824348
	pesos_i(25193) := b"0000000000000000_0000000000000000_0000010111111101_0010101110010100"; -- 0.023394321068018076
	pesos_i(25194) := b"1111111111111111_1111111111111111_1100110100001110_0101111000100011"; -- -0.19899951592911758
	pesos_i(25195) := b"1111111111111111_1111111111111111_1101010000001011_0010011110011101"; -- -0.17170479220115434
	pesos_i(25196) := b"0000000000000000_0000000000000000_0000001000111101_1010100000111100"; -- 0.008753313783376473
	pesos_i(25197) := b"0000000000000000_0000000000000000_0001010000010110_0011011011011011"; -- 0.07846396298877933
	pesos_i(25198) := b"0000000000000000_0000000000000000_0000101011100111_0010011001000001"; -- 0.04258956029893437
	pesos_i(25199) := b"0000000000000000_0000000000000000_0000110111010000_1101011110001100"; -- 0.05396792566633582
	pesos_i(25200) := b"0000000000000000_0000000000000000_0000000001010011_0011110010011110"; -- 0.0012700925632742252
	pesos_i(25201) := b"0000000000000000_0000000000000000_0001100110101010_1111011000010001"; -- 0.10026491085226397
	pesos_i(25202) := b"1111111111111111_1111111111111111_1111100001101100_0111011000110111"; -- -0.029595004707082165
	pesos_i(25203) := b"0000000000000000_0000000000000000_0010011100110101_0000010100101010"; -- 0.15315277363947963
	pesos_i(25204) := b"1111111111111111_1111111111111111_1110001001010001_1011111010101010"; -- -0.11594017366072822
	pesos_i(25205) := b"1111111111111111_1111111111111111_1110110101111111_1010100111100100"; -- -0.072270757415472
	pesos_i(25206) := b"0000000000000000_0000000000000000_0001111100011001_0111011110000011"; -- 0.12148234315998815
	pesos_i(25207) := b"1111111111111111_1111111111111111_1111110111110000_1001011011111110"; -- -0.008047640825387265
	pesos_i(25208) := b"0000000000000000_0000000000000000_0001100001000100_0101011011111011"; -- 0.09479278199939434
	pesos_i(25209) := b"0000000000000000_0000000000000000_0010110011110111_1001000110001011"; -- 0.17565259603121602
	pesos_i(25210) := b"1111111111111111_1111111111111111_1100110010100100_1100111101010100"; -- -0.20061020084681627
	pesos_i(25211) := b"1111111111111111_1111111111111111_1111100011000001_1011011000100111"; -- -0.028294196577368227
	pesos_i(25212) := b"1111111111111111_1111111111111111_1110101001101111_0010111100101001"; -- -0.0842409634648088
	pesos_i(25213) := b"1111111111111111_1111111111111111_1101000101100101_1010101010111100"; -- -0.18204243573092135
	pesos_i(25214) := b"1111111111111111_1111111111111111_1110000110100000_1001101110111111"; -- -0.11864306065587214
	pesos_i(25215) := b"1111111111111111_1111111111111111_1110100010100110_0000001111110000"; -- -0.09121680627977674
	pesos_i(25216) := b"0000000000000000_0000000000000000_0000100101101001_1100100100111011"; -- 0.036770417105138654
	pesos_i(25217) := b"0000000000000000_0000000000000000_0000000100110000_0001011101011100"; -- 0.004640064263078166
	pesos_i(25218) := b"0000000000000000_0000000000000000_0000111100101001_1110010001010101"; -- 0.0592329699942737
	pesos_i(25219) := b"0000000000000000_0000000000000000_0001110000011000_0110010011111001"; -- 0.10974722940683768
	pesos_i(25220) := b"0000000000000000_0000000000000000_0000110101101110_1100000000011000"; -- 0.05247116655960941
	pesos_i(25221) := b"1111111111111111_1111111111111111_1111000100011111_0010111110111011"; -- -0.058117882618859265
	pesos_i(25222) := b"0000000000000000_0000000000000000_0001000111110000_0010001101000000"; -- 0.07007046035393791
	pesos_i(25223) := b"1111111111111111_1111111111111111_1110111011110111_1101100100010010"; -- -0.06653064072286685
	pesos_i(25224) := b"0000000000000000_0000000000000000_0001111101010110_1111111101011100"; -- 0.1224212264630081
	pesos_i(25225) := b"1111111111111111_1111111111111111_1111101100111010_0010100001100000"; -- -0.01864383374542243
	pesos_i(25226) := b"1111111111111111_1111111111111111_1111101101011011_1101110011010010"; -- -0.01812953831509763
	pesos_i(25227) := b"0000000000000000_0000000000000000_0010010101101000_1000000111111011"; -- 0.1461259113967701
	pesos_i(25228) := b"0000000000000000_0000000000000000_0010001011100011_1010100010000110"; -- 0.13628628984294766
	pesos_i(25229) := b"0000000000000000_0000000000000000_0010011011101010_0101111101111101"; -- 0.15201374809307175
	pesos_i(25230) := b"0000000000000000_0000000000000000_0001010101110111_0110100110001101"; -- 0.08385333721573036
	pesos_i(25231) := b"0000000000000000_0000000000000000_0000101111011001_0101100000010011"; -- 0.04628515680022058
	pesos_i(25232) := b"0000000000000000_0000000000000000_0000111001011100_0101000011100001"; -- 0.0560961293896839
	pesos_i(25233) := b"1111111111111111_1111111111111111_1101110101001011_0100010000100011"; -- -0.13557027964346802
	pesos_i(25234) := b"1111111111111111_1111111111111111_1101100000010110_0100000101010111"; -- -0.15591041218065246
	pesos_i(25235) := b"1111111111111111_1111111111111111_1110101111010001_1000010011111010"; -- -0.07883423698904711
	pesos_i(25236) := b"1111111111111111_1111111111111111_1101001110101110_0111101010010111"; -- -0.17311891384381767
	pesos_i(25237) := b"0000000000000000_0000000000000000_0001101010110110_0001001101001100"; -- 0.10434074985701751
	pesos_i(25238) := b"0000000000000000_0000000000000000_0000001111000011_0001100101010101"; -- 0.014695723723706405
	pesos_i(25239) := b"1111111111111111_1111111111111111_1111011010110001_1110011011100110"; -- -0.03634793180192515
	pesos_i(25240) := b"0000000000000000_0000000000000000_0010101111110111_0101000100111110"; -- 0.17174251336920734
	pesos_i(25241) := b"0000000000000000_0000000000000000_0001111011100111_0001101111111111"; -- 0.12071394905358855
	pesos_i(25242) := b"1111111111111111_1111111111111111_1110100000100001_0110111100000000"; -- -0.09323984396108392
	pesos_i(25243) := b"0000000000000000_0000000000000000_0001101000111111_0011001100000110"; -- 0.10252684500035585
	pesos_i(25244) := b"0000000000000000_0000000000000000_0000000101011010_0000110011111001"; -- 0.005280314295531554
	pesos_i(25245) := b"1111111111111111_1111111111111111_1110010101110010_1010101110110100"; -- -0.1037190137009629
	pesos_i(25246) := b"0000000000000000_0000000000000000_0000110101111001_0111110110001100"; -- 0.052635046752604525
	pesos_i(25247) := b"0000000000000000_0000000000000000_0001011000100111_1000100101010001"; -- 0.08654077751250476
	pesos_i(25248) := b"1111111111111111_1111111111111111_1101100001010011_0110111111111010"; -- -0.1549768462172847
	pesos_i(25249) := b"0000000000000000_0000000000000000_0001000001000110_1000010111100000"; -- 0.06357609481391176
	pesos_i(25250) := b"1111111111111111_1111111111111111_1110000100110110_0011111111001111"; -- -0.12026597221453665
	pesos_i(25251) := b"1111111111111111_1111111111111111_1111011110101001_1001110101110000"; -- -0.03256813059449617
	pesos_i(25252) := b"0000000000000000_0000000000000000_0010101000110100_0010011111000100"; -- 0.16485832733563008
	pesos_i(25253) := b"1111111111111111_1111111111111111_1111100100110001_0010100100000101"; -- -0.026593624447786637
	pesos_i(25254) := b"0000000000000000_0000000000000000_0010111011100100_1100000111111001"; -- 0.18317806568687653
	pesos_i(25255) := b"1111111111111111_1111111111111111_1111110100100100_1010010000011110"; -- -0.011159651507101156
	pesos_i(25256) := b"1111111111111111_1111111111111111_1110110110101000_0111111011110011"; -- -0.07164770668640902
	pesos_i(25257) := b"1111111111111111_1111111111111111_1101101110111100_1011110000110001"; -- -0.14165138067989316
	pesos_i(25258) := b"1111111111111111_1111111111111111_1110011100010000_1010011011111011"; -- -0.09740215661981436
	pesos_i(25259) := b"1111111111111111_1111111111111111_1111110011110110_0010000001010010"; -- -0.011869411425685593
	pesos_i(25260) := b"0000000000000000_0000000000000000_0001101101010001_0111000110011111"; -- 0.10671148416782945
	pesos_i(25261) := b"1111111111111111_1111111111111111_1110010101001110_0011111110010010"; -- -0.10427477537093169
	pesos_i(25262) := b"1111111111111111_1111111111111111_1110010001111000_1000000011111101"; -- -0.10753625690096531
	pesos_i(25263) := b"0000000000000000_0000000000000000_0010101110111010_1001010111101111"; -- 0.17081582157262667
	pesos_i(25264) := b"0000000000000000_0000000000000000_0010011011110110_0011100010011101"; -- 0.15219453649965933
	pesos_i(25265) := b"0000000000000000_0000000000000000_0010010000111101_0101111100001010"; -- 0.1415614510139822
	pesos_i(25266) := b"1111111111111111_1111111111111111_1101100010111001_1100011011110101"; -- -0.15341526531864333
	pesos_i(25267) := b"0000000000000000_0000000000000000_0001011101001101_1011110001111110"; -- 0.09102991181469293
	pesos_i(25268) := b"0000000000000000_0000000000000000_0001011100001001_1010100010001010"; -- 0.08999112478631205
	pesos_i(25269) := b"1111111111111111_1111111111111111_1101001100000100_1110110111010111"; -- -0.17570603839328758
	pesos_i(25270) := b"1111111111111111_1111111111111111_1101101001000010_0111001001001101"; -- -0.14742360716770922
	pesos_i(25271) := b"1111111111111111_1111111111111111_1110000010101101_1011101110010110"; -- -0.12234904850275259
	pesos_i(25272) := b"1111111111111111_1111111111111111_1111110011110110_1111100011010000"; -- -0.011856507441747871
	pesos_i(25273) := b"1111111111111111_1111111111111111_1110001111110101_0100101100000111"; -- -0.10953837468870206
	pesos_i(25274) := b"1111111111111111_1111111111111111_1110101001001110_0101010111010001"; -- -0.08474219943037689
	pesos_i(25275) := b"1111111111111111_1111111111111111_1110111110110001_1111000110110100"; -- -0.06369103760761317
	pesos_i(25276) := b"0000000000000000_0000000000000000_0000101110010101_1011111110111100"; -- 0.045253737896937325
	pesos_i(25277) := b"1111111111111111_1111111111111111_1110110001001101_1011110100000011"; -- -0.07693880724909224
	pesos_i(25278) := b"0000000000000000_0000000000000000_0001100001001101_0101100011111001"; -- 0.09493022983016407
	pesos_i(25279) := b"0000000000000000_0000000000000000_0011001100101010_1101001111011011"; -- 0.19987224666857345
	pesos_i(25280) := b"0000000000000000_0000000000000000_0010001001111110_0010111101010010"; -- 0.1347379279995208
	pesos_i(25281) := b"1111111111111111_1111111111111111_1111111110000001_1100100101010011"; -- -0.0019258662827724188
	pesos_i(25282) := b"1111111111111111_1111111111111111_1110111110111111_0001001010111110"; -- -0.06349070413769291
	pesos_i(25283) := b"1111111111111111_1111111111111111_1110001000001000_0111001000111001"; -- -0.11705862147182397
	pesos_i(25284) := b"0000000000000000_0000000000000000_0001111010111000_1111001011011111"; -- 0.12000959334193706
	pesos_i(25285) := b"0000000000000000_0000000000000000_0011010001111100_0110110101000101"; -- 0.20502360282726806
	pesos_i(25286) := b"1111111111111111_1111111111111111_1110000000101000_1100110000000000"; -- -0.12437748908533516
	pesos_i(25287) := b"0000000000000000_0000000000000000_0010011101111010_0000000011110000"; -- 0.15420537809620707
	pesos_i(25288) := b"0000000000000000_0000000000000000_0010100011101010_1011110101100011"; -- 0.15983184505308437
	pesos_i(25289) := b"1111111111111111_1111111111111111_1101000100101100_1000000110001100"; -- -0.18291464174191022
	pesos_i(25290) := b"1111111111111111_1111111111111111_1111111000000011_1111100110111001"; -- -0.007751839043684736
	pesos_i(25291) := b"1111111111111111_1111111111111111_1111101110000111_0000110010100000"; -- -0.017470561023185515
	pesos_i(25292) := b"0000000000000000_0000000000000000_0000001100011111_1001011110001110"; -- 0.012200805762289062
	pesos_i(25293) := b"0000000000000000_0000000000000000_0010010101010110_0110100110011101"; -- 0.14584980095019845
	pesos_i(25294) := b"0000000000000000_0000000000000000_0011000001100000_0010110101010111"; -- 0.18896754616998385
	pesos_i(25295) := b"1111111111111111_1111111111111111_1110110101010010_0010011110000110"; -- -0.07296517350008525
	pesos_i(25296) := b"0000000000000000_0000000000000000_0001110010001001_1111111110001010"; -- 0.11148068532103206
	pesos_i(25297) := b"0000000000000000_0000000000000000_0000001100010011_0111110000111011"; -- 0.01201607173084727
	pesos_i(25298) := b"0000000000000000_0000000000000000_0001111000100010_0010001111101110"; -- 0.11770844033060655
	pesos_i(25299) := b"1111111111111111_1111111111111111_1111011000001011_0101011111000110"; -- -0.03888942170113478
	pesos_i(25300) := b"1111111111111111_1111111111111111_1111011010110001_0001110101111111"; -- -0.03635993611853087
	pesos_i(25301) := b"1111111111111111_1111111111111111_1111001110111101_1000000010010001"; -- -0.04788967562460281
	pesos_i(25302) := b"0000000000000000_0000000000000000_0001101011100110_0110000001000111"; -- 0.1050777599835764
	pesos_i(25303) := b"0000000000000000_0000000000000000_0010011001101101_0101000011000010"; -- 0.15010552147815234
	pesos_i(25304) := b"1111111111111111_1111111111111111_1111100101010000_1010000000100010"; -- -0.026113502137994155
	pesos_i(25305) := b"1111111111111111_1111111111111111_1111001101101100_1010010000101100"; -- -0.049123515361235964
	pesos_i(25306) := b"0000000000000000_0000000000000000_0010010010111010_0100011100101000"; -- 0.1434673759533832
	pesos_i(25307) := b"1111111111111111_1111111111111111_1101110001001100_0100111111111001"; -- -0.13946056529185258
	pesos_i(25308) := b"0000000000000000_0000000000000000_0010100101000110_1110000100000110"; -- 0.1612377776587268
	pesos_i(25309) := b"0000000000000000_0000000000000000_0000101110100011_1010110100010000"; -- 0.0454662479210279
	pesos_i(25310) := b"1111111111111111_1111111111111111_1110101010111100_1001001110101111"; -- -0.08306004513442117
	pesos_i(25311) := b"1111111111111111_1111111111111111_1111100010001001_0111011100000011"; -- -0.02915245219961888
	pesos_i(25312) := b"1111111111111111_1111111111111111_1110010001001111_1000011101010011"; -- -0.10816148965008207
	pesos_i(25313) := b"1111111111111111_1111111111111111_1110110000111110_1111000001101011"; -- -0.07716462513329585
	pesos_i(25314) := b"1111111111111111_1111111111111111_1101111101010011_0110011111001011"; -- -0.12763358391496094
	pesos_i(25315) := b"1111111111111111_1111111111111111_1110010100000010_1101010110010011"; -- -0.10542550238214451
	pesos_i(25316) := b"0000000000000000_0000000000000000_0001000011000111_0100000011101111"; -- 0.06554036926072448
	pesos_i(25317) := b"0000000000000000_0000000000000000_0001011001000010_0101010010110101"; -- 0.086949629116935
	pesos_i(25318) := b"0000000000000000_0000000000000000_0000110101011010_1011011101111001"; -- 0.052165476897756725
	pesos_i(25319) := b"0000000000000000_0000000000000000_0000101110110110_1011001011100011"; -- 0.04575651218395995
	pesos_i(25320) := b"0000000000000000_0000000000000000_0000100100110110_0101001110010101"; -- 0.03598520638850751
	pesos_i(25321) := b"0000000000000000_0000000000000000_0000001000010010_0011010001111010"; -- 0.008090286107206196
	pesos_i(25322) := b"1111111111111111_1111111111111111_1101101000101100_0100011110001010"; -- -0.14776184912445653
	pesos_i(25323) := b"1111111111111111_1111111111111111_1110110100001100_0001111111100000"; -- -0.0740337447326827
	pesos_i(25324) := b"1111111111111111_1111111111111111_1110001001100000_1101001011110100"; -- -0.11571008240842072
	pesos_i(25325) := b"1111111111111111_1111111111111111_1101011010000000_1100011110111110"; -- -0.16209746943218112
	pesos_i(25326) := b"0000000000000000_0000000000000000_0001111101110111_0101110111010000"; -- 0.12291513751196523
	pesos_i(25327) := b"0000000000000000_0000000000000000_0001111110011000_1001101110111110"; -- 0.12342236878297841
	pesos_i(25328) := b"1111111111111111_1111111111111111_1111001111011000_1111111001101111"; -- -0.04747018614669606
	pesos_i(25329) := b"0000000000000000_0000000000000000_0010000100011110_1010010011101000"; -- 0.12937384285282016
	pesos_i(25330) := b"1111111111111111_1111111111111111_1110110110100000_0100100000001001"; -- -0.07177305020366048
	pesos_i(25331) := b"0000000000000000_0000000000000000_0001011001100101_0001010110111100"; -- 0.08747993321291613
	pesos_i(25332) := b"1111111111111111_1111111111111111_1101110111110001_1011110111000010"; -- -0.133030071483543
	pesos_i(25333) := b"1111111111111111_1111111111111111_1110010000011011_1000100000110110"; -- -0.10895489393515866
	pesos_i(25334) := b"0000000000000000_0000000000000000_0000100110001110_1111111101111000"; -- 0.03733822526521307
	pesos_i(25335) := b"0000000000000000_0000000000000000_0011001011110011_1000011011111001"; -- 0.1990284307241728
	pesos_i(25336) := b"0000000000000000_0000000000000000_0000101101011100_0011101110011010"; -- 0.04437611106010198
	pesos_i(25337) := b"0000000000000000_0000000000000000_0011001101100011_1000101011001110"; -- 0.20073764362805527
	pesos_i(25338) := b"0000000000000000_0000000000000000_0010101100111010_0111111101001011"; -- 0.1688613469783928
	pesos_i(25339) := b"0000000000000000_0000000000000000_0000010110010010_0000000000000110"; -- 0.021759034584836332
	pesos_i(25340) := b"0000000000000000_0000000000000000_0000101100001001_0100101101000001"; -- 0.04311056462563149
	pesos_i(25341) := b"0000000000000000_0000000000000000_0000010011110011_0000111011110001"; -- 0.019333776266264122
	pesos_i(25342) := b"0000000000000000_0000000000000000_0010010111000010_1110010111110000"; -- 0.14750516033660535
	pesos_i(25343) := b"0000000000000000_0000000000000000_0000001011011101_0100101100000101"; -- 0.011189163928231868
	pesos_i(25344) := b"1111111111111111_1111111111111111_1111101101000110_1100011101011100"; -- -0.018451252091724858
	pesos_i(25345) := b"0000000000000000_0000000000000000_0001011110001100_0101001101011100"; -- 0.09198494909695001
	pesos_i(25346) := b"1111111111111111_1111111111111111_1101111010010011_0101100101100100"; -- -0.1305641298485282
	pesos_i(25347) := b"0000000000000000_0000000000000000_0010010010011000_0010010010101100"; -- 0.14294652168371166
	pesos_i(25348) := b"1111111111111111_1111111111111111_1110101010010110_0001110110110000"; -- -0.0836469120463661
	pesos_i(25349) := b"0000000000000000_0000000000000000_0000000001110101_1111011010101010"; -- 0.001799980731513691
	pesos_i(25350) := b"1111111111111111_1111111111111111_1110010110101001_0110000111110000"; -- -0.10288417718964357
	pesos_i(25351) := b"0000000000000000_0000000000000000_0000111110110000_1011010001011010"; -- 0.06129004667561559
	pesos_i(25352) := b"1111111111111111_1111111111111111_1111010011111001_1101010101000111"; -- -0.04306284926211905
	pesos_i(25353) := b"0000000000000000_0000000000000000_0000010100000001_0000001101000110"; -- 0.01954670379832477
	pesos_i(25354) := b"0000000000000000_0000000000000000_0000010011000010_0110011110100010"; -- 0.018591382069749415
	pesos_i(25355) := b"1111111111111111_1111111111111111_1110110110101010_0000111001110010"; -- -0.07162389496775115
	pesos_i(25356) := b"0000000000000000_0000000000000000_0001011001110001_0000000100010101"; -- 0.0876618075873479
	pesos_i(25357) := b"1111111111111111_1111111111111111_1111110001101101_1100111001010110"; -- -0.013949493330075653
	pesos_i(25358) := b"1111111111111111_1111111111111111_1101101001101110_1001111111110110"; -- -0.14674949869525572
	pesos_i(25359) := b"1111111111111111_1111111111111111_1110000000010011_1101100110101111"; -- -0.12469710799337387
	pesos_i(25360) := b"1111111111111111_1111111111111111_1110111100010011_1101010100101101"; -- -0.06610362666515548
	pesos_i(25361) := b"1111111111111111_1111111111111111_1111101001000001_1011100100000000"; -- -0.022434651893656336
	pesos_i(25362) := b"1111111111111111_1111111111111111_1101100000100110_0001001000010011"; -- -0.15566908862223514
	pesos_i(25363) := b"1111111111111111_1111111111111111_1110110001010101_1000010100011000"; -- -0.07682006983756128
	pesos_i(25364) := b"0000000000000000_0000000000000000_0001011000110111_1000110111100111"; -- 0.08678519143777959
	pesos_i(25365) := b"1111111111111111_1111111111111111_1101111001111100_0010100111011011"; -- -0.13091791545213746
	pesos_i(25366) := b"1111111111111111_1111111111111111_1101101111000101_0110111100111001"; -- -0.14151863913158041
	pesos_i(25367) := b"1111111111111111_1111111111111111_1111010010101001_1001101010010011"; -- -0.044287051254196526
	pesos_i(25368) := b"1111111111111111_1111111111111111_1101001110110011_1010000111000110"; -- -0.17304028429343818
	pesos_i(25369) := b"1111111111111111_1111111111111111_1111100111000110_1110100101101000"; -- -0.02430859765390378
	pesos_i(25370) := b"1111111111111111_1111111111111111_1101110110010111_0010100111010101"; -- -0.13441217953112364
	pesos_i(25371) := b"0000000000000000_0000000000000000_0000110100011110_1010101000101100"; -- 0.05124915677735103
	pesos_i(25372) := b"1111111111111111_1111111111111111_1101011011000010_0100100101000100"; -- -0.16109792800246164
	pesos_i(25373) := b"0000000000000000_0000000000000000_0001011011001000_1011110001011001"; -- 0.08900048420205257
	pesos_i(25374) := b"0000000000000000_0000000000000000_0011011010110111_0000010011111001"; -- 0.21373015485507482
	pesos_i(25375) := b"1111111111111111_1111111111111111_1101000000001110_0111100110111101"; -- -0.18727912089731652
	pesos_i(25376) := b"1111111111111111_1111111111111111_1111100100000101_1110011000101000"; -- -0.02725373763854575
	pesos_i(25377) := b"0000000000000000_0000000000000000_0001000010110011_0101111111001011"; -- 0.06523703301755458
	pesos_i(25378) := b"1111111111111111_1111111111111111_1111101000111111_1101110001001111"; -- -0.0224630648320649
	pesos_i(25379) := b"1111111111111111_1111111111111111_1101101001000000_1000010101110010"; -- -0.14745298364607373
	pesos_i(25380) := b"0000000000000000_0000000000000000_0010001010100010_1010111001110110"; -- 0.13529482252344224
	pesos_i(25381) := b"1111111111111111_1111111111111111_1111100010010100_0011011011110000"; -- -0.02898842471568752
	pesos_i(25382) := b"0000000000000000_0000000000000000_0001001001111111_1111010011100010"; -- 0.07226496230188376
	pesos_i(25383) := b"0000000000000000_0000000000000000_0000101110101111_0001000010101101"; -- 0.04564003201396453
	pesos_i(25384) := b"1111111111111111_1111111111111111_1110011101001110_0010110100000000"; -- -0.09646338223811624
	pesos_i(25385) := b"0000000000000000_0000000000000000_0011000001000110_1010100010110100"; -- 0.18857817077985692
	pesos_i(25386) := b"1111111111111111_1111111111111111_1110110100011110_1101010011110000"; -- -0.07374829419784652
	pesos_i(25387) := b"0000000000000000_0000000000000000_0010110101110100_1110000101011010"; -- 0.1775647014825887
	pesos_i(25388) := b"1111111111111111_1111111111111111_1110010100101000_1111101000010110"; -- -0.10484349218795908
	pesos_i(25389) := b"0000000000000000_0000000000000000_0000001100111100_1011011001010101"; -- 0.012645145095316621
	pesos_i(25390) := b"0000000000000000_0000000000000000_0010110000100010_1101000010100001"; -- 0.17240623404580202
	pesos_i(25391) := b"1111111111111111_1111111111111111_1100110100100100_0100101100101010"; -- -0.19866495355850552
	pesos_i(25392) := b"0000000000000000_0000000000000000_0011001100100001_0101101100110000"; -- 0.19972772525770263
	pesos_i(25393) := b"1111111111111111_1111111111111111_1101101001010100_0110111000010011"; -- -0.1471492008967074
	pesos_i(25394) := b"1111111111111111_1111111111111111_1101010000110010_1010100001011010"; -- -0.17110202608224317
	pesos_i(25395) := b"1111111111111111_1111111111111111_1101000100010101_0000001011011111"; -- -0.18327314421450044
	pesos_i(25396) := b"0000000000000000_0000000000000000_0000000110001101_1001111101011011"; -- 0.006067237612724124
	pesos_i(25397) := b"0000000000000000_0000000000000000_0001000111111101_0001110100001010"; -- 0.07026845459016069
	pesos_i(25398) := b"0000000000000000_0000000000000000_0010101111111001_1110101010010010"; -- 0.1717821700723169
	pesos_i(25399) := b"0000000000000000_0000000000000000_0000000101000011_0110011110110011"; -- 0.004934769787148699
	pesos_i(25400) := b"0000000000000000_0000000000000000_0000010010110000_1010011001000001"; -- 0.01832045647807279
	pesos_i(25401) := b"0000000000000000_0000000000000000_0010001001101100_1101101100111001"; -- 0.1344735159641409
	pesos_i(25402) := b"0000000000000000_0000000000000000_0010010101011100_1100011011011001"; -- 0.14594691093916767
	pesos_i(25403) := b"1111111111111111_1111111111111111_1101011111101011_0001101010101100"; -- -0.15656884484493225
	pesos_i(25404) := b"1111111111111111_1111111111111111_1101010110101111_0100101011111110"; -- -0.16529399206645878
	pesos_i(25405) := b"1111111111111111_1111111111111111_1101001000100100_1111000010000100"; -- -0.17912384780086235
	pesos_i(25406) := b"0000000000000000_0000000000000000_0010011000011000_1111110101000100"; -- 0.1488188068091291
	pesos_i(25407) := b"1111111111111111_1111111111111111_1101100010110101_1101011001010011"; -- -0.15347538439516822
	pesos_i(25408) := b"0000000000000000_0000000000000000_0000100010110111_1101000101000110"; -- 0.034054832105257976
	pesos_i(25409) := b"1111111111111111_1111111111111111_1101010000001001_0111101011010010"; -- -0.17173035015511134
	pesos_i(25410) := b"0000000000000000_0000000000000000_0001010100100001_0100110111101101"; -- 0.0825394347956951
	pesos_i(25411) := b"0000000000000000_0000000000000000_0001010011100001_0001001001000110"; -- 0.08155931678375174
	pesos_i(25412) := b"1111111111111111_1111111111111111_1100110110010010_0101111100011110"; -- -0.19698529739012138
	pesos_i(25413) := b"1111111111111111_1111111111111111_1100110000010100_0100011111011111"; -- -0.20281554028486048
	pesos_i(25414) := b"0000000000000000_0000000000000000_0011001000001001_0110010001100001"; -- 0.19545581220532512
	pesos_i(25415) := b"1111111111111111_1111111111111111_1101011011101111_1100100111000111"; -- -0.16040362254083637
	pesos_i(25416) := b"0000000000000000_0000000000000000_0000111111110001_1000001101010001"; -- 0.06227894513867831
	pesos_i(25417) := b"0000000000000000_0000000000000000_0011000000011011_0110110001011110"; -- 0.18791844649540113
	pesos_i(25418) := b"0000000000000000_0000000000000000_0001100101000100_1110001010001010"; -- 0.09870735050098638
	pesos_i(25419) := b"0000000000000000_0000000000000000_0010000001000001_0000011101000110"; -- 0.12599225481545065
	pesos_i(25420) := b"1111111111111111_1111111111111111_1101010001001000_1100010001010101"; -- -0.1707646649690852
	pesos_i(25421) := b"1111111111111111_1111111111111111_1101110111100001_0101000111011010"; -- -0.13328064375185422
	pesos_i(25422) := b"1111111111111111_1111111111111111_1110010110001101_1100011110001010"; -- -0.10330536726544015
	pesos_i(25423) := b"0000000000000000_0000000000000000_0000001101100101_0100010000110011"; -- 0.013263952716798961
	pesos_i(25424) := b"0000000000000000_0000000000000000_0001101011110011_0010011111110001"; -- 0.10527276654361052
	pesos_i(25425) := b"1111111111111111_1111111111111111_1110001000011001_0011100000110101"; -- -0.1168026801186973
	pesos_i(25426) := b"0000000000000000_0000000000000000_0000101110000111_1011011100100100"; -- 0.045039602603160214
	pesos_i(25427) := b"1111111111111111_1111111111111111_1101110001100110_0001101110100011"; -- -0.1390669562415042
	pesos_i(25428) := b"1111111111111111_1111111111111111_1111110101111100_1111100010101000"; -- -0.009811839089283169
	pesos_i(25429) := b"1111111111111111_1111111111111111_1101010000101110_0010110001111001"; -- -0.1711704448466056
	pesos_i(25430) := b"1111111111111111_1111111111111111_1101010101111111_0011100011110010"; -- -0.16602748963792233
	pesos_i(25431) := b"1111111111111111_1111111111111111_1111101001001010_1100010101111111"; -- -0.02229657787235028
	pesos_i(25432) := b"1111111111111111_1111111111111111_1101101010100001_0110001001111100"; -- -0.14597496489172967
	pesos_i(25433) := b"0000000000000000_0000000000000000_0010101001001011_0010000000001101"; -- 0.1652088196239944
	pesos_i(25434) := b"1111111111111111_1111111111111111_1101110101011010_0100011111000000"; -- -0.13534118239319615
	pesos_i(25435) := b"0000000000000000_0000000000000000_0000111011001100_1100101010010100"; -- 0.057812367479700165
	pesos_i(25436) := b"0000000000000000_0000000000000000_0010100001010010_1011100100000100"; -- 0.15751224860831053
	pesos_i(25437) := b"1111111111111111_1111111111111111_1101101111100011_0100001110000011"; -- -0.14106348091458254
	pesos_i(25438) := b"1111111111111111_1111111111111111_1110110100011011_0001111000000100"; -- -0.07380497361171304
	pesos_i(25439) := b"1111111111111111_1111111111111111_1110111101011010_1001101100100100"; -- -0.06502371197196437
	pesos_i(25440) := b"1111111111111111_1111111111111111_1110111101001101_1001001100010110"; -- -0.06522255628604268
	pesos_i(25441) := b"0000000000000000_0000000000000000_0001110010100000_1101100010010011"; -- 0.11182931500417784
	pesos_i(25442) := b"0000000000000000_0000000000000000_0010100110101010_0111011000110011"; -- 0.1627572892946818
	pesos_i(25443) := b"1111111111111111_1111111111111111_1110010011010110_1010001000000001"; -- -0.10609996292092168
	pesos_i(25444) := b"1111111111111111_1111111111111111_1110101010010100_1010111010100101"; -- -0.0836687894928687
	pesos_i(25445) := b"1111111111111111_1111111111111111_1111011101000011_0101111000111101"; -- -0.03412829400373777
	pesos_i(25446) := b"1111111111111111_1111111111111111_1110100011000101_0111011011011110"; -- -0.09073693355810049
	pesos_i(25447) := b"1111111111111111_1111111111111111_1111000100000001_1001111011100010"; -- -0.05856902101719421
	pesos_i(25448) := b"0000000000000000_0000000000000000_0000101000110111_1101011000011110"; -- 0.039914495805677755
	pesos_i(25449) := b"0000000000000000_0000000000000000_0010100110101100_0010101000110000"; -- 0.1627832763076792
	pesos_i(25450) := b"0000000000000000_0000000000000000_0011001001111001_0111110111110110"; -- 0.19716632126757425
	pesos_i(25451) := b"0000000000000000_0000000000000000_0010111101110110_1100100011011011"; -- 0.18540625914196016
	pesos_i(25452) := b"1111111111111111_1111111111111111_1110101110101100_1110110010010011"; -- -0.07939263739239208
	pesos_i(25453) := b"0000000000000000_0000000000000000_0000101001110100_0011111100110001"; -- 0.040836286141976486
	pesos_i(25454) := b"1111111111111111_1111111111111111_1110001100101111_1110101010001111"; -- -0.11255010614328932
	pesos_i(25455) := b"0000000000000000_0000000000000000_0001101101110110_0001111111100110"; -- 0.107271188446177
	pesos_i(25456) := b"0000000000000000_0000000000000000_0001101011100011_1110111011100101"; -- 0.1050404843144623
	pesos_i(25457) := b"0000000000000000_0000000000000000_0000000001000001_0101001001010101"; -- 0.0009967287054340995
	pesos_i(25458) := b"0000000000000000_0000000000000000_0010000000101110_0001000100010101"; -- 0.12570292239176326
	pesos_i(25459) := b"0000000000000000_0000000000000000_0001000110101110_1011010101011011"; -- 0.069072088874197
	pesos_i(25460) := b"1111111111111111_1111111111111111_1101101011100011_1011011000010100"; -- -0.14496290216641375
	pesos_i(25461) := b"0000000000000000_0000000000000000_0011010000101001_0100110001111011"; -- 0.20375516905446125
	pesos_i(25462) := b"0000000000000000_0000000000000000_0010000111110011_0000100111010110"; -- 0.13261472190983764
	pesos_i(25463) := b"0000000000000000_0000000000000000_0001110100101101_0001111011001010"; -- 0.11396973061792766
	pesos_i(25464) := b"0000000000000000_0000000000000000_0011000110100000_0011001111101011"; -- 0.19385075073575933
	pesos_i(25465) := b"0000000000000000_0000000000000000_0001111110000100_1110001000100001"; -- 0.12312138839162709
	pesos_i(25466) := b"0000000000000000_0000000000000000_0010010111000111_1111100110011100"; -- 0.14758262693394386
	pesos_i(25467) := b"1111111111111111_1111111111111111_1101010000011011_0000100010100100"; -- -0.1714624976091692
	pesos_i(25468) := b"1111111111111111_1111111111111111_1110010100110100_0111101111000001"; -- -0.10466791654771708
	pesos_i(25469) := b"0000000000000000_0000000000000000_0010111100010110_0000001001100100"; -- 0.1839295859486881
	pesos_i(25470) := b"0000000000000000_0000000000000000_0001100001111001_0111100001101100"; -- 0.09560349125387962
	pesos_i(25471) := b"1111111111111111_1111111111111111_1101111011110100_1010110010001110"; -- -0.12907907048979975
	pesos_i(25472) := b"1111111111111111_1111111111111111_1101001001101000_1011000110001011"; -- -0.17809000358489022
	pesos_i(25473) := b"1111111111111111_1111111111111111_1110101011110001_1000000000001101"; -- -0.08225249936900372
	pesos_i(25474) := b"0000000000000000_0000000000000000_0000011101101111_1010111011111001"; -- 0.02904790478046169
	pesos_i(25475) := b"1111111111111111_1111111111111111_1111100000001100_0100111111100011"; -- -0.031062132843193785
	pesos_i(25476) := b"0000000000000000_0000000000000000_0000100011101111_1110010101011101"; -- 0.03491052166070352
	pesos_i(25477) := b"0000000000000000_0000000000000000_0000011000000010_0010101000100000"; -- 0.02347052838141315
	pesos_i(25478) := b"1111111111111111_1111111111111111_1111100001010100_1001000101000000"; -- -0.02995960411772457
	pesos_i(25479) := b"0000000000000000_0000000000000000_0010100001011001_0001010010111000"; -- 0.15760926705807365
	pesos_i(25480) := b"0000000000000000_0000000000000000_0010010010110110_0101011111111100"; -- 0.1434073438909616
	pesos_i(25481) := b"1111111111111111_1111111111111111_1111001000100011_1011011111011111"; -- -0.05414248279375071
	pesos_i(25482) := b"1111111111111111_1111111111111111_1100100000000011_1000101000000101"; -- -0.21869599697126713
	pesos_i(25483) := b"0000000000000000_0000000000000000_0001010110110000_1001001011000001"; -- 0.08472554400353104
	pesos_i(25484) := b"1111111111111111_1111111111111111_1101111111001010_0011110111011111"; -- -0.12582028669033285
	pesos_i(25485) := b"0000000000000000_0000000000000000_0010110110001000_1001000111101101"; -- 0.1778651431530197
	pesos_i(25486) := b"0000000000000000_0000000000000000_0010010100110100_1111010110110001"; -- 0.14533935143700205
	pesos_i(25487) := b"1111111111111111_1111111111111111_1101010000011011_1010100101111011"; -- -0.17145291088112685
	pesos_i(25488) := b"1111111111111111_1111111111111111_1110001000111101_1011111100111010"; -- -0.11624531586923224
	pesos_i(25489) := b"0000000000000000_0000000000000000_0001001111000001_1111000011100101"; -- 0.07717805479191239
	pesos_i(25490) := b"0000000000000000_0000000000000000_0010000111000011_1001010100011101"; -- 0.13189060166495756
	pesos_i(25491) := b"1111111111111111_1111111111111111_1110000101100010_1011100001111011"; -- -0.11958739268535505
	pesos_i(25492) := b"1111111111111111_1111111111111111_1100111010000001_1111100011010011"; -- -0.19332928506457644
	pesos_i(25493) := b"0000000000000000_0000000000000000_0001111001101111_1001101101011100"; -- 0.11889048572434376
	pesos_i(25494) := b"1111111111111111_1111111111111111_1101001111110100_0011101100101010"; -- -0.1720545789171032
	pesos_i(25495) := b"1111111111111111_1111111111111111_1101110110111001_1010101101110011"; -- -0.13388565485566065
	pesos_i(25496) := b"1111111111111111_1111111111111111_1110011111000111_1011111100001010"; -- -0.0946083642669379
	pesos_i(25497) := b"1111111111111111_1111111111111111_1111000000100100_0010001110011110"; -- -0.06194856074871361
	pesos_i(25498) := b"1111111111111111_1111111111111111_1110010101101011_1111111110101100"; -- -0.10382082045134826
	pesos_i(25499) := b"0000000000000000_0000000000000000_0001110000111010_0011010101100100"; -- 0.11026319218583033
	pesos_i(25500) := b"0000000000000000_0000000000000000_0010111001110101_1001101110011011"; -- 0.18148205318131022
	pesos_i(25501) := b"1111111111111111_1111111111111111_1101101001011101_1100111100110110"; -- -0.14700608197479362
	pesos_i(25502) := b"0000000000000000_0000000000000000_0000100110110011_0010001010101011"; -- 0.03788963962704949
	pesos_i(25503) := b"0000000000000000_0000000000000000_0001010100010110_0101100001010111"; -- 0.08237220885717987
	pesos_i(25504) := b"1111111111111111_1111111111111111_1101011100100000_0100000001010111"; -- -0.15966413385118
	pesos_i(25505) := b"1111111111111111_1111111111111111_1111111001111000_0100100011100000"; -- -0.005977101727413699
	pesos_i(25506) := b"1111111111111111_1111111111111111_1101000000111101_1101111110110101"; -- -0.18655587982439295
	pesos_i(25507) := b"1111111111111111_1111111111111111_1101100000110110_0110111000001101"; -- -0.15541946585017066
	pesos_i(25508) := b"0000000000000000_0000000000000000_0000000110110111_0011101101100001"; -- 0.006702147714818676
	pesos_i(25509) := b"1111111111111111_1111111111111111_1101010011000101_1011001100000101"; -- -0.1688583480843404
	pesos_i(25510) := b"0000000000000000_0000000000000000_0000010110000011_1010011001110001"; -- 0.021540072031492698
	pesos_i(25511) := b"1111111111111111_1111111111111111_1101110100110001_0000101100100001"; -- -0.13597040604514354
	pesos_i(25512) := b"1111111111111111_1111111111111111_1110001110100000_1010100001010100"; -- -0.11082981050094169
	pesos_i(25513) := b"1111111111111111_1111111111111111_1101101011011111_1001011111000110"; -- -0.14502574361219514
	pesos_i(25514) := b"0000000000000000_0000000000000000_0001110001001111_1110001010010010"; -- 0.11059394899890408
	pesos_i(25515) := b"0000000000000000_0000000000000000_0010011100111010_1010101000110000"; -- 0.15323890363051615
	pesos_i(25516) := b"1111111111111111_1111111111111111_1111001010010101_1111011111111110"; -- -0.05239915902088419
	pesos_i(25517) := b"1111111111111111_1111111111111111_1111010100100000_0101010100111111"; -- -0.04247538777497555
	pesos_i(25518) := b"1111111111111111_1111111111111111_1110111111000111_1100011100100101"; -- -0.06335788097267296
	pesos_i(25519) := b"0000000000000000_0000000000000000_0001001111010101_0110100000010101"; -- 0.07747507576477589
	pesos_i(25520) := b"1111111111111111_1111111111111111_1111101100111110_0100101111111010"; -- -0.018580676467691754
	pesos_i(25521) := b"0000000000000000_0000000000000000_0001111110001101_1111011001010010"; -- 0.12325992115107008
	pesos_i(25522) := b"0000000000000000_0000000000000000_0001000010010101_0001111000111101"; -- 0.06477536193977572
	pesos_i(25523) := b"1111111111111111_1111111111111111_1110000110001011_0101100100101010"; -- -0.11896746364009461
	pesos_i(25524) := b"1111111111111111_1111111111111111_1110011100001001_0100111010111100"; -- -0.09751422801918251
	pesos_i(25525) := b"0000000000000000_0000000000000000_0000100011011110_1001110010000011"; -- 0.034646779940386715
	pesos_i(25526) := b"0000000000000000_0000000000000000_0010010111111000_0111010110010101"; -- 0.148322438208352
	pesos_i(25527) := b"1111111111111111_1111111111111111_1101000011110100_0101111011000010"; -- -0.18377120756388188
	pesos_i(25528) := b"0000000000000000_0000000000000000_0010011111001111_1000100100100100"; -- 0.15551049364851113
	pesos_i(25529) := b"1111111111111111_1111111111111111_1101111000000001_0000011110011011"; -- -0.1327967878731508
	pesos_i(25530) := b"1111111111111111_1111111111111111_1110111000000101_1011001011000101"; -- -0.07022555063872186
	pesos_i(25531) := b"1111111111111111_1111111111111111_1110000100001011_1011101011010000"; -- -0.12091476832146693
	pesos_i(25532) := b"0000000000000000_0000000000000000_0001101110111001_1111001000001110"; -- 0.10830605365404619
	pesos_i(25533) := b"0000000000000000_0000000000000000_0000111111001100_1111011100100001"; -- 0.06172127306591489
	pesos_i(25534) := b"0000000000000000_0000000000000000_0010110101111001_0100111001010101"; -- 0.17763223238803413
	pesos_i(25535) := b"0000000000000000_0000000000000000_0001010111111000_0111000000000011"; -- 0.08582210604062669
	pesos_i(25536) := b"1111111111111111_1111111111111111_1111101000101000_0010001010011101"; -- -0.02282508521105558
	pesos_i(25537) := b"1111111111111111_1111111111111111_1100111110001101_0111011001100001"; -- -0.18924770476052594
	pesos_i(25538) := b"1111111111111111_1111111111111111_1111100000001000_1111111110111011"; -- -0.031112686937044415
	pesos_i(25539) := b"0000000000000000_0000000000000000_0000110111101100_0000000001110000"; -- 0.05438235030558286
	pesos_i(25540) := b"1111111111111111_1111111111111111_1111100100110111_1101101010010100"; -- -0.026491488294971388
	pesos_i(25541) := b"0000000000000000_0000000000000000_0001110000100010_1000001110010111"; -- 0.10990164215720757
	pesos_i(25542) := b"0000000000000000_0000000000000000_0000110111000101_0111100000101111"; -- 0.053794394987263745
	pesos_i(25543) := b"1111111111111111_1111111111111111_1101001101111011_1111011101001011"; -- -0.17388967921417173
	pesos_i(25544) := b"1111111111111111_1111111111111111_1101101101010111_1110111110010001"; -- -0.14318945598187668
	pesos_i(25545) := b"1111111111111111_1111111111111111_1111111100111011_1011011000011100"; -- -0.0029951269909063976
	pesos_i(25546) := b"1111111111111111_1111111111111111_1100110101001101_1010100010110000"; -- -0.1980337687719976
	pesos_i(25547) := b"1111111111111111_1111111111111111_1101111110010010_1111001010110011"; -- -0.12666400085390697
	pesos_i(25548) := b"0000000000000000_0000000000000000_0010110110010101_1010101010101000"; -- 0.17806498135988458
	pesos_i(25549) := b"0000000000000000_0000000000000000_0001000011110011_1001010100000010"; -- 0.06621676735702052
	pesos_i(25550) := b"1111111111111111_1111111111111111_1111000101101010_1100100001110000"; -- -0.05696437141488513
	pesos_i(25551) := b"0000000000000000_0000000000000000_0001010101111101_1000101100100000"; -- 0.08394689112416416
	pesos_i(25552) := b"0000000000000000_0000000000000000_0001101100010000_0000011110011000"; -- 0.10571334336264353
	pesos_i(25553) := b"1111111111111111_1111111111111111_1101101010001000_0000110111001000"; -- -0.14636148328907825
	pesos_i(25554) := b"0000000000000000_0000000000000000_0001111000100010_0011000000111011"; -- 0.11770917362184576
	pesos_i(25555) := b"0000000000000000_0000000000000000_0001011000101101_0101111101100101"; -- 0.08662983152385165
	pesos_i(25556) := b"1111111111111111_1111111111111111_1110110010111000_1010111100010000"; -- -0.07530694834398373
	pesos_i(25557) := b"1111111111111111_1111111111111111_1111001100100101_0001001010010000"; -- -0.05021556834521783
	pesos_i(25558) := b"0000000000000000_0000000000000000_0001100011010111_1011011101011101"; -- 0.0970415690563529
	pesos_i(25559) := b"1111111111111111_1111111111111111_1111111011111001_0100101011001100"; -- -0.0040086032860780375
	pesos_i(25560) := b"1111111111111111_1111111111111111_1101011101100111_1010110011100010"; -- -0.15857429009100654
	pesos_i(25561) := b"1111111111111111_1111111111111111_1111101111110010_0011010110000000"; -- -0.015835434154369544
	pesos_i(25562) := b"0000000000000000_0000000000000000_0001011011011101_0000000001110010"; -- 0.08930971882518983
	pesos_i(25563) := b"1111111111111111_1111111111111111_1110111111111011_1010101100000010"; -- -0.06256610118025834
	pesos_i(25564) := b"0000000000000000_0000000000000000_0000000100010000_1100011010010010"; -- 0.00416222627239941
	pesos_i(25565) := b"1111111111111111_1111111111111111_1110011010111110_0100000100110111"; -- -0.09865944288482723
	pesos_i(25566) := b"0000000000000000_0000000000000000_0010100010010111_1100010011111011"; -- 0.15856581805392098
	pesos_i(25567) := b"0000000000000000_0000000000000000_0010000011011101_1100010110100011"; -- 0.12838397244592362
	pesos_i(25568) := b"1111111111111111_1111111111111111_1110111111001000_0010110001000011"; -- -0.06335185407613424
	pesos_i(25569) := b"0000000000000000_0000000000000000_0010101100111101_1110110111000011"; -- 0.16891370788566717
	pesos_i(25570) := b"0000000000000000_0000000000000000_0001101111000110_1100001000110111"; -- 0.10850156639069733
	pesos_i(25571) := b"1111111111111111_1111111111111111_1110110001000101_0010110001100110"; -- -0.07706949717330291
	pesos_i(25572) := b"0000000000000000_0000000000000000_0001110110000001_0001110001011011"; -- 0.115251323972055
	pesos_i(25573) := b"0000000000000000_0000000000000000_0001101001000010_1110010000111100"; -- 0.1025831837921749
	pesos_i(25574) := b"1111111111111111_1111111111111111_1110000011100101_1011110111011110"; -- -0.12149442040711804
	pesos_i(25575) := b"0000000000000000_0000000000000000_0000101101010110_1000000110111111"; -- 0.04428873939103827
	pesos_i(25576) := b"0000000000000000_0000000000000000_0001100111101100_1000100010001101"; -- 0.10126546322477221
	pesos_i(25577) := b"1111111111111111_1111111111111111_1110110000111110_1111110101011110"; -- -0.07716385323482976
	pesos_i(25578) := b"1111111111111111_1111111111111111_1101100000010111_1101000000111101"; -- -0.15588663591061527
	pesos_i(25579) := b"0000000000000000_0000000000000000_0000100100001001_1110100100111100"; -- 0.035307481033865926
	pesos_i(25580) := b"1111111111111111_1111111111111111_1110100110000110_1111110011001111"; -- -0.08778400360101482
	pesos_i(25581) := b"0000000000000000_0000000000000000_0010000110100010_0111011100111100"; -- 0.1313852807150036
	pesos_i(25582) := b"0000000000000000_0000000000000000_0001000010110011_0101100100100010"; -- 0.06523663607801426
	pesos_i(25583) := b"0000000000000000_0000000000000000_0001001101010100_0110110110110000"; -- 0.07550702607237186
	pesos_i(25584) := b"1111111111111111_1111111111111111_1111101001110001_1100011100010010"; -- -0.02170139124825362
	pesos_i(25585) := b"0000000000000000_0000000000000000_0010010101110000_1111100010011101"; -- 0.14625505294569627
	pesos_i(25586) := b"1111111111111111_1111111111111111_1101100011100101_1110010101011111"; -- -0.15274206571295315
	pesos_i(25587) := b"0000000000000000_0000000000000000_0010110110010100_0011001101101101"; -- 0.17804261606974517
	pesos_i(25588) := b"0000000000000000_0000000000000000_0010111001101000_1001110100101000"; -- 0.18128378125140981
	pesos_i(25589) := b"0000000000000000_0000000000000000_0010010001111011_0110100011001111"; -- 0.14250807820802108
	pesos_i(25590) := b"1111111111111111_1111111111111111_1101100000110010_1100001110001010"; -- -0.1554754054468213
	pesos_i(25591) := b"1111111111111111_1111111111111111_1110101010110111_0001100011001001"; -- -0.08314366418674816
	pesos_i(25592) := b"0000000000000000_0000000000000000_0011010000101011_0011011010000000"; -- 0.20378437644670563
	pesos_i(25593) := b"0000000000000000_0000000000000000_0000000111101100_1001011110011110"; -- 0.007516361226439719
	pesos_i(25594) := b"1111111111111111_1111111111111111_1110110100000100_0111100111001101"; -- -0.07415045498401851
	pesos_i(25595) := b"1111111111111111_1111111111111111_1101110111001000_0100111001001100"; -- -0.13366232540757486
	pesos_i(25596) := b"1111111111111111_1111111111111111_1101011000000110_1001110000011011"; -- -0.16396164262296614
	pesos_i(25597) := b"1111111111111111_1111111111111111_1111101010011100_0011111100011000"; -- -0.02105336831540282
	pesos_i(25598) := b"0000000000000000_0000000000000000_0011000110001100_0111010100000101"; -- 0.19354945529164094
	pesos_i(25599) := b"0000000000000000_0000000000000000_0001110111000100_0001101001010000"; -- 0.1162735409801205
	pesos_i(25600) := b"0000000000000000_0000000000000000_0001110010010100_0001110110100101"; -- 0.11163506769793773
	pesos_i(25601) := b"1111111111111111_1111111111111111_1110011111010010_1101100111101010"; -- -0.09443891559485142
	pesos_i(25602) := b"1111111111111111_1111111111111111_1100111011010110_1001000100101110"; -- -0.19203846564486882
	pesos_i(25603) := b"0000000000000000_0000000000000000_0001111000011001_1110000111100010"; -- 0.11758243341493213
	pesos_i(25604) := b"1111111111111111_1111111111111111_1111000011100101_1100001101011110"; -- -0.05899409242430381
	pesos_i(25605) := b"0000000000000000_0000000000000000_0010000011110011_1101000000001101"; -- 0.1287202864425659
	pesos_i(25606) := b"1111111111111111_1111111111111111_1111011011111000_1100010110110000"; -- -0.03526653728945291
	pesos_i(25607) := b"0000000000000000_0000000000000000_0010110111010110_1001111101100010"; -- 0.17905613087221878
	pesos_i(25608) := b"1111111111111111_1111111111111111_1110111000000010_1100010001110110"; -- -0.07027027232295406
	pesos_i(25609) := b"0000000000000000_0000000000000000_0000000001000110_0011100100010000"; -- 0.0010715163092965732
	pesos_i(25610) := b"1111111111111111_1111111111111111_1110011000110111_1101011101011001"; -- -0.10071043088331517
	pesos_i(25611) := b"0000000000000000_0000000000000000_0010111110001001_1110001110010100"; -- 0.1856977688351927
	pesos_i(25612) := b"1111111111111111_1111111111111111_1110110011111101_1010010000111111"; -- -0.07425473644793192
	pesos_i(25613) := b"1111111111111111_1111111111111111_1111100110010111_0101111001001010"; -- -0.025034052760380985
	pesos_i(25614) := b"1111111111111111_1111111111111111_1101011011110011_1011000010001101"; -- -0.1603440910752311
	pesos_i(25615) := b"0000000000000000_0000000000000000_0000001000110101_0011010111101110"; -- 0.008624430263436024
	pesos_i(25616) := b"0000000000000000_0000000000000000_0010100101011110_1111110110111101"; -- 0.16160570021560933
	pesos_i(25617) := b"1111111111111111_1111111111111111_1110010000100100_0100100100011110"; -- -0.10882132541495305
	pesos_i(25618) := b"0000000000000000_0000000000000000_0001100101000111_1011110111000011"; -- 0.09875093475490329
	pesos_i(25619) := b"1111111111111111_1111111111111111_1110010000000001_0101101010111010"; -- -0.10935433351920425
	pesos_i(25620) := b"0000000000000000_0000000000000000_0001000100100110_1001110001110001"; -- 0.06699540863120557
	pesos_i(25621) := b"0000000000000000_0000000000000000_0010011100010110_0001010000011101"; -- 0.15268064210759505
	pesos_i(25622) := b"0000000000000000_0000000000000000_0010100110000011_0111011000011111"; -- 0.16216219189281114
	pesos_i(25623) := b"1111111111111111_1111111111111111_1110110111100001_0011100111100100"; -- -0.07078207189920603
	pesos_i(25624) := b"0000000000000000_0000000000000000_0000010101111010_1001000010000000"; -- 0.021401435207051074
	pesos_i(25625) := b"0000000000000000_0000000000000000_0010101111110000_0111110011100010"; -- 0.17163830295830984
	pesos_i(25626) := b"0000000000000000_0000000000000000_0010001101100000_0110101011101001"; -- 0.13818996610428574
	pesos_i(25627) := b"1111111111111111_1111111111111111_1110000010100010_0101101010101010"; -- -0.12252267215644118
	pesos_i(25628) := b"1111111111111111_1111111111111111_1100111111011111_0010111100110011"; -- -0.18800072675878585
	pesos_i(25629) := b"0000000000000000_0000000000000000_0000100010100011_0001111000001000"; -- 0.03373897254918937
	pesos_i(25630) := b"1111111111111111_1111111111111111_1111100101001001_0110101100001110"; -- -0.026223477499163015
	pesos_i(25631) := b"1111111111111111_1111111111111111_1101111010110110_1000000000001101"; -- -0.13002776806147015
	pesos_i(25632) := b"1111111111111111_1111111111111111_1111011000011010_0001000010000001"; -- -0.03866478779399988
	pesos_i(25633) := b"1111111111111111_1111111111111111_1111001100001101_0001100101100011"; -- -0.05058137246486449
	pesos_i(25634) := b"1111111111111111_1111111111111111_1111000111010010_1100011001111110"; -- -0.05537757319893642
	pesos_i(25635) := b"0000000000000000_0000000000000000_0000001000010011_0111110001010011"; -- 0.008109827248122797
	pesos_i(25636) := b"0000000000000000_0000000000000000_0001100111111101_1001010101111001"; -- 0.10152563285155011
	pesos_i(25637) := b"1111111111111111_1111111111111111_1101101000011111_0001100111100111"; -- -0.14796293362671467
	pesos_i(25638) := b"1111111111111111_1111111111111111_1111000101111010_0100000010011010"; -- -0.056728327187967144
	pesos_i(25639) := b"1111111111111111_1111111111111111_1111001000011101_1111100110000010"; -- -0.05423012325185647
	pesos_i(25640) := b"0000000000000000_0000000000000000_0000100001001111_0110000111000111"; -- 0.032461272224952445
	pesos_i(25641) := b"0000000000000000_0000000000000000_0000100101101110_1100010111010111"; -- 0.03684650900508226
	pesos_i(25642) := b"0000000000000000_0000000000000000_0000100011000001_1111101100110100"; -- 0.034209919223133434
	pesos_i(25643) := b"0000000000000000_0000000000000000_0010101011110010_1001000101000110"; -- 0.16776378586452
	pesos_i(25644) := b"1111111111111111_1111111111111111_1111111001001011_0011100111001111"; -- -0.006664645103138286
	pesos_i(25645) := b"1111111111111111_1111111111111111_1111100100100001_0111001001010000"; -- -0.026833396478956172
	pesos_i(25646) := b"1111111111111111_1111111111111111_1101110000001110_1010001001100110"; -- -0.14040169718960752
	pesos_i(25647) := b"1111111111111111_1111111111111111_1101011101011001_1111101000100000"; -- -0.15878330906215624
	pesos_i(25648) := b"1111111111111111_1111111111111111_1100110011100000_1100110100111011"; -- -0.1996947985326529
	pesos_i(25649) := b"1111111111111111_1111111111111111_1110110101000110_0101001111001101"; -- -0.0731456397472757
	pesos_i(25650) := b"1111111111111111_1111111111111111_1101101010000100_1011010100001110"; -- -0.14641254808330068
	pesos_i(25651) := b"1111111111111111_1111111111111111_1110111011000100_1001000010110010"; -- -0.06731315272186271
	pesos_i(25652) := b"1111111111111111_1111111111111111_1100110111001101_1000101111101001"; -- -0.196082359033602
	pesos_i(25653) := b"0000000000000000_0000000000000000_0000110000101000_1000000000010111"; -- 0.04749298621961144
	pesos_i(25654) := b"1111111111111111_1111111111111111_1111001001101000_1011100000101000"; -- -0.05308960926266971
	pesos_i(25655) := b"1111111111111111_1111111111111111_1101101011011001_0010101110011110"; -- -0.1451237429528409
	pesos_i(25656) := b"1111111111111111_1111111111111111_1101001111000111_1000001100111010"; -- -0.1727369293441938
	pesos_i(25657) := b"1111111111111111_1111111111111111_1111100000110010_1011100101100111"; -- -0.030476009792143665
	pesos_i(25658) := b"1111111111111111_1111111111111111_1110101010111101_0101011011111111"; -- -0.08304840347106489
	pesos_i(25659) := b"1111111111111111_1111111111111111_1110010011100101_1001110000100100"; -- -0.1058714306974584
	pesos_i(25660) := b"1111111111111111_1111111111111111_1111100110110110_0110000110100101"; -- -0.024560830247890787
	pesos_i(25661) := b"1111111111111111_1111111111111111_1110011000100111_0010010010001010"; -- -0.10096522929990584
	pesos_i(25662) := b"1111111111111111_1111111111111111_1100111010011010_0010000110110001"; -- -0.1929606382546465
	pesos_i(25663) := b"1111111111111111_1111111111111111_1110001010010010_1101000000011000"; -- -0.11494731348803502
	pesos_i(25664) := b"1111111111111111_1111111111111111_1111001100101110_1000000100001101"; -- -0.05007165368277707
	pesos_i(25665) := b"1111111111111111_1111111111111111_1101010101101100_1001011111010110"; -- -0.16631175053947014
	pesos_i(25666) := b"0000000000000000_0000000000000000_0001101011010011_1100110011000110"; -- 0.10479431002215016
	pesos_i(25667) := b"0000000000000000_0000000000000000_0010100010010010_0000000110010100"; -- 0.1584778771940635
	pesos_i(25668) := b"0000000000000000_0000000000000000_0000001011100100_1010111010100010"; -- 0.011301912861851284
	pesos_i(25669) := b"1111111111111111_1111111111111111_1101011101100100_0111000101100111"; -- -0.15862361172393896
	pesos_i(25670) := b"1111111111111111_1111111111111111_1110100110101100_0010100110110000"; -- -0.08721675340254399
	pesos_i(25671) := b"0000000000000000_0000000000000000_0001111101111010_1000100100100011"; -- 0.12296349620010072
	pesos_i(25672) := b"1111111111111111_1111111111111111_1110010101000001_0101011000010100"; -- -0.10447179808294438
	pesos_i(25673) := b"0000000000000000_0000000000000000_0010000001001111_0011010001110010"; -- 0.12620857024111412
	pesos_i(25674) := b"0000000000000000_0000000000000000_0010000001101010_1110010101000111"; -- 0.1266310977043791
	pesos_i(25675) := b"0000000000000000_0000000000000000_0001100000100010_0110000001100111"; -- 0.09427454492389277
	pesos_i(25676) := b"0000000000000000_0000000000000000_0010000101010100_1010111010010101"; -- 0.13019839423328577
	pesos_i(25677) := b"1111111111111111_1111111111111111_1111010101010110_0100111011111011"; -- -0.04165178654945914
	pesos_i(25678) := b"0000000000000000_0000000000000000_0010100101000000_1001110011010011"; -- 0.16114216001190612
	pesos_i(25679) := b"1111111111111111_1111111111111111_1110011000001000_1001100110000100"; -- -0.10143127945660764
	pesos_i(25680) := b"0000000000000000_0000000000000000_0010101100101001_0011011000000100"; -- 0.16859757999975927
	pesos_i(25681) := b"1111111111111111_1111111111111111_1111101101000110_0000101011111111"; -- -0.018462479359376154
	pesos_i(25682) := b"1111111111111111_1111111111111111_1110100101000101_1110010001000110"; -- -0.08877728739138573
	pesos_i(25683) := b"0000000000000000_0000000000000000_0001111110111010_0011110010111000"; -- 0.12393550380696741
	pesos_i(25684) := b"1111111111111111_1111111111111111_1101001100100111_1011011011100100"; -- -0.17517525611394405
	pesos_i(25685) := b"1111111111111111_1111111111111111_1110110101110110_1011101110001001"; -- -0.07240703484376577
	pesos_i(25686) := b"1111111111111111_1111111111111111_1100111100111010_1000110111110111"; -- -0.19051277839615965
	pesos_i(25687) := b"0000000000000000_0000000000000000_0001001110100000_0110101011100010"; -- 0.0766665270674339
	pesos_i(25688) := b"0000000000000000_0000000000000000_0011010111101111_1010110110110000"; -- 0.21068845308855638
	pesos_i(25689) := b"0000000000000000_0000000000000000_0010000111010101_0100110110100010"; -- 0.13216099927301128
	pesos_i(25690) := b"0000000000000000_0000000000000000_0010110101000011_0111010000001000"; -- 0.17681050489745323
	pesos_i(25691) := b"1111111111111111_1111111111111111_1101110001000001_1001001100001010"; -- -0.13962441439275847
	pesos_i(25692) := b"0000000000000000_0000000000000000_0010101011001011_1010111101011011"; -- 0.1671704861828306
	pesos_i(25693) := b"0000000000000000_0000000000000000_0011000110111000_1011100000001011"; -- 0.19422483694713255
	pesos_i(25694) := b"0000000000000000_0000000000000000_0010000110111110_0001110001101101"; -- 0.13180711425293984
	pesos_i(25695) := b"0000000000000000_0000000000000000_0010110001101101_1011111110000101"; -- 0.17354962349906533
	pesos_i(25696) := b"1111111111111111_1111111111111111_1101101001101011_0100101010100011"; -- -0.14680036079702483
	pesos_i(25697) := b"1111111111111111_1111111111111111_1101001111110011_0101010010110101"; -- -0.17206831535399966
	pesos_i(25698) := b"0000000000000000_0000000000000000_0001100011000100_0101001101100111"; -- 0.0967456937558763
	pesos_i(25699) := b"1111111111111111_1111111111111111_1101011011010111_0100001010101010"; -- -0.16077788697044149
	pesos_i(25700) := b"0000000000000000_0000000000000000_0010100111000010_1101111010010011"; -- 0.16312972160178268
	pesos_i(25701) := b"0000000000000000_0000000000000000_0000110001001011_0101000111001001"; -- 0.04802428392649185
	pesos_i(25702) := b"1111111111111111_1111111111111111_1110111111000000_1011110101110101"; -- -0.06346527005706433
	pesos_i(25703) := b"1111111111111111_1111111111111111_1101101011001001_0001010110001101"; -- -0.1453691988993056
	pesos_i(25704) := b"0000000000000000_0000000000000000_0001100001101100_1011111000111100"; -- 0.09540928817632185
	pesos_i(25705) := b"1111111111111111_1111111111111111_1111100010111110_1001101001011101"; -- -0.028341629217456702
	pesos_i(25706) := b"1111111111111111_1111111111111111_1101001000000101_0111011110001101"; -- -0.1796040802490484
	pesos_i(25707) := b"1111111111111111_1111111111111111_1111101000100001_0110000000100011"; -- -0.022928229784755127
	pesos_i(25708) := b"0000000000000000_0000000000000000_0010001001011101_1011000100100100"; -- 0.13424212589933135
	pesos_i(25709) := b"0000000000000000_0000000000000000_0010101110110010_1111000100101010"; -- 0.17069918902081163
	pesos_i(25710) := b"1111111111111111_1111111111111111_1100111111010010_1010010110010001"; -- -0.1881920357262386
	pesos_i(25711) := b"1111111111111111_1111111111111111_1111111100110000_1011010001010101"; -- -0.0031630795067725996
	pesos_i(25712) := b"1111111111111111_1111111111111111_1110101000101001_1111110010101001"; -- -0.08529682984764585
	pesos_i(25713) := b"0000000000000000_0000000000000000_0000000001100001_1101101101100100"; -- 0.0014931791962061334
	pesos_i(25714) := b"0000000000000000_0000000000000000_0001001001000111_0010001001111111"; -- 0.07139793012605919
	pesos_i(25715) := b"0000000000000000_0000000000000000_0000010001001101_0000101110101100"; -- 0.016800622511983346
	pesos_i(25716) := b"1111111111111111_1111111111111111_1111101100011010_1101001001000100"; -- -0.01912198866136144
	pesos_i(25717) := b"1111111111111111_1111111111111111_1110100011001110_0001110110010010"; -- -0.09060492690750051
	pesos_i(25718) := b"0000000000000000_0000000000000000_0001111011101001_1110110100100100"; -- 0.12075693263663198
	pesos_i(25719) := b"0000000000000000_0000000000000000_0000100110100101_0011000011001111"; -- 0.03767685941352613
	pesos_i(25720) := b"1111111111111111_1111111111111111_1110110100001110_1011111101101000"; -- -0.07399371832247595
	pesos_i(25721) := b"1111111111111111_1111111111111111_1101101011110000_0010010111011011"; -- -0.14477313430465644
	pesos_i(25722) := b"0000000000000000_0000000000000000_0000010100110001_0001000010101011"; -- 0.020279924177337795
	pesos_i(25723) := b"1111111111111111_1111111111111111_1101110110011010_1000100000011000"; -- -0.1343607846347183
	pesos_i(25724) := b"1111111111111111_1111111111111111_1101100111000100_0001001101010101"; -- -0.14935187501514047
	pesos_i(25725) := b"0000000000000000_0000000000000000_0010000010100100_0111000110011001"; -- 0.12750921225508857
	pesos_i(25726) := b"0000000000000000_0000000000000000_0000111010111111_0101000000000000"; -- 0.05760669699794512
	pesos_i(25727) := b"1111111111111111_1111111111111111_1111110001001110_0111001001001001"; -- -0.014428002565069138
	pesos_i(25728) := b"1111111111111111_1111111111111111_1101001010010000_1101010101001001"; -- -0.17747752148743443
	pesos_i(25729) := b"1111111111111111_1111111111111111_1111010100101100_0010110001111001"; -- -0.04229471257567921
	pesos_i(25730) := b"0000000000000000_0000000000000000_0011000101111100_0110011011010101"; -- 0.19330446901666118
	pesos_i(25731) := b"0000000000000000_0000000000000000_0010010100011000_0011101100000100"; -- 0.1449009784293243
	pesos_i(25732) := b"1111111111111111_1111111111111111_1101100111000001_1110011000000110"; -- -0.1493850931417688
	pesos_i(25733) := b"0000000000000000_0000000000000000_0010111110010111_0001000101010010"; -- 0.18589885957464578
	pesos_i(25734) := b"1111111111111111_1111111111111111_1111000001110010_1010100110001101"; -- -0.06075039204207891
	pesos_i(25735) := b"1111111111111111_1111111111111111_1110010011001110_1010110001000111"; -- -0.10622142092162769
	pesos_i(25736) := b"0000000000000000_0000000000000000_0010111011100101_1001110000010011"; -- 0.18319106535672772
	pesos_i(25737) := b"0000000000000000_0000000000000000_0010111000000010_1101001000001010"; -- 0.17973053686963592
	pesos_i(25738) := b"1111111111111111_1111111111111111_1110101010110000_1000111101111010"; -- -0.08324340123116217
	pesos_i(25739) := b"0000000000000000_0000000000000000_0001010101001111_1110100111011111"; -- 0.08325063420149312
	pesos_i(25740) := b"1111111111111111_1111111111111111_1101000010000101_1101001111011111"; -- -0.18545795249170846
	pesos_i(25741) := b"1111111111111111_1111111111111111_1110011010101010_0010100000010101"; -- -0.09896611686359046
	pesos_i(25742) := b"0000000000000000_0000000000000000_0001100110110001_0011101110001000"; -- 0.10036060410439501
	pesos_i(25743) := b"1111111111111111_1111111111111111_1110110101010000_0010011101100110"; -- -0.0729956985635368
	pesos_i(25744) := b"1111111111111111_1111111111111111_1111001111001100_0010011111001000"; -- -0.04766608587875564
	pesos_i(25745) := b"0000000000000000_0000000000000000_0001011010010110_0100101111010000"; -- 0.08823083717444995
	pesos_i(25746) := b"0000000000000000_0000000000000000_0001111111010100_0111111111101110"; -- 0.12433623854083803
	pesos_i(25747) := b"0000000000000000_0000000000000000_0000001110111010_1010010101010110"; -- 0.014566739441863336
	pesos_i(25748) := b"0000000000000000_0000000000000000_0010001000101011_1011011011010011"; -- 0.13347952511637406
	pesos_i(25749) := b"0000000000000000_0000000000000000_0010100110000100_0100010000100110"; -- 0.16217447203443544
	pesos_i(25750) := b"1111111111111111_1111111111111111_1111100100010001_1100000000110010"; -- -0.027072894797557916
	pesos_i(25751) := b"1111111111111111_1111111111111111_1111000000111010_0111111001111101"; -- -0.06160745100314261
	pesos_i(25752) := b"1111111111111111_1111111111111111_1101000111100011_0100011110111000"; -- -0.18012573009656713
	pesos_i(25753) := b"1111111111111111_1111111111111111_1110100110101011_1101000000011010"; -- -0.08722209324336061
	pesos_i(25754) := b"1111111111111111_1111111111111111_1110001111101010_1100010000000100"; -- -0.1096990098345109
	pesos_i(25755) := b"1111111111111111_1111111111111111_1101110010101110_1001001010011010"; -- -0.1379612325236588
	pesos_i(25756) := b"1111111111111111_1111111111111111_1111111111010011_1000011110001011"; -- -0.0006785664634390381
	pesos_i(25757) := b"1111111111111111_1111111111111111_1111011000100001_1011101001000001"; -- -0.038547858258191375
	pesos_i(25758) := b"1111111111111111_1111111111111111_1111100000100011_1100010101011101"; -- -0.030704178648003785
	pesos_i(25759) := b"1111111111111111_1111111111111111_1101111100000101_1001101111101111"; -- -0.12882066170268816
	pesos_i(25760) := b"0000000000000000_0000000000000000_0000100111100001_0110000111101001"; -- 0.03859531347671728
	pesos_i(25761) := b"0000000000000000_0000000000000000_0001010011111010_0011100110100000"; -- 0.0819431319098511
	pesos_i(25762) := b"0000000000000000_0000000000000000_0000111100000111_0001000001010001"; -- 0.05870153403351829
	pesos_i(25763) := b"1111111111111111_1111111111111111_1110010000010001_1110001111111011"; -- -0.10910201197612397
	pesos_i(25764) := b"0000000000000000_0000000000000000_0010101100101001_0110001001111001"; -- 0.1686002298091767
	pesos_i(25765) := b"1111111111111111_1111111111111111_1101100001011000_1101101010111011"; -- -0.15489418917838835
	pesos_i(25766) := b"1111111111111111_1111111111111111_1110101001011010_1110011011111001"; -- -0.0845504420341525
	pesos_i(25767) := b"1111111111111111_1111111111111111_1111100001010011_1111101111110000"; -- -0.029968503860020663
	pesos_i(25768) := b"1111111111111111_1111111111111111_1111011011101101_0110100011101011"; -- -0.035439913307330435
	pesos_i(25769) := b"0000000000000000_0000000000000000_0000000111000111_1000000100110110"; -- 0.006950450620508238
	pesos_i(25770) := b"0000000000000000_0000000000000000_0000110011110101_1000110110101110"; -- 0.050621848113833814
	pesos_i(25771) := b"1111111111111111_1111111111111111_1111011001010001_0000001100010101"; -- -0.03782635445211416
	pesos_i(25772) := b"1111111111111111_1111111111111111_1101111101001001_0000101001001110"; -- -0.12779174424242248
	pesos_i(25773) := b"1111111111111111_1111111111111111_1111100100000100_1101000111001010"; -- -0.027270210446027704
	pesos_i(25774) := b"0000000000000000_0000000000000000_0010011111110111_0001010101010010"; -- 0.1561139416913305
	pesos_i(25775) := b"1111111111111111_1111111111111111_1111001000001110_0010011011111010"; -- -0.054471553760772125
	pesos_i(25776) := b"0000000000000000_0000000000000000_0000110101101100_0000000101111010"; -- 0.05242928722040674
	pesos_i(25777) := b"0000000000000000_0000000000000000_0010100111110110_0100011110000111"; -- 0.1639141753724438
	pesos_i(25778) := b"0000000000000000_0000000000000000_0001011001100100_1101110000100111"; -- 0.08747650108785203
	pesos_i(25779) := b"0000000000000000_0000000000000000_0011000011011010_1110001100100001"; -- 0.19083995406860269
	pesos_i(25780) := b"0000000000000000_0000000000000000_0000000001100010_0000100110111010"; -- 0.0014959410869569013
	pesos_i(25781) := b"1111111111111111_1111111111111111_1111000111100000_0011000101000100"; -- -0.05517284481298385
	pesos_i(25782) := b"1111111111111111_1111111111111111_1110111101011101_1001000001101010"; -- -0.06497857484575865
	pesos_i(25783) := b"1111111111111111_1111111111111111_1111111110001010_1010000101100110"; -- -0.0017909170680528697
	pesos_i(25784) := b"0000000000000000_0000000000000000_0000111100100111_1101011111100111"; -- 0.05920171144922516
	pesos_i(25785) := b"0000000000000000_0000000000000000_0000011110011010_0100000001111100"; -- 0.02969744710379995
	pesos_i(25786) := b"1111111111111111_1111111111111111_1100111000010000_0101100001101101"; -- -0.19506308871951206
	pesos_i(25787) := b"1111111111111111_1111111111111111_1110100101100111_0101010101110000"; -- -0.08826700224498416
	pesos_i(25788) := b"1111111111111111_1111111111111111_1110101100000100_0110011111100011"; -- -0.08196402272106142
	pesos_i(25789) := b"1111111111111111_1111111111111111_1101010100011101_0101000010011101"; -- -0.16752144017820822
	pesos_i(25790) := b"0000000000000000_0000000000000000_0010110111100101_0101000000111101"; -- 0.17928029517874935
	pesos_i(25791) := b"0000000000000000_0000000000000000_0000010010101110_1100111010010010"; -- 0.018292341939951877
	pesos_i(25792) := b"1111111111111111_1111111111111111_1101101010101011_0001001010010111"; -- -0.14582713911838605
	pesos_i(25793) := b"0000000000000000_0000000000000000_0011010111110011_1111011101111100"; -- 0.21075388707535117
	pesos_i(25794) := b"0000000000000000_0000000000000000_0011001001100000_1010001010011001"; -- 0.19678703528765767
	pesos_i(25795) := b"1111111111111111_1111111111111111_1111000101010000_0111110000111001"; -- -0.05736564255606066
	pesos_i(25796) := b"0000000000000000_0000000000000000_0000000010110010_1110100101001001"; -- 0.0027299692530645923
	pesos_i(25797) := b"0000000000000000_0000000000000000_0010001000111110_1101101111111111"; -- 0.13377165771215993
	pesos_i(25798) := b"1111111111111111_1111111111111111_1111010011011110_0001000010101101"; -- -0.04348655497635389
	pesos_i(25799) := b"1111111111111111_1111111111111111_1111101110100100_1000011011100101"; -- -0.01702076827265549
	pesos_i(25800) := b"0000000000000000_0000000000000000_0001001100101001_1000010101111101"; -- 0.07485231681044241
	pesos_i(25801) := b"1111111111111111_1111111111111111_1101001001110010_1110000110111101"; -- -0.17793454299172687
	pesos_i(25802) := b"0000000000000000_0000000000000000_0010101101001010_1011101000100001"; -- 0.16910899458585688
	pesos_i(25803) := b"1111111111111111_1111111111111111_1101000011111000_0000110010110110"; -- -0.18371506269111335
	pesos_i(25804) := b"1111111111111111_1111111111111111_1111010110111011_1100101011101100"; -- -0.040103261299466626
	pesos_i(25805) := b"1111111111111111_1111111111111111_1100111110101111_0100100110111001"; -- -0.18873156778226038
	pesos_i(25806) := b"1111111111111111_1111111111111111_1111000011101100_0001100010100000"; -- -0.05889745808915534
	pesos_i(25807) := b"1111111111111111_1111111111111111_1110101001001111_1011001111100001"; -- -0.08472133400463394
	pesos_i(25808) := b"0000000000000000_0000000000000000_0001111101110010_0010010111101001"; -- 0.12283551157392775
	pesos_i(25809) := b"0000000000000000_0000000000000000_0001111001110100_0011000110111001"; -- 0.11896048323911587
	pesos_i(25810) := b"0000000000000000_0000000000000000_0010010101101011_0010000000001101"; -- 0.14616585088990192
	pesos_i(25811) := b"1111111111111111_1111111111111111_1101000000101011_0111111111111010"; -- -0.1868362441546267
	pesos_i(25812) := b"0000000000000000_0000000000000000_0010100001000101_1000010001101101"; -- 0.15731074974342923
	pesos_i(25813) := b"0000000000000000_0000000000000000_0001000011010110_0101101001010011"; -- 0.06577076460989076
	pesos_i(25814) := b"0000000000000000_0000000000000000_0011000001100111_0101000011010100"; -- 0.18907647298129746
	pesos_i(25815) := b"1111111111111111_1111111111111111_1111000001101000_1100110000111001"; -- -0.06090091342547663
	pesos_i(25816) := b"0000000000000000_0000000000000000_0010011110010111_1100000001000111"; -- 0.15465928775079976
	pesos_i(25817) := b"1111111111111111_1111111111111111_1110001101101111_1001000111000001"; -- -0.11157883685446175
	pesos_i(25818) := b"1111111111111111_1111111111111111_1110010000000011_0000110010101011"; -- -0.10932846844762602
	pesos_i(25819) := b"1111111111111111_1111111111111111_1110101001100010_1100011101111001"; -- -0.08443024917989568
	pesos_i(25820) := b"0000000000000000_0000000000000000_0011000111110001_1011001101100011"; -- 0.19509431040849037
	pesos_i(25821) := b"0000000000000000_0000000000000000_0001111011010110_1011111110010101"; -- 0.12046430013066761
	pesos_i(25822) := b"0000000000000000_0000000000000000_0010110010100010_0100111001100100"; -- 0.17435159630361366
	pesos_i(25823) := b"1111111111111111_1111111111111111_1111111101000110_1011111101110011"; -- -0.0028267235047466357
	pesos_i(25824) := b"0000000000000000_0000000000000000_0000010110010101_0010111011111001"; -- 0.021807609280346807
	pesos_i(25825) := b"1111111111111111_1111111111111111_1101010000111101_1100111110011001"; -- -0.17093184013956475
	pesos_i(25826) := b"1111111111111111_1111111111111111_1100110010000101_1111111010111101"; -- -0.20108039746954684
	pesos_i(25827) := b"0000000000000000_0000000000000000_0001010111011111_0010100010100010"; -- 0.0854363818290619
	pesos_i(25828) := b"1111111111111111_1111111111111111_1111100011001110_0011010101000111"; -- -0.028103513767619815
	pesos_i(25829) := b"1111111111111111_1111111111111111_1101100000100101_1011101111111010"; -- -0.15567422044353818
	pesos_i(25830) := b"1111111111111111_1111111111111111_1101001110010101_0110111111001001"; -- -0.1735010276198534
	pesos_i(25831) := b"1111111111111111_1111111111111111_1111110111000010_0110000001110010"; -- -0.008752796335551026
	pesos_i(25832) := b"1111111111111111_1111111111111111_1100111110010010_1001100101001110"; -- -0.18916932912254453
	pesos_i(25833) := b"1111111111111111_1111111111111111_1101111011110011_0010110100001110"; -- -0.12910192883730093
	pesos_i(25834) := b"0000000000000000_0000000000000000_0010110110001011_0011100100000011"; -- 0.1779056199531423
	pesos_i(25835) := b"1111111111111111_1111111111111111_1111000000110110_1101011111001101"; -- -0.06166316260499074
	pesos_i(25836) := b"1111111111111111_1111111111111111_1101010100100100_0100110010010011"; -- -0.16741486932235236
	pesos_i(25837) := b"0000000000000000_0000000000000000_0001101010100000_0011100111101000"; -- 0.10400735779695897
	pesos_i(25838) := b"1111111111111111_1111111111111111_1111100001000001_0001001011100001"; -- -0.030257053483140176
	pesos_i(25839) := b"1111111111111111_1111111111111111_1111100000100000_0100101100100101"; -- -0.030757239860935103
	pesos_i(25840) := b"0000000000000000_0000000000000000_0011000001100101_1011011101001011"; -- 0.18905206289580406
	pesos_i(25841) := b"1111111111111111_1111111111111111_1110111001111101_0001011111110011"; -- -0.06840372399026119
	pesos_i(25842) := b"0000000000000000_0000000000000000_0001000001110111_0001110100001110"; -- 0.0643175276203425
	pesos_i(25843) := b"1111111111111111_1111111111111111_1101100101010110_1011101010001100"; -- -0.1510203750995079
	pesos_i(25844) := b"0000000000000000_0000000000000000_0011010001111101_1000000100110111"; -- 0.2050400503740019
	pesos_i(25845) := b"1111111111111111_1111111111111111_1111101101101110_0010011100010011"; -- -0.017850454192226056
	pesos_i(25846) := b"0000000000000000_0000000000000000_0010011010011111_0010111101110010"; -- 0.15086647546328802
	pesos_i(25847) := b"0000000000000000_0000000000000000_0000001000110100_1010111110111011"; -- 0.008616431402592498
	pesos_i(25848) := b"1111111111111111_1111111111111111_1111011110100000_1101010001101101"; -- -0.0327021820959186
	pesos_i(25849) := b"0000000000000000_0000000000000000_0010101000011010_0110000111110010"; -- 0.164465066398313
	pesos_i(25850) := b"1111111111111111_1111111111111111_1111001001001110_0001101011010100"; -- -0.05349571540522816
	pesos_i(25851) := b"0000000000000000_0000000000000000_0010100100110111_1010101000111111"; -- 0.1610056308874582
	pesos_i(25852) := b"1111111111111111_1111111111111111_1110111111001011_1000100100110110"; -- -0.06330053736982076
	pesos_i(25853) := b"0000000000000000_0000000000000000_0001111000100011_1101101111100101"; -- 0.11773466431859199
	pesos_i(25854) := b"1111111111111111_1111111111111111_1101010010101111_1011111011111011"; -- -0.1691933285390344
	pesos_i(25855) := b"1111111111111111_1111111111111111_1101001000000100_0101111001011010"; -- -0.17962084107644202
    return pesos_i;
    end function;
end package body mnist_weights;
    