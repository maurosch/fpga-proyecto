
-- ARCHIVO AUTOGENERADO CON generate_weights_package.py

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.perceptron_package.perceptron_input;

package matrix_weights is
    function GetWeights(Dummy: natural)
    return perceptron_input;
end package matrix_weights;

package body matrix_weights is
    function GetWeights(Dummy: natural) return perceptron_input is
        variable pesos_i : perceptron_input(17 downto 0);
    begin
	pesos_i(0) := b"0000000000000000_0000000000000000_0001100110011001_1001100110011010"; -- 0.1
	pesos_i(1) := b"0000000000000000_0000000000000000_0011001100110011_0011001100110011"; -- 0.2
	pesos_i(2) := b"0000000000000000_0000000000000000_0100110011001100_1100110011001101"; -- 0.3
	pesos_i(3) := b"0000000000000000_0000000000000000_0110011001100110_0110011001100110"; -- 0.4
	pesos_i(4) := b"0000000000000000_0000000000000000_1000000000000000_0000000000000000"; -- 0.5
	pesos_i(5) := b"0000000000000000_0000000000000000_1001100110011001_1001100110011010"; -- 0.6
	pesos_i(6) := b"1111111111111111_1111111111111111_1110011001100110_0110011001100110"; -- -0.1
	pesos_i(7) := b"1111111111111111_1111111111111111_1100110011001100_1100110011001101"; -- -0.2
	pesos_i(8) := b"1111111111111111_1111111111111111_1011001100110011_0011001100110011"; -- -0.3
	pesos_i(9) := b"1111111111111111_1111111111111111_1001100110011001_1001100110011010"; -- -0.4
	pesos_i(10) := b"1111111111111111_1111111111111111_1000000000000000_0000000000000000"; -- -0.5
	pesos_i(11) := b"1111111111111111_1111111111111111_0110011001100110_0110011001100110"; -- -0.6
	pesos_i(12) := b"1111111111111111_1111111111111111_0100110011001100_1100110011001101"; -- -0.7
	pesos_i(13) := b"1111111111111111_1111111111111111_0011001100110011_0011001100110011"; -- -0.8
	pesos_i(14) := b"1111111111111111_1111111111111111_0001100110011001_1001100110011010"; -- -0.9
	pesos_i(15) := b"0000000000000000_0000000000000001_0000000000000000_0000000000000000"; -- 1
	pesos_i(16) := b"0000000000000000_0000000000000010_0000000000000000_0000000000000000"; -- 2
	pesos_i(17) := b"0000000000000000_0000000000000011_0000000000000000_0000000000000000"; -- 3

    return pesos_i;
    end function;
end package body matrix_weights;
    