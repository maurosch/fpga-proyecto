
-- ARCHIVO AUTOGENERADO CON generate_weights_package.py

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.perceptron_package.perceptron_input;

package mnist_weights is
    function GetWeights(Dummy: natural)
    return perceptron_input;
end package mnist_weights;

package body mnist_weights is
    function GetWeights(Dummy: natural) return perceptron_input is
        variable pesos_i : perceptron_input(25855 downto 0);
    begin
	pesos_i(0) := b"1111111111111111_1111111111111111_1101100001100010_1010110111001110"; -- -0.15474427913013053
	pesos_i(1) := b"0000000000000000_0000000000000000_0010010101000011_1001111111000011"; -- 0.1455631113895911
	pesos_i(2) := b"1111111111111111_1111111111111111_1110010101100010_1110110000100011"; -- -0.10395931393041476
	pesos_i(3) := b"1111111111111111_1111111111111111_1111101100010111_1111111111001110"; -- -0.01916505075719053
	pesos_i(4) := b"1111111111111111_1111111111111111_1111001101110101_0101101000011110"; -- -0.048990600208625286
	pesos_i(5) := b"0000000000000000_0000000000000000_0000110110101100_0101011110111101"; -- 0.05341099141670477
	pesos_i(6) := b"0000000000000000_0000000000000000_0000001010110000_1111100000001110"; -- 0.010512831982210319
	pesos_i(7) := b"0000000000000000_0000000000000000_0001011001010011_0101111001111001"; -- 0.08720961039878103
	pesos_i(8) := b"1111111111111111_1111111111111111_1111000101011111_1001101001000110"; -- -0.05713496963480013
	pesos_i(9) := b"1111111111111111_1111111111111111_1110011100001010_1011001010111001"; -- -0.09749300952349603
	pesos_i(10) := b"1111111111111111_1111111111111111_1110101100100111_1111000110110000"; -- -0.08142175143561234
	pesos_i(11) := b"1111111111111111_1111111111111111_1111011100010001_0000011100111100"; -- -0.034896419495004036
	pesos_i(12) := b"0000000000000000_0000000000000000_0010010001000000_0101111011011001"; -- 0.14160721577988644
	pesos_i(13) := b"1111111111111111_1111111111111111_1101001101010001_1010000010010111"; -- -0.17453571626754683
	pesos_i(14) := b"0000000000000000_0000000000000000_0010100111011100_1110101110000000"; -- 0.16352722044597853
	pesos_i(15) := b"0000000000000000_0000000000000000_0001110111100010_0001100110011111"; -- 0.1167312635669969
	pesos_i(16) := b"0000000000000000_0000000000000000_0000101001101100_1011100100000110"; -- 0.04072147738661819
	pesos_i(17) := b"1111111111111111_1111111111111111_1111100111000001_0110101111000001"; -- -0.024392381017043475
	pesos_i(18) := b"1111111111111111_1111111111111111_1101111100101010_0101111010111010"; -- -0.12825973463903245
	pesos_i(19) := b"1111111111111111_1111111111111111_1101111010111100_0000101001000000"; -- -0.12994323666702084
	pesos_i(20) := b"1111111111111111_1111111111111111_1111101001101010_0110000011011010"; -- -0.021814295488714035
	pesos_i(21) := b"1111111111111111_1111111111111111_1110010011000101_1111100011110100"; -- -0.1063541798272583
	pesos_i(22) := b"1111111111111111_1111111111111111_1110101010001011_1010100110001100"; -- -0.08380642253752774
	pesos_i(23) := b"0000000000000000_0000000000000000_0010010101011111_0100000001010000"; -- 0.1459846683476552
	pesos_i(24) := b"0000000000000000_0000000000000000_0000010111000001_0101111101010000"; -- 0.022481877421051726
	pesos_i(25) := b"0000000000000000_0000000000000000_0010011101101000_0101100110000010"; -- 0.15393599907214392
	pesos_i(26) := b"1111111111111111_1111111111111111_1111111101011000_1001000101100010"; -- -0.0025548111771844
	pesos_i(27) := b"0000000000000000_0000000000000000_0000001000101100_1100001110011010"; -- 0.008495545517620136
	pesos_i(28) := b"1111111111111111_1111111111111111_1111100011010101_1000110100100110"; -- -0.027991464739335746
	pesos_i(29) := b"1111111111111111_1111111111111111_1110001011000111_1101001001100100"; -- -0.11413846062281013
	pesos_i(30) := b"1111111111111111_1111111111111111_1111001100001011_1010101010000011"; -- -0.0506032401063762
	pesos_i(31) := b"0000000000000000_0000000000000000_0000000010111001_1010001111000101"; -- 0.0028326373372367653
	pesos_i(32) := b"1111111111111111_1111111111111111_1101011101110111_0000010111101100"; -- -0.15834010110894653
	pesos_i(33) := b"1111111111111111_1111111111111111_1111010111011111_0110011101011011"; -- -0.03955987953063372
	pesos_i(34) := b"1111111111111111_1111111111111111_1110011101101011_0101110100111111"; -- -0.09601800161546319
	pesos_i(35) := b"1111111111111111_1111111111111111_1111100110110011_0000110000000110"; -- -0.02461171005142971
	pesos_i(36) := b"1111111111111111_1111111111111111_1111111010001110_0000001001001001"; -- -0.005645615811281775
	pesos_i(37) := b"0000000000000000_0000000000000000_0001100111111111_1010000110101001"; -- 0.1015568769173631
	pesos_i(38) := b"0000000000000000_0000000000000000_0000111111100110_0001100110011000"; -- 0.06210479690959038
	pesos_i(39) := b"1111111111111111_1111111111111111_1110101100000110_0011000110001111"; -- -0.08193674345119616
	pesos_i(40) := b"0000000000000000_0000000000000000_0000110000101001_1001010000100011"; -- 0.04750944009065072
	pesos_i(41) := b"0000000000000000_0000000000000000_0000110101100011_0001101010100110"; -- 0.052293458426997966
	pesos_i(42) := b"1111111111111111_1111111111111111_1111011100100001_0101100100111001"; -- -0.034647391842967126
	pesos_i(43) := b"1111111111111111_1111111111111111_1110001111100000_0001000010001001"; -- -0.10986229575311009
	pesos_i(44) := b"0000000000000000_0000000000000000_0001000001110011_1101001111000111"; -- 0.06426738365683018
	pesos_i(45) := b"0000000000000000_0000000000000000_0000111010011100_0011010000000100"; -- 0.05707097152322563
	pesos_i(46) := b"1111111111111111_1111111111111111_1110100101011000_1010011101100101"; -- -0.088490999078809
	pesos_i(47) := b"1111111111111111_1111111111111111_1111010101100001_0001111111010000"; -- -0.04148675124832768
	pesos_i(48) := b"0000000000000000_0000000000000000_0000011000011111_1100101011001111"; -- 0.02392261076115515
	pesos_i(49) := b"0000000000000000_0000000000000000_0010100111011010_1101100010011001"; -- 0.16349557613639462
	pesos_i(50) := b"1111111111111111_1111111111111111_1111000000011111_0001110000100011"; -- -0.06202530040775884
	pesos_i(51) := b"0000000000000000_0000000000000000_0010101101011001_0011111110000111"; -- 0.16933056866269944
	pesos_i(52) := b"0000000000000000_0000000000000000_0000011000010111_0100101100000001"; -- 0.023792922711594732
	pesos_i(53) := b"0000000000000000_0000000000000000_0001000101101111_0100110101101001"; -- 0.06810458954657223
	pesos_i(54) := b"1111111111111111_1111111111111111_1111001111010000_0000111011011011"; -- -0.047606536502442405
	pesos_i(55) := b"0000000000000000_0000000000000000_0000011100001001_0010011100111101"; -- 0.027483417995133635
	pesos_i(56) := b"1111111111111111_1111111111111111_1110000101110101_0000000000110000"; -- -0.11930846039108825
	pesos_i(57) := b"0000000000000000_0000000000000000_0010101001001011_0101110001100100"; -- 0.16521241605760922
	pesos_i(58) := b"0000000000000000_0000000000000000_0010000100000111_1100100011001111"; -- 0.12902503072852595
	pesos_i(59) := b"0000000000000000_0000000000000000_0010100110010000_0110101011010111"; -- 0.16235988384972758
	pesos_i(60) := b"0000000000000000_0000000000000000_0001110000000100_1000001001101000"; -- 0.10944380796469072
	pesos_i(61) := b"1111111111111111_1111111111111111_1111100100010101_0101100011011010"; -- -0.02701801950857455
	pesos_i(62) := b"1111111111111111_1111111111111111_1111001100101110_0101010111010000"; -- -0.050074230832606204
	pesos_i(63) := b"0000000000000000_0000000000000000_0010010000010001_0110011111000111"; -- 0.14089058496030213
	pesos_i(64) := b"1111111111111111_1111111111111111_1111111000100101_0101001110000010"; -- -0.007242947313767345
	pesos_i(65) := b"1111111111111111_1111111111111111_1111010001000110_1101011011011110"; -- -0.04579407767787791
	pesos_i(66) := b"0000000000000000_0000000000000000_0001100010010000_1010110000100010"; -- 0.09595752549374226
	pesos_i(67) := b"1111111111111111_1111111111111111_1111101110000101_1000100000111111"; -- -0.01749371022860996
	pesos_i(68) := b"0000000000000000_0000000000000000_0001000011010111_0101011010110000"; -- 0.0657858066189019
	pesos_i(69) := b"1111111111111111_1111111111111111_1110101100110010_0001010101110001"; -- -0.08126703259797076
	pesos_i(70) := b"0000000000000000_0000000000000000_0001011101100101_1011010001101100"; -- 0.0913956416363043
	pesos_i(71) := b"0000000000000000_0000000000000000_0010011011101111_1010101001010000"; -- 0.15209450194775329
	pesos_i(72) := b"0000000000000000_0000000000000000_0001111101011011_1101001101100001"; -- 0.12249489891914069
	pesos_i(73) := b"0000000000000000_0000000000000000_0001001011100111_0000111111101110"; -- 0.07383822973696107
	pesos_i(74) := b"1111111111111111_1111111111111111_1111000011010101_1101101010001001"; -- -0.05923685233525367
	pesos_i(75) := b"1111111111111111_1111111111111111_1110011101100111_0000111101010100"; -- -0.09608368121489513
	pesos_i(76) := b"0000000000000000_0000000000000000_0000111000010101_1001100101111010"; -- 0.05501708251099868
	pesos_i(77) := b"0000000000000000_0000000000000000_0001110010010001_1001010010000000"; -- 0.1115963757781782
	pesos_i(78) := b"0000000000000000_0000000000000000_0010001101011110_0101001111010010"; -- 0.13815807228685908
	pesos_i(79) := b"1111111111111111_1111111111111111_1110110011001001_0001110110011000"; -- -0.07505621944102564
	pesos_i(80) := b"1111111111111111_1111111111111111_1111110000100101_0000100011011010"; -- -0.015059897238211828
	pesos_i(81) := b"0000000000000000_0000000000000000_0000110001100001_1010000101110111"; -- 0.04836472648699808
	pesos_i(82) := b"1111111111111111_1111111111111111_1111110000001100_0000001111010001"; -- -0.015441667146472358
	pesos_i(83) := b"1111111111111111_1111111111111111_1111100110100111_1110110110110001"; -- -0.024781364684274252
	pesos_i(84) := b"1111111111111111_1111111111111111_1101110110000000_1001011010110111"; -- -0.13475664163665027
	pesos_i(85) := b"0000000000000000_0000000000000000_0010010110000101_1111110001000101"; -- 0.1465757054818761
	pesos_i(86) := b"0000000000000000_0000000000000000_0010010011100111_1010000101010111"; -- 0.14415939693849714
	pesos_i(87) := b"1111111111111111_1111111111111111_1111010110101111_1110001101010000"; -- -0.040284912959427335
	pesos_i(88) := b"1111111111111111_1111111111111111_1101001110001010_0101001110011000"; -- -0.17367055443317736
	pesos_i(89) := b"0000000000000000_0000000000000000_0000101001110101_1110010001100110"; -- 0.04086139181419998
	pesos_i(90) := b"0000000000000000_0000000000000000_0010000000111010_1011100001111000"; -- 0.12589600499827644
	pesos_i(91) := b"1111111111111111_1111111111111111_1110010010110000_0100111110010010"; -- -0.10668471033241826
	pesos_i(92) := b"1111111111111111_1111111111111111_1111011100110000_1111010111101101"; -- -0.03440916972487309
	pesos_i(93) := b"0000000000000000_0000000000000000_0010000110001010_1000111010110111"; -- 0.1310204693387015
	pesos_i(94) := b"1111111111111111_1111111111111111_1110001001010100_1101000111111011"; -- -0.11589324591777597
	pesos_i(95) := b"0000000000000000_0000000000000000_0000111101010011_0000111010100001"; -- 0.05986110145254053
	pesos_i(96) := b"0000000000000000_0000000000000000_0000100001000011_0111010101000010"; -- 0.0322793278859736
	pesos_i(97) := b"1111111111111111_1111111111111111_1110010100010011_1100111011110111"; -- -0.10516649687869767
	pesos_i(98) := b"1111111111111111_1111111111111111_1111000110110100_0111011001000111"; -- -0.05584011806802757
	pesos_i(99) := b"1111111111111111_1111111111111111_1110111101011001_0110010101100100"; -- -0.06504217431875584
	pesos_i(100) := b"1111111111111111_1111111111111111_1110111101000111_1100101110110000"; -- -0.06531073520843472
	pesos_i(101) := b"1111111111111111_1111111111111111_1110100011001010_0101010011011000"; -- -0.09066266759711435
	pesos_i(102) := b"1111111111111111_1111111111111111_1101100110110101_0111000110001111"; -- -0.1495751405601744
	pesos_i(103) := b"0000000000000000_0000000000000000_0000000000100010_1111001101011111"; -- 0.0005333048109609773
	pesos_i(104) := b"1111111111111111_1111111111111111_1101111111010000_1001100001111111"; -- -0.1257233324849441
	pesos_i(105) := b"1111111111111111_1111111111111111_1101101101101110_0111001001111011"; -- -0.14284595967224312
	pesos_i(106) := b"0000000000000000_0000000000000000_0001011010111111_1100110001100111"; -- 0.08886411193995442
	pesos_i(107) := b"0000000000000000_0000000000000000_0000010110100000_0000100101100101"; -- 0.021973216250822016
	pesos_i(108) := b"0000000000000000_0000000000000000_0001100010011111_0001001001100111"; -- 0.09617724443658979
	pesos_i(109) := b"1111111111111111_1111111111111111_1101010100001110_1000110111000100"; -- -0.16774667698165124
	pesos_i(110) := b"0000000000000000_0000000000000000_0010100001101101_1100011011000110"; -- 0.15792505578101948
	pesos_i(111) := b"0000000000000000_0000000000000000_0000001011000100_1010110111010000"; -- 0.010813582683039748
	pesos_i(112) := b"1111111111111111_1111111111111111_1111100000001100_0110100001001011"; -- -0.031060678180181156
	pesos_i(113) := b"0000000000000000_0000000000000000_0010101001101110_1110111101110011"; -- 0.1657552391307243
	pesos_i(114) := b"1111111111111111_1111111111111111_1111010101110101_0111011101000100"; -- -0.04117636278686662
	pesos_i(115) := b"1111111111111111_1111111111111111_1111001010110111_1111100001100000"; -- -0.051880337305506626
	pesos_i(116) := b"1111111111111111_1111111111111111_1111000110101001_0010010111010001"; -- -0.05601276067712278
	pesos_i(117) := b"0000000000000000_0000000000000000_0001011011010100_1101100011001000"; -- 0.08918528446653734
	pesos_i(118) := b"1111111111111111_1111111111111111_1111011100000010_1111011111011011"; -- -0.03511095900822115
	pesos_i(119) := b"0000000000000000_0000000000000000_0011000001011111_0001000101001110"; -- 0.18895061628499055
	pesos_i(120) := b"1111111111111111_1111111111111111_1101011000100110_0001100011111010"; -- -0.16348117732318684
	pesos_i(121) := b"0000000000000000_0000000000000000_0010000000000001_1111000101001111"; -- 0.12502964180393006
	pesos_i(122) := b"1111111111111111_1111111111111111_1101011111101110_0001000000011101"; -- -0.1565236976697425
	pesos_i(123) := b"1111111111111111_1111111111111111_1110010011101010_0001010100100111"; -- -0.10580318251491425
	pesos_i(124) := b"1111111111111111_1111111111111111_1111001111100101_0110000100001011"; -- -0.047281203069033606
	pesos_i(125) := b"0000000000000000_0000000000000000_0010101010000011_1000110010111001"; -- 0.16606978903928113
	pesos_i(126) := b"1111111111111111_1111111111111111_1110001100010011_0011101111100101"; -- -0.11298776299784656
	pesos_i(127) := b"1111111111111111_1111111111111111_1101010011000010_1001010001100001"; -- -0.16890595094648433
	pesos_i(128) := b"1111111111111111_1111111111111111_1110100100000001_0110111100111011"; -- -0.08982186129183585
	pesos_i(129) := b"1111111111111111_1111111111111111_1110010001100010_0010111000011111"; -- -0.1078768897425825
	pesos_i(130) := b"0000000000000000_0000000000000000_0001111111101111_1110010101001001"; -- 0.12475426714551666
	pesos_i(131) := b"0000000000000000_0000000000000000_0010100101101111_0010101101101100"; -- 0.16185256380973548
	pesos_i(132) := b"0000000000000000_0000000000000000_0001100100100110_0101111010100000"; -- 0.09824172396818584
	pesos_i(133) := b"1111111111111111_1111111111111111_1111111010011010_1111001110000010"; -- -0.005448132275870621
	pesos_i(134) := b"1111111111111111_1111111111111111_1110001001111100_0111101101101101"; -- -0.1152880533250273
	pesos_i(135) := b"1111111111111111_1111111111111111_1111110010111111_0000110000000111"; -- -0.01270985441565297
	pesos_i(136) := b"1111111111111111_1111111111111111_1111110111011111_0101101001010000"; -- -0.008310657073160779
	pesos_i(137) := b"1111111111111111_1111111111111111_1110010000001011_1011110000000110"; -- -0.10919594622609426
	pesos_i(138) := b"1111111111111111_1111111111111111_1101100100101011_0100010110001111"; -- -0.1516834760585639
	pesos_i(139) := b"1111111111111111_1111111111111111_1111110110000011_0100000000100010"; -- -0.00971602595321465
	pesos_i(140) := b"1111111111111111_1111111111111111_1111000101010111_1110100000010101"; -- -0.057252402300588805
	pesos_i(141) := b"0000000000000000_0000000000000000_0001000011110100_1001101101111011"; -- 0.06623241178753139
	pesos_i(142) := b"0000000000000000_0000000000000000_0000010001010010_1110100001110110"; -- 0.016890076482109172
	pesos_i(143) := b"0000000000000000_0000000000000000_0001100101100101_1110011110110100"; -- 0.09921119819097492
	pesos_i(144) := b"1111111111111111_1111111111111111_1110000001001110_0111011100100011"; -- -0.12380271337922452
	pesos_i(145) := b"0000000000000000_0000000000000000_0001100011010110_1111100111100110"; -- 0.09703027591872372
	pesos_i(146) := b"1111111111111111_1111111111111111_1110010000000001_0110111011010101"; -- -0.10935313512789341
	pesos_i(147) := b"1111111111111111_1111111111111111_1110110000111010_1111111010001001"; -- -0.07722481880038201
	pesos_i(148) := b"0000000000000000_0000000000000000_0001000111110000_0111001001110110"; -- 0.0700751816660594
	pesos_i(149) := b"0000000000000000_0000000000000000_0001110001111011_0011111101111000"; -- 0.11125561419039369
	pesos_i(150) := b"0000000000000000_0000000000000000_0000110010001111_1100010000011011"; -- 0.04906869553407937
	pesos_i(151) := b"1111111111111111_1111111111111111_1111110100101110_1000101111010110"; -- -0.011008510742556682
	pesos_i(152) := b"1111111111111111_1111111111111111_1110110111101110_1101100111110101"; -- -0.07057416685648175
	pesos_i(153) := b"1111111111111111_1111111111111111_1110101101110011_0110110010111001"; -- -0.08027000897762716
	pesos_i(154) := b"0000000000000000_0000000000000000_0001100011110101_1011010011001001"; -- 0.09749917884596287
	pesos_i(155) := b"1111111111111111_1111111111111111_1101100011110001_1111100111100010"; -- -0.15255773770625358
	pesos_i(156) := b"0000000000000000_0000000000000000_0000000110011110_1100101100111101"; -- 0.006329252692891979
	pesos_i(157) := b"1111111111111111_1111111111111111_1111100101101111_1101000100010110"; -- -0.02563756202030092
	pesos_i(158) := b"1111111111111111_1111111111111111_1110100000101101_0010111111111001"; -- -0.0930604950765151
	pesos_i(159) := b"0000000000000000_0000000000000000_0001010110100010_0111101011000100"; -- 0.08451049114225964
	pesos_i(160) := b"0000000000000000_0000000000000000_0010000110011100_0101100111000111"; -- 0.13129197217900876
	pesos_i(161) := b"1111111111111111_1111111111111111_1110011101100010_1010000011011101"; -- -0.09615130036426874
	pesos_i(162) := b"0000000000000000_0000000000000000_0001101100100111_1010010101010010"; -- 0.10607369654005065
	pesos_i(163) := b"1111111111111111_1111111111111111_1110011000100111_1011111011110001"; -- -0.10095602616112348
	pesos_i(164) := b"0000000000000000_0000000000000000_0000100010011001_0000110000011100"; -- 0.0335853165472436
	pesos_i(165) := b"1111111111111111_1111111111111111_1110011100111100_1111010011000010"; -- -0.09672613389331124
	pesos_i(166) := b"0000000000000000_0000000000000000_0010001001100111_0011100010011111"; -- 0.13438753025021444
	pesos_i(167) := b"0000000000000000_0000000000000000_0010010100110001_1010011101001100"; -- 0.14528890230251892
	pesos_i(168) := b"0000000000000000_0000000000000000_0000101100010000_1100111000110011"; -- 0.04322518096911196
	pesos_i(169) := b"1111111111111111_1111111111111111_1110010110111100_0110110011010011"; -- -0.10259361113243905
	pesos_i(170) := b"0000000000000000_0000000000000000_0000111001011010_0110000000011101"; -- 0.056066519873387684
	pesos_i(171) := b"0000000000000000_0000000000000000_0000101010100000_1110101011101011"; -- 0.04151790855063023
	pesos_i(172) := b"1111111111111111_1111111111111111_1110000100111011_0001010110010111"; -- -0.12019219458347075
	pesos_i(173) := b"1111111111111111_1111111111111111_1111011001000010_0101001100010111"; -- -0.038050467429098914
	pesos_i(174) := b"0000000000000000_0000000000000000_0001010011000011_0111101100100101"; -- 0.08110780395813702
	pesos_i(175) := b"0000000000000000_0000000000000000_0000111110110101_1110101100111101"; -- 0.061369612161748265
	pesos_i(176) := b"1111111111111111_1111111111111111_1110101001001101_0101111001111111"; -- -0.08475694089104654
	pesos_i(177) := b"0000000000000000_0000000000000000_0001111100101000_1110101011000100"; -- 0.12171809465652311
	pesos_i(178) := b"0000000000000000_0000000000000000_0000000010100011_1101010011110011"; -- 0.0024998754896811853
	pesos_i(179) := b"1111111111111111_1111111111111111_1101111100101111_1110010101111000"; -- -0.12817540951800938
	pesos_i(180) := b"0000000000000000_0000000000000000_0001010010001001_1001011111011111"; -- 0.08022450630379642
	pesos_i(181) := b"1111111111111111_1111111111111111_1111101011000111_0000101101000011"; -- -0.020400329759460427
	pesos_i(182) := b"1111111111111111_1111111111111111_1110111000110011_1011111110111011"; -- -0.06952287376712567
	pesos_i(183) := b"0000000000000000_0000000000000000_0000011001000101_0100010011110111"; -- 0.024494467172678894
	pesos_i(184) := b"1111111111111111_1111111111111111_1111000100110100_1100011110111000"; -- -0.05778838888489135
	pesos_i(185) := b"0000000000000000_0000000000000000_0001100000010100_0011010101001100"; -- 0.09405835262794109
	pesos_i(186) := b"0000000000000000_0000000000000000_0000010110010111_1111010010101000"; -- 0.021849909720049694
	pesos_i(187) := b"0000000000000000_0000000000000000_0000000111101011_1000000100100001"; -- 0.0074997620156546495
	pesos_i(188) := b"1111111111111111_1111111111111111_1111111111101111_0100001111101000"; -- -0.00025535179508590284
	pesos_i(189) := b"0000000000000000_0000000000000000_0010010101010010_0010100001110101"; -- 0.14578488215908494
	pesos_i(190) := b"0000000000000000_0000000000000000_0000110100111100_0000100110001101"; -- 0.051697346616227595
	pesos_i(191) := b"1111111111111111_1111111111111111_1111011000100000_1111100011001011"; -- -0.038559389422487586
	pesos_i(192) := b"0000000000000000_0000000000000000_0000010000011001_0011100101100001"; -- 0.016009889764371066
	pesos_i(193) := b"1111111111111111_1111111111111111_1110100000111011_0010101100011000"; -- -0.09284716285355878
	pesos_i(194) := b"1111111111111111_1111111111111111_1101100001111000_1010101100101110"; -- -0.15440874228038207
	pesos_i(195) := b"0000000000000000_0000000000000000_0001111000000110_1001010001001011"; -- 0.11728789164845602
	pesos_i(196) := b"1111111111111111_1111111111111111_1111110111001110_1000101000010010"; -- -0.008567209911179872
	pesos_i(197) := b"0000000000000000_0000000000000000_0010101001001101_1001000000100001"; -- 0.16524601744165598
	pesos_i(198) := b"0000000000000000_0000000000000000_0000110010101100_1100100001100011"; -- 0.04951145566270889
	pesos_i(199) := b"1111111111111111_1111111111111111_1101101000110100_0010111100001011"; -- -0.1476412390759677
	pesos_i(200) := b"0000000000000000_0000000000000000_0010011100111101_1110111110000001"; -- 0.1532888117348275
	pesos_i(201) := b"1111111111111111_1111111111111111_1111111001100111_0001110010100011"; -- -0.006239137842549845
	pesos_i(202) := b"0000000000000000_0000000000000000_0010001001101010_0001011001011011"; -- 0.13443126413237125
	pesos_i(203) := b"1111111111111111_1111111111111111_1111001001110101_0011111010001001"; -- -0.05289849440468749
	pesos_i(204) := b"1111111111111111_1111111111111111_1110010011011010_0011111111110101"; -- -0.10604477185768833
	pesos_i(205) := b"0000000000000000_0000000000000000_0000000101010101_0101001100100011"; -- 0.005208202317266477
	pesos_i(206) := b"1111111111111111_1111111111111111_1110101111101001_1111110000000100"; -- -0.07846093087785969
	pesos_i(207) := b"0000000000000000_0000000000000000_0010100000111000_1100101101100100"; -- 0.15711661512516303
	pesos_i(208) := b"1111111111111111_1111111111111111_1110001010100100_0010100101011100"; -- -0.11468259344997678
	pesos_i(209) := b"1111111111111111_1111111111111111_1111111110100111_0111110110000010"; -- -0.0013505514261706146
	pesos_i(210) := b"1111111111111111_1111111111111111_1101110000011100_1101011100001001"; -- -0.1401849369090553
	pesos_i(211) := b"0000000000000000_0000000000000000_0001110111100011_1000000100001100"; -- 0.11675268700425906
	pesos_i(212) := b"0000000000000000_0000000000000000_0010010111111101_0010101111010010"; -- 0.14839433546769806
	pesos_i(213) := b"0000000000000000_0000000000000000_0010001101000000_1011100000110110"; -- 0.13770629232854
	pesos_i(214) := b"1111111111111111_1111111111111111_1111111010110111_0011110100110000"; -- -0.005016494455593433
	pesos_i(215) := b"1111111111111111_1111111111111111_1101001010110100_1011110111100111"; -- -0.17692959892432933
	pesos_i(216) := b"1111111111111111_1111111111111111_1110101011101111_0011110000111101"; -- -0.08228705898870883
	pesos_i(217) := b"0000000000000000_0000000000000000_0010110000011100_1011101111110010"; -- 0.1723134485809633
	pesos_i(218) := b"0000000000000000_0000000000000000_0001000110001100_1100100101110100"; -- 0.06855448800535054
	pesos_i(219) := b"1111111111111111_1111111111111111_1111000000000001_1111101011011001"; -- -0.062469789639616476
	pesos_i(220) := b"1111111111111111_1111111111111111_1111010101101011_1101111000101111"; -- -0.04132281646062396
	pesos_i(221) := b"1111111111111111_1111111111111111_1110001101100111_0011111000101111"; -- -0.11170588819458592
	pesos_i(222) := b"0000000000000000_0000000000000000_0000001101100010_0100101011101100"; -- 0.013218577070978187
	pesos_i(223) := b"1111111111111111_1111111111111111_1101010011101100_0100011111100001"; -- -0.16826964156670385
	pesos_i(224) := b"1111111111111111_1111111111111111_1110000000001101_1111010001101000"; -- -0.1247870680776487
	pesos_i(225) := b"1111111111111111_1111111111111111_1110101111011100_0001100111000011"; -- -0.07867278078684586
	pesos_i(226) := b"0000000000000000_0000000000000000_0000100000000110_0010010111010011"; -- 0.03134380712701996
	pesos_i(227) := b"1111111111111111_1111111111111111_1110100010111011_1101100100101010"; -- -0.09088366255742251
	pesos_i(228) := b"0000000000000000_0000000000000000_0000010111100111_0110000111101011"; -- 0.02306186666447969
	pesos_i(229) := b"0000000000000000_0000000000000000_0000110101111011_0110100011101111"; -- 0.052664335697750156
	pesos_i(230) := b"0000000000000000_0000000000000000_0001110001110100_1111110000000010"; -- 0.11116004039946857
	pesos_i(231) := b"1111111111111111_1111111111111111_1110100010100010_1110000111011100"; -- -0.09126461392742546
	pesos_i(232) := b"1111111111111111_1111111111111111_1110000100100111_0101100011011010"; -- -0.1204933612452266
	pesos_i(233) := b"1111111111111111_1111111111111111_1101111100001001_0110100110111001"; -- -0.12876261924944477
	pesos_i(234) := b"0000000000000000_0000000000000000_0001111001110010_0010110001010111"; -- 0.11892964478650075
	pesos_i(235) := b"1111111111111111_1111111111111111_1110001011100001_0101010000111010"; -- -0.11374925223851302
	pesos_i(236) := b"1111111111111111_1111111111111111_1110101101011001_0100010100001011"; -- -0.08066910250266626
	pesos_i(237) := b"1111111111111111_1111111111111111_1111110000000000_1010101000110100"; -- -0.015614855031598629
	pesos_i(238) := b"0000000000000000_0000000000000000_0001000001100111_1000111101000110"; -- 0.06408019510505811
	pesos_i(239) := b"0000000000000000_0000000000000000_0010111101110110_0011110010111111"; -- 0.18539790782710316
	pesos_i(240) := b"0000000000000000_0000000000000000_0000011000101010_1111010110001011"; -- 0.02409300456343899
	pesos_i(241) := b"1111111111111111_1111111111111111_1110000001000010_0101110100000100"; -- -0.12398737568827643
	pesos_i(242) := b"1111111111111111_1111111111111111_1110011010100010_0101010011000100"; -- -0.0990855237919612
	pesos_i(243) := b"1111111111111111_1111111111111111_1101001100000011_1100001100011001"; -- -0.17572384495884433
	pesos_i(244) := b"0000000000000000_0000000000000000_0010011000111011_1011100011100010"; -- 0.1493487883845692
	pesos_i(245) := b"0000000000000000_0000000000000000_0010101001111101_0100110011011100"; -- 0.1659744297943291
	pesos_i(246) := b"1111111111111111_1111111111111111_1110110011111000_1011111001110110"; -- -0.07432946785722515
	pesos_i(247) := b"0000000000000000_0000000000000000_0000111010100111_1100010100010111"; -- 0.0572474652531144
	pesos_i(248) := b"0000000000000000_0000000000000000_0000101111101001_1010110110000110"; -- 0.04653439061335174
	pesos_i(249) := b"0000000000000000_0000000000000000_0010011001111001_1101111111110011"; -- 0.15029716199528476
	pesos_i(250) := b"0000000000000000_0000000000000000_0001011111101000_0011111100001000"; -- 0.093387545979588
	pesos_i(251) := b"1111111111111111_1111111111111111_1110111011011100_0000000111010111"; -- -0.06695545681311503
	pesos_i(252) := b"1111111111111111_1111111111111111_1110101110100010_0010100011000000"; -- -0.07955689726633819
	pesos_i(253) := b"0000000000000000_0000000000000000_0000110000101110_1001010111010010"; -- 0.04758583427648927
	pesos_i(254) := b"0000000000000000_0000000000000000_0010100101100100_0110010110110001"; -- 0.16168819029849427
	pesos_i(255) := b"0000000000000000_0000000000000000_0000010110001010_1000110000011011"; -- 0.021645313770284887
	pesos_i(256) := b"0000000000000000_0000000000000000_0000101111100001_0100000011110111"; -- 0.04640584964525338
	pesos_i(257) := b"1111111111111111_1111111111111111_1101001101000111_0010000000000110"; -- -0.1746959671290391
	pesos_i(258) := b"0000000000000000_0000000000000000_0000000011110011_0110011000100010"; -- 0.0037139733555769583
	pesos_i(259) := b"1111111111111111_1111111111111111_1101100001100010_0100010011100000"; -- -0.1547505334869514
	pesos_i(260) := b"1111111111111111_1111111111111111_1111101111000010_0110001111111110"; -- -0.01656508496600552
	pesos_i(261) := b"0000000000000000_0000000000000000_0010011001011011_0001100000111010"; -- 0.14982749371499784
	pesos_i(262) := b"0000000000000000_0000000000000000_0000011101101100_0100001001010000"; -- 0.028995651729948675
	pesos_i(263) := b"0000000000000000_0000000000000000_0001010111101001_1001100100111100"; -- 0.08559568144060326
	pesos_i(264) := b"1111111111111111_1111111111111111_1110010011001101_1111100010001000"; -- -0.10623213473290176
	pesos_i(265) := b"0000000000000000_0000000000000000_0001110100111011_0010001001010011"; -- 0.11418356451042308
	pesos_i(266) := b"0000000000000000_0000000000000000_0001111001100001_1000101111111110"; -- 0.11867594683559972
	pesos_i(267) := b"0000000000000000_0000000000000000_0001100110011000_1101111100011100"; -- 0.09998888430872371
	pesos_i(268) := b"1111111111111111_1111111111111111_1111110101001011_0001011001100000"; -- -0.01057300723211732
	pesos_i(269) := b"1111111111111111_1111111111111111_1110010101010100_0101111101111000"; -- -0.1041813213299396
	pesos_i(270) := b"1111111111111111_1111111111111111_1110110101000110_0011010110110100"; -- -0.07314743391464486
	pesos_i(271) := b"1111111111111111_1111111111111111_1110001011110011_1101110010101111"; -- -0.11346646045400849
	pesos_i(272) := b"1111111111111111_1111111111111111_1111001001000111_0100010000000110"; -- -0.05360007150250838
	pesos_i(273) := b"1111111111111111_1111111111111111_1101110010101101_0110001100101010"; -- -0.1379793188329046
	pesos_i(274) := b"0000000000000000_0000000000000000_0001000100110000_0100010010001101"; -- 0.06714275786222783
	pesos_i(275) := b"1111111111111111_1111111111111111_1111100100111000_1010100010101110"; -- -0.02647920374613375
	pesos_i(276) := b"1111111111111111_1111111111111111_1111011111101111_0001011010101011"; -- -0.031508048187274415
	pesos_i(277) := b"0000000000000000_0000000000000000_0010110011000010_1110110100110101"; -- 0.17484934362283897
	pesos_i(278) := b"1111111111111111_1111111111111111_1101100001101110_1011001100101110"; -- -0.1545608532410233
	pesos_i(279) := b"0000000000000000_0000000000000000_0010100010000001_0101000010011110"; -- 0.15822318889978795
	pesos_i(280) := b"1111111111111111_1111111111111111_1110000101100111_0100011011001111"; -- -0.11951787418466267
	pesos_i(281) := b"0000000000000000_0000000000000000_0001101000011001_0001100010100100"; -- 0.10194543836854969
	pesos_i(282) := b"0000000000000000_0000000000000000_0001010000000000_0110111011101011"; -- 0.07813161133838087
	pesos_i(283) := b"0000000000000000_0000000000000000_0001010010100011_1010001111001111"; -- 0.08062194641459462
	pesos_i(284) := b"1111111111111111_1111111111111111_1101110101111010_1010111111100000"; -- -0.13484669477657907
	pesos_i(285) := b"1111111111111111_1111111111111111_1110010011000101_0111100101100000"; -- -0.10636178405888988
	pesos_i(286) := b"0000000000000000_0000000000000000_0001110110100000_1001000010111111"; -- 0.11573128379433895
	pesos_i(287) := b"1111111111111111_1111111111111111_1111000110101011_0000011011011111"; -- -0.05598408748112692
	pesos_i(288) := b"0000000000000000_0000000000000000_0010100100101100_1101010010100011"; -- 0.1608403109352923
	pesos_i(289) := b"1111111111111111_1111111111111111_1110111101001001_1010100011111010"; -- -0.06528228650398907
	pesos_i(290) := b"0000000000000000_0000000000000000_0000100100010100_0010000111010101"; -- 0.03546344225769369
	pesos_i(291) := b"1111111111111111_1111111111111111_1111010001001010_1110000001000101"; -- -0.045732482062353634
	pesos_i(292) := b"1111111111111111_1111111111111111_1111010000100000_0101100011101000"; -- -0.04638141947906404
	pesos_i(293) := b"0000000000000000_0000000000000000_0000100001000100_1100001111010100"; -- 0.03229926989210122
	pesos_i(294) := b"1111111111111111_1111111111111111_1111111011100111_0000111100110010"; -- -0.004286814091942652
	pesos_i(295) := b"0000000000000000_0000000000000000_0000111101101111_0001000010001001"; -- 0.060288461098213286
	pesos_i(296) := b"0000000000000000_0000000000000000_0001111110100001_1000010110110000"; -- 0.12355838350330742
	pesos_i(297) := b"0000000000000000_0000000000000000_0001011101010110_1100011000001001"; -- 0.09116780966866671
	pesos_i(298) := b"1111111111111111_1111111111111111_1111000011001110_1100010010100010"; -- -0.05934496929369403
	pesos_i(299) := b"1111111111111111_1111111111111111_1101111111001011_1100010001000100"; -- -0.12579701738059826
	pesos_i(300) := b"0000000000000000_0000000000000000_0001000010111010_1010011001011011"; -- 0.06534805024274368
	pesos_i(301) := b"0000000000000000_0000000000000000_0001110100011100_1010110101001011"; -- 0.1137188251201214
	pesos_i(302) := b"1111111111111111_1111111111111111_1101101000000000_0111001000000000"; -- -0.1484307051560219
	pesos_i(303) := b"1111111111111111_1111111111111111_1110000010001111_0010000100111101"; -- -0.12281601204629689
	pesos_i(304) := b"1111111111111111_1111111111111111_1111000000001101_1101111101111110"; -- -0.06228831465956283
	pesos_i(305) := b"1111111111111111_1111111111111111_1111100101100001_0110001110111111"; -- -0.02585770216708162
	pesos_i(306) := b"1111111111111111_1111111111111111_1110111111110010_1100000011010101"; -- -0.06270212925024797
	pesos_i(307) := b"0000000000000000_0000000000000000_0010011000100001_0101110110010110"; -- 0.1489466182086552
	pesos_i(308) := b"1111111111111111_1111111111111111_1111001100111000_1000010100000010"; -- -0.04991882988250142
	pesos_i(309) := b"0000000000000000_0000000000000000_0001001110110110_1001000111100000"; -- 0.07700454433972623
	pesos_i(310) := b"0000000000000000_0000000000000000_0000011111011100_1100000101011100"; -- 0.0307122086872939
	pesos_i(311) := b"0000000000000000_0000000000000000_0001110100110111_0010100111011000"; -- 0.11412297756844494
	pesos_i(312) := b"0000000000000000_0000000000000000_0001101100111011_0010111010100100"; -- 0.10637179854645798
	pesos_i(313) := b"0000000000000000_0000000000000000_0000001000010001_1110001100101000"; -- 0.008085438912774419
	pesos_i(314) := b"1111111111111111_1111111111111111_1111111100010111_1101101000010010"; -- -0.0035422997610877437
	pesos_i(315) := b"1111111111111111_1111111111111111_1110100101100110_1010000011110110"; -- -0.08827775946156763
	pesos_i(316) := b"1111111111111111_1111111111111111_1110110110001010_1000001010110011"; -- -0.07210524688526632
	pesos_i(317) := b"1111111111111111_1111111111111111_1101110011011110_0110000110111110"; -- -0.13723172288467286
	pesos_i(318) := b"0000000000000000_0000000000000000_0001100110001111_1011101100101100"; -- 0.09984941315612578
	pesos_i(319) := b"1111111111111111_1111111111111111_1110100101001111_1000100111111111"; -- -0.08863008044150052
	pesos_i(320) := b"1111111111111111_1111111111111111_1110111110111001_1011000100011011"; -- -0.06357281772332757
	pesos_i(321) := b"0000000000000000_0000000000000000_0001111010101101_0100001110001010"; -- 0.11983129620392911
	pesos_i(322) := b"0000000000000000_0000000000000000_0001000011110111_0100011101011000"; -- 0.06627317323041905
	pesos_i(323) := b"0000000000000000_0000000000000000_0001010000111100_0001111101011010"; -- 0.07904239599819993
	pesos_i(324) := b"1111111111111111_1111111111111111_1110111101011110_0100101111010001"; -- -0.06496740473699035
	pesos_i(325) := b"1111111111111111_1111111111111111_1110011000001101_1101101010010101"; -- -0.10135110718318567
	pesos_i(326) := b"0000000000000000_0000000000000000_0001101110101110_0110110010100100"; -- 0.10813025485756163
	pesos_i(327) := b"1111111111111111_1111111111111111_1111100100001100_1000001010010101"; -- -0.0271528611210181
	pesos_i(328) := b"1111111111111111_1111111111111111_1110100000001110_0101000100100101"; -- -0.09353154029196172
	pesos_i(329) := b"0000000000000000_0000000000000000_0001110010111101_0101100010110010"; -- 0.11226419788114318
	pesos_i(330) := b"1111111111111111_1111111111111111_1111111011111011_0100100110011001"; -- -0.0039781571016012885
	pesos_i(331) := b"1111111111111111_1111111111111111_1111100110101101_1001111100101001"; -- -0.02469449291236025
	pesos_i(332) := b"1111111111111111_1111111111111111_1111001100100101_0100000010011001"; -- -0.050212824472708376
	pesos_i(333) := b"0000000000000000_0000000000000000_0010101010000110_1000100010001010"; -- 0.16611531608897862
	pesos_i(334) := b"1111111111111111_1111111111111111_1110101011001011_1010011110011111"; -- -0.08282997473661736
	pesos_i(335) := b"1111111111111111_1111111111111111_1110111100101001_1111010000010110"; -- -0.06576609107731916
	pesos_i(336) := b"0000000000000000_0000000000000000_0000001001100101_1010010100011000"; -- 0.009363477964486167
	pesos_i(337) := b"0000000000000000_0000000000000000_0010001110000011_0110110000101100"; -- 0.13872409896361435
	pesos_i(338) := b"1111111111111111_1111111111111111_1111110110001010_1100110111111101"; -- -0.00960075923729555
	pesos_i(339) := b"0000000000000000_0000000000000000_0010001000010010_0011010001010001"; -- 0.133090276527384
	pesos_i(340) := b"1111111111111111_1111111111111111_1110001001111011_0011000110001111"; -- -0.11530771499641523
	pesos_i(341) := b"0000000000000000_0000000000000000_0001110101001101_1100110111010100"; -- 0.11446844511685252
	pesos_i(342) := b"1111111111111111_1111111111111111_1111100000001111_0100001000111100"; -- -0.031017170313327527
	pesos_i(343) := b"0000000000000000_0000000000000000_0010110100100101_1001101011011001"; -- 0.17635505490543657
	pesos_i(344) := b"0000000000000000_0000000000000000_0010010000101001_0100110001000010"; -- 0.14125515565714794
	pesos_i(345) := b"0000000000000000_0000000000000000_0001101011001001_1000001110101111"; -- 0.10463736551073133
	pesos_i(346) := b"1111111111111111_1111111111111111_1101001011101100_0101001100010001"; -- -0.1760814746708205
	pesos_i(347) := b"0000000000000000_0000000000000000_0000001000100111_0101011001111110"; -- 0.008412748138898769
	pesos_i(348) := b"1111111111111111_1111111111111111_1101101100010111_0111010010011111"; -- -0.14417334659981307
	pesos_i(349) := b"1111111111111111_1111111111111111_1110101010111011_1111111100110000"; -- -0.08306889608866899
	pesos_i(350) := b"1111111111111111_1111111111111111_1110111011011110_1011010101000011"; -- -0.06691424468073215
	pesos_i(351) := b"1111111111111111_1111111111111111_1110111100010011_1001101100000011"; -- -0.06610709358160978
	pesos_i(352) := b"1111111111111111_1111111111111111_1110010001100000_0001101101100101"; -- -0.10790852335531534
	pesos_i(353) := b"1111111111111111_1111111111111111_1111101000101001_1111011100110110"; -- -0.02279715468714528
	pesos_i(354) := b"1111111111111111_1111111111111111_1110010011001101_0100011001001100"; -- -0.10624275832708462
	pesos_i(355) := b"1111111111111111_1111111111111111_1110100111011000_1001110100010010"; -- -0.08653848933365295
	pesos_i(356) := b"1111111111111111_1111111111111111_1110001001001010_0010100001001001"; -- -0.11605594835991709
	pesos_i(357) := b"1111111111111111_1111111111111111_1101110011111001_0100111011101000"; -- -0.13682085823233814
	pesos_i(358) := b"0000000000000000_0000000000000000_0010011110000110_1110000101101000"; -- 0.1544018630869388
	pesos_i(359) := b"1111111111111111_1111111111111111_1110100010000111_0100000010010101"; -- -0.0916862140538589
	pesos_i(360) := b"0000000000000000_0000000000000000_0001110111011110_1110110011111001"; -- 0.11668282583602932
	pesos_i(361) := b"0000000000000000_0000000000000000_0000010001111010_0010001101100000"; -- 0.017488680705044793
	pesos_i(362) := b"1111111111111111_1111111111111111_1110101100010101_0001011011011010"; -- -0.08170945343015537
	pesos_i(363) := b"0000000000000000_0000000000000000_0001010000010010_0101110100101100"; -- 0.07840521167830164
	pesos_i(364) := b"0000000000000000_0000000000000000_0001011100100111_0110110101101110"; -- 0.09044536526132295
	pesos_i(365) := b"0000000000000000_0000000000000000_0000011000011110_1010001110101000"; -- 0.023905018433114815
	pesos_i(366) := b"0000000000000000_0000000000000000_0010001010000000_0110110011011101"; -- 0.13477211372284514
	pesos_i(367) := b"0000000000000000_0000000000000000_0010000100010100_1101110010011010"; -- 0.12922457458133432
	pesos_i(368) := b"0000000000000000_0000000000000000_0010110100001101_0011011011000001"; -- 0.17598287784137454
	pesos_i(369) := b"1111111111111111_1111111111111111_1110100010110000_0111111100110011"; -- -0.09105687155425633
	pesos_i(370) := b"1111111111111111_1111111111111111_1110011000110110_1101010100100000"; -- -0.10072582219470798
	pesos_i(371) := b"0000000000000000_0000000000000000_0001111111100010_0100001011011110"; -- 0.12454622184513729
	pesos_i(372) := b"0000000000000000_0000000000000000_0000111010011111_1000010010001100"; -- 0.05712154777268234
	pesos_i(373) := b"0000000000000000_0000000000000000_0010111001011100_1101101111110110"; -- 0.1811044192785431
	pesos_i(374) := b"0000000000000000_0000000000000000_0001000110010001_0001000010001110"; -- 0.06861976109790427
	pesos_i(375) := b"0000000000000000_0000000000000000_0001011010001110_0000110111110000"; -- 0.08810507875213476
	pesos_i(376) := b"0000000000000000_0000000000000000_0010010100011001_0111111100011010"; -- 0.1449202955108221
	pesos_i(377) := b"0000000000000000_0000000000000000_0001000000100100_0110001111110101"; -- 0.06305527435803225
	pesos_i(378) := b"1111111111111111_1111111111111111_1111111001101101_0111011010010101"; -- -0.006142223924769208
	pesos_i(379) := b"1111111111111111_1111111111111111_1110001010110010_1011011011100101"; -- -0.11446053411708465
	pesos_i(380) := b"0000000000000000_0000000000000000_0010010101111101_0000101000010000"; -- 0.1464391983048644
	pesos_i(381) := b"0000000000000000_0000000000000000_0001110101101000_0011111111100010"; -- 0.1148719717082612
	pesos_i(382) := b"0000000000000000_0000000000000000_0001101000101101_1101001100011001"; -- 0.10226172786084314
	pesos_i(383) := b"1111111111111111_1111111111111111_1101010101111100_1110110010110100"; -- -0.16606255155220548
	pesos_i(384) := b"1111111111111111_1111111111111111_1101011100110001_0001000000100100"; -- -0.15940760731947123
	pesos_i(385) := b"1111111111111111_1111111111111111_1110011010101011_1010111010000010"; -- -0.09894284548151212
	pesos_i(386) := b"0000000000000000_0000000000000000_0001001100001101_1000011010000111"; -- 0.0744251327434579
	pesos_i(387) := b"0000000000000000_0000000000000000_0010100101110001_1111110011100011"; -- 0.16189556649231163
	pesos_i(388) := b"0000000000000000_0000000000000000_0010101000100000_1001001101100111"; -- 0.16455956701412086
	pesos_i(389) := b"1111111111111111_1111111111111111_1111101010100101_1000101011001110"; -- -0.020911526457499642
	pesos_i(390) := b"0000000000000000_0000000000000000_0000111101011111_0101100110001100"; -- 0.06004867240815165
	pesos_i(391) := b"0000000000000000_0000000000000000_0000101001100000_0001111011011110"; -- 0.040529183610727326
	pesos_i(392) := b"1111111111111111_1111111111111111_1101001010010000_0111001010001111"; -- -0.17748340617944708
	pesos_i(393) := b"0000000000000000_0000000000000000_0010001001111110_1000111000001111"; -- 0.13474357481578955
	pesos_i(394) := b"1111111111111111_1111111111111111_1111001000000011_0010100110010101"; -- -0.05463924519444192
	pesos_i(395) := b"0000000000000000_0000000000000000_0000110000011001_0001000000101000"; -- 0.04725743272957004
	pesos_i(396) := b"0000000000000000_0000000000000000_0000011110100000_0110110101010100"; -- 0.029791672698835175
	pesos_i(397) := b"0000000000000000_0000000000000000_0001000111101101_1010001101000001"; -- 0.07003231371339377
	pesos_i(398) := b"1111111111111111_1111111111111111_1111101100011101_1000111111110001"; -- -0.01908016548247242
	pesos_i(399) := b"0000000000000000_0000000000000000_0000111011101010_1110000111010010"; -- 0.05827151659849243
	pesos_i(400) := b"1111111111111111_1111111111111111_1110110100101000_1011111100001110"; -- -0.07359701069702332
	pesos_i(401) := b"1111111111111111_1111111111111111_1110011101110111_0100010011100011"; -- -0.09583634806192758
	pesos_i(402) := b"0000000000000000_0000000000000000_0000010110011000_1110010110111100"; -- 0.02186427905958385
	pesos_i(403) := b"0000000000000000_0000000000000000_0001100010011001_1100010010010100"; -- 0.09609631164428384
	pesos_i(404) := b"0000000000000000_0000000000000000_0001101101111011_0101000101100011"; -- 0.10735043211018218
	pesos_i(405) := b"1111111111111111_1111111111111111_1110110001000100_1000100010111001"; -- -0.07707925312144236
	pesos_i(406) := b"0000000000000000_0000000000000000_0000000110011010_1011100100100110"; -- 0.006267139188075261
	pesos_i(407) := b"1111111111111111_1111111111111111_1111111100110110_0101100101100010"; -- -0.003076947767875712
	pesos_i(408) := b"1111111111111111_1111111111111111_1111010100010000_1110111110110000"; -- -0.042710322991172826
	pesos_i(409) := b"1111111111111111_1111111111111111_1110010001010101_0000001000111011"; -- -0.10807787001279101
	pesos_i(410) := b"0000000000000000_0000000000000000_0010010011100101_0010001100011110"; -- 0.1441213557380217
	pesos_i(411) := b"0000000000000000_0000000000000000_0010001101001111_1010101101110110"; -- 0.13793441428869327
	pesos_i(412) := b"1111111111111111_1111111111111111_1110000001001010_1100011100101110"; -- -0.12385897758741837
	pesos_i(413) := b"0000000000000000_0000000000000000_0010011100100010_1111000011011000"; -- 0.15287690420620692
	pesos_i(414) := b"0000000000000000_0000000000000000_0000000110001111_1000000101010101"; -- 0.006095965608898964
	pesos_i(415) := b"0000000000000000_0000000000000000_0000000011100110_1101111111000001"; -- 0.003522858207697266
	pesos_i(416) := b"1111111111111111_1111111111111111_1110110101100000_1110110000101100"; -- -0.07273982929042111
	pesos_i(417) := b"1111111111111111_1111111111111111_1110010101110101_0000110110000110"; -- -0.10368266567554635
	pesos_i(418) := b"0000000000000000_0000000000000000_0000001101000001_0001110100001101"; -- 0.012712302954334972
	pesos_i(419) := b"0000000000000000_0000000000000000_0000011101110100_1001110011110011"; -- 0.02912312447425208
	pesos_i(420) := b"0000000000000000_0000000000000000_0010011101001010_1011001011110110"; -- 0.15348356725721085
	pesos_i(421) := b"1111111111111111_1111111111111111_1111100001011001_1110000010001000"; -- -0.029878584772387137
	pesos_i(422) := b"1111111111111111_1111111111111111_1111110001110001_1100100010011101"; -- -0.013888799302550705
	pesos_i(423) := b"1111111111111111_1111111111111111_1101111100010010_0101010111000001"; -- -0.1286264804008226
	pesos_i(424) := b"0000000000000000_0000000000000000_0010101011010110_1110000111011011"; -- 0.1673413427926362
	pesos_i(425) := b"0000000000000000_0000000000000000_0001110010010010_0110100111001010"; -- 0.1116090887378898
	pesos_i(426) := b"1111111111111111_1111111111111111_1101111100111110_1000110011001110"; -- -0.12795181236954603
	pesos_i(427) := b"1111111111111111_1111111111111111_1111100100101011_1111100100111100"; -- -0.02667276664559972
	pesos_i(428) := b"1111111111111111_1111111111111111_1111010110101111_0011000000100001"; -- -0.04029559323789816
	pesos_i(429) := b"0000000000000000_0000000000000000_0010000111101000_0111111001101000"; -- 0.13245382353281748
	pesos_i(430) := b"1111111111111111_1111111111111111_1110110110010001_1110011111110010"; -- -0.07199240066559254
	pesos_i(431) := b"1111111111111111_1111111111111111_1101111110000110_0000001010100011"; -- -0.12686141505364562
	pesos_i(432) := b"0000000000000000_0000000000000000_0001110010101011_1110101010111111"; -- 0.11199824494593577
	pesos_i(433) := b"0000000000000000_0000000000000000_0000000100000110_1011101010101000"; -- 0.0040089284156177565
	pesos_i(434) := b"1111111111111111_1111111111111111_1111100110100110_1010000000000000"; -- -0.024801254245832766
	pesos_i(435) := b"1111111111111111_1111111111111111_1101010011010000_0000110001111101"; -- -0.16870042763184265
	pesos_i(436) := b"0000000000000000_0000000000000000_0001111001101111_1010110111111001"; -- 0.11889159513262802
	pesos_i(437) := b"0000000000000000_0000000000000000_0010100110010000_1100001100011111"; -- 0.16236514575132088
	pesos_i(438) := b"1111111111111111_1111111111111111_1110011000111011_1111101010000010"; -- -0.10064730004000418
	pesos_i(439) := b"0000000000000000_0000000000000000_0000100111011101_1011011110110000"; -- 0.038539390937635615
	pesos_i(440) := b"0000000000000000_0000000000000000_0000010001000101_0011101011101111"; -- 0.016681369155181924
	pesos_i(441) := b"1111111111111111_1111111111111111_1110111011010011_0111111010010101"; -- -0.06708535059094041
	pesos_i(442) := b"0000000000000000_0000000000000000_0000101100100110_0100111100110110"; -- 0.04355330535859024
	pesos_i(443) := b"1111111111111111_1111111111111111_1111001000110011_0110001010100010"; -- -0.053903422764227986
	pesos_i(444) := b"1111111111111111_1111111111111111_1110001101100010_0100101011100000"; -- -0.11178142584134691
	pesos_i(445) := b"0000000000000000_0000000000000000_0010010010011110_1110110010111010"; -- 0.14304999856516137
	pesos_i(446) := b"0000000000000000_0000000000000000_0010011000001111_0010100110001010"; -- 0.14866885767434074
	pesos_i(447) := b"0000000000000000_0000000000000000_0000010000001110_0111011110110111"; -- 0.015845758719110942
	pesos_i(448) := b"1111111111111111_1111111111111111_1101100001011111_1111100111000001"; -- -0.1547855286127893
	pesos_i(449) := b"0000000000000000_0000000000000000_0001110001001100_0001010110011100"; -- 0.11053595592616185
	pesos_i(450) := b"0000000000000000_0000000000000000_0010010111011000_0101001010011010"; -- 0.14783207197937667
	pesos_i(451) := b"1111111111111111_1111111111111111_1101111001001110_0001111110110010"; -- -0.13162042528034507
	pesos_i(452) := b"1111111111111111_1111111111111111_1111111000010000_1010011011001010"; -- -0.007558417936643094
	pesos_i(453) := b"0000000000000000_0000000000000000_0001010110011100_1001010010001000"; -- 0.08442047434679402
	pesos_i(454) := b"0000000000000000_0000000000000000_0010000110111101_1010011110011011"; -- 0.1318001512077536
	pesos_i(455) := b"0000000000000000_0000000000000000_0000101001010011_0100101001111111"; -- 0.0403334198789215
	pesos_i(456) := b"0000000000000000_0000000000000000_0001011111000011_0010110100010110"; -- 0.09282190111753583
	pesos_i(457) := b"1111111111111111_1111111111111111_1110001101110111_1010110000010111"; -- -0.11145519673671017
	pesos_i(458) := b"0000000000000000_0000000000000000_0000110111100110_1011100011000001"; -- 0.054301783647237874
	pesos_i(459) := b"0000000000000000_0000000000000000_0010010110111111_0001010000000000"; -- 0.1474468707803997
	pesos_i(460) := b"1111111111111111_1111111111111111_1111111111001011_1011000001000000"; -- -0.0007982105385125469
	pesos_i(461) := b"1111111111111111_1111111111111111_1101100011110110_0101110110000000"; -- -0.1524907647682592
	pesos_i(462) := b"1111111111111111_1111111111111111_1111010101101011_0001111001010111"; -- -0.04133425113172055
	pesos_i(463) := b"0000000000000000_0000000000000000_0001011100000100_1111110111101010"; -- 0.08991991969070265
	pesos_i(464) := b"1111111111111111_1111111111111111_1111011110100111_1101010100001101"; -- -0.03259533332382636
	pesos_i(465) := b"0000000000000000_0000000000000000_0001001011111101_0001101010101011"; -- 0.07417456312765405
	pesos_i(466) := b"1111111111111111_1111111111111111_1110110100011000_1001000111111011"; -- -0.07384383802183012
	pesos_i(467) := b"1111111111111111_1111111111111111_1110010001011101_0101101100101110"; -- -0.10795049785205722
	pesos_i(468) := b"1111111111111111_1111111111111111_1111100111010101_0001111001011100"; -- -0.02409181846913631
	pesos_i(469) := b"1111111111111111_1111111111111111_1110001001011001_0100001110111111"; -- -0.11582542984447865
	pesos_i(470) := b"1111111111111111_1111111111111111_1110010011111000_0010010100101111"; -- -0.10558860401959302
	pesos_i(471) := b"0000000000000000_0000000000000000_0001110001001100_1111001100100011"; -- 0.1105491601286545
	pesos_i(472) := b"1111111111111111_1111111111111111_1110111001000011_1111100110100000"; -- -0.06927528225440947
	pesos_i(473) := b"1111111111111111_1111111111111111_1110010010000101_0100110010000101"; -- -0.10734102017554682
	pesos_i(474) := b"1111111111111111_1111111111111111_1101111101001010_1011011100010110"; -- -0.12776618682681798
	pesos_i(475) := b"1111111111111111_1111111111111111_1111011100001011_0100010101011111"; -- -0.03498426846722607
	pesos_i(476) := b"0000000000000000_0000000000000000_0000001011011100_1011100000101011"; -- 0.011180410945773564
	pesos_i(477) := b"1111111111111111_1111111111111111_1110100011011010_1101110011111110"; -- -0.09041041176759321
	pesos_i(478) := b"1111111111111111_1111111111111111_1110100010110000_1110011101111011"; -- -0.09105065581864313
	pesos_i(479) := b"1111111111111111_1111111111111111_1110111110001100_0100001100111000"; -- -0.06426601303260066
	pesos_i(480) := b"1111111111111111_1111111111111111_1111110110000100_1100001100101011"; -- -0.009692956888897264
	pesos_i(481) := b"0000000000000000_0000000000000000_0000000111000011_1001011110111011"; -- 0.00689075771661721
	pesos_i(482) := b"0000000000000000_0000000000000000_0010101110111101_1101011011100010"; -- 0.17086546924876642
	pesos_i(483) := b"0000000000000000_0000000000000000_0000111001000101_0010001101010111"; -- 0.055742462824480726
	pesos_i(484) := b"0000000000000000_0000000000000000_0000011101100101_1100101011110001"; -- 0.02889698400832646
	pesos_i(485) := b"0000000000000000_0000000000000000_0000010000011110_0101101101001000"; -- 0.01608820455163974
	pesos_i(486) := b"0000000000000000_0000000000000000_0000100000100101_1001000101000111"; -- 0.03182323451337561
	pesos_i(487) := b"0000000000000000_0000000000000000_0001001101100011_0011110010011101"; -- 0.07573298299870981
	pesos_i(488) := b"0000000000000000_0000000000000000_0000001000001111_1101100111101110"; -- 0.008054371426483325
	pesos_i(489) := b"0000000000000000_0000000000000000_0001010001100001_0111111001010100"; -- 0.07961263238402785
	pesos_i(490) := b"1111111111111111_1111111111111111_1111000110100100_1110100000101111"; -- -0.056077469487985275
	pesos_i(491) := b"0000000000000000_0000000000000000_0001111100111111_1111111100111110"; -- 0.12207026733572358
	pesos_i(492) := b"0000000000000000_0000000000000000_0010110011000100_0011011010010010"; -- 0.17486897535446905
	pesos_i(493) := b"1111111111111111_1111111111111111_1110000010100111_1010010100001110"; -- -0.1224419441168312
	pesos_i(494) := b"1111111111111111_1111111111111111_1110100110101111_1001101100010011"; -- -0.08716421870425854
	pesos_i(495) := b"0000000000000000_0000000000000000_0001001010111111_0100011101000110"; -- 0.07323117703327478
	pesos_i(496) := b"0000000000000000_0000000000000000_0000101010000101_0101011011101101"; -- 0.04109710010364928
	pesos_i(497) := b"1111111111111111_1111111111111111_1101111110101110_0011010011100011"; -- -0.12624806850274292
	pesos_i(498) := b"1111111111111111_1111111111111111_1110100001101100_0111110001001100"; -- -0.0920946421798213
	pesos_i(499) := b"1111111111111111_1111111111111111_1101011111101001_0001100000001111"; -- -0.15659951825596197
	pesos_i(500) := b"1111111111111111_1111111111111111_1101110000101010_0100110000101011"; -- -0.1399795909631116
	pesos_i(501) := b"1111111111111111_1111111111111111_1111010100000100_1100100001000000"; -- -0.04289577902134613
	pesos_i(502) := b"0000000000000000_0000000000000000_0000000100011000_1000110111011001"; -- 0.004280915644958536
	pesos_i(503) := b"1111111111111111_1111111111111111_1110111000011100_1111111011100000"; -- -0.06987006227498932
	pesos_i(504) := b"1111111111111111_1111111111111111_1111001110111110_1100000101010010"; -- -0.04787055729533188
	pesos_i(505) := b"1111111111111111_1111111111111111_1110101100011011_0101111101010101"; -- -0.08161358035428365
	pesos_i(506) := b"0000000000000000_0000000000000000_0001010001101111_1111010001110000"; -- 0.0798332952975451
	pesos_i(507) := b"0000000000000000_0000000000000000_0001000010111010_0100100100101111"; -- 0.06534249678763837
	pesos_i(508) := b"0000000000000000_0000000000000000_0001100011100010_0100101101011001"; -- 0.09720297739323326
	pesos_i(509) := b"0000000000000000_0000000000000000_0000111110111110_0100101100010100"; -- 0.061497394882523114
	pesos_i(510) := b"0000000000000000_0000000000000000_0001101100011101_0010100111011010"; -- 0.10591374953740862
	pesos_i(511) := b"1111111111111111_1111111111111111_1110010111011110_0001100110000100"; -- -0.10207977797779934
	pesos_i(512) := b"1111111111111111_1111111111111111_1101101001101100_0100001111100100"; -- -0.1467855042647172
	pesos_i(513) := b"1111111111111111_1111111111111111_1101111011101000_0110011011101011"; -- -0.12926632663153761
	pesos_i(514) := b"1111111111111111_1111111111111111_1111000001001010_1011100111001100"; -- -0.06135977531893874
	pesos_i(515) := b"1111111111111111_1111111111111111_1111100101110110_0001011010001101"; -- -0.025541868750453025
	pesos_i(516) := b"1111111111111111_1111111111111111_1111001010000010_1101110110001000"; -- -0.05269065314150582
	pesos_i(517) := b"0000000000000000_0000000000000000_0000000000111100_0001111001101110"; -- 0.0009173411664294939
	pesos_i(518) := b"0000000000000000_0000000000000000_0010000010110000_1101101100010101"; -- 0.12769860515348908
	pesos_i(519) := b"1111111111111111_1111111111111111_1110111100111000_1110100000010101"; -- -0.06553792453729719
	pesos_i(520) := b"0000000000000000_0000000000000000_0000001101100101_1001101111001110"; -- 0.013269174463295036
	pesos_i(521) := b"0000000000000000_0000000000000000_0001000110101000_1010000110100001"; -- 0.06897936050682361
	pesos_i(522) := b"0000000000000000_0000000000000000_0000010010000001_1111111100100110"; -- 0.017608591749571956
	pesos_i(523) := b"1111111111111111_1111111111111111_1111100011010101_1011000010011100"; -- -0.027989351101863832
	pesos_i(524) := b"1111111111111111_1111111111111111_1101010000100000_0000000000100010"; -- -0.17138671085185186
	pesos_i(525) := b"1111111111111111_1111111111111111_1111110100011111_0101110111111010"; -- -0.011240126057702228
	pesos_i(526) := b"0000000000000000_0000000000000000_0001000001100100_1101110011101111"; -- 0.06403904748361441
	pesos_i(527) := b"0000000000000000_0000000000000000_0001000001110001_0001100110001110"; -- 0.06422576626080553
	pesos_i(528) := b"1111111111111111_1111111111111111_1111000100001011_0000100011111011"; -- -0.058425368154483986
	pesos_i(529) := b"1111111111111111_1111111111111111_1110101111001011_0000100101110111"; -- -0.07893315157474573
	pesos_i(530) := b"1111111111111111_1111111111111111_1101110100011110_0101010011101011"; -- -0.13625592481107257
	pesos_i(531) := b"1111111111111111_1111111111111111_1101111011001001_1010110110100000"; -- -0.12973513454438293
	pesos_i(532) := b"0000000000000000_0000000000000000_0000101001110011_1001110101000100"; -- 0.04082663455117994
	pesos_i(533) := b"1111111111111111_1111111111111111_1110100010101011_0111110001011000"; -- -0.09113333555008954
	pesos_i(534) := b"0000000000000000_0000000000000000_0001000010101101_1101000000001101"; -- 0.06515217133932626
	pesos_i(535) := b"1111111111111111_1111111111111111_1110101110100101_1011100001100001"; -- -0.07950255991459496
	pesos_i(536) := b"1111111111111111_1111111111111111_1111110010111100_0111010011001001"; -- -0.012749386684036268
	pesos_i(537) := b"1111111111111111_1111111111111111_1110110011111001_0111000100101000"; -- -0.07431881693304067
	pesos_i(538) := b"1111111111111111_1111111111111111_1110111111110010_1000010100010101"; -- -0.0627056906922364
	pesos_i(539) := b"0000000000000000_0000000000000000_0000100011010101_0110011001101000"; -- 0.034506225884029615
	pesos_i(540) := b"1111111111111111_1111111111111111_1110011011011010_0011101000001100"; -- -0.09823262403377521
	pesos_i(541) := b"0000000000000000_0000000000000000_0010010110101011_1000111111001100"; -- 0.1471490739352665
	pesos_i(542) := b"1111111111111111_1111111111111111_1110111111101010_0011111101100011"; -- -0.06283191513409692
	pesos_i(543) := b"1111111111111111_1111111111111111_1110111110111100_1001101101010100"; -- -0.0635283392817023
	pesos_i(544) := b"1111111111111111_1111111111111111_1101001101000111_1001011001101111"; -- -0.17468890937677864
	pesos_i(545) := b"0000000000000000_0000000000000000_0001010000011100_1111001011110110"; -- 0.07856672759128715
	pesos_i(546) := b"1111111111111111_1111111111111111_1111101001011100_0100011101101000"; -- -0.02202943529323978
	pesos_i(547) := b"1111111111111111_1111111111111111_1111100101000101_0010110111000111"; -- -0.02628816500651653
	pesos_i(548) := b"0000000000000000_0000000000000000_0000001001100000_0011111101100011"; -- 0.00928112184249869
	pesos_i(549) := b"1111111111111111_1111111111111111_1111111110000001_1101000100001011"; -- -0.0019254062214281672
	pesos_i(550) := b"0000000000000000_0000000000000000_0000001001101111_0100011000001010"; -- 0.009510400131147281
	pesos_i(551) := b"0000000000000000_0000000000000000_0000000010001000_0100111100111001"; -- 0.0020799172482235673
	pesos_i(552) := b"1111111111111111_1111111111111111_1111001001101110_1001000001000010"; -- -0.05300043482858724
	pesos_i(553) := b"1111111111111111_1111111111111111_1111101010010011_1000001101111110"; -- -0.021186620524544585
	pesos_i(554) := b"1111111111111111_1111111111111111_1101010010010110_1100000010010111"; -- -0.16957470232980207
	pesos_i(555) := b"1111111111111111_1111111111111111_1101101000010111_1001111100101110"; -- -0.14807705992114134
	pesos_i(556) := b"1111111111111111_1111111111111111_1101110000000001_1111101110001001"; -- -0.14059474855940732
	pesos_i(557) := b"1111111111111111_1111111111111111_1110100110011001_0100110101011001"; -- -0.08750454506719604
	pesos_i(558) := b"1111111111111111_1111111111111111_1111100010001010_0111011001110110"; -- -0.0291372262261329
	pesos_i(559) := b"1111111111111111_1111111111111111_1110000101100100_1011011101001011"; -- -0.1195569459379613
	pesos_i(560) := b"1111111111111111_1111111111111111_1110100100101111_1100001000101011"; -- -0.08911501363695222
	pesos_i(561) := b"1111111111111111_1111111111111111_1110100011010111_0111110110001001"; -- -0.0904618778110664
	pesos_i(562) := b"1111111111111111_1111111111111111_1111000010110010_1001110011010110"; -- -0.05977458749282203
	pesos_i(563) := b"0000000000000000_0000000000000000_0010100101010110_0011001001100011"; -- 0.1614715092104108
	pesos_i(564) := b"1111111111111111_1111111111111111_1111111101010010_1010001011110000"; -- -0.0026453173571489466
	pesos_i(565) := b"1111111111111111_1111111111111111_1110101101011010_0110001001100101"; -- -0.08065209416845909
	pesos_i(566) := b"0000000000000000_0000000000000000_0000011001011100_1101001100101110"; -- 0.024853895846472445
	pesos_i(567) := b"0000000000000000_0000000000000000_0010000001011110_1000111100011001"; -- 0.126442855495957
	pesos_i(568) := b"0000000000000000_0000000000000000_0001100101000101_1111010110010010"; -- 0.0987237435158195
	pesos_i(569) := b"0000000000000000_0000000000000000_0000010001011011_1000101101111111"; -- 0.017021864493069402
	pesos_i(570) := b"0000000000000000_0000000000000000_0001101101011000_1101000011110101"; -- 0.10682397824266601
	pesos_i(571) := b"1111111111111111_1111111111111111_1111000100111101_0111111111000010"; -- -0.05765534888535404
	pesos_i(572) := b"0000000000000000_0000000000000000_0010010011111001_1000000101000110"; -- 0.1444321437807051
	pesos_i(573) := b"1111111111111111_1111111111111111_1111011111111111_1101100110111000"; -- -0.031252281657342035
	pesos_i(574) := b"0000000000000000_0000000000000000_0000111110111101_0100011101101010"; -- 0.06148191776217262
	pesos_i(575) := b"1111111111111111_1111111111111111_1110011010011100_0000011010111110"; -- -0.09918172713760756
	pesos_i(576) := b"0000000000000000_0000000000000000_0001011110011001_0010110110111111"; -- 0.09218107151650659
	pesos_i(577) := b"0000000000000000_0000000000000000_0000100101100001_0001100011101111"; -- 0.036637838805157114
	pesos_i(578) := b"0000000000000000_0000000000000000_0000101011001000_0001101100111010"; -- 0.042115880569898984
	pesos_i(579) := b"0000000000000000_0000000000000000_0001110001100100_0100111011110001"; -- 0.11090558419750761
	pesos_i(580) := b"0000000000000000_0000000000000000_0001100101110111_1111001000111111"; -- 0.09948648479386951
	pesos_i(581) := b"0000000000000000_0000000000000000_0001110111100100_1111010111111001"; -- 0.11677491493391493
	pesos_i(582) := b"0000000000000000_0000000000000000_0001100000100110_1101110101100000"; -- 0.09434302891809049
	pesos_i(583) := b"1111111111111111_1111111111111111_1111001000001100_0000110111111101"; -- -0.05450356080045829
	pesos_i(584) := b"0000000000000000_0000000000000000_0000100001001110_0100110100100000"; -- 0.03244478257463834
	pesos_i(585) := b"0000000000000000_0000000000000000_0001110011000101_0000011000000101"; -- 0.11238134023393095
	pesos_i(586) := b"0000000000000000_0000000000000000_0010100000111110_1101011101110001"; -- 0.15720888614777234
	pesos_i(587) := b"0000000000000000_0000000000000000_0000101011011000_1100111000010000"; -- 0.04237068075691585
	pesos_i(588) := b"1111111111111111_1111111111111111_1110011101100100_1111111010001110"; -- -0.0961151984339132
	pesos_i(589) := b"0000000000000000_0000000000000000_0001001100011011_1111101110011110"; -- 0.07464573489312536
	pesos_i(590) := b"0000000000000000_0000000000000000_0001001100101010_0010111110011011"; -- 0.07486245667711905
	pesos_i(591) := b"0000000000000000_0000000000000000_0010010001110010_0011110110010001"; -- 0.14236817150228598
	pesos_i(592) := b"1111111111111111_1111111111111111_1110101011100010_0100011101100011"; -- -0.08248475874022507
	pesos_i(593) := b"0000000000000000_0000000000000000_0010000111100010_0110001110011011"; -- 0.1323606732649876
	pesos_i(594) := b"0000000000000000_0000000000000000_0001010110111010_0001101010111111"; -- 0.08487097899252823
	pesos_i(595) := b"0000000000000000_0000000000000000_0001101011001010_0011001010100110"; -- 0.10464779420954586
	pesos_i(596) := b"1111111111111111_1111111111111111_1101110111000001_0110010011101000"; -- -0.13376778932384895
	pesos_i(597) := b"1111111111111111_1111111111111111_1111111111001101_1100110111111101"; -- -0.0007659204077666541
	pesos_i(598) := b"0000000000000000_0000000000000000_0010001100000011_0001000010000011"; -- 0.13676551044386692
	pesos_i(599) := b"1111111111111111_1111111111111111_1101001100010001_0111010011011011"; -- -0.17551488538513038
	pesos_i(600) := b"1111111111111111_1111111111111111_1100100000000000_0111100110100010"; -- -0.21874275013880887
	pesos_i(601) := b"1111111111111111_1111111111111111_1101011000011110_0100000111001100"; -- -0.1636008145168789
	pesos_i(602) := b"0000000000000000_0000000000000000_0001010011110101_0110100111111111"; -- 0.0818697211760018
	pesos_i(603) := b"0000000000000000_0000000000000000_0001011110110000_1000001011010110"; -- 0.09253709534722872
	pesos_i(604) := b"0000000000000000_0000000000000000_0000110101110100_0010010001001110"; -- 0.05255343338999171
	pesos_i(605) := b"0000000000000000_0000000000000000_0000111010000010_0101011101100110"; -- 0.05667635189975874
	pesos_i(606) := b"1111111111111111_1111111111111111_1111000111000011_1001000011001001"; -- -0.05560965617716906
	pesos_i(607) := b"0000000000000000_0000000000000000_0010011010010010_1010001010010001"; -- 0.15067497300814817
	pesos_i(608) := b"1111111111111111_1111111111111111_1101111010110011_1110000001111011"; -- -0.13006779675757515
	pesos_i(609) := b"0000000000000000_0000000000000000_0000100000001110_0101101111110011"; -- 0.03146910363986294
	pesos_i(610) := b"1111111111111111_1111111111111111_1101001000110100_0010110100100000"; -- -0.17889135335224474
	pesos_i(611) := b"0000000000000000_0000000000000000_0000000001111101_0100001011101111"; -- 0.0019113381796248133
	pesos_i(612) := b"1111111111111111_1111111111111111_1111101010100110_0000100101111110"; -- -0.02090397533547577
	pesos_i(613) := b"1111111111111111_1111111111111111_1101101111101100_1010101011111001"; -- -0.14091998511383602
	pesos_i(614) := b"1111111111111111_1111111111111111_1110110111010110_1101001111011010"; -- -0.0709407417625665
	pesos_i(615) := b"0000000000000000_0000000000000000_0001000100001101_0001011010100010"; -- 0.06660596326256904
	pesos_i(616) := b"1111111111111111_1111111111111111_1110010101001000_1010010100100011"; -- -0.1043602742268615
	pesos_i(617) := b"1111111111111111_1111111111111111_1111110010010110_1011101011001000"; -- -0.0133250485467273
	pesos_i(618) := b"0000000000000000_0000000000000000_0010001101010010_1111011001011100"; -- 0.13798465487416472
	pesos_i(619) := b"1111111111111111_1111111111111111_1101110010010010_1101011100000101"; -- -0.13838440062769924
	pesos_i(620) := b"1111111111111111_1111111111111111_1110101110001010_0100010000011101"; -- -0.07992147729130555
	pesos_i(621) := b"0000000000000000_0000000000000000_0010001111001001_1100010000010010"; -- 0.1397974533179754
	pesos_i(622) := b"0000000000000000_0000000000000000_0000001101011100_0011100110101000"; -- 0.013125995059488908
	pesos_i(623) := b"0000000000000000_0000000000000000_0001001100111101_1011110010001001"; -- 0.07516077376111335
	pesos_i(624) := b"1111111111111111_1111111111111111_1110011111100100_0010100110110100"; -- -0.09417476032538004
	pesos_i(625) := b"1111111111111111_1111111111111111_1110110101011111_0110100001000110"; -- -0.07276294990260536
	pesos_i(626) := b"1111111111111111_1111111111111111_1111001010001011_0110110010100101"; -- -0.05256005259781067
	pesos_i(627) := b"0000000000000000_0000000000000000_0001011000001010_1111110010101101"; -- 0.08610514851606561
	pesos_i(628) := b"1111111111111111_1111111111111111_1101011111001001_0111110011100101"; -- -0.15708178903392847
	pesos_i(629) := b"0000000000000000_0000000000000000_0001000001100011_0010101110010011"; -- 0.06401321734275442
	pesos_i(630) := b"0000000000000000_0000000000000000_0000111001111101_1101110111100100"; -- 0.05660807424985115
	pesos_i(631) := b"1111111111111111_1111111111111111_1110100001100000_0101111101101011"; -- -0.09227946900222339
	pesos_i(632) := b"1111111111111111_1111111111111111_1111110110011000_0101101010100001"; -- -0.009394012243079147
	pesos_i(633) := b"1111111111111111_1111111111111111_1101110010111000_1110100011000001"; -- -0.13780350955054557
	pesos_i(634) := b"1111111111111111_1111111111111111_1111001110010001_1110010110101001"; -- -0.04855503683398945
	pesos_i(635) := b"0000000000000000_0000000000000000_0001011011101110_1110110101001001"; -- 0.08958323502488602
	pesos_i(636) := b"1111111111111111_1111111111111111_1110100111101111_0010010110100100"; -- -0.08619465580122236
	pesos_i(637) := b"0000000000000000_0000000000000000_0000001010111011_1010111010010101"; -- 0.010676299407353372
	pesos_i(638) := b"1111111111111111_1111111111111111_1110000111001001_0010001100101111"; -- -0.11802463639800152
	pesos_i(639) := b"1111111111111111_1111111111111111_1111110111101110_1001100001011111"; -- -0.008078076147435009
	pesos_i(640) := b"1111111111111111_1111111111111111_1110000111010010_0110110010101111"; -- -0.11788292619039466
	pesos_i(641) := b"0000000000000000_0000000000000000_0000011010111001_0111111010001100"; -- 0.026267918650297005
	pesos_i(642) := b"1111111111111111_1111111111111111_1101110111111100_0001101010101110"; -- -0.132871944944185
	pesos_i(643) := b"1111111111111111_1111111111111111_1101010100110100_0000001101100111"; -- -0.16717509028005845
	pesos_i(644) := b"0000000000000000_0000000000000000_0001110010001011_1011000000001011"; -- 0.11150646473389034
	pesos_i(645) := b"0000000000000000_0000000000000000_0001110011101000_1000100011001010"; -- 0.11292319232932217
	pesos_i(646) := b"0000000000000000_0000000000000000_0001010001001000_0110111110101101"; -- 0.07923028921963304
	pesos_i(647) := b"0000000000000000_0000000000000000_0001100010111010_0011111001110111"; -- 0.0965918579053571
	pesos_i(648) := b"0000000000000000_0000000000000000_0000000100001110_0100100111011011"; -- 0.0041242752477173026
	pesos_i(649) := b"1111111111111111_1111111111111111_1110110110101011_0000011010111000"; -- -0.07160909658879022
	pesos_i(650) := b"1111111111111111_1111111111111111_1101011011110110_1001100110010010"; -- -0.16029968446939927
	pesos_i(651) := b"1111111111111111_1111111111111111_1101110111001011_0011001101000000"; -- -0.13361816107449895
	pesos_i(652) := b"1111111111111111_1111111111111111_1110111010000110_0101110010001000"; -- -0.06826230687690157
	pesos_i(653) := b"0000000000000000_0000000000000000_0010101000010011_1000101110111101"; -- 0.16436074599294095
	pesos_i(654) := b"0000000000000000_0000000000000000_0001000101010110_0111011101000110"; -- 0.06772561512928371
	pesos_i(655) := b"1111111111111111_1111111111111111_1111100101101110_1010110110011001"; -- -0.025654935874821306
	pesos_i(656) := b"0000000000000000_0000000000000000_0001101010100101_0111100011000100"; -- 0.10408739832528466
	pesos_i(657) := b"0000000000000000_0000000000000000_0001000110011011_0011010001111001"; -- 0.06877448986654869
	pesos_i(658) := b"1111111111111111_1111111111111111_1111001010110110_0100011010001001"; -- -0.051906196109856105
	pesos_i(659) := b"0000000000000000_0000000000000000_0010100100001010_0110101001011001"; -- 0.16031517664573774
	pesos_i(660) := b"1111111111111111_1111111111111111_1110001111001010_0011011111001100"; -- -0.11019564877886322
	pesos_i(661) := b"1111111111111111_1111111111111111_1111011010011101_1011111011111111"; -- -0.03665548593577314
	pesos_i(662) := b"1111111111111111_1111111111111111_1101010110101111_1000010111000111"; -- -0.16529048807124708
	pesos_i(663) := b"1111111111111111_1111111111111111_1110101100011101_1010010010111010"; -- -0.0815789265695909
	pesos_i(664) := b"1111111111111111_1111111111111111_1110011101010011_1111110010101110"; -- -0.09637470971452403
	pesos_i(665) := b"1111111111111111_1111111111111111_1110000001111001_1101100001100100"; -- -0.12314078862061993
	pesos_i(666) := b"0000000000000000_0000000000000000_0000111111000110_1100011011101100"; -- 0.061626846879996734
	pesos_i(667) := b"0000000000000000_0000000000000000_0001100111111110_1000101001111001"; -- 0.10154023595666369
	pesos_i(668) := b"0000000000000000_0000000000000000_0001110101000010_1001010010001110"; -- 0.11429718464427015
	pesos_i(669) := b"0000000000000000_0000000000000000_0001100100111101_1100000011110101"; -- 0.09859853724033812
	pesos_i(670) := b"0000000000000000_0000000000000000_0010001101100011_0010001010000101"; -- 0.13823142772868108
	pesos_i(671) := b"1111111111111111_1111111111111111_1110001110101110_0101010010100100"; -- -0.11062117564916361
	pesos_i(672) := b"1111111111111111_1111111111111111_1110010011000111_1001001110100110"; -- -0.10632970045784032
	pesos_i(673) := b"1111111111111111_1111111111111111_1101010111010000_1110011101110011"; -- -0.16478112647292587
	pesos_i(674) := b"0000000000000000_0000000000000000_0001100000101101_1101111011001011"; -- 0.09444992508046125
	pesos_i(675) := b"1111111111111111_1111111111111111_1111010101100011_1001100100001011"; -- -0.041449007776505904
	pesos_i(676) := b"1111111111111111_1111111111111111_1111000101000011_1011000011111111"; -- -0.05756086141542242
	pesos_i(677) := b"1111111111111111_1111111111111111_1111101100011110_1100010001110101"; -- -0.019061776629993945
	pesos_i(678) := b"0000000000000000_0000000000000000_0001001000100000_0000101101110000"; -- 0.07080146302492958
	pesos_i(679) := b"0000000000000000_0000000000000000_0010011010010011_1001010011101111"; -- 0.1506894192323837
	pesos_i(680) := b"1111111111111111_1111111111111111_1101011001010010_1110100000010111"; -- -0.162797445730527
	pesos_i(681) := b"0000000000000000_0000000000000000_0000001010001010_0010110010000111"; -- 0.009920866901778111
	pesos_i(682) := b"0000000000000000_0000000000000000_0000010100001110_1111110111100001"; -- 0.019760005428681678
	pesos_i(683) := b"0000000000000000_0000000000000000_0000001011111110_1001010011111010"; -- 0.011697112079924046
	pesos_i(684) := b"0000000000000000_0000000000000000_0001001010010011_1011010101001110"; -- 0.0725663485511953
	pesos_i(685) := b"0000000000000000_0000000000000000_0010011000110001_0010100010001011"; -- 0.14918759728251568
	pesos_i(686) := b"1111111111111111_1111111111111111_1110101001000110_0000000100010111"; -- -0.08486931984357646
	pesos_i(687) := b"0000000000000000_0000000000000000_0000111100101010_0010010100001001"; -- 0.05923682664329342
	pesos_i(688) := b"0000000000000000_0000000000000000_0000110110111010_1010111011111011"; -- 0.05362981433913991
	pesos_i(689) := b"1111111111111111_1111111111111111_1111111101111100_0010010111111010"; -- -0.0020118966563967664
	pesos_i(690) := b"0000000000000000_0000000000000000_0010011000100000_0011001000000110"; -- 0.14892876278465153
	pesos_i(691) := b"1111111111111111_1111111111111111_1110110111011000_0101101000111000"; -- -0.07091747415269874
	pesos_i(692) := b"0000000000000000_0000000000000000_0000110110111100_0100010001011010"; -- 0.053653976529592314
	pesos_i(693) := b"1111111111111111_1111111111111111_1110000110010101_1111101011101011"; -- -0.11880523460303175
	pesos_i(694) := b"1111111111111111_1111111111111111_1110110000101011_0010111111010101"; -- -0.07746602115753938
	pesos_i(695) := b"1111111111111111_1111111111111111_1101111110110101_1111010010111110"; -- -0.12612982130635805
	pesos_i(696) := b"1111111111111111_1111111111111111_1111010110001001_1111000010010100"; -- -0.04086395623394207
	pesos_i(697) := b"1111111111111111_1111111111111111_1111111100101011_0000100000101111"; -- -0.003249634288691343
	pesos_i(698) := b"0000000000000000_0000000000000000_0000100011001010_1011000110011000"; -- 0.03434286087998387
	pesos_i(699) := b"0000000000000000_0000000000000000_0001011101101000_1110011001110010"; -- 0.09144439978079993
	pesos_i(700) := b"1111111111111111_1111111111111111_1110011101111010_1001000011000010"; -- -0.09578604944770384
	pesos_i(701) := b"1111111111111111_1111111111111111_1110101111101000_1001111100110000"; -- -0.07848172268861185
	pesos_i(702) := b"1111111111111111_1111111111111111_1110000000010110_1010110000110100"; -- -0.12465404250368275
	pesos_i(703) := b"0000000000000000_0000000000000000_0000100001100010_0001111000100110"; -- 0.03274715837560119
	pesos_i(704) := b"1111111111111111_1111111111111111_1111001110001100_0010011011101001"; -- -0.048642700218213625
	pesos_i(705) := b"0000000000000000_0000000000000000_0000111101101110_0100011111111111"; -- 0.06027650808261179
	pesos_i(706) := b"1111111111111111_1111111111111111_1101101100111011_0110011101010111"; -- -0.14362482191783002
	pesos_i(707) := b"0000000000000000_0000000000000000_0001010011010011_0000111001111011"; -- 0.08134546755772382
	pesos_i(708) := b"0000000000000000_0000000000000000_0010010010010001_0010011110010000"; -- 0.1428398824966119
	pesos_i(709) := b"1111111111111111_1111111111111111_1101101011000100_1001001100010110"; -- -0.1454380102310973
	pesos_i(710) := b"0000000000000000_0000000000000000_0010001101111011_0000110100010010"; -- 0.13859636010747878
	pesos_i(711) := b"1111111111111111_1111111111111111_1110001010000000_0110000101111101"; -- -0.11522856419015716
	pesos_i(712) := b"1111111111111111_1111111111111111_1111011110111101_1001011011000010"; -- -0.032263352985465746
	pesos_i(713) := b"1111111111111111_1111111111111111_1111001100010010_0001110111111011"; -- -0.050504804932735216
	pesos_i(714) := b"1111111111111111_1111111111111111_1111101000000010_0010000011101011"; -- -0.02340502034202097
	pesos_i(715) := b"1111111111111111_1111111111111111_1110001001100001_1101000010010011"; -- -0.11569496546522161
	pesos_i(716) := b"0000000000000000_0000000000000000_0000100001110011_1000111001000001"; -- 0.033013239677142
	pesos_i(717) := b"0000000000000000_0000000000000000_0010001011010010_0111100100110111"; -- 0.13602407055891375
	pesos_i(718) := b"1111111111111111_1111111111111111_1111101001000011_1001110110111001"; -- -0.02240576021551759
	pesos_i(719) := b"0000000000000000_0000000000000000_0001000011111111_1101100101111110"; -- 0.06640395472260413
	pesos_i(720) := b"0000000000000000_0000000000000000_0000010111110000_0111111110011110"; -- 0.023200965950176955
	pesos_i(721) := b"1111111111111111_1111111111111111_1110111101000010_0010010101101001"; -- -0.06539694002803252
	pesos_i(722) := b"1111111111111111_1111111111111111_1101100100101110_1101110000100000"; -- -0.1516287252327105
	pesos_i(723) := b"1111111111111111_1111111111111111_1110010010110110_1000001000010101"; -- -0.10659014690806184
	pesos_i(724) := b"1111111111111111_1111111111111111_1111111101010001_1110011111110011"; -- -0.0026564628680601737
	pesos_i(725) := b"1111111111111111_1111111111111111_1110110011101101_0001100010001111"; -- -0.0745072031591057
	pesos_i(726) := b"0000000000000000_0000000000000000_0000110101111100_0001000010110100"; -- 0.05267433549449989
	pesos_i(727) := b"1111111111111111_1111111111111111_1110011110000101_0010110001011101"; -- -0.0956241867905778
	pesos_i(728) := b"1111111111111111_1111111111111111_1110100110110111_0101000110110011"; -- -0.08704652198293286
	pesos_i(729) := b"0000000000000000_0000000000000000_0000001000010100_0011001010100001"; -- 0.008120693553469898
	pesos_i(730) := b"1111111111111111_1111111111111111_1101101000110101_0001010001110111"; -- -0.14762756429548693
	pesos_i(731) := b"1111111111111111_1111111111111111_1101011110101101_1110110010110101"; -- -0.15750237075722257
	pesos_i(732) := b"1111111111111111_1111111111111111_1111101000010101_1000111001111101"; -- -0.023108572408034284
	pesos_i(733) := b"1111111111111111_1111111111111111_1101101101110110_1000110010111111"; -- -0.14272232371823262
	pesos_i(734) := b"0000000000000000_0000000000000000_0001000001101000_1001110001001010"; -- 0.06409622972646113
	pesos_i(735) := b"0000000000000000_0000000000000000_0000001100100000_1000101000001010"; -- 0.012215259071398143
	pesos_i(736) := b"0000000000000000_0000000000000000_0010100110000011_0000110001001101"; -- 0.16215588448149046
	pesos_i(737) := b"1111111111111111_1111111111111111_1110011001111100_0011110100101001"; -- -0.09966676474338393
	pesos_i(738) := b"1111111111111111_1111111111111111_1110001011001001_1011111010110100"; -- -0.1141091167119519
	pesos_i(739) := b"1111111111111111_1111111111111111_1110010100100011_1011111101111001"; -- -0.10492327960819146
	pesos_i(740) := b"0000000000000000_0000000000000000_0001000110110010_0110100101111111"; -- 0.06912860244844636
	pesos_i(741) := b"0000000000000000_0000000000000000_0001001110100110_1110001100111101"; -- 0.07676525345404872
	pesos_i(742) := b"0000000000000000_0000000000000000_0000000101101001_0001100101101001"; -- 0.005509937432759739
	pesos_i(743) := b"1111111111111111_1111111111111111_1111001100011110_1000100110001011"; -- -0.05031528817487699
	pesos_i(744) := b"0000000000000000_0000000000000000_0001110000100100_0100001101100111"; -- 0.10992833394470322
	pesos_i(745) := b"0000000000000000_0000000000000000_0010011100011000_0000001110010010"; -- 0.15271017371616158
	pesos_i(746) := b"0000000000000000_0000000000000000_0010011111010111_0001100001000010"; -- 0.15562583550760034
	pesos_i(747) := b"1111111111111111_1111111111111111_1101011000001001_0001000001000111"; -- -0.1639242006856534
	pesos_i(748) := b"1111111111111111_1111111111111111_1101101010101001_0110010111011100"; -- -0.14585269341652166
	pesos_i(749) := b"0000000000000000_0000000000000000_0010100110111000_1000110110010000"; -- 0.16297230492948528
	pesos_i(750) := b"1111111111111111_1111111111111111_1111000101001111_1111011110110100"; -- -0.057373541399587766
	pesos_i(751) := b"0000000000000000_0000000000000000_0000111011000010_0011101100111010"; -- 0.05765123516921208
	pesos_i(752) := b"1111111111111111_1111111111111111_1111101111101010_1101011011110100"; -- -0.015947881097979733
	pesos_i(753) := b"1111111111111111_1111111111111111_1111000001010110_0010101100110110"; -- -0.061185168676039674
	pesos_i(754) := b"0000000000000000_0000000000000000_0001101001000011_0111101111110010"; -- 0.10259222646850347
	pesos_i(755) := b"1111111111111111_1111111111111111_1111001101111010_1110010001110001"; -- -0.0489060614881914
	pesos_i(756) := b"1111111111111111_1111111111111111_1111100100001000_1000000000010110"; -- -0.027214045126740617
	pesos_i(757) := b"1111111111111111_1111111111111111_1110010100110100_0010011011000010"; -- -0.10467298272291901
	pesos_i(758) := b"1111111111111111_1111111111111111_1101110011011011_1011101000110111"; -- -0.13727222582348417
	pesos_i(759) := b"1111111111111111_1111111111111111_1110001001011001_1010100011000111"; -- -0.11581940789541746
	pesos_i(760) := b"1111111111111111_1111111111111111_1110010010110100_1101111101110110"; -- -0.10661509863888854
	pesos_i(761) := b"1111111111111111_1111111111111111_1111010101111001_0010001001010100"; -- -0.04112039045902019
	pesos_i(762) := b"0000000000000000_0000000000000000_0001100001100001_0111110111110111"; -- 0.0952376105648045
	pesos_i(763) := b"0000000000000000_0000000000000000_0001000111101110_0110111110110010"; -- 0.07004449943489251
	pesos_i(764) := b"0000000000000000_0000000000000000_0000011000001010_1011101111001001"; -- 0.02360128083138042
	pesos_i(765) := b"0000000000000000_0000000000000000_0010110110010001_0001101110110011"; -- 0.17799542552193856
	pesos_i(766) := b"0000000000000000_0000000000000000_0001000100000001_1111100111100100"; -- 0.06643640338604018
	pesos_i(767) := b"0000000000000000_0000000000000000_0010011011110001_0100011001111010"; -- 0.15211906883087062
	pesos_i(768) := b"0000000000000000_0000000000000000_0001100111101010_0100110110110111"; -- 0.10123143891352113
	pesos_i(769) := b"0000000000000000_0000000000000000_0000101011101101_1110000000101111"; -- 0.04269219533142286
	pesos_i(770) := b"0000000000000000_0000000000000000_0010010011100011_1010000011101111"; -- 0.1440983374874874
	pesos_i(771) := b"1111111111111111_1111111111111111_1110001001111011_0010000111010111"; -- -0.11530865189506538
	pesos_i(772) := b"0000000000000000_0000000000000000_0000101100001011_1100000101110000"; -- 0.04314812640409229
	pesos_i(773) := b"0000000000000000_0000000000000000_0001011000100101_1001000001100011"; -- 0.08651068127385986
	pesos_i(774) := b"0000000000000000_0000000000000000_0010001100111101_0111101101100000"; -- 0.13765688985209404
	pesos_i(775) := b"1111111111111111_1111111111111111_1111101111111110_0100110110011110"; -- -0.015650891149165833
	pesos_i(776) := b"0000000000000000_0000000000000000_0001110010101100_1011010011001011"; -- 0.11201028785998712
	pesos_i(777) := b"1111111111111111_1111111111111111_1101110011111100_0011011000000011"; -- -0.1367765658479749
	pesos_i(778) := b"0000000000000000_0000000000000000_0001011111111010_1000010110001110"; -- 0.09366640773236273
	pesos_i(779) := b"0000000000000000_0000000000000000_0000010110000100_1110000000001111"; -- 0.02155876508826595
	pesos_i(780) := b"0000000000000000_0000000000000000_0000010100111000_1100001111100000"; -- 0.020397417141956132
	pesos_i(781) := b"0000000000000000_0000000000000000_0000011010010111_1001001001110001"; -- 0.02575030585170747
	pesos_i(782) := b"1111111111111111_1111111111111111_1111101011100100_0100100001111110"; -- -0.019954175170643528
	pesos_i(783) := b"0000000000000000_0000000000000000_0000011011111001_1001101110001111"; -- 0.02724621049033008
	pesos_i(784) := b"1111111111111111_1111111111111111_1111000100101110_1110100001100101"; -- -0.057877993875661615
	pesos_i(785) := b"0000000000000000_0000000000000000_0001111110101001_0000011010101110"; -- 0.1236728835660868
	pesos_i(786) := b"0000000000000000_0000000000000000_0000011010011111_1111101100010010"; -- 0.025878612387488745
	pesos_i(787) := b"0000000000000000_0000000000000000_0001100110000101_0000001110011100"; -- 0.09968588397051477
	pesos_i(788) := b"0000000000000000_0000000000000000_0000101001110011_0110000000000101"; -- 0.04082298391680804
	pesos_i(789) := b"0000000000000000_0000000000000000_0010011001011110_0011100110010001"; -- 0.14987525736442567
	pesos_i(790) := b"1111111111111111_1111111111111111_1111110101101011_0010001010100101"; -- -0.01008399467302579
	pesos_i(791) := b"1111111111111111_1111111111111111_1101100101000011_1111011100100110"; -- -0.1513066800460513
	pesos_i(792) := b"1111111111111111_1111111111111111_1101111110001111_1110111010110100"; -- -0.12671001542057136
	pesos_i(793) := b"0000000000000000_0000000000000000_0000111000000101_0010010111100001"; -- 0.054766051629243834
	pesos_i(794) := b"0000000000000000_0000000000000000_0010011000010001_0111000110000011"; -- 0.14870366523650147
	pesos_i(795) := b"0000000000000000_0000000000000000_0001000010011001_1011000000000101"; -- 0.06484508620672577
	pesos_i(796) := b"1111111111111111_1111111111111111_1111001000001000_1011101101011110"; -- -0.05455426174985817
	pesos_i(797) := b"1111111111111111_1111111111111111_1101111011011110_1010111100011001"; -- -0.1294146121385083
	pesos_i(798) := b"1111111111111111_1111111111111111_1101110001101101_0000000110110001"; -- -0.13896169115463977
	pesos_i(799) := b"0000000000000000_0000000000000000_0010101110001110_0000000111110100"; -- 0.17013561435554272
	pesos_i(800) := b"0000000000000000_0000000000000000_0010000111110001_1111101001101001"; -- 0.13259854377823024
	pesos_i(801) := b"1111111111111111_1111111111111111_1111010001101000_0111111111001010"; -- -0.045280469124948416
	pesos_i(802) := b"0000000000000000_0000000000000000_0000010100111010_0010110110101010"; -- 0.02041898166763824
	pesos_i(803) := b"0000000000000000_0000000000000000_0000101010101101_0111110010110110"; -- 0.04170970386051803
	pesos_i(804) := b"1111111111111111_1111111111111111_1110000100101010_0110011111000101"; -- -0.1204466956023502
	pesos_i(805) := b"0000000000000000_0000000000000000_0010100011100001_0100111010010101"; -- 0.15968791134865198
	pesos_i(806) := b"0000000000000000_0000000000000000_0000111111010010_1001011111101101"; -- 0.06180715115999831
	pesos_i(807) := b"0000000000000000_0000000000000000_0001001010010100_1101001100000111"; -- 0.07258337895761763
	pesos_i(808) := b"0000000000000000_0000000000000000_0001101111100011_0011111001010001"; -- 0.1089362094084397
	pesos_i(809) := b"0000000000000000_0000000000000000_0000010010111010_0010001101110010"; -- 0.018465247390866413
	pesos_i(810) := b"1111111111111111_1111111111111111_1111110111011001_1000011001110000"; -- -0.008399579667631172
	pesos_i(811) := b"1111111111111111_1111111111111111_1110010111100110_1010110011000000"; -- -0.10194893179002287
	pesos_i(812) := b"1111111111111111_1111111111111111_1101101101111000_1001111110010000"; -- -0.14269068466628942
	pesos_i(813) := b"1111111111111111_1111111111111111_1111111111011000_1011011011011001"; -- -0.0005994531069677728
	pesos_i(814) := b"1111111111111111_1111111111111111_1110000001110000_0001111001110111"; -- -0.1232891996932219
	pesos_i(815) := b"0000000000000000_0000000000000000_0000111000000110_0000011111011100"; -- 0.05477952109750873
	pesos_i(816) := b"1111111111111111_1111111111111111_1110000000110011_0111001111100011"; -- -0.12421489432033328
	pesos_i(817) := b"1111111111111111_1111111111111111_1110011110100001_0000000100001110"; -- -0.09519952217631242
	pesos_i(818) := b"0000000000000000_0000000000000000_0000011111000000_0010000100010010"; -- 0.030275408633993965
	pesos_i(819) := b"0000000000000000_0000000000000000_0001010010001110_0111011001011000"; -- 0.08029880192070402
	pesos_i(820) := b"1111111111111111_1111111111111111_1101100101101110_0001010111101010"; -- -0.15066397692013103
	pesos_i(821) := b"1111111111111111_1111111111111111_1111101101100001_0111110111110111"; -- -0.01804363944588249
	pesos_i(822) := b"1111111111111111_1111111111111111_1111011001011100_1001101100110101"; -- -0.0376494403002018
	pesos_i(823) := b"1111111111111111_1111111111111111_1101100000011000_1011110000101000"; -- -0.15587257416581438
	pesos_i(824) := b"0000000000000000_0000000000000000_0001101010000110_1011101010001000"; -- 0.10361829591450292
	pesos_i(825) := b"1111111111111111_1111111111111111_1111000011000111_1101100001001101"; -- -0.059450608418494005
	pesos_i(826) := b"1111111111111111_1111111111111111_1111000100111110_0000001111110100"; -- -0.057647469384336784
	pesos_i(827) := b"1111111111111111_1111111111111111_1110100011010010_1101011101000110"; -- -0.09053282310696484
	pesos_i(828) := b"1111111111111111_1111111111111111_1101011100110101_1001101101010100"; -- -0.15933827596186084
	pesos_i(829) := b"0000000000000000_0000000000000000_0000110001111101_0001000100101101"; -- 0.04878337234808197
	pesos_i(830) := b"1111111111111111_1111111111111111_1110110111110100_1010011001100010"; -- -0.07048568826841611
	pesos_i(831) := b"0000000000000000_0000000000000000_0000000111010111_1100110000000101"; -- 0.007199050154283548
	pesos_i(832) := b"1111111111111111_1111111111111111_1101100000110010_0011100110101101"; -- -0.1554836227428243
	pesos_i(833) := b"1111111111111111_1111111111111111_1111111101001010_0101110110110011"; -- -0.002771514673822089
	pesos_i(834) := b"1111111111111111_1111111111111111_1110000010011111_1001110011001011"; -- -0.12256450692094044
	pesos_i(835) := b"0000000000000000_0000000000000000_0010100000000111_1101111000000010"; -- 0.1563700441166806
	pesos_i(836) := b"0000000000000000_0000000000000000_0000001001000110_1010111100110111"; -- 0.008891058797588523
	pesos_i(837) := b"0000000000000000_0000000000000000_0000000001011010_0011000111011100"; -- 0.0013762629034033322
	pesos_i(838) := b"0000000000000000_0000000000000000_0001011010010011_0101101000001111"; -- 0.08818590985001183
	pesos_i(839) := b"1111111111111111_1111111111111111_1110100010101001_1011000001011000"; -- -0.09116075380854607
	pesos_i(840) := b"0000000000000000_0000000000000000_0010010111001000_0110101110010111"; -- 0.14758942071138234
	pesos_i(841) := b"0000000000000000_0000000000000000_0001110001110001_1100101000000000"; -- 0.11111128322419353
	pesos_i(842) := b"0000000000000000_0000000000000000_0000010110110100_0111000000001110"; -- 0.02228451089764708
	pesos_i(843) := b"1111111111111111_1111111111111111_1101100010001011_0100111101111011"; -- -0.15412429094885396
	pesos_i(844) := b"0000000000000000_0000000000000000_0000110101010010_1001001100110110"; -- 0.0520412451208641
	pesos_i(845) := b"1111111111111111_1111111111111111_1111101001101111_1011000111111001"; -- -0.02173316632823178
	pesos_i(846) := b"1111111111111111_1111111111111111_1111001000001110_1011000001100001"; -- -0.05446336406706381
	pesos_i(847) := b"1111111111111111_1111111111111111_1110101111100001_0000110101011000"; -- -0.07859722714488566
	pesos_i(848) := b"1111111111111111_1111111111111111_1101001100011100_1010011100001011"; -- -0.1753440474737514
	pesos_i(849) := b"0000000000000000_0000000000000000_0001011111100111_0011010010000100"; -- 0.09337166046352766
	pesos_i(850) := b"1111111111111111_1111111111111111_1110100011110101_1010101011011101"; -- -0.09000141249160727
	pesos_i(851) := b"1111111111111111_1111111111111111_1111111001101011_1001000000110000"; -- -0.006171215411176681
	pesos_i(852) := b"0000000000000000_0000000000000000_0010001111001111_1011000110101000"; -- 0.1398879085371876
	pesos_i(853) := b"0000000000000000_0000000000000000_0000110010011000_1100111101111000"; -- 0.04920670195180029
	pesos_i(854) := b"0000000000000000_0000000000000000_0001100011111011_1001000110000010"; -- 0.09758862899835713
	pesos_i(855) := b"1111111111111111_1111111111111111_1110111111110010_1001001001011110"; -- -0.06270489878272228
	pesos_i(856) := b"0000000000000000_0000000000000000_0010110001111001_0000001101101110"; -- 0.17372151780924863
	pesos_i(857) := b"1111111111111111_1111111111111111_1111000000001111_1111110011000011"; -- -0.06225605243326878
	pesos_i(858) := b"0000000000000000_0000000000000000_0010011010011111_1111111110111111"; -- 0.15087889111804242
	pesos_i(859) := b"0000000000000000_0000000000000000_0010101011000110_1000101101111100"; -- 0.16709205416335696
	pesos_i(860) := b"0000000000000000_0000000000000000_0000110001101110_1100110100000111"; -- 0.04856568749309406
	pesos_i(861) := b"0000000000000000_0000000000000000_0010010010111110_1010000100101101"; -- 0.14353377676826728
	pesos_i(862) := b"0000000000000000_0000000000000000_0010010010010011_0101000011101100"; -- 0.14287286522652595
	pesos_i(863) := b"0000000000000000_0000000000000000_0001000000001000_0010011100101110"; -- 0.06262440569953401
	pesos_i(864) := b"0000000000000000_0000000000000000_0010010111001110_1001101001011011"; -- 0.14768376073965436
	pesos_i(865) := b"1111111111111111_1111111111111111_1101010110001111_0110110011111111"; -- -0.16578024646343867
	pesos_i(866) := b"0000000000000000_0000000000000000_0001011101010011_0110111011000100"; -- 0.09111683170128883
	pesos_i(867) := b"0000000000000000_0000000000000000_0010010001001001_1011001101111101"; -- 0.1417495899674546
	pesos_i(868) := b"1111111111111111_1111111111111111_1101110010010111_0100010010010100"; -- -0.1383168351878537
	pesos_i(869) := b"0000000000000000_0000000000000000_0001111010010110_1111111111110010"; -- 0.11949157387302535
	pesos_i(870) := b"1111111111111111_1111111111111111_1110100011000011_0100111110110110"; -- -0.09076978508692062
	pesos_i(871) := b"1111111111111111_1111111111111111_1110011000100110_1000110011001000"; -- -0.10097427470442098
	pesos_i(872) := b"0000000000000000_0000000000000000_0000000101101010_0010111100101001"; -- 0.0055264926982744045
	pesos_i(873) := b"1111111111111111_1111111111111111_1111110011001111_1110011100110101"; -- -0.012452649761955915
	pesos_i(874) := b"1111111111111111_1111111111111111_1111100001101001_0010100110101011"; -- -0.029645343438564526
	pesos_i(875) := b"1111111111111111_1111111111111111_1110111011100100_0110110101111101"; -- -0.06682696999489393
	pesos_i(876) := b"1111111111111111_1111111111111111_1110000100101011_1100000010111100"; -- -0.12042613419922348
	pesos_i(877) := b"1111111111111111_1111111111111111_1111111111100101_1010000001010101"; -- -0.0004024308335276978
	pesos_i(878) := b"0000000000000000_0000000000000000_0000010101100011_1010110110011001"; -- 0.021052217267345276
	pesos_i(879) := b"1111111111111111_1111111111111111_1101110011110111_1010000011001101"; -- -0.1368464946074729
	pesos_i(880) := b"1111111111111111_1111111111111111_1111110100001101_1001110010110110"; -- -0.011511044992317698
	pesos_i(881) := b"0000000000000000_0000000000000000_0010011111000100_1001001100101000"; -- 0.15534324374391767
	pesos_i(882) := b"0000000000000000_0000000000000000_0010010010111011_1101010010100010"; -- 0.14349106756354355
	pesos_i(883) := b"1111111111111111_1111111111111111_1101011110101101_1010010101101010"; -- -0.1575066200502935
	pesos_i(884) := b"0000000000000000_0000000000000000_0010010010110110_0001011111000011"; -- 0.14340351597658177
	pesos_i(885) := b"1111111111111111_1111111111111111_1101011000001010_0000110111000100"; -- -0.16390909163702855
	pesos_i(886) := b"0000000000000000_0000000000000000_0010001011000010_1100110000001100"; -- 0.13578486711433885
	pesos_i(887) := b"1111111111111111_1111111111111111_1111001011001010_1100111100111110"; -- -0.05159287195062949
	pesos_i(888) := b"1111111111111111_1111111111111111_1101110011100011_0110100110111110"; -- -0.13715495204952688
	pesos_i(889) := b"1111111111111111_1111111111111111_1101001100010100_1101011110010110"; -- -0.1754632244040598
	pesos_i(890) := b"0000000000000000_0000000000000000_0010100100101100_1001100001100101"; -- 0.16083672023202436
	pesos_i(891) := b"1111111111111111_1111111111111111_1111110110010011_0001010110011001"; -- -0.009474420742318912
	pesos_i(892) := b"1111111111111111_1111111111111111_1101011000111000_0110110110111000"; -- -0.16320146795567259
	pesos_i(893) := b"1111111111111111_1111111111111111_1111101000001010_1111101110101100"; -- -0.02326991130893088
	pesos_i(894) := b"0000000000000000_0000000000000000_0000001001000101_1000000000011010"; -- 0.00887299193454915
	pesos_i(895) := b"0000000000000000_0000000000000000_0001010111111111_1110010001011111"; -- 0.08593585324911139
	pesos_i(896) := b"0000000000000000_0000000000000000_0000111100011111_0100101101000011"; -- 0.05907125835725449
	pesos_i(897) := b"1111111111111111_1111111111111111_1101010010100100_1101100000100100"; -- -0.1693596756587596
	pesos_i(898) := b"0000000000000000_0000000000000000_0000011101111011_0011011111001010"; -- 0.029223906342966635
	pesos_i(899) := b"1111111111111111_1111111111111111_1111101110011111_1001101000101011"; -- -0.017095913305277877
	pesos_i(900) := b"1111111111111111_1111111111111111_1110101100100000_1000011000110101"; -- -0.0815349694991317
	pesos_i(901) := b"1111111111111111_1111111111111111_1111001001111101_0000010010010001"; -- -0.05277987911795069
	pesos_i(902) := b"1111111111111111_1111111111111111_1101101110001101_1101111000111001"; -- -0.14236651517277493
	pesos_i(903) := b"0000000000000000_0000000000000000_0010101000100100_1101001110101100"; -- 0.1646244330346119
	pesos_i(904) := b"0000000000000000_0000000000000000_0011101011000110_0010100111010101"; -- 0.22958623358574146
	pesos_i(905) := b"1111111111111111_1111111111111111_1111010110010010_0110010001100011"; -- -0.04073498320381372
	pesos_i(906) := b"0000000000000000_0000000000000000_0001110111100101_1100010001000001"; -- 0.11678721032116132
	pesos_i(907) := b"1111111111111111_1111111111111111_1110010111011010_1101110110010000"; -- -0.1021291278731253
	pesos_i(908) := b"1111111111111111_1111111111111111_1111010011000000_1110001000000111"; -- -0.043931840204365
	pesos_i(909) := b"0000000000000000_0000000000000000_0010010101010011_1011110110011000"; -- 0.1458090302453925
	pesos_i(910) := b"1111111111111111_1111111111111111_1110110000010110_0100011011001001"; -- -0.07778508747274657
	pesos_i(911) := b"0000000000000000_0000000000000000_0000000111010100_1100010011011111"; -- 0.007152847807281601
	pesos_i(912) := b"1111111111111111_1111111111111111_1101111100111010_0010111001100001"; -- -0.1280184759493489
	pesos_i(913) := b"0000000000000000_0000000000000000_0010001000111111_1110011000110110"; -- 0.13378752524267293
	pesos_i(914) := b"1111111111111111_1111111111111111_1111011101001101_0100001110110010"; -- -0.03397728836042645
	pesos_i(915) := b"0000000000000000_0000000000000000_0000111000101110_0001101011101011"; -- 0.055391008712254
	pesos_i(916) := b"0000000000000000_0000000000000000_0000001001101110_0111000111011011"; -- 0.009497753128699582
	pesos_i(917) := b"0000000000000000_0000000000000000_0010001000001110_1101110011100111"; -- 0.13303928974559748
	pesos_i(918) := b"0000000000000000_0000000000000000_0010010100000000_0000111000011001"; -- 0.1445320901779372
	pesos_i(919) := b"1111111111111111_1111111111111111_1101110011011001_0010110000110000"; -- -0.13731120909463465
	pesos_i(920) := b"0000000000000000_0000000000000000_0000010001001011_1111000000100100"; -- 0.016783722773346495
	pesos_i(921) := b"0000000000000000_0000000000000000_0000101001111001_0001111101011011"; -- 0.04091068232420833
	pesos_i(922) := b"0000000000000000_0000000000000000_0001011100111110_1000111110100000"; -- 0.09079835563881261
	pesos_i(923) := b"1111111111111111_1111111111111111_1110011100011010_1010011110001100"; -- -0.09724953498151825
	pesos_i(924) := b"0000000000000000_0000000000000000_0001101110010111_1001010110011100"; -- 0.10778174465027257
	pesos_i(925) := b"0000000000000000_0000000000000000_0010010000110110_1110011000100100"; -- 0.14146269208971138
	pesos_i(926) := b"1111111111111111_1111111111111111_1111001100100001_1011000001110011"; -- -0.05026719266297107
	pesos_i(927) := b"0000000000000000_0000000000000000_0000110011000001_1000010111101100"; -- 0.04982792858192803
	pesos_i(928) := b"0000000000000000_0000000000000000_0000110111000101_1111110010110001"; -- 0.05380229295949729
	pesos_i(929) := b"1111111111111111_1111111111111111_1111110001100001_1101010100111001"; -- -0.01413218839382919
	pesos_i(930) := b"0000000000000000_0000000000000000_0010011111100000_1110100100001001"; -- 0.15577560884203054
	pesos_i(931) := b"0000000000000000_0000000000000000_0001000001000000_0110010000111001"; -- 0.0634825361825713
	pesos_i(932) := b"0000000000000000_0000000000000000_0001110111001110_0101001111101111"; -- 0.11642956336614231
	pesos_i(933) := b"0000000000000000_0000000000000000_0001100111011101_1001001100011110"; -- 0.10103721129080441
	pesos_i(934) := b"0000000000000000_0000000000000000_0010001101111000_1110010011011111"; -- 0.13856344651798091
	pesos_i(935) := b"1111111111111111_1111111111111111_1110100001011010_0111101000110010"; -- -0.0923694255552706
	pesos_i(936) := b"0000000000000000_0000000000000000_0001001000001110_0001101000000100"; -- 0.07052767370506591
	pesos_i(937) := b"0000000000000000_0000000000000000_0010010110010111_1000100111110101"; -- 0.1468435499226162
	pesos_i(938) := b"1111111111111111_1111111111111111_1111101011100111_1010110111000010"; -- -0.019902362969685703
	pesos_i(939) := b"1111111111111111_1111111111111111_1110011100111000_1001010111011111"; -- -0.09679282475180707
	pesos_i(940) := b"1111111111111111_1111111111111111_1111011000100000_1110100011100011"; -- -0.03856033761641765
	pesos_i(941) := b"1111111111111111_1111111111111111_1101101100100111_0111110000000010"; -- -0.14392876572199018
	pesos_i(942) := b"0000000000000000_0000000000000000_0000100101110110_0010000000100100"; -- 0.03695870273751159
	pesos_i(943) := b"0000000000000000_0000000000000000_0001111110111101_0001000110110100"; -- 0.12397871632306058
	pesos_i(944) := b"0000000000000000_0000000000000000_0001001011101101_0100010000111000"; -- 0.07393289913185233
	pesos_i(945) := b"1111111111111111_1111111111111111_1110111011010110_1000011010111000"; -- -0.067039089341505
	pesos_i(946) := b"0000000000000000_0000000000000000_0000111000100010_1111011111000100"; -- 0.055221066785211444
	pesos_i(947) := b"0000000000000000_0000000000000000_0000110011011011_0100101011110100"; -- 0.05022114226281256
	pesos_i(948) := b"1111111111111111_1111111111111111_1101101000110010_1001000000100101"; -- -0.14766596892247888
	pesos_i(949) := b"0000000000000000_0000000000000000_0000111101001100_1011111011011011"; -- 0.05976479372814357
	pesos_i(950) := b"1111111111111111_1111111111111111_1111011100101000_1001110011000100"; -- -0.034536554583689094
	pesos_i(951) := b"0000000000000000_0000000000000000_0001000101011110_1010111000000101"; -- 0.06785094858538078
	pesos_i(952) := b"1111111111111111_1111111111111111_1111000100111010_0100100000010011"; -- -0.05770444421669482
	pesos_i(953) := b"1111111111111111_1111111111111111_1111000100001110_1010101011110011"; -- -0.05836993754036631
	pesos_i(954) := b"1111111111111111_1111111111111111_1111010001001000_0010010011001000"; -- -0.04577417488246389
	pesos_i(955) := b"0000000000000000_0000000000000000_0001101001001111_0111100001011100"; -- 0.10277511837839459
	pesos_i(956) := b"1111111111111111_1111111111111111_1111110000011000_0110010100101001"; -- -0.015252759516385014
	pesos_i(957) := b"1111111111111111_1111111111111111_1110010101011110_0000010100011011"; -- -0.1040341194401163
	pesos_i(958) := b"1111111111111111_1111111111111111_1111000000001001_0010100110011011"; -- -0.06236019104817243
	pesos_i(959) := b"1111111111111111_1111111111111111_1110110111100010_1011001100101000"; -- -0.07075958520891974
	pesos_i(960) := b"1111111111111111_1111111111111111_1111001011101110_1111000001100000"; -- -0.05104158084982549
	pesos_i(961) := b"0000000000000000_0000000000000000_0000011001101001_1001111111100111"; -- 0.025049203730892793
	pesos_i(962) := b"1111111111111111_1111111111111111_1101110100100000_1111010110011111"; -- -0.13621582854718584
	pesos_i(963) := b"0000000000000000_0000000000000000_0001011110111010_1011000010010001"; -- 0.09269240883297475
	pesos_i(964) := b"1111111111111111_1111111111111111_1110111001001011_0000110100100100"; -- -0.06916730754443284
	pesos_i(965) := b"0000000000000000_0000000000000000_0000010011010101_0110010101100110"; -- 0.018881165803933394
	pesos_i(966) := b"0000000000000000_0000000000000000_0000000000000101_0001111111000010"; -- 7.818686160492831e-05
	pesos_i(967) := b"1111111111111111_1111111111111111_1110010111011011_0001000011111010"; -- -0.1021260632130975
	pesos_i(968) := b"0000000000000000_0000000000000000_0001111010000001_0111100100010010"; -- 0.11916310025579001
	pesos_i(969) := b"1111111111111111_1111111111111111_1111011110101000_0111110010100010"; -- -0.03258534479611099
	pesos_i(970) := b"1111111111111111_1111111111111111_1110101100100101_1010100010111101"; -- -0.08145661724887733
	pesos_i(971) := b"0000000000000000_0000000000000000_0000011011011000_1000010101101111"; -- 0.026741351627518766
	pesos_i(972) := b"0000000000000000_0000000000000000_0000111101000010_0010110010010100"; -- 0.05960348713865025
	pesos_i(973) := b"0000000000000000_0000000000000000_0001101101101111_1101111101111001"; -- 0.10717579550240319
	pesos_i(974) := b"0000000000000000_0000000000000000_0001111111011011_1010101101010000"; -- 0.12444563583633116
	pesos_i(975) := b"1111111111111111_1111111111111111_1101111111011101_1100101100111110"; -- -0.12552194334543113
	pesos_i(976) := b"0000000000000000_0000000000000000_0001001111111010_0001100100110111"; -- 0.07803495019983334
	pesos_i(977) := b"0000000000000000_0000000000000000_0010101110000010_1011100010001110"; -- 0.16996339283787126
	pesos_i(978) := b"0000000000000000_0000000000000000_0001110110101101_1110110010111010"; -- 0.11593513043204315
	pesos_i(979) := b"1111111111111111_1111111111111111_1101010110010001_0011001011100100"; -- -0.1657531923406096
	pesos_i(980) := b"0000000000000000_0000000000000000_0001110100101111_0100011110010010"; -- 0.11400267901054799
	pesos_i(981) := b"0000000000000000_0000000000000000_0010000101000001_0001100010100111"; -- 0.1298995406527615
	pesos_i(982) := b"1111111111111111_1111111111111111_1111001011100010_1100111111001100"; -- -0.051226627987835116
	pesos_i(983) := b"1111111111111111_1111111111111111_1111111100010010_1011001110000001"; -- -0.0036208925793164933
	pesos_i(984) := b"1111111111111111_1111111111111111_1111101001101110_0000111111110000"; -- -0.021758083247520266
	pesos_i(985) := b"0000000000000000_0000000000000000_0000101001000100_1010001100110110"; -- 0.04010982574881817
	pesos_i(986) := b"0000000000000000_0000000000000000_0000101001000101_1001110001001110"; -- 0.04012467298079332
	pesos_i(987) := b"0000000000000000_0000000000000000_0001000111101010_0110111110000010"; -- 0.06998345291089733
	pesos_i(988) := b"0000000000000000_0000000000000000_0001001101010010_0110001110011111"; -- 0.07547590846664082
	pesos_i(989) := b"0000000000000000_0000000000000000_0000001010100000_0100101000001110"; -- 0.010258320151366643
	pesos_i(990) := b"0000000000000000_0000000000000000_0000001011101000_1011010100101111"; -- 0.01136333843813914
	pesos_i(991) := b"1111111111111111_1111111111111111_1111011010110010_1101110110110101"; -- -0.03633322075317261
	pesos_i(992) := b"1111111111111111_1111111111111111_1101110011011100_0010000011010011"; -- -0.13726610981558343
	pesos_i(993) := b"1111111111111111_1111111111111111_1110011011101101_1001011110001000"; -- -0.09793713512499742
	pesos_i(994) := b"1111111111111111_1111111111111111_1111000011110111_0011110001001111"; -- -0.05872748448924108
	pesos_i(995) := b"1111111111111111_1111111111111111_1110101110100001_0000010111101001"; -- -0.0795742326205354
	pesos_i(996) := b"0000000000000000_0000000000000000_0001000010101001_1101110110110100"; -- 0.06509194987009745
	pesos_i(997) := b"0000000000000000_0000000000000000_0000011100101110_0111101001000010"; -- 0.028052941408019266
	pesos_i(998) := b"1111111111111111_1111111111111111_1110110001100101_0101111100010101"; -- -0.07657819507452159
	pesos_i(999) := b"0000000000000000_0000000000000000_0000111011011101_1100000000111101"; -- 0.05807115071968194
	pesos_i(1000) := b"1111111111111111_1111111111111111_1111101101100110_0010100101111111"; -- -0.017972380163748164
	pesos_i(1001) := b"1111111111111111_1111111111111111_1101111010011000_0011100101101110"; -- -0.13048974103366678
	pesos_i(1002) := b"0000000000000000_0000000000000000_0000010000010001_0011110101101100"; -- 0.015888060330745975
	pesos_i(1003) := b"1111111111111111_1111111111111111_1111010010001110_1001000111101101"; -- -0.04469955408610918
	pesos_i(1004) := b"1111111111111111_1111111111111111_1110110001110000_1001000000111010"; -- -0.07640741909050845
	pesos_i(1005) := b"0000000000000000_0000000000000000_0001000100111010_1001100111001100"; -- 0.06730042686297186
	pesos_i(1006) := b"1111111111111111_1111111111111111_1110011111110101_1010000100000000"; -- -0.09390825041858286
	pesos_i(1007) := b"1111111111111111_1111111111111111_1111101111000000_1111010101110010"; -- -0.016586932770919587
	pesos_i(1008) := b"0000000000000000_0000000000000000_0001100001110100_1001111111100100"; -- 0.09552954976220338
	pesos_i(1009) := b"0000000000000000_0000000000000000_0000100010111000_1001001100100110"; -- 0.034066387882523926
	pesos_i(1010) := b"0000000000000000_0000000000000000_0010100000100010_0001111011000110"; -- 0.1567706329555089
	pesos_i(1011) := b"0000000000000000_0000000000000000_0001101101110110_1010011010110101"; -- 0.10727922359509139
	pesos_i(1012) := b"0000000000000000_0000000000000000_0001001001001100_0100001111111010"; -- 0.07147621980186639
	pesos_i(1013) := b"1111111111111111_1111111111111111_1111110010010011_0001111111101100"; -- -0.013380055372536904
	pesos_i(1014) := b"0000000000000000_0000000000000000_0001101111101000_0001001011110101"; -- 0.10900991888074382
	pesos_i(1015) := b"1111111111111111_1111111111111111_1110101110100101_1101111000000100"; -- -0.07950031663965579
	pesos_i(1016) := b"1111111111111111_1111111111111111_1101110010000000_1001111001101101"; -- -0.1386624320717042
	pesos_i(1017) := b"1111111111111111_1111111111111111_1110011000011010_0100010110110111"; -- -0.10116161615546149
	pesos_i(1018) := b"0000000000000000_0000000000000000_0001101010101101_0001011101100110"; -- 0.10420366511876526
	pesos_i(1019) := b"1111111111111111_1111111111111111_1111100000110100_1001101011011000"; -- -0.030447313471769873
	pesos_i(1020) := b"0000000000000000_0000000000000000_0000010001111111_0001101000001100"; -- 0.01756441865098776
	pesos_i(1021) := b"0000000000000000_0000000000000000_0000100101110011_1010010010101000"; -- 0.03692082504086008
	pesos_i(1022) := b"1111111111111111_1111111111111111_1101101101011110_0101011001111110"; -- -0.14309176841430668
	pesos_i(1023) := b"1111111111111111_1111111111111111_1101101110001100_1001110010101001"; -- -0.1423856818768858
	pesos_i(1024) := b"1111111111111111_1111111111111111_1110100011100000_0011101000101010"; -- -0.09032856443692557
	pesos_i(1025) := b"1111111111111111_1111111111111111_1111000011000010_0000000110011001"; -- -0.05953969969478208
	pesos_i(1026) := b"0000000000000000_0000000000000000_0000111010000110_1000000000111100"; -- 0.05673982108794779
	pesos_i(1027) := b"0000000000000000_0000000000000000_0000001001100111_0000010110110000"; -- 0.00938449435600445
	pesos_i(1028) := b"1111111111111111_1111111111111111_1110011011101100_0010001100011111"; -- -0.09795933231164061
	pesos_i(1029) := b"1111111111111111_1111111111111111_1101011010010011_0011000100001100"; -- -0.16181653470059468
	pesos_i(1030) := b"1111111111111111_1111111111111111_1110010010100110_0000000001000001"; -- -0.10684202596001706
	pesos_i(1031) := b"1111111111111111_1111111111111111_1101111110100100_1111001101001101"; -- -0.12638930670362866
	pesos_i(1032) := b"0000000000000000_0000000000000000_0001001100011011_0111110001011111"; -- 0.07463815038123162
	pesos_i(1033) := b"0000000000000000_0000000000000000_0000010100111101_0001011010000110"; -- 0.020463378574377914
	pesos_i(1034) := b"1111111111111111_1111111111111111_1110011011111100_0100011011110010"; -- -0.09771305643199066
	pesos_i(1035) := b"1111111111111111_1111111111111111_1110101110101100_0101001001110000"; -- -0.07940182473022697
	pesos_i(1036) := b"1111111111111111_1111111111111111_1111100010110011_1111110010100001"; -- -0.02850361897157706
	pesos_i(1037) := b"1111111111111111_1111111111111111_1111100111111111_1110011011110001"; -- -0.023438993705064824
	pesos_i(1038) := b"0000000000000000_0000000000000000_0010101101101100_0011000100110011"; -- 0.16961963179774062
	pesos_i(1039) := b"0000000000000000_0000000000000000_0000100111100110_0010010010001000"; -- 0.03866794899689739
	pesos_i(1040) := b"1111111111111111_1111111111111111_1111111111110001_1100011000011111"; -- -0.00021707279336258267
	pesos_i(1041) := b"0000000000000000_0000000000000000_0010000100100100_1110101001100011"; -- 0.1294695369744795
	pesos_i(1042) := b"0000000000000000_0000000000000000_0010100110001100_0101111000010100"; -- 0.16229808794117895
	pesos_i(1043) := b"0000000000000000_0000000000000000_0010001101110000_1100010000101111"; -- 0.13843942782942786
	pesos_i(1044) := b"1111111111111111_1111111111111111_1111111100010010_0001111111101001"; -- -0.003629689849513825
	pesos_i(1045) := b"1111111111111111_1111111111111111_1110101010100010_1001111010101100"; -- -0.08345611857137936
	pesos_i(1046) := b"1111111111111111_1111111111111111_1101110010110010_0001001001000110"; -- -0.13790784638393988
	pesos_i(1047) := b"0000000000000000_0000000000000000_0000001101111010_1010111000111000"; -- 0.01359070642947646
	pesos_i(1048) := b"1111111111111111_1111111111111111_1101010001010010_1111011100011001"; -- -0.1706090511694843
	pesos_i(1049) := b"1111111111111111_1111111111111111_1110100110110000_1101000100011010"; -- -0.08714573976832792
	pesos_i(1050) := b"0000000000000000_0000000000000000_0000100000100011_0010001110100100"; -- 0.03178618192288777
	pesos_i(1051) := b"1111111111111111_1111111111111111_1101111010111110_0010000110100001"; -- -0.12991132559639343
	pesos_i(1052) := b"1111111111111111_1111111111111111_1101101110001110_0100010011101110"; -- -0.14236039344061782
	pesos_i(1053) := b"1111111111111111_1111111111111111_1111101011001111_1001000100100101"; -- -0.020270279396039384
	pesos_i(1054) := b"0000000000000000_0000000000000000_0001110010101010_0111101011111100"; -- 0.11197632461384245
	pesos_i(1055) := b"0000000000000000_0000000000000000_0000101101111100_1010000000110100"; -- 0.04487038859002951
	pesos_i(1056) := b"1111111111111111_1111111111111111_1110000111000111_1000001001011111"; -- -0.11804948019166725
	pesos_i(1057) := b"0000000000000000_0000000000000000_0001001100011100_0000100101110011"; -- 0.07464655936587491
	pesos_i(1058) := b"0000000000000000_0000000000000000_0010110100100111_0001011011010011"; -- 0.17637770309937786
	pesos_i(1059) := b"1111111111111111_1111111111111111_1101100100011000_1111010010000111"; -- -0.15196296401535708
	pesos_i(1060) := b"1111111111111111_1111111111111111_1101010101101101_0011101111100001"; -- -0.16630197294041765
	pesos_i(1061) := b"1111111111111111_1111111111111111_1111100111010011_0000000011111110"; -- -0.024124086343003188
	pesos_i(1062) := b"0000000000000000_0000000000000000_0000011101101000_1111010101110001"; -- 0.02894529344272202
	pesos_i(1063) := b"0000000000000000_0000000000000000_0010011101110101_0111001100101111"; -- 0.15413589387328527
	pesos_i(1064) := b"0000000000000000_0000000000000000_0001001001011011_1111010100110110"; -- 0.07171566557662035
	pesos_i(1065) := b"1111111111111111_1111111111111111_1101011010111101_0011111111101001"; -- -0.1611747794869651
	pesos_i(1066) := b"1111111111111111_1111111111111111_1111010010101000_0101100010110101"; -- -0.04430623606269351
	pesos_i(1067) := b"0000000000000000_0000000000000000_0001111001001011_0111000010001111"; -- 0.11833861821181754
	pesos_i(1068) := b"1111111111111111_1111111111111111_1101010001111111_0100001111000100"; -- -0.1699330945918244
	pesos_i(1069) := b"0000000000000000_0000000000000000_0001000000011111_0010110100011110"; -- 0.0629757117182275
	pesos_i(1070) := b"0000000000000000_0000000000000000_0010001101101011_1111111101110110"; -- 0.13836666709842182
	pesos_i(1071) := b"1111111111111111_1111111111111111_1100111111001001_1010101000011011"; -- -0.18832909428882977
	pesos_i(1072) := b"0000000000000000_0000000000000000_0001110011110001_0100011101101011"; -- 0.11305662493593491
	pesos_i(1073) := b"1111111111111111_1111111111111111_1111101111000101_1010001010100010"; -- -0.01651557481434249
	pesos_i(1074) := b"0000000000000000_0000000000000000_0010001111000011_0001111010010100"; -- 0.13969603656439078
	pesos_i(1075) := b"0000000000000000_0000000000000000_0000010001001100_1101110111100111"; -- 0.016797894386653148
	pesos_i(1076) := b"1111111111111111_1111111111111111_1110010100111011_0111001011111111"; -- -0.10456162708916245
	pesos_i(1077) := b"1111111111111111_1111111111111111_1110101111001010_1001101010000110"; -- -0.0789397643608438
	pesos_i(1078) := b"1111111111111111_1111111111111111_1111110011100001_1100000011110011"; -- -0.012180271777680291
	pesos_i(1079) := b"1111111111111111_1111111111111111_1110010100000110_0101110000001010"; -- -0.10537171134108889
	pesos_i(1080) := b"1111111111111111_1111111111111111_1110011000010001_1000011111011110"; -- -0.1012950021787031
	pesos_i(1081) := b"1111111111111111_1111111111111111_1111001001010001_1111100001100010"; -- -0.05343673342248135
	pesos_i(1082) := b"0000000000000000_0000000000000000_0001010010111010_0001100100101100"; -- 0.08096463518134084
	pesos_i(1083) := b"0000000000000000_0000000000000000_0001111010100011_1100100011111110"; -- 0.11968666259697604
	pesos_i(1084) := b"1111111111111111_1111111111111111_1111100001111110_0011100111110001"; -- -0.029323938981289793
	pesos_i(1085) := b"1111111111111111_1111111111111111_1110001110110000_0000001000010000"; -- -0.1105955801120072
	pesos_i(1086) := b"1111111111111111_1111111111111111_1110000010000010_0011110111000011"; -- -0.12301267621247923
	pesos_i(1087) := b"1111111111111111_1111111111111111_1111011101010100_0111001100011110"; -- -0.0338676501390177
	pesos_i(1088) := b"1111111111111111_1111111111111111_1111100100100111_0011101111010001"; -- -0.026745091796410908
	pesos_i(1089) := b"1111111111111111_1111111111111111_1111001010111011_1000011100011100"; -- -0.05182605318907886
	pesos_i(1090) := b"0000000000000000_0000000000000000_0001111100011110_1000000010011101"; -- 0.12155917960349656
	pesos_i(1091) := b"0000000000000000_0000000000000000_0000101001101100_1111011100100001"; -- 0.04072517917325051
	pesos_i(1092) := b"1111111111111111_1111111111111111_1101110000000110_1001100110010000"; -- -0.14052429415402032
	pesos_i(1093) := b"1111111111111111_1111111111111111_1101011111001101_1011011100011110"; -- -0.15701728362481115
	pesos_i(1094) := b"0000000000000000_0000000000000000_0000101011011010_1001010010111100"; -- 0.04239778133736867
	pesos_i(1095) := b"0000000000000000_0000000000000000_0001011100100101_1100111110110100"; -- 0.09042070523636037
	pesos_i(1096) := b"0000000000000000_0000000000000000_0011000101010001_0111101100111101"; -- 0.1926495574938786
	pesos_i(1097) := b"1111111111111111_1111111111111111_1110101111111001_1110110100100110"; -- -0.07821767643781058
	pesos_i(1098) := b"0000000000000000_0000000000000000_0000100111110010_0000010000110000"; -- 0.038849126455651126
	pesos_i(1099) := b"0000000000000000_0000000000000000_0000000010111000_0111111111101111"; -- 0.0028152426581372976
	pesos_i(1100) := b"0000000000000000_0000000000000000_0010001110010110_1111100110100001"; -- 0.13902244743325945
	pesos_i(1101) := b"1111111111111111_1111111111111111_1111110000111101_1100110001001001"; -- -0.014682037527355436
	pesos_i(1102) := b"1111111111111111_1111111111111111_1111110101110010_1110011001001101"; -- -0.009965521072980257
	pesos_i(1103) := b"1111111111111111_1111111111111111_1101110110110011_0000110010010110"; -- -0.13398667666061104
	pesos_i(1104) := b"0000000000000000_0000000000000000_0001001010011100_0100100010010011"; -- 0.07269719678306302
	pesos_i(1105) := b"1111111111111111_1111111111111111_1110000011101010_0011100101010110"; -- -0.12142602584053395
	pesos_i(1106) := b"0000000000000000_0000000000000000_0010001101010011_1000101101010010"; -- 0.1379935335568405
	pesos_i(1107) := b"0000000000000000_0000000000000000_0001110011100110_0110010101011001"; -- 0.11289056231194741
	pesos_i(1108) := b"1111111111111111_1111111111111111_1110111011011000_1101010011000110"; -- -0.06700391933014202
	pesos_i(1109) := b"1111111111111111_1111111111111111_1101111101101010_1110001111011101"; -- -0.12727523667100019
	pesos_i(1110) := b"1111111111111111_1111111111111111_1101100010101110_1111101010010001"; -- -0.15358003576826418
	pesos_i(1111) := b"0000000000000000_0000000000000000_0000001111010110_0010011110001110"; -- 0.014986488570928429
	pesos_i(1112) := b"1111111111111111_1111111111111111_1111001001010011_1100010110101111"; -- -0.05340923754245091
	pesos_i(1113) := b"0000000000000000_0000000000000000_0000000000110101_0010011111011001"; -- 0.0008110910342101219
	pesos_i(1114) := b"1111111111111111_1111111111111111_1110101110111001_1100011011111100"; -- -0.07919651356009637
	pesos_i(1115) := b"0000000000000000_0000000000000000_0000110011001111_0000100100010010"; -- 0.05003410992858616
	pesos_i(1116) := b"1111111111111111_1111111111111111_1111100000011010_0010110101110100"; -- -0.030850562252847883
	pesos_i(1117) := b"0000000000000000_0000000000000000_0001011001111101_0011000100010110"; -- 0.0878477744383165
	pesos_i(1118) := b"1111111111111111_1111111111111111_1110101001010111_1000110010011001"; -- -0.08460160516069896
	pesos_i(1119) := b"1111111111111111_1111111111111111_1101010101011101_1100100000010100"; -- -0.166537756968651
	pesos_i(1120) := b"0000000000000000_0000000000000000_0001101111011111_0000011100111101"; -- 0.10887189129332633
	pesos_i(1121) := b"0000000000000000_0000000000000000_0010111000101000_1110011010110011"; -- 0.18031160232529828
	pesos_i(1122) := b"1111111111111111_1111111111111111_1101001111111110_0010100100100111"; -- -0.17190306467607094
	pesos_i(1123) := b"1111111111111111_1111111111111111_1110110001001011_1100000101111110"; -- -0.07696905769042084
	pesos_i(1124) := b"1111111111111111_1111111111111111_1101010001101111_0010010110111100"; -- -0.17017902518814015
	pesos_i(1125) := b"0000000000000000_0000000000000000_0001101011011011_0100111111110001"; -- 0.10490893974346173
	pesos_i(1126) := b"0000000000000000_0000000000000000_0000000110100001_1010000000011111"; -- 0.006372458922348944
	pesos_i(1127) := b"0000000000000000_0000000000000000_0000111110111100_0110000000111100"; -- 0.06146813828500147
	pesos_i(1128) := b"0000000000000000_0000000000000000_0000100110101110_0111101101011100"; -- 0.037818632159293625
	pesos_i(1129) := b"0000000000000000_0000000000000000_0010000110101000_1011000110011010"; -- 0.1314803125047912
	pesos_i(1130) := b"0000000000000000_0000000000000000_0001000111110100_1010001110101111"; -- 0.07013915088006886
	pesos_i(1131) := b"0000000000000000_0000000000000000_0001001010001101_1011010110000111"; -- 0.07247480921086225
	pesos_i(1132) := b"0000000000000000_0000000000000000_0010110001001001_1010100110101001"; -- 0.17299900418476505
	pesos_i(1133) := b"1111111111111111_1111111111111111_1111110001000000_0010111100110011"; -- -0.01464562411768379
	pesos_i(1134) := b"1111111111111111_1111111111111111_1110010100110100_0001110011001100"; -- -0.10467357662665841
	pesos_i(1135) := b"1111111111111111_1111111111111111_1110000111100101_0011011100100101"; -- -0.11759620053103195
	pesos_i(1136) := b"1111111111111111_1111111111111111_1111001010111111_1011011001001001"; -- -0.05176220624740499
	pesos_i(1137) := b"0000000000000000_0000000000000000_0010001010010010_1110100100110011"; -- 0.1350541830636096
	pesos_i(1138) := b"0000000000000000_0000000000000000_0010011000111011_1111000011000001"; -- 0.1493521187030535
	pesos_i(1139) := b"1111111111111111_1111111111111111_1111010001111111_0111010111101111"; -- -0.044930104412139245
	pesos_i(1140) := b"0000000000000000_0000000000000000_0010011100000000_0111100001000111"; -- 0.15235091913087748
	pesos_i(1141) := b"1111111111111111_1111111111111111_1110001100110100_0101001010000011"; -- -0.11248287492695369
	pesos_i(1142) := b"1111111111111111_1111111111111111_1111010001000011_1011100100010011"; -- -0.045841629819462125
	pesos_i(1143) := b"1111111111111111_1111111111111111_1111000001111000_0100000110001010"; -- -0.060665038922627035
	pesos_i(1144) := b"0000000000000000_0000000000000000_0000110101101110_1010011110001110"; -- 0.052469703802084544
	pesos_i(1145) := b"1111111111111111_1111111111111111_1110010011011101_1110011001101110"; -- -0.1059890730161087
	pesos_i(1146) := b"0000000000000000_0000000000000000_0001001000111011_1101000010110010"; -- 0.0712252077413672
	pesos_i(1147) := b"0000000000000000_0000000000000000_0001110100101101_1010000110011111"; -- 0.11397752897390326
	pesos_i(1148) := b"1111111111111111_1111111111111111_1110011111111101_1101111111010001"; -- -0.09378243585348502
	pesos_i(1149) := b"1111111111111111_1111111111111111_1110001101101000_1010100100101000"; -- -0.11168425354795819
	pesos_i(1150) := b"1111111111111111_1111111111111111_1111110100110111_1000000111101010"; -- -0.010871773058921945
	pesos_i(1151) := b"0000000000000000_0000000000000000_0001101100011011_1000111111110001"; -- 0.10588931687143607
	pesos_i(1152) := b"1111111111111111_1111111111111111_1101100100101000_1010000101011011"; -- -0.151723781006828
	pesos_i(1153) := b"1111111111111111_1111111111111111_1101111101001011_1100100100000011"; -- -0.1277498596692663
	pesos_i(1154) := b"1111111111111111_1111111111111111_1101101111101100_0100101100100010"; -- -0.1409256976234094
	pesos_i(1155) := b"0000000000000000_0000000000000000_0010101101010010_1000001000010010"; -- 0.16922772348600176
	pesos_i(1156) := b"0000000000000000_0000000000000000_0000101001111011_0010111001110010"; -- 0.040942099381396445
	pesos_i(1157) := b"0000000000000000_0000000000000000_0010100110010011_0110000001010010"; -- 0.16240503309528392
	pesos_i(1158) := b"0000000000000000_0000000000000000_0001010110000100_1000011100101100"; -- 0.08405346694007342
	pesos_i(1159) := b"1111111111111111_1111111111111111_1110010000110111_1011011010000000"; -- -0.10852488879528924
	pesos_i(1160) := b"0000000000000000_0000000000000000_0010110001010011_0010001110111101"; -- 0.17314360957602207
	pesos_i(1161) := b"0000000000000000_0000000000000000_0001100001011100_0011100101010000"; -- 0.09515722458217998
	pesos_i(1162) := b"1111111111111111_1111111111111111_1111101100001001_1000011000100111"; -- -0.01938592483532288
	pesos_i(1163) := b"0000000000000000_0000000000000000_0000111100101111_0001001111011001"; -- 0.05931209612128081
	pesos_i(1164) := b"1111111111111111_1111111111111111_1111100001000000_0101110100101110"; -- -0.03026788350758984
	pesos_i(1165) := b"0000000000000000_0000000000000000_0010000011000100_1101011100101111"; -- 0.1280035486629998
	pesos_i(1166) := b"1111111111111111_1111111111111111_1110111010001010_0000111010100011"; -- -0.06820591474137168
	pesos_i(1167) := b"1111111111111111_1111111111111111_1111001001111101_0110110110010000"; -- -0.05277362095540221
	pesos_i(1168) := b"1111111111111111_1111111111111111_1110010101111111_1110111100101101"; -- -0.10351662780193693
	pesos_i(1169) := b"0000000000000000_0000000000000000_0010011000110000_1111010111111011"; -- 0.14918458353402483
	pesos_i(1170) := b"1111111111111111_1111111111111111_1111110001001101_1010100100001110"; -- -0.014439996912870345
	pesos_i(1171) := b"1111111111111111_1111111111111111_1111000100011111_1011001000000000"; -- -0.05811011782494319
	pesos_i(1172) := b"1111111111111111_1111111111111111_1101001101011110_1001010100010000"; -- -0.17433803889697153
	pesos_i(1173) := b"0000000000000000_0000000000000000_0000011011000010_1001111011001011"; -- 0.026407169902539076
	pesos_i(1174) := b"1111111111111111_1111111111111111_1101111101010101_1011110000111001"; -- -0.1275980340413998
	pesos_i(1175) := b"0000000000000000_0000000000000000_0000000111010011_0101010011011001"; -- 0.0071309118900866495
	pesos_i(1176) := b"0000000000000000_0000000000000000_0000011110100000_0110011010001100"; -- 0.029791268472834653
	pesos_i(1177) := b"0000000000000000_0000000000000000_0001000000110111_0100000010011100"; -- 0.06334308447432767
	pesos_i(1178) := b"1111111111111111_1111111111111111_1101110101100110_1111010011000010"; -- -0.13514776487863878
	pesos_i(1179) := b"0000000000000000_0000000000000000_0010010010011001_0100110110111010"; -- 0.14296422764606942
	pesos_i(1180) := b"1111111111111111_1111111111111111_1110000111111010_0010011100000100"; -- -0.11727672716140945
	pesos_i(1181) := b"1111111111111111_1111111111111111_1110111000111111_1001000001001101"; -- -0.06934259522212757
	pesos_i(1182) := b"0000000000000000_0000000000000000_0010111000001000_0011111100110100"; -- 0.17981333748431655
	pesos_i(1183) := b"1111111111111111_1111111111111111_1111001000110000_1011100000101101"; -- -0.05394410034485857
	pesos_i(1184) := b"1111111111111111_1111111111111111_1110110011110000_1011101001011010"; -- -0.07445178317997757
	pesos_i(1185) := b"1111111111111111_1111111111111111_1101100011100100_1110001111000001"; -- -0.15275742079850893
	pesos_i(1186) := b"1111111111111111_1111111111111111_1111000010100111_0001111111010111"; -- -0.05994988440734834
	pesos_i(1187) := b"1111111111111111_1111111111111111_1101010100010000_0110101110010011"; -- -0.16771819737017454
	pesos_i(1188) := b"1111111111111111_1111111111111111_1111101011001001_1110101010110001"; -- -0.020356494654439165
	pesos_i(1189) := b"1111111111111111_1111111111111111_1111000111000101_1000100111110111"; -- -0.055579545177170495
	pesos_i(1190) := b"0000000000000000_0000000000000000_0000000111000011_0000010110100110"; -- 0.006882050466636599
	pesos_i(1191) := b"0000000000000000_0000000000000000_0001010011001111_0001111010010010"; -- 0.0812853915426546
	pesos_i(1192) := b"0000000000000000_0000000000000000_0001000111010010_1011110010010100"; -- 0.06962183593117544
	pesos_i(1193) := b"1111111111111111_1111111111111111_1110110100110001_1110101011101100"; -- -0.07345706688726078
	pesos_i(1194) := b"0000000000000000_0000000000000000_0000001100100110_0111100011011111"; -- 0.01230578838827447
	pesos_i(1195) := b"0000000000000000_0000000000000000_0000011011011100_1101101001000101"; -- 0.026807443436267852
	pesos_i(1196) := b"0000000000000000_0000000000000000_0000010111110001_0111110100101111"; -- 0.023216079696937963
	pesos_i(1197) := b"0000000000000000_0000000000000000_0001101000111100_1111010001000101"; -- 0.10249258699486885
	pesos_i(1198) := b"0000000000000000_0000000000000000_0010010111010001_0011100001100111"; -- 0.14772369885715564
	pesos_i(1199) := b"1111111111111111_1111111111111111_1101100001010010_1000010101110001"; -- -0.15499082564813044
	pesos_i(1200) := b"0000000000000000_0000000000000000_0000101100010010_0101000001101100"; -- 0.043248201756958815
	pesos_i(1201) := b"1111111111111111_1111111111111111_1111001101111110_1111011100101000"; -- -0.04884391087751025
	pesos_i(1202) := b"0000000000000000_0000000000000000_0001110110110100_1101101110111100"; -- 0.11604092929092265
	pesos_i(1203) := b"1111111111111111_1111111111111111_1101001011100100_0010011001010101"; -- -0.17620621130896605
	pesos_i(1204) := b"0000000000000000_0000000000000000_0001011010010101_1101000111101001"; -- 0.0882235711423614
	pesos_i(1205) := b"1111111111111111_1111111111111111_1111111000000001_0011001100110010"; -- -0.007794189725503582
	pesos_i(1206) := b"1111111111111111_1111111111111111_1111100010001110_0011100010110000"; -- -0.0290798731881738
	pesos_i(1207) := b"0000000000000000_0000000000000000_0000111000101000_1011100001001010"; -- 0.05530883604318467
	pesos_i(1208) := b"1111111111111111_1111111111111111_1110110101001101_0101110101011100"; -- -0.07303825861391411
	pesos_i(1209) := b"1111111111111111_1111111111111111_1111101001111010_0100111101101011"; -- -0.021571194115815873
	pesos_i(1210) := b"1111111111111111_1111111111111111_1111101111110001_0100001000010001"; -- -0.015849943947757354
	pesos_i(1211) := b"0000000000000000_0000000000000000_0001101011000011_1110110001001110"; -- 0.10455204862427508
	pesos_i(1212) := b"1111111111111111_1111111111111111_1101111001100110_1001001011111111"; -- -0.13124734186819473
	pesos_i(1213) := b"0000000000000000_0000000000000000_0010001100100110_0001111100010000"; -- 0.13730043541987783
	pesos_i(1214) := b"0000000000000000_0000000000000000_0000011000010000_0011001011000011"; -- 0.023684666343298064
	pesos_i(1215) := b"0000000000000000_0000000000000000_0001001001110011_0001001100000111"; -- 0.07206839484018134
	pesos_i(1216) := b"0000000000000000_0000000000000000_0001110011100111_0101110111001100"; -- 0.1129053710758022
	pesos_i(1217) := b"0000000000000000_0000000000000000_0000101000111100_0101000000000010"; -- 0.039982796133509996
	pesos_i(1218) := b"0000000000000000_0000000000000000_0010101100101101_1110110000111000"; -- 0.16866947530554297
	pesos_i(1219) := b"1111111111111111_1111111111111111_1110011101110010_0110011001000110"; -- -0.09591065210547678
	pesos_i(1220) := b"1111111111111111_1111111111111111_1101010101001000_0011100101111000"; -- -0.16686669178942692
	pesos_i(1221) := b"1111111111111111_1111111111111111_1111010011000111_1001110010001010"; -- -0.043829170603470906
	pesos_i(1222) := b"1111111111111111_1111111111111111_1101101010111011_0101000011111000"; -- -0.1455792803147857
	pesos_i(1223) := b"0000000000000000_0000000000000000_0000001100011001_1100110010001000"; -- 0.012112410661401462
	pesos_i(1224) := b"1111111111111111_1111111111111111_1110000111110111_0111111011001001"; -- -0.11731727200113405
	pesos_i(1225) := b"1111111111111111_1111111111111111_1101111100011111_0101101101011010"; -- -0.12842778262564103
	pesos_i(1226) := b"1111111111111111_1111111111111111_1110111010110011_0100110011000111"; -- -0.06757660038356617
	pesos_i(1227) := b"1111111111111111_1111111111111111_1111101100001010_0110110110100101"; -- -0.01937212674771055
	pesos_i(1228) := b"0000000000000000_0000000000000000_0010001110011010_1001010001100100"; -- 0.13907744830884744
	pesos_i(1229) := b"1111111111111111_1111111111111111_1101101001101101_0001010010100100"; -- -0.14677306163830914
	pesos_i(1230) := b"1111111111111111_1111111111111111_1110010101101001_1011101110100101"; -- -0.1038553927394253
	pesos_i(1231) := b"1111111111111111_1111111111111111_1101110000000100_1100001000000001"; -- -0.14055240141461833
	pesos_i(1232) := b"0000000000000000_0000000000000000_0000001110001000_0111111100010110"; -- 0.013801520233640174
	pesos_i(1233) := b"0000000000000000_0000000000000000_0000001010001001_1000101010000001"; -- 0.00991120956303264
	pesos_i(1234) := b"1111111111111111_1111111111111111_1101011111010010_1001001100100011"; -- -0.15694313416902128
	pesos_i(1235) := b"0000000000000000_0000000000000000_0000110001010111_0010011000011000"; -- 0.04820478525520279
	pesos_i(1236) := b"1111111111111111_1111111111111111_1111101101111000_1001101001010001"; -- -0.01769099728216546
	pesos_i(1237) := b"1111111111111111_1111111111111111_1111010111100001_0111100101111010"; -- -0.03952828187345579
	pesos_i(1238) := b"0000000000000000_0000000000000000_0001011110110000_1001111001010000"; -- 0.09253873309221182
	pesos_i(1239) := b"0000000000000000_0000000000000000_0001110100110000_1111011110010110"; -- 0.11402842905516264
	pesos_i(1240) := b"0000000000000000_0000000000000000_0001010111100110_0011011000100001"; -- 0.08554399770934355
	pesos_i(1241) := b"1111111111111111_1111111111111111_1101011101000100_0110011110110100"; -- -0.15911247104702023
	pesos_i(1242) := b"1111111111111111_1111111111111111_1110011001011110_1111100001111000"; -- -0.10011336397023364
	pesos_i(1243) := b"0000000000000000_0000000000000000_0001001100110011_0110111011001110"; -- 0.07500355282870753
	pesos_i(1244) := b"1111111111111111_1111111111111111_1101111011100110_0000100111010110"; -- -0.1293023921584605
	pesos_i(1245) := b"0000000000000000_0000000000000000_0001011010110010_1110011101101001"; -- 0.0886673576561329
	pesos_i(1246) := b"0000000000000000_0000000000000000_0000001000100001_0111101010010111"; -- 0.00832334702405672
	pesos_i(1247) := b"0000000000000000_0000000000000000_0010001011100001_1110011101100110"; -- 0.13625951987445298
	pesos_i(1248) := b"0000000000000000_0000000000000000_0000011111110000_0011100010110000"; -- 0.031009238195292776
	pesos_i(1249) := b"0000000000000000_0000000000000000_0000000001101011_0101000110100101"; -- 0.0016375569131573042
	pesos_i(1250) := b"0000000000000000_0000000000000000_0010001010000110_1000000000101110"; -- 0.13486481785730384
	pesos_i(1251) := b"1111111111111111_1111111111111111_1110011101010100_1101011001101101"; -- -0.09636173103048243
	pesos_i(1252) := b"1111111111111111_1111111111111111_1111110000101111_0000111000101100"; -- -0.014906992240111314
	pesos_i(1253) := b"1111111111111111_1111111111111111_1101010010011100_1101110010001001"; -- -0.16948148387748024
	pesos_i(1254) := b"1111111111111111_1111111111111111_1110011100000111_0010111110010101"; -- -0.09754660227422497
	pesos_i(1255) := b"0000000000000000_0000000000000000_0001010110011101_0011111011111101"; -- 0.08443063422026778
	pesos_i(1256) := b"0000000000000000_0000000000000000_0010000010101010_1000110000000001"; -- 0.12760233894918985
	pesos_i(1257) := b"0000000000000000_0000000000000000_0001011100001011_1010010011010001"; -- 0.09002142043660265
	pesos_i(1258) := b"1111111111111111_1111111111111111_1110001010001100_1110011011101100"; -- -0.1150375054544097
	pesos_i(1259) := b"1111111111111111_1111111111111111_1110111000000101_1011111101000100"; -- -0.07022480573127574
	pesos_i(1260) := b"1111111111111111_1111111111111111_1111010111011001_0101011000001011"; -- -0.03965246431951158
	pesos_i(1261) := b"1111111111111111_1111111111111111_1101100101101110_0011100000101000"; -- -0.15066193613457385
	pesos_i(1262) := b"0000000000000000_0000000000000000_0001111101010001_0001000100110110"; -- 0.12233073783660817
	pesos_i(1263) := b"1111111111111111_1111111111111111_1110011000100011_1111010010111011"; -- -0.10101385522737687
	pesos_i(1264) := b"1111111111111111_1111111111111111_1110000111110010_1110100111000001"; -- -0.11738719030565287
	pesos_i(1265) := b"0000000000000000_0000000000000000_0000011101010011_1101011110001101"; -- 0.02862307735566378
	pesos_i(1266) := b"1111111111111111_1111111111111111_1101101111100110_0000001111101101"; -- -0.14102149459302413
	pesos_i(1267) := b"0000000000000000_0000000000000000_0000000100101010_1111000000110000"; -- 0.004561435468633754
	pesos_i(1268) := b"1111111111111111_1111111111111111_1110110000010110_0110011101100111"; -- -0.07778314332064559
	pesos_i(1269) := b"0000000000000000_0000000000000000_0010110011000111_1001011001010101"; -- 0.17492045952412777
	pesos_i(1270) := b"0000000000000000_0000000000000000_0010100001110011_1101101110111101"; -- 0.1580178581485789
	pesos_i(1271) := b"1111111111111111_1111111111111111_1101111101100110_1000111010101100"; -- -0.12734134970858493
	pesos_i(1272) := b"0000000000000000_0000000000000000_0010110001010011_0011010011000000"; -- 0.1731446236556615
	pesos_i(1273) := b"0000000000000000_0000000000000000_0001011011000101_0110101101011001"; -- 0.08894987992287491
	pesos_i(1274) := b"0000000000000000_0000000000000000_0000101000011000_1000110000001000"; -- 0.039437057458793945
	pesos_i(1275) := b"1111111111111111_1111111111111111_1110010110100010_0111100110010110"; -- -0.10298957908630646
	pesos_i(1276) := b"1111111111111111_1111111111111111_1101011000101101_0010011000011101"; -- -0.16337358282572909
	pesos_i(1277) := b"1111111111111111_1111111111111111_1111001000011110_1001000000100110"; -- -0.05422114436287571
	pesos_i(1278) := b"0000000000000000_0000000000000000_0001101000011101_0101111110111110"; -- 0.10201071152830316
	pesos_i(1279) := b"0000000000000000_0000000000000000_0010101111000011_1000000101000110"; -- 0.1709519191517062
	pesos_i(1280) := b"0000000000000000_0000000000000000_0000100100110110_1010011101010110"; -- 0.03599019869803635
	pesos_i(1281) := b"1111111111111111_1111111111111111_1101111011000111_1110001111000101"; -- -0.12976242491850584
	pesos_i(1282) := b"0000000000000000_0000000000000000_0010011101110111_1101110000110011"; -- 0.1541726708518937
	pesos_i(1283) := b"1111111111111111_1111111111111111_1111100001000111_1000111001110111"; -- -0.030158134511613123
	pesos_i(1284) := b"0000000000000000_0000000000000000_0000010100001110_1001001010100110"; -- 0.019753613872627845
	pesos_i(1285) := b"1111111111111111_1111111111111111_1101011010111110_1000000011010011"; -- -0.16115565155264625
	pesos_i(1286) := b"1111111111111111_1111111111111111_1111101100000011_1100011101101000"; -- -0.01947358803701382
	pesos_i(1287) := b"1111111111111111_1111111111111111_1101110010100111_0100000100100000"; -- -0.13807290055687013
	pesos_i(1288) := b"0000000000000000_0000000000000000_0010100100001010_0110010011100000"; -- 0.16031485051536262
	pesos_i(1289) := b"1111111111111111_1111111111111111_1111001001100110_1001001101110011"; -- -0.05312231490125276
	pesos_i(1290) := b"0000000000000000_0000000000000000_0001000111111011_1111001111001010"; -- 0.07025073712012767
	pesos_i(1291) := b"0000000000000000_0000000000000000_0000000111001101_0010000001111111"; -- 0.007036238773467475
	pesos_i(1292) := b"1111111111111111_1111111111111111_1111101010101011_1001000100101000"; -- -0.020819594978071992
	pesos_i(1293) := b"1111111111111111_1111111111111111_1111101010001010_1101111111001000"; -- -0.02131844864783698
	pesos_i(1294) := b"1111111111111111_1111111111111111_1111101101111001_0000011101110100"; -- -0.017684492274516787
	pesos_i(1295) := b"1111111111111111_1111111111111111_1111100111101011_1011001101111011"; -- -0.023747236737874374
	pesos_i(1296) := b"1111111111111111_1111111111111111_1101010000000101_0111101110110110"; -- -0.17179133228249288
	pesos_i(1297) := b"0000000000000000_0000000000000000_0010011000110100_1000000100101110"; -- 0.14923865669395628
	pesos_i(1298) := b"1111111111111111_1111111111111111_1101111110110110_0001101101111101"; -- -0.12612751185959167
	pesos_i(1299) := b"1111111111111111_1111111111111111_1111000011000010_0011100100100100"; -- -0.05953638916500203
	pesos_i(1300) := b"1111111111111111_1111111111111111_1111110010001010_1100100010001101"; -- -0.013507333241960986
	pesos_i(1301) := b"0000000000000000_0000000000000000_0010000100000100_1111000011101110"; -- 0.12898164560927908
	pesos_i(1302) := b"0000000000000000_0000000000000000_0001010010011000_0010000011010000"; -- 0.08044629167274137
	pesos_i(1303) := b"0000000000000000_0000000000000000_0001010111001100_0010101111100111"; -- 0.0851466598020833
	pesos_i(1304) := b"0000000000000000_0000000000000000_0001110101011110_0001111001011011"; -- 0.11471738554538974
	pesos_i(1305) := b"0000000000000000_0000000000000000_0001001111110011_1011010111110111"; -- 0.07793748165390219
	pesos_i(1306) := b"0000000000000000_0000000000000000_0010000110000101_0010000010110000"; -- 0.13093761725953906
	pesos_i(1307) := b"0000000000000000_0000000000000000_0001100000011111_0001111001011001"; -- 0.09422483139570892
	pesos_i(1308) := b"1111111111111111_1111111111111111_1101010010111101_0101101110011100"; -- -0.16898562846755794
	pesos_i(1309) := b"0000000000000000_0000000000000000_0000111011110101_1010101000011010"; -- 0.05843604222895698
	pesos_i(1310) := b"0000000000000000_0000000000000000_0000110000000011_1110111010111110"; -- 0.04693500640665751
	pesos_i(1311) := b"1111111111111111_1111111111111111_1101010110100111_0011101110100000"; -- -0.16541697833524785
	pesos_i(1312) := b"1111111111111111_1111111111111111_1110101001001000_1101001111000000"; -- -0.08482624591947902
	pesos_i(1313) := b"0000000000000000_0000000000000000_0000011100010101_0101110000100011"; -- 0.027669676456799516
	pesos_i(1314) := b"1111111111111111_1111111111111111_1101100111101100_1010110111010100"; -- -0.14873231492026684
	pesos_i(1315) := b"1111111111111111_1111111111111111_1110011110110011_1100111111001000"; -- -0.09491254202256028
	pesos_i(1316) := b"0000000000000000_0000000000000000_0001010110011001_1111101110110100"; -- 0.08438084747502486
	pesos_i(1317) := b"1111111111111111_1111111111111111_1101010010001001_1110010011011001"; -- -0.16977090560556607
	pesos_i(1318) := b"1111111111111111_1111111111111111_1111001000100011_1111101010100000"; -- -0.054138504064155546
	pesos_i(1319) := b"1111111111111111_1111111111111111_1101111100011001_0111101111011000"; -- -0.12851739860897377
	pesos_i(1320) := b"1111111111111111_1111111111111111_1110011001101110_1101111011110111"; -- -0.09987074340475931
	pesos_i(1321) := b"1111111111111111_1111111111111111_1111101111100101_0010100011111010"; -- -0.016034544843744485
	pesos_i(1322) := b"1111111111111111_1111111111111111_1110100110100011_0110101000111100"; -- -0.08735023531000466
	pesos_i(1323) := b"1111111111111111_1111111111111111_1101100000110011_0100000010100011"; -- -0.15546794921457296
	pesos_i(1324) := b"0000000000000000_0000000000000000_0010001111110000_1010110110000001"; -- 0.14039120094150453
	pesos_i(1325) := b"0000000000000000_0000000000000000_0000100001111011_1110001001101111"; -- 0.03314032757727479
	pesos_i(1326) := b"0000000000000000_0000000000000000_0001100101010010_0110101000111010"; -- 0.09891380221045941
	pesos_i(1327) := b"1111111111111111_1111111111111111_1111111101001101_1100011011000011"; -- -0.00271947606250983
	pesos_i(1328) := b"1111111111111111_1111111111111111_1110100010111101_0101000101111111"; -- -0.09086123124839478
	pesos_i(1329) := b"0000000000000000_0000000000000000_0010001001010001_0011110100110110"; -- 0.13405211033115674
	pesos_i(1330) := b"1111111111111111_1111111111111111_1110011101000100_1001110101000110"; -- -0.0966092781282703
	pesos_i(1331) := b"0000000000000000_0000000000000000_0010001010100101_0111010111110001"; -- 0.13533723013527496
	pesos_i(1332) := b"1111111111111111_1111111111111111_1101100101001011_0100110001100000"; -- -0.15119478847504889
	pesos_i(1333) := b"0000000000000000_0000000000000000_0001010011010100_0010111010011010"; -- 0.0813626409853532
	pesos_i(1334) := b"0000000000000000_0000000000000000_0001111101111000_1110001001101011"; -- 0.12293830035443416
	pesos_i(1335) := b"1111111111111111_1111111111111111_1111011000101101_0100001101011010"; -- -0.03837183998093153
	pesos_i(1336) := b"1111111111111111_1111111111111111_1110010000011100_1101001101001011"; -- -0.10893515979524199
	pesos_i(1337) := b"0000000000000000_0000000000000000_0000001000010011_0111010110110011"; -- 0.008109432420244235
	pesos_i(1338) := b"0000000000000000_0000000000000000_0001100011101000_1010101100101101"; -- 0.09730024183275163
	pesos_i(1339) := b"1111111111111111_1111111111111111_1111000100010000_1010110000011010"; -- -0.05833935136545004
	pesos_i(1340) := b"1111111111111111_1111111111111111_1111000001000110_1000100001100101"; -- -0.06142375501957999
	pesos_i(1341) := b"1111111111111111_1111111111111111_1110011010001001_0000110111111111"; -- -0.09947121168333815
	pesos_i(1342) := b"1111111111111111_1111111111111111_1111100011101011_1111101100000000"; -- -0.027649223872235975
	pesos_i(1343) := b"1111111111111111_1111111111111111_1110111101101010_1000110110000110"; -- -0.0647803829591472
	pesos_i(1344) := b"1111111111111111_1111111111111111_1111001010111010_0010100110010101"; -- -0.05184688685105891
	pesos_i(1345) := b"1111111111111111_1111111111111111_1110001011011000_0010010100001111"; -- -0.1138893927465605
	pesos_i(1346) := b"0000000000000000_0000000000000000_0001011101010000_1100000010011111"; -- 0.09107593424072385
	pesos_i(1347) := b"1111111111111111_1111111111111111_1110000010100111_0100101100010000"; -- -0.12244730822942688
	pesos_i(1348) := b"0000000000000000_0000000000000000_0001010011101000_0101100010010010"; -- 0.08167031821231484
	pesos_i(1349) := b"1111111111111111_1111111111111111_1110100000000110_1011101010111111"; -- -0.0936473163779239
	pesos_i(1350) := b"0000000000000000_0000000000000000_0001011110001001_1111110011010101"; -- 0.0919492739635515
	pesos_i(1351) := b"1111111111111111_1111111111111111_1111011011101110_1001011011111101"; -- -0.035421908513081295
	pesos_i(1352) := b"0000000000000000_0000000000000000_0000001000100111_1000010101110100"; -- 0.00841554731027673
	pesos_i(1353) := b"1111111111111111_1111111111111111_1110111010101111_1100101010000010"; -- -0.06763014157477427
	pesos_i(1354) := b"0000000000000000_0000000000000000_0000110010101111_1000000011001000"; -- 0.04955296406422515
	pesos_i(1355) := b"0000000000000000_0000000000000000_0010001111111110_0111110001111100"; -- 0.1406019023241885
	pesos_i(1356) := b"0000000000000000_0000000000000000_0010101000011101_0101111001110000"; -- 0.1645106337469802
	pesos_i(1357) := b"1111111111111111_1111111111111111_1111100101111010_0101111000001111"; -- -0.025476571409065285
	pesos_i(1358) := b"1111111111111111_1111111111111111_1110100111000000_1011000010111110"; -- -0.08690352783676566
	pesos_i(1359) := b"0000000000000000_0000000000000000_0010001110000000_1110010001000100"; -- 0.13868548075262732
	pesos_i(1360) := b"0000000000000000_0000000000000000_0010101100001101_0000011001010111"; -- 0.16816749213378943
	pesos_i(1361) := b"0000000000000000_0000000000000000_0001011100101011_0001111000010011"; -- 0.09050167050210965
	pesos_i(1362) := b"0000000000000000_0000000000000000_0000110100001110_1001001111110011"; -- 0.05100369141179089
	pesos_i(1363) := b"0000000000000000_0000000000000000_0010101101010000_0001001110100111"; -- 0.16919062440263544
	pesos_i(1364) := b"0000000000000000_0000000000000000_0000111010001010_1100000011001111"; -- 0.056804705154028086
	pesos_i(1365) := b"0000000000000000_0000000000000000_0001010101000101_1000111100010011"; -- 0.08309263427288477
	pesos_i(1366) := b"0000000000000000_0000000000000000_0010000000111011_1000011110000011"; -- 0.1259083455820374
	pesos_i(1367) := b"0000000000000000_0000000000000000_0001001000100010_0111001101111011"; -- 0.07083818190593165
	pesos_i(1368) := b"1111111111111111_1111111111111111_1111001011101010_0000000000011101"; -- -0.0511169366906058
	pesos_i(1369) := b"1111111111111111_1111111111111111_1110010011000111_0010000011111101"; -- -0.10633653479378087
	pesos_i(1370) := b"1111111111111111_1111111111111111_1110001000110011_0111110111110010"; -- -0.11640179491254393
	pesos_i(1371) := b"1111111111111111_1111111111111111_1110000010100001_0001101011100110"; -- -0.12254173157783219
	pesos_i(1372) := b"0000000000000000_0000000000000000_0010100010101010_0111111111000011"; -- 0.15885160942439078
	pesos_i(1373) := b"1111111111111111_1111111111111111_1111001000010111_1101110101101001"; -- -0.05432335081521976
	pesos_i(1374) := b"0000000000000000_0000000000000000_0000010101110001_0101110100111001"; -- 0.02126104977307298
	pesos_i(1375) := b"1111111111111111_1111111111111111_1110010000111100_1110100111111000"; -- -0.10844552699112375
	pesos_i(1376) := b"1111111111111111_1111111111111111_1101111100100011_1110000001010000"; -- -0.1283588223083884
	pesos_i(1377) := b"1111111111111111_1111111111111111_1111010111010100_1101110011111011"; -- -0.0397207151844078
	pesos_i(1378) := b"1111111111111111_1111111111111111_1111001011100001_0101000110011001"; -- -0.05124940893715792
	pesos_i(1379) := b"1111111111111111_1111111111111111_1110101101101111_0111100001100110"; -- -0.08033034820102732
	pesos_i(1380) := b"0000000000000000_0000000000000000_0010000100000001_0101110101111011"; -- 0.12892708067439002
	pesos_i(1381) := b"1111111111111111_1111111111111111_1101111000110010_1111011000000100"; -- -0.13203489691869494
	pesos_i(1382) := b"1111111111111111_1111111111111111_1110101011010010_0101011001011011"; -- -0.08272800717188243
	pesos_i(1383) := b"1111111111111111_1111111111111111_1110001001001101_0111101101110000"; -- -0.11600521577068018
	pesos_i(1384) := b"1111111111111111_1111111111111111_1101001111110011_1100001010001100"; -- -0.17206176825377384
	pesos_i(1385) := b"1111111111111111_1111111111111111_1111100101001001_1001111111101101"; -- -0.026220326086445072
	pesos_i(1386) := b"0000000000000000_0000000000000000_0010010101011101_1111000011110111"; -- 0.14596468010877128
	pesos_i(1387) := b"0000000000000000_0000000000000000_0000010001100100_0011110110001111"; -- 0.017154548069065707
	pesos_i(1388) := b"1111111111111111_1111111111111111_1101100100010111_0011100001010001"; -- -0.15198944118394211
	pesos_i(1389) := b"1111111111111111_1111111111111111_1110011001001000_0010010110101110"; -- -0.10046162141690132
	pesos_i(1390) := b"0000000000000000_0000000000000000_0000010010001011_1010110000001110"; -- 0.01775622705454051
	pesos_i(1391) := b"1111111111111111_1111111111111111_1110010101110111_0001011110101110"; -- -0.10365154260075143
	pesos_i(1392) := b"0000000000000000_0000000000000000_0001000111001101_0010110101000010"; -- 0.0695369992876455
	pesos_i(1393) := b"0000000000000000_0000000000000000_0000110000111010_0101100100011000"; -- 0.04776532014533355
	pesos_i(1394) := b"1111111111111111_1111111111111111_1111010010010000_1011011100101010"; -- -0.04466681686215042
	pesos_i(1395) := b"1111111111111111_1111111111111111_1110000011010101_0000001011110110"; -- -0.12174970136502924
	pesos_i(1396) := b"0000000000000000_0000000000000000_0001011110010001_0110011000000110"; -- 0.0920623554959106
	pesos_i(1397) := b"1111111111111111_1111111111111111_1111000010101110_0100000100011000"; -- -0.059841090726647
	pesos_i(1398) := b"1111111111111111_1111111111111111_1111110110011101_1001010101101010"; -- -0.009314214438436134
	pesos_i(1399) := b"0000000000000000_0000000000000000_0001100110011001_1111111001001110"; -- 0.10000600243263945
	pesos_i(1400) := b"0000000000000000_0000000000000000_0000011010110011_1101001110010001"; -- 0.026181433593127912
	pesos_i(1401) := b"1111111111111111_1111111111111111_1111100101110010_1010001100001000"; -- -0.02559453060484616
	pesos_i(1402) := b"0000000000000000_0000000000000000_0000110011101100_0111100001000100"; -- 0.050483242538528504
	pesos_i(1403) := b"1111111111111111_1111111111111111_1110111001100110_1011101111101110"; -- -0.06874490211831022
	pesos_i(1404) := b"0000000000000000_0000000000000000_0001011011000101_0011010111100111"; -- 0.08894669419560605
	pesos_i(1405) := b"1111111111111111_1111111111111111_1111001001010110_0001110111111000"; -- -0.05337345786692766
	pesos_i(1406) := b"1111111111111111_1111111111111111_1111101101000000_0001101100000111"; -- -0.018553076563938026
	pesos_i(1407) := b"0000000000000000_0000000000000000_0001000010100001_0110100001101110"; -- 0.06496288942275665
	pesos_i(1408) := b"0000000000000000_0000000000000000_0001010011011111_1001010011011000"; -- 0.08153658175707143
	pesos_i(1409) := b"0000000000000000_0000000000000000_0000111101000010_0100001100100100"; -- 0.059604832031064876
	pesos_i(1410) := b"0000000000000000_0000000000000000_0001001010101011_0001110010010111"; -- 0.07292345708337289
	pesos_i(1411) := b"1111111111111111_1111111111111111_1111000111111100_0100001011100101"; -- -0.05474454785054922
	pesos_i(1412) := b"1111111111111111_1111111111111111_1111010010001000_0100100010110100"; -- -0.044795471295766484
	pesos_i(1413) := b"1111111111111111_1111111111111111_1110001110000101_1000100011000111"; -- -0.1112436784679165
	pesos_i(1414) := b"1111111111111111_1111111111111111_1110111100110111_1100001010110110"; -- -0.06555541081978272
	pesos_i(1415) := b"0000000000000000_0000000000000000_0010010111101010_1011111101001001"; -- 0.14811320822486268
	pesos_i(1416) := b"0000000000000000_0000000000000000_0001011010001011_0110000110000110"; -- 0.08806428456552434
	pesos_i(1417) := b"1111111111111111_1111111111111111_1101011000101110_0000101011010101"; -- -0.16335995001653666
	pesos_i(1418) := b"1111111111111111_1111111111111111_1110001101000010_1000001110100111"; -- -0.11226632287252135
	pesos_i(1419) := b"1111111111111111_1111111111111111_1101101001001111_0011010000001111"; -- -0.14722895282220247
	pesos_i(1420) := b"0000000000000000_0000000000000000_0001101011001001_1110000010011111"; -- 0.10464290498156445
	pesos_i(1421) := b"0000000000000000_0000000000000000_0010110011011011_1101101001010000"; -- 0.17522968734955488
	pesos_i(1422) := b"0000000000000000_0000000000000000_0000101100001000_1000101101011101"; -- 0.043099126897747496
	pesos_i(1423) := b"0000000000000000_0000000000000000_0000010010000100_1011110101111010"; -- 0.017650453836960123
	pesos_i(1424) := b"1111111111111111_1111111111111111_1110000001001100_1110001000111100"; -- -0.1238268474130263
	pesos_i(1425) := b"1111111111111111_1111111111111111_1110010111110011_0000011011010001"; -- -0.10176045800713616
	pesos_i(1426) := b"0000000000000000_0000000000000000_0001100100011010_1101001111000001"; -- 0.09806560000292194
	pesos_i(1427) := b"0000000000000000_0000000000000000_0010001001111100_0101000001001110"; -- 0.1347093764660063
	pesos_i(1428) := b"0000000000000000_0000000000000000_0001100000101010_1111101110011110"; -- 0.09440586661675926
	pesos_i(1429) := b"1111111111111111_1111111111111111_1101101100010010_0111100011101101"; -- -0.14424938412224642
	pesos_i(1430) := b"1111111111111111_1111111111111111_1111101111100111_1000110110001111"; -- -0.01599803212135101
	pesos_i(1431) := b"0000000000000000_0000000000000000_0010100101101001_1101110010010111"; -- 0.16177157108716558
	pesos_i(1432) := b"0000000000000000_0000000000000000_0001010110100011_1111111001011000"; -- 0.08453359274826072
	pesos_i(1433) := b"0000000000000000_0000000000000000_0010001000010110_0111100110111111"; -- 0.13315545000529871
	pesos_i(1434) := b"1111111111111111_1111111111111111_1110000001000011_1010011111100001"; -- -0.12396765467233523
	pesos_i(1435) := b"1111111111111111_1111111111111111_1101011101000011_0010000100101111"; -- -0.1591319332182632
	pesos_i(1436) := b"1111111111111111_1111111111111111_1110100011110001_1001110101000011"; -- -0.09006325839440552
	pesos_i(1437) := b"0000000000000000_0000000000000000_0001010011010001_1100011110000000"; -- 0.08132597811971187
	pesos_i(1438) := b"1111111111111111_1111111111111111_1111000001100011_1011010100010000"; -- -0.060978587609581685
	pesos_i(1439) := b"0000000000000000_0000000000000000_0000011101101101_0001000101100010"; -- 0.0290079940269157
	pesos_i(1440) := b"0000000000000000_0000000000000000_0001111011011101_0001100110111010"; -- 0.12056122576405184
	pesos_i(1441) := b"0000000000000000_0000000000000000_0000011000010101_0001111001100110"; -- 0.023759746564010868
	pesos_i(1442) := b"1111111111111111_1111111111111111_1110001000110001_0000110000111101"; -- -0.1164390899285697
	pesos_i(1443) := b"1111111111111111_1111111111111111_1110111101100000_1000110011011001"; -- -0.06493301112016303
	pesos_i(1444) := b"0000000000000000_0000000000000000_0010111010010110_0001011000100100"; -- 0.18197763800685612
	pesos_i(1445) := b"0000000000000000_0000000000000000_0010101010101011_1101101101000000"; -- 0.16668482134766818
	pesos_i(1446) := b"0000000000000000_0000000000000000_0001000000010100_0111001111001101"; -- 0.06281207798019033
	pesos_i(1447) := b"0000000000000000_0000000000000000_0001011100111010_1111101011000100"; -- 0.09074370661837469
	pesos_i(1448) := b"1111111111111111_1111111111111111_1111010001010100_1000011000111001"; -- -0.04558526151057851
	pesos_i(1449) := b"0000000000000000_0000000000000000_0000110010011100_1010000111101111"; -- 0.049265023188817605
	pesos_i(1450) := b"1111111111111111_1111111111111111_1111101100100011_0101011110000010"; -- -0.018991976567794368
	pesos_i(1451) := b"1111111111111111_1111111111111111_1111011100101100_0000100101001101"; -- -0.03448430895743523
	pesos_i(1452) := b"0000000000000000_0000000000000000_0001001101010000_0100100110101000"; -- 0.07544384331688771
	pesos_i(1453) := b"0000000000000000_0000000000000000_0000010100110111_1001000110111111"; -- 0.02037917047373899
	pesos_i(1454) := b"1111111111111111_1111111111111111_1111011110000010_1111100011011100"; -- -0.0331577741559749
	pesos_i(1455) := b"0000000000000000_0000000000000000_0001101111011001_1100000111110110"; -- 0.10879146819764203
	pesos_i(1456) := b"0000000000000000_0000000000000000_0010010000100011_1111011100010001"; -- 0.14117378390263383
	pesos_i(1457) := b"0000000000000000_0000000000000000_0010001111010000_0110001010100001"; -- 0.13989845680989774
	pesos_i(1458) := b"1111111111111111_1111111111111111_1111110011001010_1100110100010010"; -- -0.012530501580487453
	pesos_i(1459) := b"0000000000000000_0000000000000000_0001100111101111_0001111001100010"; -- 0.10130491157150442
	pesos_i(1460) := b"1111111111111111_1111111111111111_1110000000001010_0110110101101101"; -- -0.12484088970819869
	pesos_i(1461) := b"1111111111111111_1111111111111111_1111100101100111_0100111011101001"; -- -0.025767391430557174
	pesos_i(1462) := b"0000000000000000_0000000000000000_0001110110010111_0010111010110001"; -- 0.11558811017437966
	pesos_i(1463) := b"0000000000000000_0000000000000000_0000010101001110_0101010011100110"; -- 0.02072649590514797
	pesos_i(1464) := b"1111111111111111_1111111111111111_1111010110011001_0101110111010001"; -- -0.04062856340478013
	pesos_i(1465) := b"1111111111111111_1111111111111111_1101110010111000_1011100101011011"; -- -0.13780633470612352
	pesos_i(1466) := b"1111111111111111_1111111111111111_1110010011101000_1110011010011011"; -- -0.10582121569901462
	pesos_i(1467) := b"1111111111111111_1111111111111111_1111111111111001_0111111101010100"; -- -9.922209268195539e-05
	pesos_i(1468) := b"1111111111111111_1111111111111111_1101110101001111_1011001010100010"; -- -0.1355026583212973
	pesos_i(1469) := b"0000000000000000_0000000000000000_0001000001100111_1111100101000010"; -- 0.06408651220991064
	pesos_i(1470) := b"0000000000000000_0000000000000000_0000001010001001_0010100101110010"; -- 0.009905424347016446
	pesos_i(1471) := b"1111111111111111_1111111111111111_1110001100111101_1000010000001110"; -- -0.11234259268795888
	pesos_i(1472) := b"0000000000000000_0000000000000000_0000110101010110_0110101010010101"; -- 0.05209985867652775
	pesos_i(1473) := b"1111111111111111_1111111111111111_1110010011001110_0101001000010010"; -- -0.10622679763056123
	pesos_i(1474) := b"0000000000000000_0000000000000000_0010011111000000_0100010011000011"; -- 0.15527753590202223
	pesos_i(1475) := b"0000000000000000_0000000000000000_0010100011011101_1111011001000010"; -- 0.15963687044980188
	pesos_i(1476) := b"0000000000000000_0000000000000000_0000100001110110_1110110010000111"; -- 0.03306463526976255
	pesos_i(1477) := b"0000000000000000_0000000000000000_0000001000010100_1001101010111011"; -- 0.008126898510377036
	pesos_i(1478) := b"0000000000000000_0000000000000000_0010000110000101_1001010101001101"; -- 0.13094456789903863
	pesos_i(1479) := b"1111111111111111_1111111111111111_1101110011100010_0000100011001010"; -- -0.13717598976060205
	pesos_i(1480) := b"0000000000000000_0000000000000000_0001001101100110_0110100001101101"; -- 0.07578137067433857
	pesos_i(1481) := b"0000000000000000_0000000000000000_0000110010111010_1110110000100010"; -- 0.049727209418769326
	pesos_i(1482) := b"0000000000000000_0000000000000000_0001100010110001_0001001111010110"; -- 0.09645198797489205
	pesos_i(1483) := b"1111111111111111_1111111111111111_1111100100100101_1110111011110000"; -- -0.026764933126669516
	pesos_i(1484) := b"1111111111111111_1111111111111111_1110001110101111_0100000111001011"; -- -0.11060704041175795
	pesos_i(1485) := b"0000000000000000_0000000000000000_0001010010011000_1001010011100101"; -- 0.0804532107713789
	pesos_i(1486) := b"1111111111111111_1111111111111111_1111010000110101_1111101011111110"; -- -0.046051323906760394
	pesos_i(1487) := b"1111111111111111_1111111111111111_1110010000001110_1011110101011110"; -- -0.1091500898159115
	pesos_i(1488) := b"1111111111111111_1111111111111111_1111000101100101_1001011100100011"; -- -0.05704360394666763
	pesos_i(1489) := b"0000000000000000_0000000000000000_0010000001001000_0010011010010110"; -- 0.12610093267277353
	pesos_i(1490) := b"0000000000000000_0000000000000000_0001010100111001_1101010010001011"; -- 0.08291366944513515
	pesos_i(1491) := b"1111111111111111_1111111111111111_1101001001010000_0111000111010111"; -- -0.1784600114908428
	pesos_i(1492) := b"1111111111111111_1111111111111111_1110100011001101_0101100111010011"; -- -0.09061659421926148
	pesos_i(1493) := b"1111111111111111_1111111111111111_1110011001010111_1100001000000011"; -- -0.10022342143504373
	pesos_i(1494) := b"0000000000000000_0000000000000000_0000101001100111_0010001011011000"; -- 0.040636232022014565
	pesos_i(1495) := b"0000000000000000_0000000000000000_0010110111111110_1101000001100001"; -- 0.17966940280608693
	pesos_i(1496) := b"1111111111111111_1111111111111111_1101101111100111_0100010111000011"; -- -0.14100231157193813
	pesos_i(1497) := b"1111111111111111_1111111111111111_1111001110110011_1100111001011000"; -- -0.048037627681543585
	pesos_i(1498) := b"1111111111111111_1111111111111111_1101100011100111_1100111110100111"; -- -0.15271284276883415
	pesos_i(1499) := b"0000000000000000_0000000000000000_0010000010000010_0111100100101101"; -- 0.12699086531213516
	pesos_i(1500) := b"0000000000000000_0000000000000000_0001100000000001_1000100001110111"; -- 0.09377339263466955
	pesos_i(1501) := b"1111111111111111_1111111111111111_1110101010011000_0100010110010111"; -- -0.08361401617966974
	pesos_i(1502) := b"1111111111111111_1111111111111111_1110101000000001_1001001001100111"; -- -0.08591351498832847
	pesos_i(1503) := b"1111111111111111_1111111111111111_1111001000001001_0101100000010010"; -- -0.05454492160794276
	pesos_i(1504) := b"0000000000000000_0000000000000000_0001110001110010_1010000100111010"; -- 0.1111241118745653
	pesos_i(1505) := b"1111111111111111_1111111111111111_1111011011110110_1001001011111101"; -- -0.03530007679470348
	pesos_i(1506) := b"0000000000000000_0000000000000000_0001001110100000_1111011010010100"; -- 0.07667485334706305
	pesos_i(1507) := b"1111111111111111_1111111111111111_1111111000111100_0010111110100010"; -- -0.006894133542286785
	pesos_i(1508) := b"0000000000000000_0000000000000000_0000011011111010_0100111010000010"; -- 0.02725687660174034
	pesos_i(1509) := b"1111111111111111_1111111111111111_1110011001100111_1110000001101011"; -- -0.09997746831472891
	pesos_i(1510) := b"0000000000000000_0000000000000000_0000101111110001_1001010010100111"; -- 0.04665497845538884
	pesos_i(1511) := b"0000000000000000_0000000000000000_0000111100100100_1011000101100010"; -- 0.059153639282883586
	pesos_i(1512) := b"1111111111111111_1111111111111111_1110010100000100_0101101010000010"; -- -0.1054023201328656
	pesos_i(1513) := b"0000000000000000_0000000000000000_0010100000100110_1100000101001010"; -- 0.1568413548205878
	pesos_i(1514) := b"0000000000000000_0000000000000000_0001001110110011_0000111000110001"; -- 0.07695091907685339
	pesos_i(1515) := b"1111111111111111_1111111111111111_1101111000111101_1010010101100000"; -- -0.13187185684201255
	pesos_i(1516) := b"1111111111111111_1111111111111111_1110001010100111_0011111111101100"; -- -0.11463547221768938
	pesos_i(1517) := b"1111111111111111_1111111111111111_1110100111000101_1101100110100111"; -- -0.08682479557396071
	pesos_i(1518) := b"0000000000000000_0000000000000000_0010001100101001_1011111000100100"; -- 0.1373556935966369
	pesos_i(1519) := b"1111111111111111_1111111111111111_1110001000011100_1100111111011101"; -- -0.1167478642911726
	pesos_i(1520) := b"0000000000000000_0000000000000000_0001011010101101_0111101001111111"; -- 0.08858457188354654
	pesos_i(1521) := b"0000000000000000_0000000000000000_0000011101010110_1101000110101010"; -- 0.028668502906158876
	pesos_i(1522) := b"1111111111111111_1111111111111111_1110001001110010_0010011000000001"; -- -0.11544573278738146
	pesos_i(1523) := b"1111111111111111_1111111111111111_1101001011011010_1101111100000000"; -- -0.1763477921282215
	pesos_i(1524) := b"1111111111111111_1111111111111111_1111100001011011_0101100000110011"; -- -0.02985619303294265
	pesos_i(1525) := b"0000000000000000_0000000000000000_0000110011101111_0101101000010110"; -- 0.05052722017283235
	pesos_i(1526) := b"1111111111111111_1111111111111111_1101111000010010_1001010011000101"; -- -0.13252897454852688
	pesos_i(1527) := b"1111111111111111_1111111111111111_1100101111101011_0001101100100001"; -- -0.20344381754057705
	pesos_i(1528) := b"0000000000000000_0000000000000000_0001100011000101_0100110001111110"; -- 0.09676054075736237
	pesos_i(1529) := b"1111111111111111_1111111111111111_1111100101000101_0101011101011011"; -- -0.02628568667875834
	pesos_i(1530) := b"0000000000000000_0000000000000000_0001011011100111_1110000011110010"; -- 0.08947568801703101
	pesos_i(1531) := b"1111111111111111_1111111111111111_1111100001111110_1110101000100100"; -- -0.02931343676654939
	pesos_i(1532) := b"1111111111111111_1111111111111111_1110101001110011_1001001000111000"; -- -0.08417402403146591
	pesos_i(1533) := b"1111111111111111_1111111111111111_1111010010110110_0000011010000100"; -- -0.04409751195619033
	pesos_i(1534) := b"1111111111111111_1111111111111111_1111000110000101_1000010000010000"; -- -0.05655645941564435
	pesos_i(1535) := b"0000000000000000_0000000000000000_0001011111100000_0100101100100001"; -- 0.09326619676753514
	pesos_i(1536) := b"0000000000000000_0000000000000000_0001010000101001_0010100100001101"; -- 0.07875305716876277
	pesos_i(1537) := b"0000000000000000_0000000000000000_0000111011011001_0111000011000010"; -- 0.0580053782135321
	pesos_i(1538) := b"1111111111111111_1111111111111111_1111011111000010_0010001111001111"; -- -0.032193910537671684
	pesos_i(1539) := b"0000000000000000_0000000000000000_0010000100101111_0011011000110011"; -- 0.1296266435703927
	pesos_i(1540) := b"1111111111111111_1111111111111111_1110110001111000_0111011010101111"; -- -0.07628687127298353
	pesos_i(1541) := b"0000000000000000_0000000000000000_0000111011101111_1001111001110110"; -- 0.05834379551942117
	pesos_i(1542) := b"0000000000000000_0000000000000000_0001101110001001_1111001000101000"; -- 0.107573637780285
	pesos_i(1543) := b"1111111111111111_1111111111111111_1111110101100010_1000001110111100"; -- -0.010215536608337968
	pesos_i(1544) := b"1111111111111111_1111111111111111_1111110010001001_1011111001100110"; -- -0.013523197320801858
	pesos_i(1545) := b"0000000000000000_0000000000000000_0010010000000100_0011011011101101"; -- 0.1406893089838368
	pesos_i(1546) := b"1111111111111111_1111111111111111_1110110001011111_0110111110110101"; -- -0.07666875685055441
	pesos_i(1547) := b"1111111111111111_1111111111111111_1110111011011110_0110111010001011"; -- -0.06691845983876822
	pesos_i(1548) := b"0000000000000000_0000000000000000_0000111000001010_1110101011000011"; -- 0.054854080709576196
	pesos_i(1549) := b"0000000000000000_0000000000000000_0001101110100101_1100000010101001"; -- 0.10799793367726865
	pesos_i(1550) := b"1111111111111111_1111111111111111_1101101011100011_1010111111010101"; -- -0.1449632745624653
	pesos_i(1551) := b"1111111111111111_1111111111111111_1111001010001111_1100111100111111"; -- -0.05249314041483817
	pesos_i(1552) := b"1111111111111111_1111111111111111_1111000100111110_0011001001000011"; -- -0.057644709283098824
	pesos_i(1553) := b"0000000000000000_0000000000000000_0010100001100101_0000011100100001"; -- 0.15779156259413496
	pesos_i(1554) := b"1111111111111111_1111111111111111_1110101001011011_1100100000111001"; -- -0.08453701607001639
	pesos_i(1555) := b"1111111111111111_1111111111111111_1101100010111011_1010101011010000"; -- -0.15338642519533466
	pesos_i(1556) := b"1111111111111111_1111111111111111_1101010110101110_1111011001010101"; -- -0.16529903814513808
	pesos_i(1557) := b"1111111111111111_1111111111111111_1111111010111100_1010011010001010"; -- -0.0049339210912089405
	pesos_i(1558) := b"0000000000000000_0000000000000000_0000101010011111_1110111111000101"; -- 0.04150293880810471
	pesos_i(1559) := b"1111111111111111_1111111111111111_1100100111101111_1111000110101010"; -- -0.2111824950927349
	pesos_i(1560) := b"0000000000000000_0000000000000000_0001111110100110_0010111011110100"; -- 0.1236295076098436
	pesos_i(1561) := b"0000000000000000_0000000000000000_0001000000110101_1110100001111011"; -- 0.06332257263949494
	pesos_i(1562) := b"1111111111111111_1111111111111111_1110001010111001_0111011010100011"; -- -0.11435755268575681
	pesos_i(1563) := b"0000000000000000_0000000000000000_0000100010111010_0011101010000110"; -- 0.03409162313669589
	pesos_i(1564) := b"1111111111111111_1111111111111111_1111010101101111_1001111101111110"; -- -0.04126551786183622
	pesos_i(1565) := b"1111111111111111_1111111111111111_1101010011000010_1010110101111011"; -- -0.168904454731855
	pesos_i(1566) := b"1111111111111111_1111111111111111_1110001111001010_0110111111001000"; -- -0.11019231198140333
	pesos_i(1567) := b"0000000000000000_0000000000000000_0001100011100010_0111010011111000"; -- 0.09720545819269868
	pesos_i(1568) := b"1111111111111111_1111111111111111_1111010011000010_1110001010000100"; -- -0.043901293652104434
	pesos_i(1569) := b"0000000000000000_0000000000000000_0010010010001101_1110010110011100"; -- 0.14279017495952698
	pesos_i(1570) := b"0000000000000000_0000000000000000_0010100011111000_0110000011001001"; -- 0.16003994860786414
	pesos_i(1571) := b"0000000000000000_0000000000000000_0001110110011010_0100111001001001"; -- 0.11563576956067494
	pesos_i(1572) := b"0000000000000000_0000000000000000_0000110000001101_0110000111101111"; -- 0.04707920148486307
	pesos_i(1573) := b"0000000000000000_0000000000000000_0010011110111001_0001111001111100"; -- 0.15516844291258033
	pesos_i(1574) := b"1111111111111111_1111111111111111_1110111011000011_1011011000101110"; -- -0.0673261773837968
	pesos_i(1575) := b"0000000000000000_0000000000000000_0010001110011101_1111100111111010"; -- 0.139129279628921
	pesos_i(1576) := b"0000000000000000_0000000000000000_0001011101001010_1000011010100001"; -- 0.09098092487894502
	pesos_i(1577) := b"0000000000000000_0000000000000000_0001111101011001_1000010010010001"; -- 0.12245968380588429
	pesos_i(1578) := b"1111111111111111_1111111111111111_1111101011010101_1000010001010110"; -- -0.020179490074773567
	pesos_i(1579) := b"0000000000000000_0000000000000000_0001110000011110_1001100110010010"; -- 0.10984191726669619
	pesos_i(1580) := b"0000000000000000_0000000000000000_0000110001011110_0011101110010110"; -- 0.048312877765939524
	pesos_i(1581) := b"1111111111111111_1111111111111111_1110001010110001_1111111010011110"; -- -0.11447151792835655
	pesos_i(1582) := b"0000000000000000_0000000000000000_0001100101100100_0010110100101101"; -- 0.09918482163640106
	pesos_i(1583) := b"0000000000000000_0000000000000000_0001011110001111_1011010110111011"; -- 0.09203658873353612
	pesos_i(1584) := b"0000000000000000_0000000000000000_0000110110011010_1111001101100010"; -- 0.05314561022338243
	pesos_i(1585) := b"0000000000000000_0000000000000000_0010100111001000_0111011110101011"; -- 0.1632151405562986
	pesos_i(1586) := b"1111111111111111_1111111111111111_1110000111011111_0011010100000011"; -- -0.11768788039149114
	pesos_i(1587) := b"0000000000000000_0000000000000000_0001110000000110_0100100010010110"; -- 0.10947087923195338
	pesos_i(1588) := b"0000000000000000_0000000000000000_0000010011101100_0010100001101111"; -- 0.019228484155004093
	pesos_i(1589) := b"1111111111111111_1111111111111111_1110111000110001_1011101110011011"; -- -0.06955363717578847
	pesos_i(1590) := b"1111111111111111_1111111111111111_1110101011110011_0100110011000100"; -- -0.08222503860921825
	pesos_i(1591) := b"1111111111111111_1111111111111111_1111110101011011_1000011100111110"; -- -0.010322139218010288
	pesos_i(1592) := b"0000000000000000_0000000000000000_0001001011000101_1100011111000110"; -- 0.0733303888084342
	pesos_i(1593) := b"1111111111111111_1111111111111111_1101111001011101_0011110000101111"; -- -0.13138984550375837
	pesos_i(1594) := b"1111111111111111_1111111111111111_1101010011010001_0111001000100111"; -- -0.1686791090560417
	pesos_i(1595) := b"0000000000000000_0000000000000000_0001001000011100_0000111110101001"; -- 0.07074067940064169
	pesos_i(1596) := b"0000000000000000_0000000000000000_0000000110100010_0001001010001101"; -- 0.006379279496273894
	pesos_i(1597) := b"1111111111111111_1111111111111111_1110100110111000_1011011111111110"; -- -0.08702516612971786
	pesos_i(1598) := b"1111111111111111_1111111111111111_1111010000010110_1100010001100011"; -- -0.04652760111105383
	pesos_i(1599) := b"1111111111111111_1111111111111111_1111010110011000_1011001111101001"; -- -0.04063869056847848
	pesos_i(1600) := b"1111111111111111_1111111111111111_1111011001001011_0010101010011110"; -- -0.03791555053159343
	pesos_i(1601) := b"0000000000000000_0000000000000000_0001111010001101_0101101010100101"; -- 0.11934439212118467
	pesos_i(1602) := b"1111111111111111_1111111111111111_1101010011101110_1001100000001001"; -- -0.16823434616906294
	pesos_i(1603) := b"1111111111111111_1111111111111111_1101111111110110_0110101001011011"; -- -0.1251462486455685
	pesos_i(1604) := b"1111111111111111_1111111111111111_1101011110001010_0000011010111011"; -- -0.15805013590492656
	pesos_i(1605) := b"1111111111111111_1111111111111111_1111101101101001_0011011110110011"; -- -0.017925757258927543
	pesos_i(1606) := b"1111111111111111_1111111111111111_1111000110100001_0001110011001000"; -- -0.05613536943603127
	pesos_i(1607) := b"1111111111111111_1111111111111111_1100101101101001_0111110010110110"; -- -0.2054216437135523
	pesos_i(1608) := b"1111111111111111_1111111111111111_1111001101111001_0010000110111010"; -- -0.04893292618101163
	pesos_i(1609) := b"1111111111111111_1111111111111111_1111111100001010_0001101011001111"; -- -0.00375206417276508
	pesos_i(1610) := b"1111111111111111_1111111111111111_1111000001100110_0000000011010111"; -- -0.060943553437935505
	pesos_i(1611) := b"0000000000000000_0000000000000000_0001110011101101_1010101011000100"; -- 0.11300151142211093
	pesos_i(1612) := b"0000000000000000_0000000000000000_0010100000001001_1111111100101000"; -- 0.15640253766575593
	pesos_i(1613) := b"0000000000000000_0000000000000000_0000101010001011_0101111011100011"; -- 0.04118912729385195
	pesos_i(1614) := b"0000000000000000_0000000000000000_0000100100100001_0100110101100010"; -- 0.03566440236453552
	pesos_i(1615) := b"0000000000000000_0000000000000000_0010000010101100_1100011100110100"; -- 0.12763638510387573
	pesos_i(1616) := b"0000000000000000_0000000000000000_0001100010000110_0110011100111100"; -- 0.09580083091952621
	pesos_i(1617) := b"0000000000000000_0000000000000000_0000111010101110_0001110111011101"; -- 0.057344309255067734
	pesos_i(1618) := b"1111111111111111_1111111111111111_1111110000010110_1100011010001111"; -- -0.015277471525326504
	pesos_i(1619) := b"0000000000000000_0000000000000000_0001000011001110_0101111100000100"; -- 0.06564897389170629
	pesos_i(1620) := b"1111111111111111_1111111111111111_1110110011001001_1001010000100000"; -- -0.07504915457298732
	pesos_i(1621) := b"0000000000000000_0000000000000000_0010100011000111_1000100100111011"; -- 0.15929467851709186
	pesos_i(1622) := b"0000000000000000_0000000000000000_0001110001101000_0010111001011001"; -- 0.1109646765009698
	pesos_i(1623) := b"0000000000000000_0000000000000000_0000101111100110_0001010110101011"; -- 0.04647956310917177
	pesos_i(1624) := b"0000000000000000_0000000000000000_0010100111000111_1001100101010100"; -- 0.163201888061936
	pesos_i(1625) := b"0000000000000000_0000000000000000_0001111000101000_1101101011111001"; -- 0.11781090346018694
	pesos_i(1626) := b"0000000000000000_0000000000000000_0000111110001001_0100110001010001"; -- 0.06068875286694574
	pesos_i(1627) := b"1111111111111111_1111111111111111_1101011000000010_0110101110001101"; -- -0.16402557196148143
	pesos_i(1628) := b"1111111111111111_1111111111111111_1110110011100101_1101000100100001"; -- -0.07461827226275508
	pesos_i(1629) := b"1111111111111111_1111111111111111_1111001110101010_1010000111001010"; -- -0.048177612562211966
	pesos_i(1630) := b"1111111111111111_1111111111111111_1101001110001111_1010110111010110"; -- -0.1735888817409888
	pesos_i(1631) := b"1111111111111111_1111111111111111_1110000001011101_0101010100110100"; -- -0.12357585423025796
	pesos_i(1632) := b"0000000000000000_0000000000000000_0001001010010010_0001101111101101"; -- 0.07254194767369446
	pesos_i(1633) := b"0000000000000000_0000000000000000_0001000000101100_1000001100011011"; -- 0.0631792012058485
	pesos_i(1634) := b"1111111111111111_1111111111111111_1101011100001000_1010100011111001"; -- -0.16002410819230303
	pesos_i(1635) := b"1111111111111111_1111111111111111_1111010000001100_0111001011010101"; -- -0.04668504996812945
	pesos_i(1636) := b"1111111111111111_1111111111111111_1101100011110011_1111110001101000"; -- -0.15252706958854756
	pesos_i(1637) := b"1111111111111111_1111111111111111_1110000111001000_0010001001101100"; -- -0.11803994053216046
	pesos_i(1638) := b"1111111111111111_1111111111111111_1110111001100001_0011101000110111"; -- -0.06882892768015651
	pesos_i(1639) := b"1111111111111111_1111111111111111_1111011001001101_0010010111110000"; -- -0.037885311928785
	pesos_i(1640) := b"1111111111111111_1111111111111111_1111100011001001_1000011100010000"; -- -0.028174932951804593
	pesos_i(1641) := b"0000000000000000_0000000000000000_0000111000001001_1110111110000001"; -- 0.05483910469342127
	pesos_i(1642) := b"1111111111111111_1111111111111111_1111110100111101_0110111100000011"; -- -0.010781347161920245
	pesos_i(1643) := b"1111111111111111_1111111111111111_1110110101001111_0101110011101111"; -- -0.07300776631931116
	pesos_i(1644) := b"0000000000000000_0000000000000000_0010101000001000_0011010000101010"; -- 0.16418767953383315
	pesos_i(1645) := b"0000000000000000_0000000000000000_0000100001010101_1011010101000100"; -- 0.03255780136825506
	pesos_i(1646) := b"1111111111111111_1111111111111111_1110011101011100_0010011000101000"; -- -0.09625016710263873
	pesos_i(1647) := b"1111111111111111_1111111111111111_1101010001011001_1110111010010110"; -- -0.17050274682921437
	pesos_i(1648) := b"0000000000000000_0000000000000000_0010001000001110_1101100100010010"; -- 0.133039061392529
	pesos_i(1649) := b"1111111111111111_1111111111111111_1110100110100001_0111110000000111"; -- -0.08737969232939878
	pesos_i(1650) := b"0000000000000000_0000000000000000_0001110110111100_0001101101010001"; -- 0.11615153044964276
	pesos_i(1651) := b"0000000000000000_0000000000000000_0010010010110010_0010000010100011"; -- 0.14334300982287815
	pesos_i(1652) := b"0000000000000000_0000000000000000_0010001001101100_1000010000111101"; -- 0.13446833118974802
	pesos_i(1653) := b"1111111111111111_1111111111111111_1110111100011101_1101001111101110"; -- -0.06595111313218935
	pesos_i(1654) := b"1111111111111111_1111111111111111_1111010101111011_0101011001111111"; -- -0.04108676335418267
	pesos_i(1655) := b"1111111111111111_1111111111111111_1111101001001001_1000110011000001"; -- -0.02231521877404631
	pesos_i(1656) := b"1111111111111111_1111111111111111_1111010100101010_0000101101010001"; -- -0.042327206289176744
	pesos_i(1657) := b"1111111111111111_1111111111111111_1111110111111111_1001010101100001"; -- -0.007818855065611661
	pesos_i(1658) := b"1111111111111111_1111111111111111_1101011110100011_0011010111001110"; -- -0.15766586046849085
	pesos_i(1659) := b"0000000000000000_0000000000000000_0010000111010011_1011000101101101"; -- 0.13213642992362
	pesos_i(1660) := b"0000000000000000_0000000000000000_0001111101011100_1000011101110111"; -- 0.1225056329845741
	pesos_i(1661) := b"0000000000000000_0000000000000000_0010011001001011_1100010111111011"; -- 0.14959370978713862
	pesos_i(1662) := b"1111111111111111_1111111111111111_1101100010110000_1000100100110111"; -- -0.15355627438000352
	pesos_i(1663) := b"1111111111111111_1111111111111111_1110100010110001_0100100011011010"; -- -0.09104485198273449
	pesos_i(1664) := b"1111111111111111_1111111111111111_1110010111101100_1101011110110110"; -- -0.10185481834056198
	pesos_i(1665) := b"1111111111111111_1111111111111111_1110110000110000_1101011100101010"; -- -0.07737975339387451
	pesos_i(1666) := b"1111111111111111_1111111111111111_1111101101011111_1010100010101011"; -- -0.01807161162565645
	pesos_i(1667) := b"0000000000000000_0000000000000000_0001011100110000_0011110110110111"; -- 0.0905798503758528
	pesos_i(1668) := b"0000000000000000_0000000000000000_0010001011001011_0110000001000001"; -- 0.13591577137217753
	pesos_i(1669) := b"1111111111111111_1111111111111111_1110110100010000_0101010101000011"; -- -0.07396952746497856
	pesos_i(1670) := b"1111111111111111_1111111111111111_1111001010010111_1000011001101101"; -- -0.052375410441100397
	pesos_i(1671) := b"1111111111111111_1111111111111111_1110101010111100_0010000110100110"; -- -0.08306684198237764
	pesos_i(1672) := b"0000000000000000_0000000000000000_0000111001111101_1011010111000111"; -- 0.056605683386763694
	pesos_i(1673) := b"1111111111111111_1111111111111111_1111110010010110_0110000111000100"; -- -0.013330354457523655
	pesos_i(1674) := b"0000000000000000_0000000000000000_0001101110111101_0111101101111110"; -- 0.10836002178569566
	pesos_i(1675) := b"0000000000000000_0000000000000000_0010001111111011_0111101110110110"; -- 0.14055607983481402
	pesos_i(1676) := b"1111111111111111_1111111111111111_1111100100110001_0111010111010000"; -- -0.026589047245872906
	pesos_i(1677) := b"1111111111111111_1111111111111111_1101001100011101_0110010000000010"; -- -0.17533278408692776
	pesos_i(1678) := b"1111111111111111_1111111111111111_1101011000101111_1000011011101101"; -- -0.16333729465893085
	pesos_i(1679) := b"0000000000000000_0000000000000000_0000111011000101_1001001000100100"; -- 0.05770219207675224
	pesos_i(1680) := b"0000000000000000_0000000000000000_0000111000001101_1001100000001001"; -- 0.05489492620415287
	pesos_i(1681) := b"0000000000000000_0000000000000000_0001010010000010_1001100000110011"; -- 0.08011771444499177
	pesos_i(1682) := b"0000000000000000_0000000000000000_0010000000000100_1110101110110001"; -- 0.12507508352212388
	pesos_i(1683) := b"0000000000000000_0000000000000000_0001000000111000_1100111100001101"; -- 0.0633668333671856
	pesos_i(1684) := b"0000000000000000_0000000000000000_0001011010001001_1111111011001111"; -- 0.08804314185014792
	pesos_i(1685) := b"1111111111111111_1111111111111111_1111010000010101_1111100000001001"; -- -0.04653978142197135
	pesos_i(1686) := b"0000000000000000_0000000000000000_0001010101001111_1111001000000011"; -- 0.08325111929109663
	pesos_i(1687) := b"1111111111111111_1111111111111111_1101101101111111_1111011001001100"; -- -0.14257870340537976
	pesos_i(1688) := b"0000000000000000_0000000000000000_0000110001110100_1110010001010001"; -- 0.0486586282069459
	pesos_i(1689) := b"1111111111111111_1111111111111111_1111011011001001_1001011100001100"; -- -0.035986480368497796
	pesos_i(1690) := b"0000000000000000_0000000000000000_0001011100111010_1100001010001110"; -- 0.09074035620074791
	pesos_i(1691) := b"0000000000000000_0000000000000000_0000001011100000_0111110100101001"; -- 0.011237928967255199
	pesos_i(1692) := b"1111111111111111_1111111111111111_1111001111000010_1110111011110010"; -- -0.0478068027778893
	pesos_i(1693) := b"0000000000000000_0000000000000000_0010001011001111_0101001011101101"; -- 0.13597601208926646
	pesos_i(1694) := b"1111111111111111_1111111111111111_1110101110000011_1010101001011101"; -- -0.08002219421705177
	pesos_i(1695) := b"0000000000000000_0000000000000000_0010000111001101_0100011100011011"; -- 0.13203853987149047
	pesos_i(1696) := b"0000000000000000_0000000000000000_0000100000110101_1011010111001110"; -- 0.032069552257142614
	pesos_i(1697) := b"0000000000000000_0000000000000000_0000011011010100_0011010100001011"; -- 0.026675524888257866
	pesos_i(1698) := b"1111111111111111_1111111111111111_1111001111001111_0010100111100100"; -- -0.047620183684983795
	pesos_i(1699) := b"0000000000000000_0000000000000000_0000100011001111_0101100110000100"; -- 0.03441390495705051
	pesos_i(1700) := b"0000000000000000_0000000000000000_0010010011000000_0101000100100110"; -- 0.14355952440412592
	pesos_i(1701) := b"0000000000000000_0000000000000000_0001111000111010_1010000010101010"; -- 0.11808208605921078
	pesos_i(1702) := b"1111111111111111_1111111111111111_1101100100010110_1101000001010010"; -- -0.1519956397895736
	pesos_i(1703) := b"0000000000000000_0000000000000000_0000111010010011_1111111000001000"; -- 0.056945683453306584
	pesos_i(1704) := b"0000000000000000_0000000000000000_0000000110001110_1000010001110100"; -- 0.0060808928661237605
	pesos_i(1705) := b"1111111111111111_1111111111111111_1110011011101001_0100110111000000"; -- -0.0980025679354762
	pesos_i(1706) := b"0000000000000000_0000000000000000_0010001110111000_0000111011100100"; -- 0.13952725480692227
	pesos_i(1707) := b"1111111111111111_1111111111111111_1110011110011011_0100100001000010"; -- -0.09528683077578444
	pesos_i(1708) := b"0000000000000000_0000000000000000_0001100111010101_0101001010011110"; -- 0.10091129633489736
	pesos_i(1709) := b"1111111111111111_1111111111111111_1111000011101000_1001110001011011"; -- -0.058950641321679535
	pesos_i(1710) := b"1111111111111111_1111111111111111_1100100101110001_0010011101000110"; -- -0.21311716586204182
	pesos_i(1711) := b"0000000000000000_0000000000000000_0010101000010100_1011010110000101"; -- 0.16437849507856872
	pesos_i(1712) := b"1111111111111111_1111111111111111_1111011101011011_1000001100000010"; -- -0.03375989146525557
	pesos_i(1713) := b"0000000000000000_0000000000000000_0000000010110001_0011011110000011"; -- 0.002704114369737234
	pesos_i(1714) := b"0000000000000000_0000000000000000_0000100111110110_0101110000101010"; -- 0.03891540559289184
	pesos_i(1715) := b"1111111111111111_1111111111111111_1110011010100000_1101001101101101"; -- -0.09910849168886154
	pesos_i(1716) := b"1111111111111111_1111111111111111_1101100001011110_0001110110011111"; -- -0.15481390830546882
	pesos_i(1717) := b"0000000000000000_0000000000000000_0010101001100101_0101100000111010"; -- 0.1656088963158975
	pesos_i(1718) := b"1111111111111111_1111111111111111_1111111001010011_1111001111011011"; -- -0.006531485640636406
	pesos_i(1719) := b"1111111111111111_1111111111111111_1101111010101101_1101011110010111"; -- -0.13015987922195316
	pesos_i(1720) := b"1111111111111111_1111111111111111_1111011010001011_1011101101100010"; -- -0.036930359517664824
	pesos_i(1721) := b"0000000000000000_0000000000000000_0000111010010110_0110000011111000"; -- 0.056982098199756005
	pesos_i(1722) := b"1111111111111111_1111111111111111_1101111001111110_0101111101011001"; -- -0.1308842095121119
	pesos_i(1723) := b"0000000000000000_0000000000000000_0000110111001101_0101011101010101"; -- 0.05391450725513755
	pesos_i(1724) := b"1111111111111111_1111111111111111_1101100101000100_0101110100001101"; -- -0.15130060619125554
	pesos_i(1725) := b"1111111111111111_1111111111111111_1110100110111001_1110110010001010"; -- -0.0870067753007816
	pesos_i(1726) := b"0000000000000000_0000000000000000_0001111011101000_1111110111000010"; -- 0.12074266424436585
	pesos_i(1727) := b"1111111111111111_1111111111111111_1101000110000011_0101110001000101"; -- -0.18158934892271583
	pesos_i(1728) := b"1111111111111111_1111111111111111_1111001011000000_0000111110010101"; -- -0.051756883733360154
	pesos_i(1729) := b"0000000000000000_0000000000000000_0001111100100100_0111110100001011"; -- 0.12165051957052374
	pesos_i(1730) := b"1111111111111111_1111111111111111_1101110001011111_1011011011001010"; -- -0.13916451995857715
	pesos_i(1731) := b"0000000000000000_0000000000000000_0001100101011111_1110001111011010"; -- 0.0991194158622606
	pesos_i(1732) := b"1111111111111111_1111111111111111_1111001111011100_0000101011101010"; -- -0.0474236659678067
	pesos_i(1733) := b"1111111111111111_1111111111111111_1111000110001001_1011110011011000"; -- -0.05649203983432021
	pesos_i(1734) := b"1111111111111111_1111111111111111_1110110101101010_0011011011011101"; -- -0.07259804834311752
	pesos_i(1735) := b"0000000000000000_0000000000000000_0000111110110000_0101000010000010"; -- 0.061284095610344334
	pesos_i(1736) := b"0000000000000000_0000000000000000_0001100000101011_0001001100011110"; -- 0.09440726744407565
	pesos_i(1737) := b"1111111111111111_1111111111111111_1110000110100000_1001001110001101"; -- -0.11864354909383407
	pesos_i(1738) := b"0000000000000000_0000000000000000_0000100111010011_1011011111001000"; -- 0.0383868086407304
	pesos_i(1739) := b"0000000000000000_0000000000000000_0000101111100110_1111000000010100"; -- 0.04649258130142464
	pesos_i(1740) := b"1111111111111111_1111111111111111_1111101110110101_1110011010110110"; -- -0.016755657625607254
	pesos_i(1741) := b"0000000000000000_0000000000000000_0010100001101100_0001111101000111"; -- 0.15789981352891855
	pesos_i(1742) := b"0000000000000000_0000000000000000_0001011111011000_1110111110011110"; -- 0.0931539308230333
	pesos_i(1743) := b"0000000000000000_0000000000000000_0010010011001001_1011100111010000"; -- 0.1437030918281923
	pesos_i(1744) := b"1111111111111111_1111111111111111_1111000100001101_0000001111101000"; -- -0.058395152873382775
	pesos_i(1745) := b"1111111111111111_1111111111111111_1111100000111011_1001100011000010"; -- -0.030340626476127473
	pesos_i(1746) := b"1111111111111111_1111111111111111_1111001111010010_1010101111011011"; -- -0.04756666089316749
	pesos_i(1747) := b"1111111111111111_1111111111111111_1110011000010110_0110101010101101"; -- -0.10122044835778295
	pesos_i(1748) := b"0000000000000000_0000000000000000_0010110011000001_1010111010100000"; -- 0.17483035481266831
	pesos_i(1749) := b"1111111111111111_1111111111111111_1110101000101001_1111111011110100"; -- -0.08529669336043749
	pesos_i(1750) := b"0000000000000000_0000000000000000_0001110111110101_0010110111010100"; -- 0.11702238483326122
	pesos_i(1751) := b"1111111111111111_1111111111111111_1111100110110001_1011101111001110"; -- -0.024631750203090393
	pesos_i(1752) := b"0000000000000000_0000000000000000_0000001101111101_0111000111100101"; -- 0.01363288734355629
	pesos_i(1753) := b"0000000000000000_0000000000000000_0000011101101110_1110110110010111"; -- 0.02903637824498213
	pesos_i(1754) := b"1111111111111111_1111111111111111_1110000001010001_1001000000100011"; -- -0.12375544681196728
	pesos_i(1755) := b"0000000000000000_0000000000000000_0000111101000000_1100101101000011"; -- 0.05958242774767805
	pesos_i(1756) := b"0000000000000000_0000000000000000_0000111110101110_0100101001010111"; -- 0.0612532104051584
	pesos_i(1757) := b"1111111111111111_1111111111111111_1110001000111000_1101011101100011"; -- -0.11632016986079587
	pesos_i(1758) := b"1111111111111111_1111111111111111_1111000001011001_1100001000101100"; -- -0.06113039413552518
	pesos_i(1759) := b"0000000000000000_0000000000000000_0010110100100000_0100000011100010"; -- 0.17627339860956273
	pesos_i(1760) := b"1111111111111111_1111111111111111_1101101101110110_1000010011000111"; -- -0.1427227988583812
	pesos_i(1761) := b"0000000000000000_0000000000000000_0001000001110011_0101000111010100"; -- 0.06425963818796207
	pesos_i(1762) := b"1111111111111111_1111111111111111_1111010011100000_0110000011010010"; -- -0.04345126041234408
	pesos_i(1763) := b"1111111111111111_1111111111111111_1101111001101010_0100010010011000"; -- -0.13119097977970676
	pesos_i(1764) := b"0000000000000000_0000000000000000_0001011110101001_0111001000000011"; -- 0.09242928089037808
	pesos_i(1765) := b"1111111111111111_1111111111111111_1110110010000000_1100011010100000"; -- -0.07616003597286385
	pesos_i(1766) := b"0000000000000000_0000000000000000_0001001111100110_0110001010000100"; -- 0.07773414358454067
	pesos_i(1767) := b"0000000000000000_0000000000000000_0001110011101011_0111101010000101"; -- 0.11296811812493238
	pesos_i(1768) := b"0000000000000000_0000000000000000_0001110111000100_1110011111101011"; -- 0.11628579595069291
	pesos_i(1769) := b"0000000000000000_0000000000000000_0000111010011011_1100010010111110"; -- 0.05706433912479368
	pesos_i(1770) := b"0000000000000000_0000000000000000_0010010011010100_0100001001011101"; -- 0.14386381878754861
	pesos_i(1771) := b"1111111111111111_1111111111111111_1101010110110101_0110010110100001"; -- -0.16520085162430942
	pesos_i(1772) := b"1111111111111111_1111111111111111_1110000111001110_0010101010010111"; -- -0.11794790094970632
	pesos_i(1773) := b"1111111111111111_1111111111111111_1111100011000111_1110111101011011"; -- -0.028199234207080055
	pesos_i(1774) := b"0000000000000000_0000000000000000_0000000111000111_0000101010110011"; -- 0.00694338676239888
	pesos_i(1775) := b"0000000000000000_0000000000000000_0001110110010110_1100001010110110"; -- 0.11558167415146547
	pesos_i(1776) := b"0000000000000000_0000000000000000_0001010100011000_0110110000111000"; -- 0.0824039113463392
	pesos_i(1777) := b"0000000000000000_0000000000000000_0010000111010110_0100011111111011"; -- 0.13217592133849587
	pesos_i(1778) := b"1111111111111111_1111111111111111_1110110011010010_0101011010111111"; -- -0.07491548383670915
	pesos_i(1779) := b"1111111111111111_1111111111111111_1101111101000001_1011011011001010"; -- -0.12790353363635937
	pesos_i(1780) := b"0000000000000000_0000000000000000_0010001111011001_0101101110110111"; -- 0.1400353737875712
	pesos_i(1781) := b"1111111111111111_1111111111111111_1110000010101001_1011100100111111"; -- -0.12241022300495176
	pesos_i(1782) := b"1111111111111111_1111111111111111_1101111001010010_1111010001101100"; -- -0.13154671052121686
	pesos_i(1783) := b"0000000000000000_0000000000000000_0000011001111100_1000100101001101"; -- 0.02533777355891842
	pesos_i(1784) := b"1111111111111111_1111111111111111_1101100101101110_0100101111001101"; -- -0.15066076506171416
	pesos_i(1785) := b"0000000000000000_0000000000000000_0001110111011010_1111100000011000"; -- 0.1166224534691417
	pesos_i(1786) := b"1111111111111111_1111111111111111_1111000101110011_1100001110010000"; -- -0.056827332881397505
	pesos_i(1787) := b"1111111111111111_1111111111111111_1111111001101100_0101110010100010"; -- -0.006159029489122067
	pesos_i(1788) := b"0000000000000000_0000000000000000_0000001010111000_1101011001001101"; -- 0.010632890624867206
	pesos_i(1789) := b"0000000000000000_0000000000000000_0001010000100001_1111010000001000"; -- 0.07864308546287312
	pesos_i(1790) := b"1111111111111111_1111111111111111_1101011010000010_0001101011011110"; -- -0.16207725593014483
	pesos_i(1791) := b"0000000000000000_0000000000000000_0000011110100011_0000111010011111"; -- 0.02983180415600135
	pesos_i(1792) := b"0000000000000000_0000000000000000_0000111110101010_0011001011101101"; -- 0.06119077955630331
	pesos_i(1793) := b"1111111111111111_1111111111111111_1101100111001000_1100001000010101"; -- -0.1492804239709488
	pesos_i(1794) := b"0000000000000000_0000000000000000_0010100100001100_0001100010110111"; -- 0.16034082863472268
	pesos_i(1795) := b"0000000000000000_0000000000000000_0001110101000011_0011101100000000"; -- 0.1143071055934564
	pesos_i(1796) := b"0000000000000000_0000000000000000_0000110101100101_1000011111001001"; -- 0.05233048101121252
	pesos_i(1797) := b"0000000000000000_0000000000000000_0010010100111100_1111011100010000"; -- 0.14546150351366496
	pesos_i(1798) := b"0000000000000000_0000000000000000_0000001100000101_0001010100001010"; -- 0.011796297939214419
	pesos_i(1799) := b"0000000000000000_0000000000000000_0000010101111011_1100101010110110"; -- 0.021420163473970362
	pesos_i(1800) := b"0000000000000000_0000000000000000_0000110100001010_1010100111011111"; -- 0.0509439630596992
	pesos_i(1801) := b"1111111111111111_1111111111111111_1111010111010111_1111010110111000"; -- -0.03967346441911802
	pesos_i(1802) := b"1111111111111111_1111111111111111_1111100100000011_0001000001011001"; -- -0.027296999286341276
	pesos_i(1803) := b"0000000000000000_0000000000000000_0000110001110011_0000000100011010"; -- 0.04862982630894419
	pesos_i(1804) := b"1111111111111111_1111111111111111_1101101111011000_0110000101100011"; -- -0.14122954682358224
	pesos_i(1805) := b"1111111111111111_1111111111111111_1101010101100000_1111101110111111"; -- -0.16648890112015768
	pesos_i(1806) := b"1111111111111111_1111111111111111_1101001010011010_1111101100101011"; -- -0.17732267578363067
	pesos_i(1807) := b"0000000000000000_0000000000000000_0001110010001101_0011010000111011"; -- 0.11152960247695169
	pesos_i(1808) := b"0000000000000000_0000000000000000_0000111110110000_1110000111010101"; -- 0.06129275744996873
	pesos_i(1809) := b"1111111111111111_1111111111111111_1110000001011110_0101011100110101"; -- -0.1235604758922434
	pesos_i(1810) := b"1111111111111111_1111111111111111_1110010111001110_1001101011111000"; -- -0.10231620251591253
	pesos_i(1811) := b"0000000000000000_0000000000000000_0001100010010011_0111011100111000"; -- 0.0960001480378336
	pesos_i(1812) := b"0000000000000000_0000000000000000_0000000011110010_0010110111100010"; -- 0.003695361666452725
	pesos_i(1813) := b"0000000000000000_0000000000000000_0001010101000100_0010110100101111"; -- 0.08307154089419663
	pesos_i(1814) := b"0000000000000000_0000000000000000_0000100000111111_0011011011110111"; -- 0.03221457984559153
	pesos_i(1815) := b"0000000000000000_0000000000000000_0001110101110000_1011001011100001"; -- 0.11500089629622037
	pesos_i(1816) := b"0000000000000000_0000000000000000_0000100001011110_1011110000010001"; -- 0.03269553589788615
	pesos_i(1817) := b"1111111111111111_1111111111111111_1111010011010011_1101001101000111"; -- -0.04364280248209123
	pesos_i(1818) := b"0000000000000000_0000000000000000_0010010011001110_1011111100101011"; -- 0.14377970501958293
	pesos_i(1819) := b"0000000000000000_0000000000000000_0000111110110010_0010100101000101"; -- 0.061312274254473526
	pesos_i(1820) := b"0000000000000000_0000000000000000_0010010111000100_1100000011010010"; -- 0.14753346571976167
	pesos_i(1821) := b"0000000000000000_0000000000000000_0001110001000110_0000110011010101"; -- 0.11044388012751175
	pesos_i(1822) := b"0000000000000000_0000000000000000_0001101000101101_1010101101110000"; -- 0.10225936392172764
	pesos_i(1823) := b"1111111111111111_1111111111111111_1101101110001111_1100110000110010"; -- -0.14233707208148072
	pesos_i(1824) := b"1111111111111111_1111111111111111_1111111001001101_1010000000001000"; -- -0.006628034691788992
	pesos_i(1825) := b"1111111111111111_1111111111111111_1111101001101100_1011001100011010"; -- -0.021778875485434973
	pesos_i(1826) := b"0000000000000000_0000000000000000_0010000100000001_0110100101000110"; -- 0.12892778347945696
	pesos_i(1827) := b"0000000000000000_0000000000000000_0000101101111001_0100101111001010"; -- 0.04481958077550599
	pesos_i(1828) := b"0000000000000000_0000000000000000_0010001101101010_1000011110110000"; -- 0.13834426922831294
	pesos_i(1829) := b"0000000000000000_0000000000000000_0000101000100001_1000000000100110"; -- 0.03957367831490843
	pesos_i(1830) := b"1111111111111111_1111111111111111_1110111011111000_1000110010011010"; -- -0.06651993980089303
	pesos_i(1831) := b"0000000000000000_0000000000000000_0001101001011110_1111111100001110"; -- 0.10301202862071482
	pesos_i(1832) := b"0000000000000000_0000000000000000_0010011010110111_0010010111111011"; -- 0.15123212213273493
	pesos_i(1833) := b"0000000000000000_0000000000000000_0010100010010111_1110000010001000"; -- 0.15856746029399468
	pesos_i(1834) := b"1111111111111111_1111111111111111_1101011111111010_1011111010001000"; -- -0.15633019625567499
	pesos_i(1835) := b"1111111111111111_1111111111111111_1101101011111110_0110011100001010"; -- -0.1445556258895361
	pesos_i(1836) := b"1111111111111111_1111111111111111_1101001001111010_0000000100011111"; -- -0.17782586081103668
	pesos_i(1837) := b"1111111111111111_1111111111111111_1101100011101101_0011110010000000"; -- -0.152630060796031
	pesos_i(1838) := b"0000000000000000_0000000000000000_0000101100001110_1111111110111100"; -- 0.04319761601792568
	pesos_i(1839) := b"1111111111111111_1111111111111111_1100111101000010_1110000010111011"; -- -0.19038577492186456
	pesos_i(1840) := b"0000000000000000_0000000000000000_0000100101001101_1000110011000110"; -- 0.03633956762165666
	pesos_i(1841) := b"1111111111111111_1111111111111111_1101100000010100_1101000010010001"; -- -0.1559323926631963
	pesos_i(1842) := b"1111111111111111_1111111111111111_1111110001111010_1001011001100110"; -- -0.013754463403941975
	pesos_i(1843) := b"0000000000000000_0000000000000000_0010000100111011_1100111010011000"; -- 0.12981883260019245
	pesos_i(1844) := b"0000000000000000_0000000000000000_0010100110101101_0111001100110101"; -- 0.16280288735032414
	pesos_i(1845) := b"0000000000000000_0000000000000000_0000001100001100_1010011010101001"; -- 0.011911789225761592
	pesos_i(1846) := b"0000000000000000_0000000000000000_0010010000111001_0010111110011100"; -- 0.14149758862772635
	pesos_i(1847) := b"1111111111111111_1111111111111111_1110110001011001_0110001011111100"; -- -0.07676106780893528
	pesos_i(1848) := b"1111111111111111_1111111111111111_1111000000111110_0000010110001101"; -- -0.0615536243209857
	pesos_i(1849) := b"1111111111111111_1111111111111111_1111110011100000_0010100110011110"; -- -0.012204550590462028
	pesos_i(1850) := b"1111111111111111_1111111111111111_1101010000011101_0101100111111010"; -- -0.17142713211883062
	pesos_i(1851) := b"0000000000000000_0000000000000000_0000100111110001_1000000000000101"; -- 0.0388412486768172
	pesos_i(1852) := b"0000000000000000_0000000000000000_0000000000010001_1111011001000000"; -- 0.00027407711663866266
	pesos_i(1853) := b"0000000000000000_0000000000000000_0000100000000110_1101001010001010"; -- 0.03135410173710482
	pesos_i(1854) := b"1111111111111111_1111111111111111_1110000011100110_1101101100011010"; -- -0.12147741914350935
	pesos_i(1855) := b"1111111111111111_1111111111111111_1110111100111100_0000000010110010"; -- -0.06549068128300745
	pesos_i(1856) := b"0000000000000000_0000000000000000_0000100110000110_0000101001111100"; -- 0.03720155265717237
	pesos_i(1857) := b"0000000000000000_0000000000000000_0001000111010000_0111010101110111"; -- 0.06958707963116925
	pesos_i(1858) := b"0000000000000000_0000000000000000_0000111010101111_0000010100111000"; -- 0.0573580990944305
	pesos_i(1859) := b"1111111111111111_1111111111111111_1111011101000100_0101101000010000"; -- -0.03411328424301386
	pesos_i(1860) := b"0000000000000000_0000000000000000_0000100110010001_1100011111101011"; -- 0.0373806904823338
	pesos_i(1861) := b"1111111111111111_1111111111111111_1110000100111000_1000111110001111"; -- -0.12023070102145797
	pesos_i(1862) := b"0000000000000000_0000000000000000_0001100101000111_1101001000000001"; -- 0.0987521411876143
	pesos_i(1863) := b"0000000000000000_0000000000000000_0001001000101000_0011000010100010"; -- 0.07092575019579185
	pesos_i(1864) := b"1111111111111111_1111111111111111_1110110101101011_0001011100100101"; -- -0.07258468009748631
	pesos_i(1865) := b"1111111111111111_1111111111111111_1111000001100011_1101000000010011"; -- -0.060976977615506085
	pesos_i(1866) := b"1111111111111111_1111111111111111_1110011010100100_0111011000000100"; -- -0.09905302423797137
	pesos_i(1867) := b"0000000000000000_0000000000000000_0000011001001101_1101001000101001"; -- 0.024624953185633965
	pesos_i(1868) := b"1111111111111111_1111111111111111_1110000000110111_1011001001100100"; -- -0.1241501337885814
	pesos_i(1869) := b"1111111111111111_1111111111111111_1110010100010011_0101111000100010"; -- -0.10517322222713313
	pesos_i(1870) := b"1111111111111111_1111111111111111_1101011010110010_1000001000010111"; -- -0.16133868154424147
	pesos_i(1871) := b"0000000000000000_0000000000000000_0000011010100001_0010101011000011"; -- 0.025896713863470575
	pesos_i(1872) := b"1111111111111111_1111111111111111_1101010101101010_1001100001110000"; -- -0.16634223233729256
	pesos_i(1873) := b"1111111111111111_1111111111111111_1101100000101000_1001110000010011"; -- -0.15563034567381986
	pesos_i(1874) := b"1111111111111111_1111111111111111_1101111011001000_1110100110001110"; -- -0.12974682123031128
	pesos_i(1875) := b"1111111111111111_1111111111111111_1101110101100011_0111110000111111"; -- -0.1352007242737983
	pesos_i(1876) := b"1111111111111111_1111111111111111_1110000010010101_0111011010010100"; -- -0.12271937263644242
	pesos_i(1877) := b"1111111111111111_1111111111111111_1110000001001010_1010010011011110"; -- -0.12386102272963968
	pesos_i(1878) := b"0000000000000000_0000000000000000_0010011010101101_0010001100101010"; -- 0.15107936650429624
	pesos_i(1879) := b"0000000000000000_0000000000000000_0001001001000101_0010100011010001"; -- 0.0713677893339084
	pesos_i(1880) := b"0000000000000000_0000000000000000_0001010010110100_0001000101001100"; -- 0.08087261302248581
	pesos_i(1881) := b"1111111111111111_1111111111111111_1111110010111000_1100110000001010"; -- -0.012805221086686093
	pesos_i(1882) := b"1111111111111111_1111111111111111_1101010110110000_0001111100110001"; -- -0.165281343918724
	pesos_i(1883) := b"0000000000000000_0000000000000000_0001000011000010_0010100110111000"; -- 0.06546269178014481
	pesos_i(1884) := b"1111111111111111_1111111111111111_1101100100110000_1100011010011101"; -- -0.15159948991322544
	pesos_i(1885) := b"0000000000000000_0000000000000000_0001111100100101_1111110111111010"; -- 0.12167346340822095
	pesos_i(1886) := b"0000000000000000_0000000000000000_0000100111001110_1001001011110011"; -- 0.03830831929765845
	pesos_i(1887) := b"1111111111111111_1111111111111111_1111110101111100_1110101110101110"; -- -0.00981261263447017
	pesos_i(1888) := b"0000000000000000_0000000000000000_0000101000101010_1111000000001101"; -- 0.03971767718060379
	pesos_i(1889) := b"0000000000000000_0000000000000000_0001000101011111_0010110101111101"; -- 0.06785854627837043
	pesos_i(1890) := b"1111111111111111_1111111111111111_1111010010001010_1010011001011001"; -- -0.04475937203514719
	pesos_i(1891) := b"0000000000000000_0000000000000000_0010100000110011_0010001010100011"; -- 0.15703026269924927
	pesos_i(1892) := b"1111111111111111_1111111111111111_1111100010110010_1111001010110101"; -- -0.028519469169573014
	pesos_i(1893) := b"0000000000000000_0000000000000000_0001000011101000_0001000100001010"; -- 0.06604105458159307
	pesos_i(1894) := b"0000000000000000_0000000000000000_0010001101001111_1000010001100001"; -- 0.1379320848242947
	pesos_i(1895) := b"0000000000000000_0000000000000000_0010010011110110_0101011000101011"; -- 0.14438379815738636
	pesos_i(1896) := b"0000000000000000_0000000000000000_0000000001100110_0100001000111001"; -- 0.0015603437333068793
	pesos_i(1897) := b"0000000000000000_0000000000000000_0000000011110100_0110010001001011"; -- 0.0037291224447702728
	pesos_i(1898) := b"1111111111111111_1111111111111111_1101011101100101_0011010100110001"; -- -0.158611941944477
	pesos_i(1899) := b"1111111111111111_1111111111111111_1101101110010011_1010100111111101"; -- -0.1422780758267724
	pesos_i(1900) := b"0000000000000000_0000000000000000_0000111100011111_0001101000111101"; -- 0.05906833637795175
	pesos_i(1901) := b"1111111111111111_1111111111111111_1101111100010000_1110101001101010"; -- -0.12864813726716598
	pesos_i(1902) := b"1111111111111111_1111111111111111_1110110011011011_1100001010110011"; -- -0.07477172033386648
	pesos_i(1903) := b"1111111111111111_1111111111111111_1110001011000100_0110010100001000"; -- -0.11419075539515258
	pesos_i(1904) := b"0000000000000000_0000000000000000_0000110101011100_1011001100011001"; -- 0.05219573372200256
	pesos_i(1905) := b"0000000000000000_0000000000000000_0000000100101001_1101111001010001"; -- 0.004545111383155448
	pesos_i(1906) := b"0000000000000000_0000000000000000_0001001000010111_0011011100001101"; -- 0.07066673341756784
	pesos_i(1907) := b"0000000000000000_0000000000000000_0010100011111010_0101100011000111"; -- 0.16006998881935403
	pesos_i(1908) := b"0000000000000000_0000000000000000_0000000110101100_1110001110101101"; -- 0.00654433233660492
	pesos_i(1909) := b"0000000000000000_0000000000000000_0000000110001111_1010101110000111"; -- 0.00609848073266072
	pesos_i(1910) := b"0000000000000000_0000000000000000_0000101011111011_1100000001010001"; -- 0.042903919051431476
	pesos_i(1911) := b"0000000000000000_0000000000000000_0010100000100000_0001101111001100"; -- 0.1567399381038998
	pesos_i(1912) := b"0000000000000000_0000000000000000_0001110110111011_0001111011100001"; -- 0.11613648418663738
	pesos_i(1913) := b"0000000000000000_0000000000000000_0000100000101011_0010010101110010"; -- 0.03190835986945847
	pesos_i(1914) := b"1111111111111111_1111111111111111_1111000100010100_0011100101101111"; -- -0.0582851509051261
	pesos_i(1915) := b"0000000000000000_0000000000000000_0001101011111011_0110111010011101"; -- 0.10539904901604225
	pesos_i(1916) := b"1111111111111111_1111111111111111_1110001100101100_0110011110100100"; -- -0.1126036859099877
	pesos_i(1917) := b"0000000000000000_0000000000000000_0001011100001110_1111000100000011"; -- 0.09007173854983992
	pesos_i(1918) := b"1111111111111111_1111111111111111_1110001000001001_0110011100011000"; -- -0.11704402592665639
	pesos_i(1919) := b"0000000000000000_0000000000000000_0000001110100000_1111110111111001"; -- 0.01417529412800856
	pesos_i(1920) := b"1111111111111111_1111111111111111_1101010000111011_1101111011101111"; -- -0.1709614434863065
	pesos_i(1921) := b"1111111111111111_1111111111111111_1101100110101000_1000101111111110"; -- -0.14977192923650934
	pesos_i(1922) := b"1111111111111111_1111111111111111_1111100001110001_0001100101010001"; -- -0.02952424782076006
	pesos_i(1923) := b"0000000000000000_0000000000000000_0001100100011001_0001101000100101"; -- 0.09803927811861518
	pesos_i(1924) := b"0000000000000000_0000000000000000_0001101000100111_1101000110100011"; -- 0.102170088136012
	pesos_i(1925) := b"0000000000000000_0000000000000000_0010100001100111_1001000010111011"; -- 0.15783028190179602
	pesos_i(1926) := b"1111111111111111_1111111111111111_1111100011011110_1010010001111000"; -- -0.027852745689684946
	pesos_i(1927) := b"0000000000000000_0000000000000000_0010001001010011_1000000010100001"; -- 0.13408664641723333
	pesos_i(1928) := b"0000000000000000_0000000000000000_0000010010000100_0101110010111001"; -- 0.01764468692629294
	pesos_i(1929) := b"0000000000000000_0000000000000000_0001001100110111_1101101110110010"; -- 0.07507107814681112
	pesos_i(1930) := b"1111111111111111_1111111111111111_1111111110001010_0111110000011111"; -- -0.0017931388753282104
	pesos_i(1931) := b"1111111111111111_1111111111111111_1101100000100101_0010110000011110"; -- -0.15568279522670972
	pesos_i(1932) := b"1111111111111111_1111111111111111_1101101111001111_1101011111111000"; -- -0.1413598078452596
	pesos_i(1933) := b"1111111111111111_1111111111111111_1101101010101110_1000110110110111"; -- -0.14577402378847532
	pesos_i(1934) := b"1111111111111111_1111111111111111_1101111010101011_0010101001101111"; -- -0.13020071788926935
	pesos_i(1935) := b"1111111111111111_1111111111111111_1110011000000101_0010000110100000"; -- -0.10148420181222359
	pesos_i(1936) := b"1111111111111111_1111111111111111_1101110001110000_1101001001100100"; -- -0.1389034753750053
	pesos_i(1937) := b"0000000000000000_0000000000000000_0001101100000100_0010111110100001"; -- 0.1055326240700306
	pesos_i(1938) := b"0000000000000000_0000000000000000_0000001000011110_1101000100010100"; -- 0.008282725592324817
	pesos_i(1939) := b"0000000000000000_0000000000000000_0000100111101111_0110111000001000"; -- 0.038809658881462546
	pesos_i(1940) := b"0000000000000000_0000000000000000_0001000001100011_1110101110010100"; -- 0.06402466166581022
	pesos_i(1941) := b"0000000000000000_0000000000000000_0010001011010101_1000110100100011"; -- 0.1360710345410395
	pesos_i(1942) := b"0000000000000000_0000000000000000_0001101011010000_0001001001000110"; -- 0.10473741739193951
	pesos_i(1943) := b"1111111111111111_1111111111111111_1111001101001011_0011101010011111"; -- -0.04963334681118704
	pesos_i(1944) := b"0000000000000000_0000000000000000_0010000011000110_1000100100110111"; -- 0.12802941895590098
	pesos_i(1945) := b"0000000000000000_0000000000000000_0000001100111101_1010001111101000"; -- 0.01265930579391574
	pesos_i(1946) := b"0000000000000000_0000000000000000_0001111010011100_1011101110010100"; -- 0.11957905151847639
	pesos_i(1947) := b"0000000000000000_0000000000000000_0001010111000100_1110011110101101"; -- 0.08503578161879696
	pesos_i(1948) := b"0000000000000000_0000000000000000_0001110111101110_1100000101000000"; -- 0.11692436036712667
	pesos_i(1949) := b"0000000000000000_0000000000000000_0001000010111011_0110100110110000"; -- 0.06535969300615711
	pesos_i(1950) := b"0000000000000000_0000000000000000_0010100110010000_1110010110010110"; -- 0.16236720007626343
	pesos_i(1951) := b"0000000000000000_0000000000000000_0010110000000101_0101100101101110"; -- 0.17195662434045902
	pesos_i(1952) := b"1111111111111111_1111111111111111_1101101101100100_1000110000111110"; -- -0.14299701206352924
	pesos_i(1953) := b"1111111111111111_1111111111111111_1111110101011101_0101101111100111"; -- -0.010294204724308559
	pesos_i(1954) := b"1111111111111111_1111111111111111_1111110100010111_1101100001011101"; -- -0.011354901539933404
	pesos_i(1955) := b"0000000000000000_0000000000000000_0010001100110101_1110101101101010"; -- 0.13754149761291073
	pesos_i(1956) := b"1111111111111111_1111111111111111_1110110111000110_0111100010110100"; -- -0.07119031518944222
	pesos_i(1957) := b"1111111111111111_1111111111111111_1111001111001110_0011011110001011"; -- -0.04763462892015347
	pesos_i(1958) := b"1111111111111111_1111111111111111_1110100111000110_0011101110001001"; -- -0.08681896125196553
	pesos_i(1959) := b"1111111111111111_1111111111111111_1111000110100100_0101110001001000"; -- -0.056085808312091825
	pesos_i(1960) := b"0000000000000000_0000000000000000_0010001010000110_0111100000101111"; -- 0.1348643412008297
	pesos_i(1961) := b"1111111111111111_1111111111111111_1110100010110110_1110111111101001"; -- -0.09095860074170582
	pesos_i(1962) := b"0000000000000000_0000000000000000_0010101100000100_1110101010111110"; -- 0.16804377690386127
	pesos_i(1963) := b"0000000000000000_0000000000000000_0001110001110111_1101001000110011"; -- 0.11120332480538792
	pesos_i(1964) := b"1111111111111111_1111111111111111_1111011011111110_0111000100010011"; -- -0.035180027880060145
	pesos_i(1965) := b"1111111111111111_1111111111111111_1110010001011101_1100011110011111"; -- -0.10794403423110915
	pesos_i(1966) := b"1111111111111111_1111111111111111_1101011111000100_0000111100111101"; -- -0.1571646191361238
	pesos_i(1967) := b"0000000000000000_0000000000000000_0010001110111111_0001101100011111"; -- 0.13963479514488367
	pesos_i(1968) := b"1111111111111111_1111111111111111_1111000101011010_0000010001000111"; -- -0.0572202039549346
	pesos_i(1969) := b"1111111111111111_1111111111111111_1101001001010000_1110101111000000"; -- -0.17845274500471564
	pesos_i(1970) := b"0000000000000000_0000000000000000_0001101101110010_0111100010110000"; -- 0.10721544544812497
	pesos_i(1971) := b"1111111111111111_1111111111111111_1110111001101111_1110001011001010"; -- -0.06860525676463115
	pesos_i(1972) := b"0000000000000000_0000000000000000_0001101011100101_0000110011111111"; -- 0.10505753740153415
	pesos_i(1973) := b"1111111111111111_1111111111111111_1111110110110111_1111001010100010"; -- -0.00891192957614535
	pesos_i(1974) := b"1111111111111111_1111111111111111_1111010010101111_1011101011100001"; -- -0.04419357300874172
	pesos_i(1975) := b"0000000000000000_0000000000000000_0001101100011100_0011101100001100"; -- 0.10589951550975152
	pesos_i(1976) := b"0000000000000000_0000000000000000_0010010001111101_1001111000100000"; -- 0.1425417736453616
	pesos_i(1977) := b"0000000000000000_0000000000000000_0001101110100111_1101100111110111"; -- 0.10802995949875356
	pesos_i(1978) := b"1111111111111111_1111111111111111_1111001000110110_1010111100101001"; -- -0.05385308506283718
	pesos_i(1979) := b"1111111111111111_1111111111111111_1110101111011000_1110101001101000"; -- -0.07872137987792391
	pesos_i(1980) := b"0000000000000000_0000000000000000_0000010101100110_0001011111101011"; -- 0.021089071992896526
	pesos_i(1981) := b"1111111111111111_1111111111111111_1111111000000110_1100101011010011"; -- -0.007708858045407788
	pesos_i(1982) := b"0000000000000000_0000000000000000_0000100111011101_1111100100000000"; -- 0.03854328383742032
	pesos_i(1983) := b"1111111111111111_1111111111111111_1101100101000111_0111000111110111"; -- -0.15125358321020388
	pesos_i(1984) := b"0000000000000000_0000000000000000_0000101101001111_1000011011000010"; -- 0.044182226472737424
	pesos_i(1985) := b"0000000000000000_0000000000000000_0010010001110100_0010111011101000"; -- 0.142397815246552
	pesos_i(1986) := b"0000000000000000_0000000000000000_0001010111111100_1100110000111101"; -- 0.08588863834987057
	pesos_i(1987) := b"1111111111111111_1111111111111111_1101111100010011_1110010101111000"; -- -0.12860265565295317
	pesos_i(1988) := b"1111111111111111_1111111111111111_1101101010100000_0101101000010111"; -- -0.14599072393801474
	pesos_i(1989) := b"0000000000000000_0000000000000000_0010101001010111_1100001000010101"; -- 0.16540158284022427
	pesos_i(1990) := b"0000000000000000_0000000000000000_0000011010010100_0110110101001010"; -- 0.025702315030700053
	pesos_i(1991) := b"0000000000000000_0000000000000000_0001101101001101_1010000111001100"; -- 0.10665332063136305
	pesos_i(1992) := b"1111111111111111_1111111111111111_1111000011011101_1101110110110000"; -- -0.05911459398829604
	pesos_i(1993) := b"1111111111111111_1111111111111111_1110111110111111_0110110000001111"; -- -0.0634853804426586
	pesos_i(1994) := b"0000000000000000_0000000000000000_0000111100110101_0110000001101000"; -- 0.059408212020515175
	pesos_i(1995) := b"1111111111111111_1111111111111111_1110100111001011_1111000000111101"; -- -0.08673189655174939
	pesos_i(1996) := b"1111111111111111_1111111111111111_1101110001110001_1111001100111000"; -- -0.13888625981356237
	pesos_i(1997) := b"0000000000000000_0000000000000000_0001110010000100_1101110111100000"; -- 0.11140238482602322
	pesos_i(1998) := b"1111111111111111_1111111111111111_1101101110101011_0100101010111101"; -- -0.14191754228269013
	pesos_i(1999) := b"1111111111111111_1111111111111111_1111111101011100_1100001111010001"; -- -0.002490769751525604
	pesos_i(2000) := b"0000000000000000_0000000000000000_0000000000110100_0011100110100001"; -- 0.000796891883658446
	pesos_i(2001) := b"0000000000000000_0000000000000000_0010001111101111_1100001001110000"; -- 0.1403771899237435
	pesos_i(2002) := b"0000000000000000_0000000000000000_0000001011111101_0011101100111101"; -- 0.011676504394961392
	pesos_i(2003) := b"1111111111111111_1111111111111111_1101110011000001_0011001100111011"; -- -0.13767700021217988
	pesos_i(2004) := b"1111111111111111_1111111111111111_1110010110000010_1100000101100101"; -- -0.10347358023659078
	pesos_i(2005) := b"1111111111111111_1111111111111111_1110111101011000_0101010001110000"; -- -0.06505844370225962
	pesos_i(2006) := b"1111111111111111_1111111111111111_1111101101010011_1100001110010011"; -- -0.018253113316455086
	pesos_i(2007) := b"0000000000000000_0000000000000000_0001101101111111_1011001001000011"; -- 0.10741724146803236
	pesos_i(2008) := b"0000000000000000_0000000000000000_0010101001000000_0000000100000000"; -- 0.16503912217425795
	pesos_i(2009) := b"0000000000000000_0000000000000000_0000000110101111_0101100101010011"; -- 0.00658186224414315
	pesos_i(2010) := b"1111111111111111_1111111111111111_1101100110111001_1100110011101001"; -- -0.14950866032431187
	pesos_i(2011) := b"1111111111111111_1111111111111111_1110010110111101_1111010010100001"; -- -0.10257025790107724
	pesos_i(2012) := b"1111111111111111_1111111111111111_1101101111010010_0110011110110101"; -- -0.14132072280180494
	pesos_i(2013) := b"0000000000000000_0000000000000000_0000011110010001_0000010111000111"; -- 0.02955661886799816
	pesos_i(2014) := b"0000000000000000_0000000000000000_0001101100101010_0010011011000000"; -- 0.10611192880955671
	pesos_i(2015) := b"0000000000000000_0000000000000000_0010001010011101_0110110011010000"; -- 0.13521461572566526
	pesos_i(2016) := b"0000000000000000_0000000000000000_0001110010101010_1010101110010010"; -- 0.11197922062152224
	pesos_i(2017) := b"0000000000000000_0000000000000000_0001001001010011_1000111111100000"; -- 0.07158755519522214
	pesos_i(2018) := b"1111111111111111_1111111111111111_1111000111000011_1110001101100110"; -- -0.0556047321503933
	pesos_i(2019) := b"1111111111111111_1111111111111111_1101100010101101_0100110100011001"; -- -0.15360563416692835
	pesos_i(2020) := b"1111111111111111_1111111111111111_1111111001010100_0101100111000110"; -- -0.006525410809821995
	pesos_i(2021) := b"0000000000000000_0000000000000000_0000011011100000_1111100010011110"; -- 0.02687028754969759
	pesos_i(2022) := b"0000000000000000_0000000000000000_0000110000100100_0011001011100010"; -- 0.0474273493239212
	pesos_i(2023) := b"0000000000000000_0000000000000000_0010001010000010_0001110011001110"; -- 0.1347978595062115
	pesos_i(2024) := b"1111111111111111_1111111111111111_1111001110001110_0111100110011001"; -- -0.048607254273453804
	pesos_i(2025) := b"1111111111111111_1111111111111111_1101111101110010_1111101100110111"; -- -0.12715177437430478
	pesos_i(2026) := b"1111111111111111_1111111111111111_1110010001010000_0011010000011111"; -- -0.10815119028240179
	pesos_i(2027) := b"0000000000000000_0000000000000000_0010000110000101_0101110011010101"; -- 0.1309412022438188
	pesos_i(2028) := b"1111111111111111_1111111111111111_1110011011001000_1001101000101001"; -- -0.09850155358162764
	pesos_i(2029) := b"0000000000000000_0000000000000000_0000100111110100_1110001110100011"; -- 0.03889296282979481
	pesos_i(2030) := b"1111111111111111_1111111111111111_1101010011000111_1011110010000011"; -- -0.1688272647634254
	pesos_i(2031) := b"0000000000000000_0000000000000000_0001111000001001_1111010111111001"; -- 0.11733949027672679
	pesos_i(2032) := b"0000000000000000_0000000000000000_0001111011001111_1111100101000001"; -- 0.12036092593395123
	pesos_i(2033) := b"1111111111111111_1111111111111111_1111110110001111_1000010000000001"; -- -0.009528875079574407
	pesos_i(2034) := b"0000000000000000_0000000000000000_0001011001001101_0001110101000011"; -- 0.08711417090822321
	pesos_i(2035) := b"1111111111111111_1111111111111111_1111111000111001_0110001110101000"; -- -0.0069368089759813505
	pesos_i(2036) := b"0000000000000000_0000000000000000_0000101010111111_0011001010110000"; -- 0.04197994997173429
	pesos_i(2037) := b"1111111111111111_1111111111111111_1101100000101010_0101001010011011"; -- -0.15560420709551617
	pesos_i(2038) := b"0000000000000000_0000000000000000_0001111110111000_0011010100010101"; -- 0.12390453118819873
	pesos_i(2039) := b"1111111111111111_1111111111111111_1110100011101001_1010000011001111"; -- -0.09018511722181898
	pesos_i(2040) := b"0000000000000000_0000000000000000_0001110000000100_1011000101110101"; -- 0.10944661238339728
	pesos_i(2041) := b"1111111111111111_1111111111111111_1110100100101001_1001111111001100"; -- -0.08920861501376615
	pesos_i(2042) := b"0000000000000000_0000000000000000_0010001101111111_1100001111111101"; -- 0.13866829792403965
	pesos_i(2043) := b"0000000000000000_0000000000000000_0010001100100010_1110010100100011"; -- 0.13725120642946545
	pesos_i(2044) := b"0000000000000000_0000000000000000_0001110010011000_1101000110110111"; -- 0.11170683591239454
	pesos_i(2045) := b"1111111111111111_1111111111111111_1110000110000000_0110000100101101"; -- -0.11913483298058633
	pesos_i(2046) := b"0000000000000000_0000000000000000_0010000100011000_0001001110011110"; -- 0.12927363017935684
	pesos_i(2047) := b"0000000000000000_0000000000000000_0000100011000111_1110000000011110"; -- 0.0342998575377427
	pesos_i(2048) := b"0000000000000000_0000000000000000_0010001010011111_0101001100100001"; -- 0.13524360232807972
	pesos_i(2049) := b"1111111111111111_1111111111111111_1111011110011111_1000001000001101"; -- -0.03272235096040199
	pesos_i(2050) := b"0000000000000000_0000000000000000_0010010010100110_0110000001100011"; -- 0.14316370415384888
	pesos_i(2051) := b"0000000000000000_0000000000000000_0000001001000011_1101010101000000"; -- 0.008847549443828965
	pesos_i(2052) := b"1111111111111111_1111111111111111_1110011111100001_0101000111010000"; -- -0.09421814597079889
	pesos_i(2053) := b"0000000000000000_0000000000000000_0000011101101100_1101100011100101"; -- 0.029004627081689743
	pesos_i(2054) := b"0000000000000000_0000000000000000_0001101010010111_0001000000110010"; -- 0.10386754246019951
	pesos_i(2055) := b"0000000000000000_0000000000000000_0001010101000111_0110111000011000"; -- 0.08312118609549458
	pesos_i(2056) := b"0000000000000000_0000000000000000_0001100011110101_0001100011000110"; -- 0.09748987998542981
	pesos_i(2057) := b"1111111111111111_1111111111111111_1101001010111010_0001001100011101"; -- -0.17684822596403513
	pesos_i(2058) := b"0000000000000000_0000000000000000_0010011001000101_1011101011001110"; -- 0.1495014908197393
	pesos_i(2059) := b"1111111111111111_1111111111111111_1101010010011010_0011000100011011"; -- -0.16952221966337416
	pesos_i(2060) := b"0000000000000000_0000000000000000_0001010110001110_1000001000100010"; -- 0.08420575451680606
	pesos_i(2061) := b"0000000000000000_0000000000000000_0010101101010000_0011001001100100"; -- 0.1691924565816401
	pesos_i(2062) := b"0000000000000000_0000000000000000_0010101110001011_1000000101011001"; -- 0.17009743143966005
	pesos_i(2063) := b"0000000000000000_0000000000000000_0001001101101101_0001001011111010"; -- 0.07588308914074876
	pesos_i(2064) := b"0000000000000000_0000000000000000_0001111110111011_0101001101011100"; -- 0.12395211223085487
	pesos_i(2065) := b"0000000000000000_0000000000000000_0010100001110110_0110000001001011"; -- 0.1580562766846676
	pesos_i(2066) := b"1111111111111111_1111111111111111_1110001111101010_1111000100110001"; -- -0.10969631732751615
	pesos_i(2067) := b"1111111111111111_1111111111111111_1110010000111100_1100011011010010"; -- -0.10844762210164323
	pesos_i(2068) := b"1111111111111111_1111111111111111_1111001010110101_0001010111011111"; -- -0.05192435547997167
	pesos_i(2069) := b"1111111111111111_1111111111111111_1110001001111010_0101010001000101"; -- -0.11532090487298678
	pesos_i(2070) := b"0000000000000000_0000000000000000_0001000010001100_1010110001100000"; -- 0.06464650477529217
	pesos_i(2071) := b"1111111111111111_1111111111111111_1111001101000011_1011001011100000"; -- -0.04974824933152517
	pesos_i(2072) := b"1111111111111111_1111111111111111_1101010011001101_1011001100011010"; -- -0.16873627300484814
	pesos_i(2073) := b"0000000000000000_0000000000000000_0010001101011110_0110001001101010"; -- 0.13815894200047843
	pesos_i(2074) := b"1111111111111111_1111111111111111_1111011010001100_1000010000101000"; -- -0.03691839242286105
	pesos_i(2075) := b"1111111111111111_1111111111111111_1110100111011000_0001110100101011"; -- -0.08654611297928042
	pesos_i(2076) := b"0000000000000000_0000000000000000_0001101001010000_1001110110100011"; -- 0.10279259891146508
	pesos_i(2077) := b"0000000000000000_0000000000000000_0010001110100101_1111000100101111"; -- 0.1392508258723814
	pesos_i(2078) := b"0000000000000000_0000000000000000_0000111100111011_1110110001010101"; -- 0.059508105142526135
	pesos_i(2079) := b"1111111111111111_1111111111111111_1110011110010100_1011111001010100"; -- -0.09538660486650867
	pesos_i(2080) := b"0000000000000000_0000000000000000_0000011111010001_1100101011000110"; -- 0.030544923074623642
	pesos_i(2081) := b"0000000000000000_0000000000000000_0010011101001011_1011101010110010"; -- 0.1534992871726246
	pesos_i(2082) := b"0000000000000000_0000000000000000_0000000010011001_1110110111111100"; -- 0.0023487796912701094
	pesos_i(2083) := b"0000000000000000_0000000000000000_0000101100110010_0001100001101010"; -- 0.04373314473443421
	pesos_i(2084) := b"0000000000000000_0000000000000000_0000011010111000_1100001111111110"; -- 0.026256799166647818
	pesos_i(2085) := b"1111111111111111_1111111111111111_1110111000100011_1101110111011100"; -- -0.06976521864060403
	pesos_i(2086) := b"1111111111111111_1111111111111111_1101101000110000_0101011100101111"; -- -0.14769988156299677
	pesos_i(2087) := b"1111111111111111_1111111111111111_1111000001010111_1110110010010110"; -- -0.06115838375705443
	pesos_i(2088) := b"0000000000000000_0000000000000000_0000110100000011_1011001101001111"; -- 0.05083771390046868
	pesos_i(2089) := b"1111111111111111_1111111111111111_1111100010110000_0111100000010111"; -- -0.028557295261208017
	pesos_i(2090) := b"0000000000000000_0000000000000000_0001011111111111_0101010101101010"; -- 0.09373983235017275
	pesos_i(2091) := b"0000000000000000_0000000000000000_0010100011001101_1001101001010000"; -- 0.15938724941072688
	pesos_i(2092) := b"1111111111111111_1111111111111111_1111001100000100_0011100000010011"; -- -0.05071687248935781
	pesos_i(2093) := b"1111111111111111_1111111111111111_1101111100000001_0100000110000101"; -- -0.12888708587881526
	pesos_i(2094) := b"0000000000000000_0000000000000000_0010001011101000_1011011011110010"; -- 0.1363634434870649
	pesos_i(2095) := b"0000000000000000_0000000000000000_0001111000001010_0010111101111101"; -- 0.11734291832376903
	pesos_i(2096) := b"1111111111111111_1111111111111111_1110010111111011_1011010110011101"; -- -0.10162796897904625
	pesos_i(2097) := b"0000000000000000_0000000000000000_0001110001100101_0001110000110111"; -- 0.11091781951252581
	pesos_i(2098) := b"1111111111111111_1111111111111111_1101001100101111_1011010111110001"; -- -0.17505324244771273
	pesos_i(2099) := b"0000000000000000_0000000000000000_0001000010011100_1110001001110110"; -- 0.06489386921552592
	pesos_i(2100) := b"0000000000000000_0000000000000000_0001010100111000_0100100101000011"; -- 0.08289010899369911
	pesos_i(2101) := b"1111111111111111_1111111111111111_1101111111110100_0100001000101110"; -- -0.1251791608655727
	pesos_i(2102) := b"0000000000000000_0000000000000000_0000011010000000_1101010000111110"; -- 0.025403275682876487
	pesos_i(2103) := b"1111111111111111_1111111111111111_1111000111111000_1010011101001110"; -- -0.054799598063621315
	pesos_i(2104) := b"0000000000000000_0000000000000000_0000011010101101_0010001011010010"; -- 0.02607934587622049
	pesos_i(2105) := b"1111111111111111_1111111111111111_1111110110001010_0001010111110010"; -- -0.009611729144448258
	pesos_i(2106) := b"0000000000000000_0000000000000000_0001100110011011_1001111111011011"; -- 0.10003089048003125
	pesos_i(2107) := b"0000000000000000_0000000000000000_0000010110101100_1010100101111001"; -- 0.022165863162147227
	pesos_i(2108) := b"0000000000000000_0000000000000000_0010100110100010_0101100011100000"; -- 0.16263347115190702
	pesos_i(2109) := b"1111111111111111_1111111111111111_1101110110101100_0000100110100100"; -- -0.1340936636186268
	pesos_i(2110) := b"0000000000000000_0000000000000000_0010001010111011_1010100000100011"; -- 0.1356759152878016
	pesos_i(2111) := b"1111111111111111_1111111111111111_1101101100001100_0010010001111111"; -- -0.1443459692885682
	pesos_i(2112) := b"0000000000000000_0000000000000000_0001101001010011_0110000010111110"; -- 0.10283474573450038
	pesos_i(2113) := b"0000000000000000_0000000000000000_0000111101101011_1010101001100100"; -- 0.06023659642730035
	pesos_i(2114) := b"1111111111111111_1111111111111111_1111111010101001_0110000100100100"; -- -0.005227974662522913
	pesos_i(2115) := b"1111111111111111_1111111111111111_1111101010101011_1110101000101000"; -- -0.0208142902115775
	pesos_i(2116) := b"0000000000000000_0000000000000000_0010000101011010_1101111110110101"; -- 0.13029287507698709
	pesos_i(2117) := b"1111111111111111_1111111111111111_1101100100000111_1010001111110000"; -- -0.15222716698807381
	pesos_i(2118) := b"0000000000000000_0000000000000000_0000010000001110_0000010001011000"; -- 0.015838881889797023
	pesos_i(2119) := b"0000000000000000_0000000000000000_0000110010100011_1101001010110111"; -- 0.04937474229942058
	pesos_i(2120) := b"1111111111111111_1111111111111111_1101101111101110_1111011100100111"; -- -0.1408849268440321
	pesos_i(2121) := b"1111111111111111_1111111111111111_1111011000111111_0000001010101001"; -- -0.03810103763618672
	pesos_i(2122) := b"0000000000000000_0000000000000000_0001110100100110_0011101101100110"; -- 0.11386462441453674
	pesos_i(2123) := b"1111111111111111_1111111111111111_1111111000010000_1011011110001101"; -- -0.007557418923614498
	pesos_i(2124) := b"1111111111111111_1111111111111111_1111000011100001_0110010101000011"; -- -0.05906073682468613
	pesos_i(2125) := b"0000000000000000_0000000000000000_0000011110101001_0011011110000101"; -- 0.029925794660346842
	pesos_i(2126) := b"0000000000000000_0000000000000000_0010101010100101_1110110110101010"; -- 0.16659436613737072
	pesos_i(2127) := b"0000000000000000_0000000000000000_0001010010001110_1000010110010010"; -- 0.08029970955380021
	pesos_i(2128) := b"1111111111111111_1111111111111111_1110100111111101_1011001110101001"; -- -0.08597256772146078
	pesos_i(2129) := b"1111111111111111_1111111111111111_1111011101111110_1001100001010000"; -- -0.03322456395020112
	pesos_i(2130) := b"0000000000000000_0000000000000000_0000011111101011_1010110010101100"; -- 0.03093985741817683
	pesos_i(2131) := b"0000000000000000_0000000000000000_0000001111100101_1111111100000000"; -- 0.015228211949553877
	pesos_i(2132) := b"1111111111111111_1111111111111111_1101111010111011_0100101001101000"; -- -0.12995467149694684
	pesos_i(2133) := b"1111111111111111_1111111111111111_1111110101000100_0110011100000111"; -- -0.010675011539998369
	pesos_i(2134) := b"1111111111111111_1111111111111111_1111001111100110_0100110010001111"; -- -0.04726716528264983
	pesos_i(2135) := b"0000000000000000_0000000000000000_0000001010111010_0111000101000011"; -- 0.010657385699267049
	pesos_i(2136) := b"0000000000000000_0000000000000000_0010111110010100_1010010000000100"; -- 0.18586182688674405
	pesos_i(2137) := b"0000000000000000_0000000000000000_0000111110010101_0000100101111000"; -- 0.06086787400969976
	pesos_i(2138) := b"0000000000000000_0000000000000000_0010000100101001_1000101010111010"; -- 0.12954012912261653
	pesos_i(2139) := b"0000000000000000_0000000000000000_0000001101011011_0011010101000000"; -- 0.013110473779611222
	pesos_i(2140) := b"0000000000000000_0000000000000000_0001010110111011_0100000101011000"; -- 0.08488853831514302
	pesos_i(2141) := b"0000000000000000_0000000000000000_0001011001010111_1101101110011100"; -- 0.08727810427651532
	pesos_i(2142) := b"1111111111111111_1111111111111111_1111100010010001_1101100001100101"; -- -0.029024577469646443
	pesos_i(2143) := b"0000000000000000_0000000000000000_0000011010100111_0100100001011011"; -- 0.025990030474924708
	pesos_i(2144) := b"0000000000000000_0000000000000000_0000110111110110_0011110010011101"; -- 0.05453852493125941
	pesos_i(2145) := b"1111111111111111_1111111111111111_1110001000000010_0000010010111000"; -- -0.11715670121425519
	pesos_i(2146) := b"1111111111111111_1111111111111111_1110010000110100_1001111001101011"; -- -0.10857210050683119
	pesos_i(2147) := b"0000000000000000_0000000000000000_0001000000010111_0101110001000001"; -- 0.0628564508177845
	pesos_i(2148) := b"1111111111111111_1111111111111111_1110000101110011_1111100100111111"; -- -0.11932413297342274
	pesos_i(2149) := b"1111111111111111_1111111111111111_1111011111101010_1101000000010000"; -- -0.031573291759887934
	pesos_i(2150) := b"1111111111111111_1111111111111111_1111111000000000_1111101011011100"; -- -0.007797547650203024
	pesos_i(2151) := b"1111111111111111_1111111111111111_1110000011011010_0011011001100100"; -- -0.12167034209048608
	pesos_i(2152) := b"1111111111111111_1111111111111111_1110110001100110_0000100000000000"; -- -0.07656812669513181
	pesos_i(2153) := b"1111111111111111_1111111111111111_1101000000001010_1011010010010011"; -- -0.1873366490036946
	pesos_i(2154) := b"1111111111111111_1111111111111111_1111000110011111_0011000100000111"; -- -0.05616468036542009
	pesos_i(2155) := b"1111111111111111_1111111111111111_1110010010100100_0100010101111111"; -- -0.10686841634778194
	pesos_i(2156) := b"1111111111111111_1111111111111111_1110111101000001_1000001011011011"; -- -0.06540662921475811
	pesos_i(2157) := b"0000000000000000_0000000000000000_0000100001011010_0100100110110010"; -- 0.03262768362391273
	pesos_i(2158) := b"1111111111111111_1111111111111111_1111110000011000_0101111010101111"; -- -0.01525314558293137
	pesos_i(2159) := b"0000000000000000_0000000000000000_0000001111001010_1100011110111101"; -- 0.014812930798054768
	pesos_i(2160) := b"1111111111111111_1111111111111111_1110010000110010_0100001000101010"; -- -0.108608116806836
	pesos_i(2161) := b"1111111111111111_1111111111111111_1111000010010100_0000000110111111"; -- -0.060241595212335616
	pesos_i(2162) := b"0000000000000000_0000000000000000_0010010011111110_0110000101010110"; -- 0.14450653420918097
	pesos_i(2163) := b"1111111111111111_1111111111111111_1110001101101110_0110101111010001"; -- -0.1115963567854876
	pesos_i(2164) := b"0000000000000000_0000000000000000_0001000000011011_1100111110010111"; -- 0.0629243606384586
	pesos_i(2165) := b"1111111111111111_1111111111111111_1111011101000101_0010100011010101"; -- -0.034100959691329036
	pesos_i(2166) := b"1111111111111111_1111111111111111_1111101110000011_0101011100010111"; -- -0.017527157680532705
	pesos_i(2167) := b"1111111111111111_1111111111111111_1101101100011101_1000001110011111"; -- -0.14408089992863382
	pesos_i(2168) := b"1111111111111111_1111111111111111_1101111011100111_0000000001010000"; -- -0.12928770099628384
	pesos_i(2169) := b"1111111111111111_1111111111111111_1110001001001101_1100011011110010"; -- -0.1160007152072679
	pesos_i(2170) := b"1111111111111111_1111111111111111_1101110011100111_1010011010010100"; -- -0.13709029096768727
	pesos_i(2171) := b"1111111111111111_1111111111111111_1111100101011010_0000101001100100"; -- -0.02596983965381081
	pesos_i(2172) := b"1111111111111111_1111111111111111_1101011110110110_0110011000010100"; -- -0.15737306611106577
	pesos_i(2173) := b"1111111111111111_1111111111111111_1101100010110110_0111001011010001"; -- -0.15346605684548728
	pesos_i(2174) := b"1111111111111111_1111111111111111_1111100011110001_1011000111001111"; -- -0.02756203371538738
	pesos_i(2175) := b"0000000000000000_0000000000000000_0000011010000100_0001011100110100"; -- 0.025453043226012335
	pesos_i(2176) := b"1111111111111111_1111111111111111_1111011101100010_0011010110000010"; -- -0.03365769925928622
	pesos_i(2177) := b"1111111111111111_1111111111111111_1101111110011110_0011111001110110"; -- -0.1264916383988321
	pesos_i(2178) := b"0000000000000000_0000000000000000_0000001011010100_1110000010010000"; -- 0.011060748328837364
	pesos_i(2179) := b"0000000000000000_0000000000000000_0010101000110010_1111110011001110"; -- 0.1648405078055516
	pesos_i(2180) := b"1111111111111111_1111111111111111_1101110001100010_0101010110100001"; -- -0.13912453480181272
	pesos_i(2181) := b"0000000000000000_0000000000000000_0000101000110101_1000011101100010"; -- 0.03987928518956163
	pesos_i(2182) := b"0000000000000000_0000000000000000_0000101011000110_1000001000011010"; -- 0.04209149486537079
	pesos_i(2183) := b"1111111111111111_1111111111111111_1111000000010100_1000100111100010"; -- -0.062186605699397345
	pesos_i(2184) := b"0000000000000000_0000000000000000_0001000100010011_1001010001011001"; -- 0.06670500926880293
	pesos_i(2185) := b"0000000000000000_0000000000000000_0010000100101001_0011000100010111"; -- 0.12953478631994705
	pesos_i(2186) := b"0000000000000000_0000000000000000_0000111000100010_1010101110101010"; -- 0.055216530824455046
	pesos_i(2187) := b"1111111111111111_1111111111111111_1101100011011101_0010000100100000"; -- -0.15287583325900592
	pesos_i(2188) := b"1111111111111111_1111111111111111_1100111000010100_1111010100011010"; -- -0.19499271508396482
	pesos_i(2189) := b"1111111111111111_1111111111111111_1101110100001111_0010100010110011"; -- -0.13648744236841784
	pesos_i(2190) := b"1111111111111111_1111111111111111_1101101000011111_1000010001110110"; -- -0.14795658223266941
	pesos_i(2191) := b"0000000000000000_0000000000000000_0010100001011111_0100101101111101"; -- 0.1577040843181504
	pesos_i(2192) := b"1111111111111111_1111111111111111_1101100011011100_0111110011001001"; -- -0.15288562872755626
	pesos_i(2193) := b"0000000000000000_0000000000000000_0010000010011000_0000111101110000"; -- 0.12732025612693604
	pesos_i(2194) := b"1111111111111111_1111111111111111_1101001111101000_0101010010110111"; -- -0.17223616146864681
	pesos_i(2195) := b"0000000000000000_0000000000000000_0001010001111111_0010010000111000"; -- 0.08006502495233914
	pesos_i(2196) := b"0000000000000000_0000000000000000_0000000110111001_0100000111011000"; -- 0.006733050639479783
	pesos_i(2197) := b"0000000000000000_0000000000000000_0000011101111110_1110001000010001"; -- 0.029279831913605843
	pesos_i(2198) := b"1111111111111111_1111111111111111_1111001000100001_1111111110010010"; -- -0.05416872673327706
	pesos_i(2199) := b"0000000000000000_0000000000000000_0001101001100001_0001101001100100"; -- 0.10304417562132116
	pesos_i(2200) := b"1111111111111111_1111111111111111_1110101010110001_1111010100111110"; -- -0.08322207669643727
	pesos_i(2201) := b"1111111111111111_1111111111111111_1110011101101110_1101010001100010"; -- -0.09596512417475393
	pesos_i(2202) := b"0000000000000000_0000000000000000_0001111000000101_0110000011001100"; -- 0.11726956349845924
	pesos_i(2203) := b"1111111111111111_1111111111111111_1111111111101011_0100011111110101"; -- -0.00031614556686876806
	pesos_i(2204) := b"1111111111111111_1111111111111111_1111110010011011_1100011100010010"; -- -0.013248022077443362
	pesos_i(2205) := b"1111111111111111_1111111111111111_1111000000110101_0110100101101010"; -- -0.06168500097467782
	pesos_i(2206) := b"1111111111111111_1111111111111111_1101111110100111_1001011101110110"; -- -0.12634900447667313
	pesos_i(2207) := b"0000000000000000_0000000000000000_0010001000000010_1001111001001001"; -- 0.13285245206736454
	pesos_i(2208) := b"0000000000000000_0000000000000000_0000011101100111_0011111001101001"; -- 0.028919125195579265
	pesos_i(2209) := b"0000000000000000_0000000000000000_0001000000000001_1000100001110011"; -- 0.06252339185649076
	pesos_i(2210) := b"0000000000000000_0000000000000000_0000110010000100_1001101010010100"; -- 0.048898373743832005
	pesos_i(2211) := b"1111111111111111_1111111111111111_1111100111111101_0010010010101010"; -- -0.02348109104066658
	pesos_i(2212) := b"0000000000000000_0000000000000000_0000100011010101_0010111010001011"; -- 0.03450289623810007
	pesos_i(2213) := b"0000000000000000_0000000000000000_0001010101110110_1010001110101000"; -- 0.08384154170605435
	pesos_i(2214) := b"1111111111111111_1111111111111111_1101110001010010_1111011100010111"; -- -0.1393590515699545
	pesos_i(2215) := b"0000000000000000_0000000000000000_0000001100011010_0001001101110010"; -- 0.012116637499582084
	pesos_i(2216) := b"0000000000000000_0000000000000000_0001110100101111_0100111000011000"; -- 0.11400306780608718
	pesos_i(2217) := b"1111111111111111_1111111111111111_1111100011101101_0100011100100111"; -- -0.027629425966574795
	pesos_i(2218) := b"0000000000000000_0000000000000000_0000100010110101_0010000101111100"; -- 0.03401383674160754
	pesos_i(2219) := b"0000000000000000_0000000000000000_0001101101011100_1100000111111010"; -- 0.1068841206028208
	pesos_i(2220) := b"0000000000000000_0000000000000000_0000010101111011_1000100101000110"; -- 0.021416263106121932
	pesos_i(2221) := b"1111111111111111_1111111111111111_1111100001011100_1100011110111011"; -- -0.02983428665175347
	pesos_i(2222) := b"0000000000000000_0000000000000000_0001111101001000_1101101110111011"; -- 0.12220547977993333
	pesos_i(2223) := b"0000000000000000_0000000000000000_0000110011110001_0011001111110010"; -- 0.05055546430232744
	pesos_i(2224) := b"0000000000000000_0000000000000000_0010001010101110_1001110000100101"; -- 0.13547683614609676
	pesos_i(2225) := b"0000000000000000_0000000000000000_0001010111011001_1000111101100011"; -- 0.08535095385158381
	pesos_i(2226) := b"1111111111111111_1111111111111111_1101110110111110_0101110111010010"; -- -0.13381398792995755
	pesos_i(2227) := b"0000000000000000_0000000000000000_0010011000011101_1001001111011100"; -- 0.14888881807383433
	pesos_i(2228) := b"0000000000000000_0000000000000000_0000110011101111_0001110001010011"; -- 0.05052353877157223
	pesos_i(2229) := b"0000000000000000_0000000000000000_0000101010110011_0100011101011011"; -- 0.041798076474055555
	pesos_i(2230) := b"1111111111111111_1111111111111111_1111000000001101_0001110111011101"; -- -0.06229985581567853
	pesos_i(2231) := b"1111111111111111_1111111111111111_1110010000101101_0101000100000111"; -- -0.10868352488541941
	pesos_i(2232) := b"1111111111111111_1111111111111111_1111000110001001_0010001000101001"; -- -0.05650125990584297
	pesos_i(2233) := b"1111111111111111_1111111111111111_1110110010100000_1011101010000011"; -- -0.07567247668195763
	pesos_i(2234) := b"0000000000000000_0000000000000000_0001100100011111_1111010011011110"; -- 0.09814386777550058
	pesos_i(2235) := b"0000000000000000_0000000000000000_0000111000101111_1011010111001000"; -- 0.05541549815550746
	pesos_i(2236) := b"0000000000000000_0000000000000000_0000010001110011_0000101100100001"; -- 0.017380424145026753
	pesos_i(2237) := b"0000000000000000_0000000000000000_0010001111100000_0110100110001010"; -- 0.14014300927521456
	pesos_i(2238) := b"0000000000000000_0000000000000000_0001001111101101_0110110001111000"; -- 0.07784154816975196
	pesos_i(2239) := b"1111111111111111_1111111111111111_1101100101001011_0111101110001101"; -- -0.15119197668683015
	pesos_i(2240) := b"1111111111111111_1111111111111111_1110010010101011_1010000001100101"; -- -0.10675618671184232
	pesos_i(2241) := b"1111111111111111_1111111111111111_1111011111110100_0010000101011111"; -- -0.031431116314261424
	pesos_i(2242) := b"0000000000000000_0000000000000000_0001110011001010_0001110101100000"; -- 0.11245902616986479
	pesos_i(2243) := b"0000000000000000_0000000000000000_0000000110010101_1010000001011110"; -- 0.006189368234019214
	pesos_i(2244) := b"1111111111111111_1111111111111111_1101111100110100_1010101101000110"; -- -0.12810258422104448
	pesos_i(2245) := b"1111111111111111_1111111111111111_1111001100101000_0111001001101011"; -- -0.050164078608087054
	pesos_i(2246) := b"0000000000000000_0000000000000000_0000100110110010_0000011100101100"; -- 0.0378727418737193
	pesos_i(2247) := b"1111111111111111_1111111111111111_1111000001011101_1100000010010001"; -- -0.06106945476484196
	pesos_i(2248) := b"1111111111111111_1111111111111111_1101110101000010_1011100000011111"; -- -0.13570069545918975
	pesos_i(2249) := b"0000000000000000_0000000000000000_0010011001111010_1111011110110101"; -- 0.15031383671895723
	pesos_i(2250) := b"1111111111111111_1111111111111111_1111101111000000_1110100011101011"; -- -0.016587679456325246
	pesos_i(2251) := b"0000000000000000_0000000000000000_0010001000110110_1101011011001111"; -- 0.13364927819762287
	pesos_i(2252) := b"0000000000000000_0000000000000000_0010010010101011_0111001011010000"; -- 0.14324109634783153
	pesos_i(2253) := b"0000000000000000_0000000000000000_0010011100100010_1000011100010100"; -- 0.15287060022249
	pesos_i(2254) := b"0000000000000000_0000000000000000_0001110110110111_0010100001100100"; -- 0.11607601586214131
	pesos_i(2255) := b"0000000000000000_0000000000000000_0001101011110110_0101100010110001"; -- 0.10532144861125171
	pesos_i(2256) := b"0000000000000000_0000000000000000_0010100110011110_0111000010110001"; -- 0.16257385559139056
	pesos_i(2257) := b"0000000000000000_0000000000000000_0010100111010001_1010101011110010"; -- 0.16335552596955288
	pesos_i(2258) := b"1111111111111111_1111111111111111_1111010001010101_1110010011000101"; -- -0.0455643673018638
	pesos_i(2259) := b"0000000000000000_0000000000000000_0000000011001101_0011011110010011"; -- 0.0031313642889132013
	pesos_i(2260) := b"0000000000000000_0000000000000000_0000111101001101_1000010110000111"; -- 0.0597766356382305
	pesos_i(2261) := b"1111111111111111_1111111111111111_1111010000100111_0000011101111111"; -- -0.046279460496375956
	pesos_i(2262) := b"1111111111111111_1111111111111111_1111101010011001_1010110100100110"; -- -0.02109258486370364
	pesos_i(2263) := b"1111111111111111_1111111111111111_1110010110010011_0110100101011010"; -- -0.10321942855208484
	pesos_i(2264) := b"1111111111111111_1111111111111111_1111010011111001_1011001000001000"; -- -0.043064950102288606
	pesos_i(2265) := b"0000000000000000_0000000000000000_0001011100000011_1100001100110000"; -- 0.08990116044745612
	pesos_i(2266) := b"1111111111111111_1111111111111111_1111110010100001_0001110111111110"; -- -0.013166547262885587
	pesos_i(2267) := b"1111111111111111_1111111111111111_1110001110010101_0101101111000011"; -- -0.11100222098822607
	pesos_i(2268) := b"1111111111111111_1111111111111111_1111001000001010_0110101010000110"; -- -0.05452856279413938
	pesos_i(2269) := b"1111111111111111_1111111111111111_1110110011010100_0011011010011011"; -- -0.07488688194335867
	pesos_i(2270) := b"0000000000000000_0000000000000000_0000010101111001_1011100111001010"; -- 0.021388637308533562
	pesos_i(2271) := b"1111111111111111_1111111111111111_1101011111011100_1001100111111001"; -- -0.15679013893424323
	pesos_i(2272) := b"0000000000000000_0000000000000000_0001111100110001_1011101011001011"; -- 0.12185256445004441
	pesos_i(2273) := b"1111111111111111_1111111111111111_1111110000100001_1100100110010001"; -- -0.015109445596480857
	pesos_i(2274) := b"1111111111111111_1111111111111111_1110011010011111_0010001001101000"; -- -0.09913430177182127
	pesos_i(2275) := b"0000000000000000_0000000000000000_0010110101001001_0110111100000100"; -- 0.1769017587233738
	pesos_i(2276) := b"0000000000000000_0000000000000000_0001000011110010_1101101000111111"; -- 0.06620563539188518
	pesos_i(2277) := b"0000000000000000_0000000000000000_0000101010111010_1011010110110011"; -- 0.04191146497872821
	pesos_i(2278) := b"0000000000000000_0000000000000000_0000010110111110_0010100101110110"; -- 0.022432891073266202
	pesos_i(2279) := b"1111111111111111_1111111111111111_1111000010101000_1010100110110001"; -- -0.0599264089766373
	pesos_i(2280) := b"0000000000000000_0000000000000000_0000101000000010_1010011011101110"; -- 0.03910296743331085
	pesos_i(2281) := b"1111111111111111_1111111111111111_1101111101000001_0001011110111011"; -- -0.12791301419009332
	pesos_i(2282) := b"0000000000000000_0000000000000000_0010100101101000_1001001111001101"; -- 0.1617519736070923
	pesos_i(2283) := b"1111111111111111_1111111111111111_1110110111011111_0110010111100000"; -- -0.07080996784687672
	pesos_i(2284) := b"1111111111111111_1111111111111111_1111010110010010_1101010101110000"; -- -0.040728244987489684
	pesos_i(2285) := b"1111111111111111_1111111111111111_1111100110000100_0100000011100110"; -- -0.02532572155471062
	pesos_i(2286) := b"1111111111111111_1111111111111111_1110100011100100_0000011000010110"; -- -0.09027063339911393
	pesos_i(2287) := b"0000000000000000_0000000000000000_0001111101101110_1101110010101010"; -- 0.12278536934055537
	pesos_i(2288) := b"0000000000000000_0000000000000000_0000101000010001_1111011011100011"; -- 0.039336614981157814
	pesos_i(2289) := b"0000000000000000_0000000000000000_0010100011110011_1001100010010011"; -- 0.15996697986193936
	pesos_i(2290) := b"0000000000000000_0000000000000000_0001001000000100_1111101111001011"; -- 0.07038854328371794
	pesos_i(2291) := b"0000000000000000_0000000000000000_0001110001100001_1001000001010110"; -- 0.11086370568485063
	pesos_i(2292) := b"1111111111111111_1111111111111111_1110001111110010_0011110101100111"; -- -0.10958496314972682
	pesos_i(2293) := b"1111111111111111_1111111111111111_1110001000001100_0001001011101011"; -- -0.1170032668651334
	pesos_i(2294) := b"0000000000000000_0000000000000000_0000100100000100_1101000010001000"; -- 0.035229714516474796
	pesos_i(2295) := b"0000000000000000_0000000000000000_0001010101010110_1111011110001100"; -- 0.0833582608685116
	pesos_i(2296) := b"0000000000000000_0000000000000000_0000101101111110_0111001110100110"; -- 0.044898250611748014
	pesos_i(2297) := b"0000000000000000_0000000000000000_0001010001010001_0000111010001110"; -- 0.07936182951933689
	pesos_i(2298) := b"0000000000000000_0000000000000000_0010011011001011_0111000110001111"; -- 0.1515418028041764
	pesos_i(2299) := b"1111111111111111_1111111111111111_1110011000111101_1110010100001011"; -- -0.1006180619209773
	pesos_i(2300) := b"1111111111111111_1111111111111111_1101011001101011_0100100010110110"; -- -0.1624254756644745
	pesos_i(2301) := b"0000000000000000_0000000000000000_0010000100000000_1110001101100110"; -- 0.12891980389396746
	pesos_i(2302) := b"0000000000000000_0000000000000000_0000000001001001_0100011010000100"; -- 0.0011180946006764114
	pesos_i(2303) := b"0000000000000000_0000000000000000_0001001011001110_1111010110011010"; -- 0.07347044965203751
	pesos_i(2304) := b"1111111111111111_1111111111111111_1110100011100100_0111111000110111"; -- -0.09026347300785574
	pesos_i(2305) := b"0000000000000000_0000000000000000_0000101011100010_1001101001000011"; -- 0.0425201811040926
	pesos_i(2306) := b"0000000000000000_0000000000000000_0010010100011001_1110001001110110"; -- 0.14492621785308651
	pesos_i(2307) := b"1111111111111111_1111111111111111_1101111110011011_1111011110101011"; -- -0.12652637556281288
	pesos_i(2308) := b"0000000000000000_0000000000000000_0000111101110011_1101010001001101"; -- 0.060361164832355436
	pesos_i(2309) := b"0000000000000000_0000000000000000_0001011010000000_0111000011001011"; -- 0.08789734792218924
	pesos_i(2310) := b"0000000000000000_0000000000000000_0000110111011100_0110100110001110"; -- 0.05414447505295451
	pesos_i(2311) := b"1111111111111111_1111111111111111_1111011111100101_0100000000001110"; -- -0.03165816925857021
	pesos_i(2312) := b"1111111111111111_1111111111111111_1111000000110111_1111100011010111"; -- -0.0616459345647633
	pesos_i(2313) := b"1111111111111111_1111111111111111_1101100001001100_0111110001110100"; -- -0.1550829140529897
	pesos_i(2314) := b"0000000000000000_0000000000000000_0010001111100011_0110000111111111"; -- 0.14018833608763934
	pesos_i(2315) := b"0000000000000000_0000000000000000_0000001101010011_0101011011000111"; -- 0.012990401766572028
	pesos_i(2316) := b"1111111111111111_1111111111111111_1110110111011110_1011011101111111"; -- -0.07082036150584292
	pesos_i(2317) := b"0000000000000000_0000000000000000_0000110110111011_0001011100100111"; -- 0.05363602345222458
	pesos_i(2318) := b"1111111111111111_1111111111111111_1101110010100110_1101000100000111"; -- -0.1380795819202567
	pesos_i(2319) := b"0000000000000000_0000000000000000_0010001111000111_0011001100010100"; -- 0.1397582934027241
	pesos_i(2320) := b"1111111111111111_1111111111111111_1111011011010000_0000111111011110"; -- -0.03588772602543955
	pesos_i(2321) := b"1111111111111111_1111111111111111_1111110110101111_1111101100000000"; -- -0.009033501129999696
	pesos_i(2322) := b"1111111111111111_1111111111111111_1110111001001111_1011011111000010"; -- -0.06909610282936637
	pesos_i(2323) := b"1111111111111111_1111111111111111_1111000111011101_0111010001011111"; -- -0.05521462133363295
	pesos_i(2324) := b"0000000000000000_0000000000000000_0001011110110000_1000100101010100"; -- 0.09253748224162044
	pesos_i(2325) := b"0000000000000000_0000000000000000_0001100000111111_1001000101101011"; -- 0.09471997139047393
	pesos_i(2326) := b"0000000000000000_0000000000000000_0001100000000001_1100001010101101"; -- 0.09377686237379301
	pesos_i(2327) := b"1111111111111111_1111111111111111_1101101101100100_1110110101111000"; -- -0.14299121680046054
	pesos_i(2328) := b"1111111111111111_1111111111111111_1110001001010001_0111011110111101"; -- -0.11594440105142474
	pesos_i(2329) := b"0000000000000000_0000000000000000_0001001010001010_0000110011010011"; -- 0.07241897733824178
	pesos_i(2330) := b"1111111111111111_1111111111111111_1110000101111010_0100010001000010"; -- -0.11922810924544257
	pesos_i(2331) := b"0000000000000000_0000000000000000_0010001010100100_1110100011101101"; -- 0.1353288248765596
	pesos_i(2332) := b"0000000000000000_0000000000000000_0000100100111101_0111001101011100"; -- 0.0360939121879765
	pesos_i(2333) := b"0000000000000000_0000000000000000_0001011101010110_0001010011000011"; -- 0.09115724342680177
	pesos_i(2334) := b"0000000000000000_0000000000000000_0000011001100010_1111010101111000"; -- 0.024947492345985933
	pesos_i(2335) := b"0000000000000000_0000000000000000_0010001000011111_1010111001011001"; -- 0.1332959142895014
	pesos_i(2336) := b"1111111111111111_1111111111111111_1101110111001011_0011001100101011"; -- -0.13361816592033607
	pesos_i(2337) := b"1111111111111111_1111111111111111_1110111001111100_1110000001001010"; -- -0.06840704156293893
	pesos_i(2338) := b"0000000000000000_0000000000000000_0010001011111101_0110011101101101"; -- 0.1366791383179454
	pesos_i(2339) := b"1111111111111111_1111111111111111_1110100010100111_0010000000110101"; -- -0.09119986248549618
	pesos_i(2340) := b"0000000000000000_0000000000000000_0001011000101000_1011010101110000"; -- 0.08655866613940431
	pesos_i(2341) := b"0000000000000000_0000000000000000_0000001010001001_0110111110000110"; -- 0.009909601409799986
	pesos_i(2342) := b"1111111111111111_1111111111111111_1110001001001110_1011111100001010"; -- -0.11598592757031786
	pesos_i(2343) := b"0000000000000000_0000000000000000_0001111001010001_0100110010100101"; -- 0.11842803039194902
	pesos_i(2344) := b"0000000000000000_0000000000000000_0001000010101100_1010111101010101"; -- 0.06513496223395007
	pesos_i(2345) := b"1111111111111111_1111111111111111_1101110001100010_1100101000001110"; -- -0.1391175953468415
	pesos_i(2346) := b"1111111111111111_1111111111111111_1111111110100010_0001011110101011"; -- -0.001432915500067466
	pesos_i(2347) := b"0000000000000000_0000000000000000_0001111011100000_1110111110101000"; -- 0.12061975348906918
	pesos_i(2348) := b"1111111111111111_1111111111111111_1101011010000011_0100111000000100"; -- -0.16205894848144853
	pesos_i(2349) := b"1111111111111111_1111111111111111_1101011110000101_0010101110000010"; -- -0.1581242378081672
	pesos_i(2350) := b"1111111111111111_1111111111111111_1101010000100011_0010111100110011"; -- -0.17133812902286738
	pesos_i(2351) := b"0000000000000000_0000000000000000_0000111101111011_0111111011101010"; -- 0.06047814576974223
	pesos_i(2352) := b"1111111111111111_1111111111111111_1101101011001000_1101000101110011"; -- -0.14537325795546557
	pesos_i(2353) := b"0000000000000000_0000000000000000_0010000101100010_1101110101110000"; -- 0.13041480997557695
	pesos_i(2354) := b"0000000000000000_0000000000000000_0001000010111000_1000110010100000"; -- 0.06531599916269301
	pesos_i(2355) := b"0000000000000000_0000000000000000_0000011011001101_0010000001111010"; -- 0.026567487523363853
	pesos_i(2356) := b"0000000000000000_0000000000000000_0010010100101010_1011000110000101"; -- 0.1451827000411632
	pesos_i(2357) := b"1111111111111111_1111111111111111_1111101001100001_0110100000000110"; -- -0.02195119728932479
	pesos_i(2358) := b"0000000000000000_0000000000000000_0010000011010000_0110101110000011"; -- 0.12818023641962123
	pesos_i(2359) := b"0000000000000000_0000000000000000_0001101101011010_0000111100100110"; -- 0.1068429439619297
	pesos_i(2360) := b"1111111111111111_1111111111111111_1110010101010000_1001111001100101"; -- -0.10423860589887149
	pesos_i(2361) := b"1111111111111111_1111111111111111_1110011000010111_0001110110011000"; -- -0.10120978381291804
	pesos_i(2362) := b"0000000000000000_0000000000000000_0001001000000101_0111110001001001"; -- 0.07039620197024216
	pesos_i(2363) := b"1111111111111111_1111111111111111_1111101110101001_0110101010101010"; -- -0.016946156881982873
	pesos_i(2364) := b"1111111111111111_1111111111111111_1110100011110011_0101000010101011"; -- -0.09003730614404722
	pesos_i(2365) := b"0000000000000000_0000000000000000_0001111111100101_1100000111010110"; -- 0.12459956620173131
	pesos_i(2366) := b"0000000000000000_0000000000000000_0001011101011100_1000011110011010"; -- 0.09125564098699364
	pesos_i(2367) := b"1111111111111111_1111111111111111_1111010010101001_1101101011000100"; -- -0.04428322512275106
	pesos_i(2368) := b"1111111111111111_1111111111111111_1111110000101101_1110101111000000"; -- -0.014924302613048335
	pesos_i(2369) := b"0000000000000000_0000000000000000_0001000101000111_1000100101100001"; -- 0.0674978123848221
	pesos_i(2370) := b"1111111111111111_1111111111111111_1111110100011011_0010110011001010"; -- -0.011304092971406665
	pesos_i(2371) := b"1111111111111111_1111111111111111_1111011001010111_1011111011010100"; -- -0.03772361110967663
	pesos_i(2372) := b"0000000000000000_0000000000000000_0000101110100011_0001110001100001"; -- 0.04545762415307839
	pesos_i(2373) := b"0000000000000000_0000000000000000_0010001000011001_0100011010011100"; -- 0.1331981782858722
	pesos_i(2374) := b"1111111111111111_1111111111111111_1111101110111010_1011101011000001"; -- -0.016681983884718064
	pesos_i(2375) := b"0000000000000000_0000000000000000_0000101110000010_0001110011110101"; -- 0.04495411844122509
	pesos_i(2376) := b"0000000000000000_0000000000000000_0001000111011111_1110010010011111"; -- 0.0698225868892641
	pesos_i(2377) := b"0000000000000000_0000000000000000_0000010111101101_0111010001111111"; -- 0.02315452666317336
	pesos_i(2378) := b"1111111111111111_1111111111111111_1110100010100001_1111110010001111"; -- -0.09127828138897931
	pesos_i(2379) := b"0000000000000000_0000000000000000_0010100100011110_0110001010100000"; -- 0.16061989217391476
	pesos_i(2380) := b"0000000000000000_0000000000000000_0010011010100011_0110111011111011"; -- 0.15093129749268713
	pesos_i(2381) := b"1111111111111111_1111111111111111_1110111001110100_1000101100000111"; -- -0.06853419389940264
	pesos_i(2382) := b"0000000000000000_0000000000000000_0001001110011110_1011011100011111"; -- 0.07664055364482879
	pesos_i(2383) := b"1111111111111111_1111111111111111_1111010111011100_0111100010000000"; -- -0.039604633967551435
	pesos_i(2384) := b"0000000000000000_0000000000000000_0000101111001011_1001010110011010"; -- 0.04607520113177416
	pesos_i(2385) := b"0000000000000000_0000000000000000_0001100110111001_0101100000101001"; -- 0.1004843806732334
	pesos_i(2386) := b"0000000000000000_0000000000000000_0000011000011000_0110100001000001"; -- 0.02380992501003587
	pesos_i(2387) := b"0000000000000000_0000000000000000_0000001100111010_0000000010010110"; -- 0.012603794789769486
	pesos_i(2388) := b"0000000000000000_0000000000000000_0010100101110011_0000110010000001"; -- 0.1619117561481104
	pesos_i(2389) := b"0000000000000000_0000000000000000_0010011111100111_1010001010000100"; -- 0.15587821700768778
	pesos_i(2390) := b"0000000000000000_0000000000000000_0001011001110001_1101101001010100"; -- 0.08767475658335618
	pesos_i(2391) := b"1111111111111111_1111111111111111_1111101110100101_0001001011011010"; -- -0.0170124262444615
	pesos_i(2392) := b"0000000000000000_0000000000000000_0001101011011000_1010001000111100"; -- 0.10486806830264848
	pesos_i(2393) := b"0000000000000000_0000000000000000_0001001110010111_1011000110001010"; -- 0.07653340923680012
	pesos_i(2394) := b"1111111111111111_1111111111111111_1111000011100111_1101100101111111"; -- -0.058962255948379824
	pesos_i(2395) := b"0000000000000000_0000000000000000_0001100100000001_1011010100010100"; -- 0.09768230197010502
	pesos_i(2396) := b"1111111111111111_1111111111111111_1110010010001001_1101101111111010"; -- -0.10727143438377791
	pesos_i(2397) := b"0000000000000000_0000000000000000_0010001111111011_1100001111011101"; -- 0.14056038046217428
	pesos_i(2398) := b"1111111111111111_1111111111111111_1111111011111100_0101101111010110"; -- -0.003961811328204062
	pesos_i(2399) := b"0000000000000000_0000000000000000_0000111111100000_1000010010001000"; -- 0.0620196182860909
	pesos_i(2400) := b"1111111111111111_1111111111111111_1111001010001000_0011000101000000"; -- -0.052609369061281025
	pesos_i(2401) := b"0000000000000000_0000000000000000_0000101111110101_1111101111101111"; -- 0.04672216970884489
	pesos_i(2402) := b"0000000000000000_0000000000000000_0000001110101011_1101111101100101"; -- 0.014341318321299467
	pesos_i(2403) := b"0000000000000000_0000000000000000_0000010011111101_1110000000000100"; -- 0.01949882606473052
	pesos_i(2404) := b"0000000000000000_0000000000000000_0000001000101010_1111011000100010"; -- 0.008468039804325238
	pesos_i(2405) := b"1111111111111111_1111111111111111_1110011000000111_1100100100110010"; -- -0.10144369622214891
	pesos_i(2406) := b"0000000000000000_0000000000000000_0001100110000010_1010101011010100"; -- 0.09965007470081898
	pesos_i(2407) := b"0000000000000000_0000000000000000_0000011011010011_0000110011110011"; -- 0.026657876386475043
	pesos_i(2408) := b"1111111111111111_1111111111111111_1101010110000101_0101111111101100"; -- -0.16593361370652557
	pesos_i(2409) := b"0000000000000000_0000000000000000_0001000010110110_0100000110101100"; -- 0.06528101385817674
	pesos_i(2410) := b"0000000000000000_0000000000000000_0001010001010000_1010100101001010"; -- 0.07935579361781166
	pesos_i(2411) := b"1111111111111111_1111111111111111_1111101111010111_1111100100000010"; -- -0.016235768376706056
	pesos_i(2412) := b"0000000000000000_0000000000000000_0000101000100110_0110001111111101"; -- 0.039648293843676526
	pesos_i(2413) := b"0000000000000000_0000000000000000_0001000101101111_1001111001011001"; -- 0.06810941391710916
	pesos_i(2414) := b"0000000000000000_0000000000000000_0010011010111010_1101101111000110"; -- 0.15128873424005496
	pesos_i(2415) := b"1111111111111111_1111111111111111_1110011011110110_1011011011000111"; -- -0.09779794356723297
	pesos_i(2416) := b"1111111111111111_1111111111111111_1110101000101111_1101011111000010"; -- -0.0852074766730872
	pesos_i(2417) := b"1111111111111111_1111111111111111_1111111101001010_1011000000111011"; -- -0.0027665953868315084
	pesos_i(2418) := b"0000000000000000_0000000000000000_0010100111100110_0001110111010010"; -- 0.16366754901977862
	pesos_i(2419) := b"0000000000000000_0000000000000000_0001010000110101_1010100101011110"; -- 0.07894381099719293
	pesos_i(2420) := b"0000000000000000_0000000000000000_0001001110110000_0111010110000001"; -- 0.0769113006687931
	pesos_i(2421) := b"1111111111111111_1111111111111111_1111000100111001_0111110100001100"; -- -0.05771654573181137
	pesos_i(2422) := b"1111111111111111_1111111111111111_1110010100111000_0101000110010011"; -- -0.10460939555318581
	pesos_i(2423) := b"0000000000000000_0000000000000000_0001100000101001_0010100110100100"; -- 0.0943780922611759
	pesos_i(2424) := b"1111111111111111_1111111111111111_1110101111011110_0000111000010001"; -- -0.07864296050118547
	pesos_i(2425) := b"0000000000000000_0000000000000000_0010100111001100_0010001100001110"; -- 0.16327113235171042
	pesos_i(2426) := b"1111111111111111_1111111111111111_1101101111110110_1001000101111011"; -- -0.14076891649339443
	pesos_i(2427) := b"0000000000000000_0000000000000000_0010000000110110_0101001101111110"; -- 0.1258289510847107
	pesos_i(2428) := b"1111111111111111_1111111111111111_1101101110000000_1001100110000110"; -- -0.14256897431871168
	pesos_i(2429) := b"0000000000000000_0000000000000000_0000110010110000_1010011010011011"; -- 0.049570477339498424
	pesos_i(2430) := b"1111111111111111_1111111111111111_1111000011111010_1000110010010011"; -- -0.05867692375412119
	pesos_i(2431) := b"0000000000000000_0000000000000000_0000100111110111_0011111010100000"; -- 0.03892890375048988
	pesos_i(2432) := b"0000000000000000_0000000000000000_0001011000011110_1111001011100010"; -- 0.08640974058170811
	pesos_i(2433) := b"0000000000000000_0000000000000000_0001101110111001_0010110001111111"; -- 0.1082942780462266
	pesos_i(2434) := b"1111111111111111_1111111111111111_1101101011110100_1010110110101111"; -- -0.14470400302989242
	pesos_i(2435) := b"0000000000000000_0000000000000000_0000110110011101_1111100110010110"; -- 0.05319175639683956
	pesos_i(2436) := b"1111111111111111_1111111111111111_1110010000001010_1011111101011100"; -- -0.1092110060872152
	pesos_i(2437) := b"0000000000000000_0000000000000000_0000111110000000_0000100011000011"; -- 0.06054739735085173
	pesos_i(2438) := b"0000000000000000_0000000000000000_0010011100100101_0110111100011001"; -- 0.15291494709562564
	pesos_i(2439) := b"1111111111111111_1111111111111111_1111000100010111_1111010001111011"; -- -0.058228225769505565
	pesos_i(2440) := b"0000000000000000_0000000000000000_0011010111011010_1000001110000010"; -- 0.2103655044129282
	pesos_i(2441) := b"1111111111111111_1111111111111111_1110000110011000_1111111011101000"; -- -0.11875922053915307
	pesos_i(2442) := b"1111111111111111_1111111111111111_1111011010011000_0110111101110000"; -- -0.03673652192066379
	pesos_i(2443) := b"0000000000000000_0000000000000000_0001000000110100_1011001010010101"; -- 0.06330410143662027
	pesos_i(2444) := b"0000000000000000_0000000000000000_0001000000110011_0011010010011000"; -- 0.06328133310820525
	pesos_i(2445) := b"0000000000000000_0000000000000000_0001100001101000_1000000011011110"; -- 0.09534459513168167
	pesos_i(2446) := b"0000000000000000_0000000000000000_0000001111001001_0010011011010001"; -- 0.014788080135688532
	pesos_i(2447) := b"0000000000000000_0000000000000000_0000000100110010_1011010001111001"; -- 0.004679946362217294
	pesos_i(2448) := b"1111111111111111_1111111111111111_1110100111001001_0111111100001000"; -- -0.08676916174654709
	pesos_i(2449) := b"0000000000000000_0000000000000000_0010011111101000_1111101111111010"; -- 0.15589880805153702
	pesos_i(2450) := b"0000000000000000_0000000000000000_0001100001010000_0000100010011110"; -- 0.09497121674880542
	pesos_i(2451) := b"0000000000000000_0000000000000000_0001110100001100_1000011101001010"; -- 0.11347241938792263
	pesos_i(2452) := b"0000000000000000_0000000000000000_0001010100010011_0110111111100110"; -- 0.08232783667726398
	pesos_i(2453) := b"1111111111111111_1111111111111111_1110111011000110_1001001101110011"; -- -0.06728247102561448
	pesos_i(2454) := b"0000000000000000_0000000000000000_0000000110100101_0000000111100011"; -- 0.006424062741350294
	pesos_i(2455) := b"1111111111111111_1111111111111111_1101111111111001_1010001101000111"; -- -0.12509707945273418
	pesos_i(2456) := b"0000000000000000_0000000000000000_0001110001100101_0100111100010000"; -- 0.11092085016988129
	pesos_i(2457) := b"0000000000000000_0000000000000000_0001110100001000_0000001000010101"; -- 0.11340344439275192
	pesos_i(2458) := b"1111111111111111_1111111111111111_1110101010100001_1110110001010101"; -- -0.08346674856452019
	pesos_i(2459) := b"0000000000000000_0000000000000000_0000110100110100_0111100100001111"; -- 0.05158192267868992
	pesos_i(2460) := b"0000000000000000_0000000000000000_0000001100011101_1100111101000110"; -- 0.01217360924482657
	pesos_i(2461) := b"1111111111111111_1111111111111111_1110110000110011_1111110101000101"; -- -0.07733170576434943
	pesos_i(2462) := b"0000000000000000_0000000000000000_0010010010000100_0101100111011111"; -- 0.14264451693717167
	pesos_i(2463) := b"1111111111111111_1111111111111111_1111111000111001_1100110001001001"; -- -0.00693057269433045
	pesos_i(2464) := b"0000000000000000_0000000000000000_0000010001001110_1100010101101111"; -- 0.016826953405915834
	pesos_i(2465) := b"0000000000000000_0000000000000000_0001010011101010_1001101010000110"; -- 0.08170476692313534
	pesos_i(2466) := b"1111111111111111_1111111111111111_1110011001011101_1101001100011001"; -- -0.10013085033137538
	pesos_i(2467) := b"0000000000000000_0000000000000000_0001000100111011_0001010010100101"; -- 0.06730774904465955
	pesos_i(2468) := b"0000000000000000_0000000000000000_0010000011011000_1101011000101110"; -- 0.12830866449675873
	pesos_i(2469) := b"1111111111111111_1111111111111111_1101110100011011_0011101101110111"; -- -0.136303218264186
	pesos_i(2470) := b"1111111111111111_1111111111111111_1101001001110010_1001000110011010"; -- -0.17793931946402008
	pesos_i(2471) := b"1111111111111111_1111111111111111_1111000100100011_0111101100000010"; -- -0.05805236043553666
	pesos_i(2472) := b"1111111111111111_1111111111111111_1111000110101101_0100011100010100"; -- -0.05594974279685459
	pesos_i(2473) := b"1111111111111111_1111111111111111_1110111000110100_0111111001101101"; -- -0.06951150733927908
	pesos_i(2474) := b"0000000000000000_0000000000000000_0000010011101100_1111001001101100"; -- 0.019240523731193622
	pesos_i(2475) := b"1111111111111111_1111111111111111_1110111110001011_0101010001010010"; -- -0.06428025240335943
	pesos_i(2476) := b"0000000000000000_0000000000000000_0000111011010101_0011000000110001"; -- 0.057940494462674165
	pesos_i(2477) := b"1111111111111111_1111111111111111_1101111001100001_0110111110111000"; -- -0.1313257385561056
	pesos_i(2478) := b"0000000000000000_0000000000000000_0001011000110100_0111110011010111"; -- 0.08673839807106394
	pesos_i(2479) := b"1111111111111111_1111111111111111_1100101101001111_1101100010010000"; -- -0.20581289757911045
	pesos_i(2480) := b"1111111111111111_1111111111111111_1101101101011011_0111010011000110"; -- -0.14313573985017078
	pesos_i(2481) := b"1111111111111111_1111111111111111_1101100001011111_0010001110011100"; -- -0.15479829262205239
	pesos_i(2482) := b"1111111111111111_1111111111111111_1111011111001111_1000000100100011"; -- -0.03198998349648388
	pesos_i(2483) := b"1111111111111111_1111111111111111_1110101111100110_0111101111111001"; -- -0.07851433914279438
	pesos_i(2484) := b"0000000000000000_0000000000000000_0000100101001001_0100011111100110"; -- 0.036274427145006664
	pesos_i(2485) := b"1111111111111111_1111111111111111_1111010001010100_0111011111110110"; -- -0.04558611157431835
	pesos_i(2486) := b"0000000000000000_0000000000000000_0010101101100100_0011000011000110"; -- 0.16949753607322907
	pesos_i(2487) := b"0000000000000000_0000000000000000_0001101011110111_1001111100010010"; -- 0.10534090224181786
	pesos_i(2488) := b"1111111111111111_1111111111111111_1110111010101100_0011001101101001"; -- -0.06768492392965943
	pesos_i(2489) := b"1111111111111111_1111111111111111_1110000000011011_1011101011101101"; -- -0.12457687110543705
	pesos_i(2490) := b"1111111111111111_1111111111111111_1111101101110101_0110111000000011"; -- -0.01773941456265938
	pesos_i(2491) := b"0000000000000000_0000000000000000_0001000010101011_1000011100110011"; -- 0.06511731154331381
	pesos_i(2492) := b"1111111111111111_1111111111111111_1101100000010100_0011011010100101"; -- -0.1559415671396384
	pesos_i(2493) := b"1111111111111111_1111111111111111_1111001101011101_0101101101110000"; -- -0.0493567325947901
	pesos_i(2494) := b"1111111111111111_1111111111111111_1110101100100110_1101100011000100"; -- -0.08143849578093232
	pesos_i(2495) := b"1111111111111111_1111111111111111_1110010110001011_1101000001011010"; -- -0.10333535956933022
	pesos_i(2496) := b"1111111111111111_1111111111111111_1101101001011101_0010011010101111"; -- -0.14701612681409204
	pesos_i(2497) := b"1111111111111111_1111111111111111_1111000011000101_1110001010110001"; -- -0.05948050661948582
	pesos_i(2498) := b"0000000000000000_0000000000000000_0010101010010101_1110101110100010"; -- 0.16635010433079728
	pesos_i(2499) := b"1111111111111111_1111111111111111_1111100001111001_0011010110010110"; -- -0.029400492471202935
	pesos_i(2500) := b"1111111111111111_1111111111111111_1111111110101101_1101110000000000"; -- -0.0012533663749924005
	pesos_i(2501) := b"0000000000000000_0000000000000000_0000111111110010_1100010100111111"; -- 0.06229813362467926
	pesos_i(2502) := b"0000000000000000_0000000000000000_0000000010101011_1110100110010001"; -- 0.002623174468634587
	pesos_i(2503) := b"1111111111111111_1111111111111111_1110001001010010_1100101010001100"; -- -0.11592420654565873
	pesos_i(2504) := b"1111111111111111_1111111111111111_1101011011011100_1001001011101011"; -- -0.16069680942406275
	pesos_i(2505) := b"1111111111111111_1111111111111111_1110001111101101_1111001101010101"; -- -0.10965041323442895
	pesos_i(2506) := b"1111111111111111_1111111111111111_1111010000011111_0100000100000000"; -- -0.0463981031967143
	pesos_i(2507) := b"1111111111111111_1111111111111111_1111110101111111_1110010101010000"; -- -0.009767215763244437
	pesos_i(2508) := b"1111111111111111_1111111111111111_1110011001111101_0010001100100011"; -- -0.09965305710868537
	pesos_i(2509) := b"1111111111111111_1111111111111111_1110000010010010_1111011100000011"; -- -0.12275749366674972
	pesos_i(2510) := b"0000000000000000_0000000000000000_0001001001011001_1000001110011001"; -- 0.07167837616013113
	pesos_i(2511) := b"1111111111111111_1111111111111111_1111100010110101_0101011101001010"; -- -0.02848295641693359
	pesos_i(2512) := b"0000000000000000_0000000000000000_0010000000100101_0000011111101111"; -- 0.12556504806514565
	pesos_i(2513) := b"1111111111111111_1111111111111111_1110010011100011_0000010010111100"; -- -0.1059109727636675
	pesos_i(2514) := b"1111111111111111_1111111111111111_1110001000111110_0100101001101100"; -- -0.1162370190883691
	pesos_i(2515) := b"0000000000000000_0000000000000000_0001001110010000_0010010100100100"; -- 0.07641822934668473
	pesos_i(2516) := b"0000000000000000_0000000000000000_0001011100100011_1011110000011001"; -- 0.09038901901471644
	pesos_i(2517) := b"0000000000000000_0000000000000000_0010010010110111_1100110000111110"; -- 0.14342953210750511
	pesos_i(2518) := b"0000000000000000_0000000000000000_0000101000000010_0100001111001110"; -- 0.03909705901577192
	pesos_i(2519) := b"0000000000000000_0000000000000000_0010011011111101_1001011100001011"; -- 0.1523069765047831
	pesos_i(2520) := b"0000000000000000_0000000000000000_0000100001010010_1000110001010101"; -- 0.03250958524045785
	pesos_i(2521) := b"1111111111111111_1111111111111111_1101101010001110_0111001100111010"; -- -0.14626388394271497
	pesos_i(2522) := b"1111111111111111_1111111111111111_1111110010100011_1011011100000010"; -- -0.013126909179211055
	pesos_i(2523) := b"0000000000000000_0000000000000000_0001000000000011_0100001101110101"; -- 0.06254979722952937
	pesos_i(2524) := b"0000000000000000_0000000000000000_0000100101001010_1010010110101000"; -- 0.03629527420647516
	pesos_i(2525) := b"0000000000000000_0000000000000000_0000100100101101_1000001010101011"; -- 0.03585068390171331
	pesos_i(2526) := b"1111111111111111_1111111111111111_1111111010000100_0111101111010101"; -- -0.005790958802879203
	pesos_i(2527) := b"0000000000000000_0000000000000000_0001011011111111_1010010110111101"; -- 0.08983836995412423
	pesos_i(2528) := b"0000000000000000_0000000000000000_0000110101010110_1000111000111110"; -- 0.05210198419090087
	pesos_i(2529) := b"0000000000000000_0000000000000000_0000111100001110_1100110101100011"; -- 0.05881961506344331
	pesos_i(2530) := b"0000000000000000_0000000000000000_0001101001101111_0111110010000000"; -- 0.10326364643885548
	pesos_i(2531) := b"1111111111111111_1111111111111111_1101111100000110_1000011001100100"; -- -0.12880668688706215
	pesos_i(2532) := b"1111111111111111_1111111111111111_1101111000001001_0011000100101001"; -- -0.1326722406333486
	pesos_i(2533) := b"1111111111111111_1111111111111111_1101100111010011_1100010110110111"; -- -0.14911236082397344
	pesos_i(2534) := b"1111111111111111_1111111111111111_1110110011001110_1100111111100110"; -- -0.07496929775824747
	pesos_i(2535) := b"1111111111111111_1111111111111111_1111100001100011_1111100000011000"; -- -0.029724592279859213
	pesos_i(2536) := b"1111111111111111_1111111111111111_1110111101001110_0010010111010100"; -- -0.06521380967428139
	pesos_i(2537) := b"1111111111111111_1111111111111111_1111101000011011_1110110010110100"; -- -0.023011404199783512
	pesos_i(2538) := b"1111111111111111_1111111111111111_1111001110111010_0110010101101011"; -- -0.04793707026724813
	pesos_i(2539) := b"0000000000000000_0000000000000000_0000101100001101_0111001000010100"; -- 0.043173913770429666
	pesos_i(2540) := b"1111111111111111_1111111111111111_1111011101010001_0010011111001101"; -- -0.03391791580847021
	pesos_i(2541) := b"0000000000000000_0000000000000000_0000010000100110_0110110000110110"; -- 0.01621128383045661
	pesos_i(2542) := b"1111111111111111_1111111111111111_1110100100101001_0000101111000010"; -- -0.08921743884445055
	pesos_i(2543) := b"0000000000000000_0000000000000000_0010101000101101_0001010111100111"; -- 0.16475045103717043
	pesos_i(2544) := b"1111111111111111_1111111111111111_1111001010110111_0110101111101010"; -- -0.05188870940280725
	pesos_i(2545) := b"1111111111111111_1111111111111111_1110111110001010_0110101100000000"; -- -0.06429415940479488
	pesos_i(2546) := b"0000000000000000_0000000000000000_0001001010111010_1011001000001101"; -- 0.07316124740834153
	pesos_i(2547) := b"1111111111111111_1111111111111111_1101111111100110_1101010101100101"; -- -0.1253840091808809
	pesos_i(2548) := b"0000000000000000_0000000000000000_0000111110101110_1111111001110001"; -- 0.06126394527999182
	pesos_i(2549) := b"1111111111111111_1111111111111111_1111110110001000_1101110110110010"; -- -0.00963034066995174
	pesos_i(2550) := b"0000000000000000_0000000000000000_0010101010010010_0000000111101110"; -- 0.16629039822269698
	pesos_i(2551) := b"1111111111111111_1111111111111111_1101111010110010_1110110110000111"; -- -0.1300822778539497
	pesos_i(2552) := b"0000000000000000_0000000000000000_0000011010100011_0100101011100011"; -- 0.025929146212573445
	pesos_i(2553) := b"1111111111111111_1111111111111111_1101100000010100_1100001101010011"; -- -0.15593318198457556
	pesos_i(2554) := b"1111111111111111_1111111111111111_1110101110111111_1010010000001000"; -- -0.07910704435305027
	pesos_i(2555) := b"0000000000000000_0000000000000000_0000110000001000_0000101111000011"; -- 0.046997771291505785
	pesos_i(2556) := b"0000000000000000_0000000000000000_0001011010001000_0011110110100000"; -- 0.0880163684301261
	pesos_i(2557) := b"0000000000000000_0000000000000000_0010011101011101_0000100011111001"; -- 0.15376335218230144
	pesos_i(2558) := b"1111111111111111_1111111111111111_1111001001010000_0101001100110110"; -- -0.05346183713812694
	pesos_i(2559) := b"1111111111111111_1111111111111111_1111100001001111_1101101111110110"; -- -0.030031444922828197
	pesos_i(2560) := b"0000000000000000_0000000000000000_0000111010111010_0110100101011000"; -- 0.05753191369524363
	pesos_i(2561) := b"0000000000000000_0000000000000000_0010000111011100_0110010010111110"; -- 0.13226918824167108
	pesos_i(2562) := b"1111111111111111_1111111111111111_1111110011010110_1110010100110111"; -- -0.012345956948622692
	pesos_i(2563) := b"0000000000000000_0000000000000000_0001000010110110_1010011100001100"; -- 0.06528705642450564
	pesos_i(2564) := b"1111111111111111_1111111111111111_1110100000110100_1111101011010000"; -- -0.09294159337513655
	pesos_i(2565) := b"1111111111111111_1111111111111111_1111011100010000_0000001110000110"; -- -0.034911899291558274
	pesos_i(2566) := b"1111111111111111_1111111111111111_1111111111001000_1111101000101110"; -- -0.0008395802489116942
	pesos_i(2567) := b"1111111111111111_1111111111111111_1110101000100101_1110010110100111"; -- -0.08535923644189705
	pesos_i(2568) := b"1111111111111111_1111111111111111_1110111000011101_1111101010000011"; -- -0.06985506336486337
	pesos_i(2569) := b"1111111111111111_1111111111111111_1101101100100111_1110100101010011"; -- -0.14392224999095102
	pesos_i(2570) := b"0000000000000000_0000000000000000_0000000111111010_1001001011010111"; -- 0.007729699491053174
	pesos_i(2571) := b"1111111111111111_1111111111111111_1101111011000010_1111101011110010"; -- -0.1298373375094841
	pesos_i(2572) := b"0000000000000000_0000000000000000_0010101001111011_1101100000110111"; -- 0.16595221851509984
	pesos_i(2573) := b"0000000000000000_0000000000000000_0001101101000000_1101100010001110"; -- 0.10645822020396901
	pesos_i(2574) := b"0000000000000000_0000000000000000_0000100011000011_0110110100100111"; -- 0.03423196985881158
	pesos_i(2575) := b"0000000000000000_0000000000000000_0010000111100010_0100000001011101"; -- 0.1323585726046538
	pesos_i(2576) := b"1111111111111111_1111111111111111_1111111001101011_0101011010000100"; -- -0.006174652868502523
	pesos_i(2577) := b"1111111111111111_1111111111111111_1101110110001101_0000100010100010"; -- -0.13456674627576348
	pesos_i(2578) := b"1111111111111111_1111111111111111_1101100001010001_0110101111110110"; -- -0.1550076031612932
	pesos_i(2579) := b"1111111111111111_1111111111111111_1101100010001100_1110000001101100"; -- -0.15410039287368069
	pesos_i(2580) := b"1111111111111111_1111111111111111_1110110111010100_0100010110110000"; -- -0.0709797329202937
	pesos_i(2581) := b"1111111111111111_1111111111111111_1110000100101100_0011011101001011"; -- -0.12041906760597756
	pesos_i(2582) := b"1111111111111111_1111111111111111_1111100000101100_1001010001110010"; -- -0.030569765261537495
	pesos_i(2583) := b"0000000000000000_0000000000000000_0000111110010001_0011100010111110"; -- 0.06080965658749575
	pesos_i(2584) := b"0000000000000000_0000000000000000_0000111010111101_1101101010101111"; -- 0.05758444573131387
	pesos_i(2585) := b"0000000000000000_0000000000000000_0001000111011110_1000010101011011"; -- 0.06980164986962034
	pesos_i(2586) := b"0000000000000000_0000000000000000_0000111101010010_0010011101010100"; -- 0.05984731477796528
	pesos_i(2587) := b"1111111111111111_1111111111111111_1101101010000111_1011101101000010"; -- -0.1463664021267296
	pesos_i(2588) := b"0000000000000000_0000000000000000_0010011010111111_0000011111100110"; -- 0.15135239938221265
	pesos_i(2589) := b"0000000000000000_0000000000000000_0010010110001110_1100010011100000"; -- 0.14670973264579215
	pesos_i(2590) := b"0000000000000000_0000000000000000_0001011011100110_1001101011000010"; -- 0.08945624588520065
	pesos_i(2591) := b"0000000000000000_0000000000000000_0001000001001101_0000101101010001"; -- 0.06367560126256214
	pesos_i(2592) := b"0000000000000000_0000000000000000_0000111010101001_0001110000101010"; -- 0.05726791416669086
	pesos_i(2593) := b"1111111111111111_1111111111111111_1111010011101010_0101001000011001"; -- -0.0432995499986443
	pesos_i(2594) := b"1111111111111111_1111111111111111_1111101111001111_1100110000110011"; -- -0.016360509392226257
	pesos_i(2595) := b"1111111111111111_1111111111111111_1110111011010000_1101100111000010"; -- -0.06712569246781616
	pesos_i(2596) := b"0000000000000000_0000000000000000_0000010001101001_0111110111111011"; -- 0.01723468191693971
	pesos_i(2597) := b"1111111111111111_1111111111111111_1111001100010101_0101001001001101"; -- -0.05045590999497575
	pesos_i(2598) := b"0000000000000000_0000000000000000_0010011000000000_0100000101101000"; -- 0.1484413986004414
	pesos_i(2599) := b"1111111111111111_1111111111111111_1110110110000110_0010110001100110"; -- -0.07217142584183223
	pesos_i(2600) := b"1111111111111111_1111111111111111_1101111001101001_1010101010110010"; -- -0.13120015286531644
	pesos_i(2601) := b"1111111111111111_1111111111111111_1111011100010101_0100011010011111"; -- -0.03483160606605336
	pesos_i(2602) := b"1111111111111111_1111111111111111_1111110011000111_1001011011101000"; -- -0.012579506350230732
	pesos_i(2603) := b"1111111111111111_1111111111111111_1110100100011001_1010100011101010"; -- -0.08945221217156152
	pesos_i(2604) := b"0000000000000000_0000000000000000_0001111101011001_0110111100110010"; -- 0.12245841006943226
	pesos_i(2605) := b"1111111111111111_1111111111111111_1111001010110111_0100011011111110"; -- -0.05189091005638276
	pesos_i(2606) := b"0000000000000000_0000000000000000_0001011001101100_0011101010001111"; -- 0.08758893957889131
	pesos_i(2607) := b"0000000000000000_0000000000000000_0001000011011000_0000001111001110"; -- 0.06579612518090468
	pesos_i(2608) := b"0000000000000000_0000000000000000_0001000001110010_1110110001111101"; -- 0.06425359771185268
	pesos_i(2609) := b"0000000000000000_0000000000000000_0000000110001000_1000110011001000"; -- 0.005989836473052549
	pesos_i(2610) := b"0000000000000000_0000000000000000_0001001011001111_0010101001111111"; -- 0.07347360227475151
	pesos_i(2611) := b"1111111111111111_1111111111111111_1111001001111111_1101001000110100"; -- -0.05273710475658762
	pesos_i(2612) := b"1111111111111111_1111111111111111_1110000011001100_1100001010000011"; -- -0.12187561323089346
	pesos_i(2613) := b"0000000000000000_0000000000000000_0001110000101011_1100010101010000"; -- 0.11004288877608562
	pesos_i(2614) := b"0000000000000000_0000000000000000_0000001000000010_1101101110111101"; -- 0.007856114987874955
	pesos_i(2615) := b"0000000000000000_0000000000000000_0001010001110101_1101101010010110"; -- 0.07992330702637761
	pesos_i(2616) := b"0000000000000000_0000000000000000_0000101010000011_1110001001000100"; -- 0.041074887792914155
	pesos_i(2617) := b"1111111111111111_1111111111111111_1111000001100101_0011001001001111"; -- -0.060955863793090086
	pesos_i(2618) := b"0000000000000000_0000000000000000_0000001100110010_0011100101010010"; -- 0.012485106009266448
	pesos_i(2619) := b"0000000000000000_0000000000000000_0001001110000100_1100111101000011"; -- 0.07624526394657259
	pesos_i(2620) := b"1111111111111111_1111111111111111_1101011011111101_0000111100000010"; -- -0.16020113175920261
	pesos_i(2621) := b"0000000000000000_0000000000000000_0001101000110100_1101101101111011"; -- 0.10236903914406287
	pesos_i(2622) := b"1111111111111111_1111111111111111_1110011101011010_1010011010110110"; -- -0.09627302223619372
	pesos_i(2623) := b"1111111111111111_1111111111111111_1101110110110001_1011010000101001"; -- -0.13400720596772434
	pesos_i(2624) := b"0000000000000000_0000000000000000_0010001111110001_0101000011100110"; -- 0.1404009400792582
	pesos_i(2625) := b"1111111111111111_1111111111111111_1110000001100011_1000110100100010"; -- -0.12348096778163532
	pesos_i(2626) := b"0000000000000000_0000000000000000_0010010111100011_0011111110000110"; -- 0.14799878141695227
	pesos_i(2627) := b"1111111111111111_1111111111111111_1111010101101000_1000001011101111"; -- -0.04137403159675013
	pesos_i(2628) := b"0000000000000000_0000000000000000_0001100011100001_0110011100100110"; -- 0.09718937555477372
	pesos_i(2629) := b"1111111111111111_1111111111111111_1110001100111000_1010011000010111"; -- -0.11241685813657701
	pesos_i(2630) := b"0000000000000000_0000000000000000_0001011010000011_0101001001100100"; -- 0.0879413121852928
	pesos_i(2631) := b"1111111111111111_1111111111111111_1110011100101111_0010110011010110"; -- -0.09693641439449842
	pesos_i(2632) := b"1111111111111111_1111111111111111_1100111000000001_1100001110001111"; -- -0.19528558507581018
	pesos_i(2633) := b"1111111111111111_1111111111111111_1111111100101111_0110000000100001"; -- -0.0031833572373535903
	pesos_i(2634) := b"1111111111111111_1111111111111111_1101010011000101_0000001010001010"; -- -0.16886886728672013
	pesos_i(2635) := b"1111111111111111_1111111111111111_1111100011111010_1111111111001100"; -- -0.027420056155270912
	pesos_i(2636) := b"0000000000000000_0000000000000000_0000110111000011_1001010110010011"; -- 0.05376562930091888
	pesos_i(2637) := b"0000000000000000_0000000000000000_0000000111101101_1101101101110100"; -- 0.007535663389033881
	pesos_i(2638) := b"0000000000000000_0000000000000000_0001001110111001_0001101010101001"; -- 0.07704321499630874
	pesos_i(2639) := b"1111111111111111_1111111111111111_1110100000110010_0001100100101011"; -- -0.09298556050519209
	pesos_i(2640) := b"0000000000000000_0000000000000000_0000111000110010_1011011011011011"; -- 0.05546133841275899
	pesos_i(2641) := b"1111111111111111_1111111111111111_1101111001110101_1001110010001000"; -- -0.1310178917334423
	pesos_i(2642) := b"1111111111111111_1111111111111111_1111011101101011_1101000011101011"; -- -0.0335111070843321
	pesos_i(2643) := b"0000000000000000_0000000000000000_0001000010100011_1111001001010111"; -- 0.06500162720142819
	pesos_i(2644) := b"0000000000000000_0000000000000000_0001100011001011_1001010010111011"; -- 0.09685639932181632
	pesos_i(2645) := b"0000000000000000_0000000000000000_0010000000101100_1010011010101101"; -- 0.12568132137200438
	pesos_i(2646) := b"1111111111111111_1111111111111111_1110100110001111_0110001111111100"; -- -0.08765578367020425
	pesos_i(2647) := b"1111111111111111_1111111111111111_1110101100000011_1111110001111010"; -- -0.08197042485868826
	pesos_i(2648) := b"0000000000000000_0000000000000000_0010110011111111_1110011110110100"; -- 0.17577980178802854
	pesos_i(2649) := b"1111111111111111_1111111111111111_1101101110111110_1000100110100101"; -- -0.14162387576670937
	pesos_i(2650) := b"0000000000000000_0000000000000000_0001011011110011_1111100000110101"; -- 0.0896601799344872
	pesos_i(2651) := b"1111111111111111_1111111111111111_1110110101001110_0110101101011000"; -- -0.07302216627306732
	pesos_i(2652) := b"0000000000000000_0000000000000000_0001010000000010_0011011000010001"; -- 0.07815874011788944
	pesos_i(2653) := b"1111111111111111_1111111111111111_1101101101101101_1011010101100011"; -- -0.14285723058938452
	pesos_i(2654) := b"1111111111111111_1111111111111111_1101110010111001_0001010001101100"; -- -0.13780090670557052
	pesos_i(2655) := b"1111111111111111_1111111111111111_1110101011010100_0100110000110001"; -- -0.08269809546435465
	pesos_i(2656) := b"1111111111111111_1111111111111111_1101010101010111_1101111011110010"; -- -0.16662794673323572
	pesos_i(2657) := b"1111111111111111_1111111111111111_1111101110101100_1101010001100011"; -- -0.016894078991372855
	pesos_i(2658) := b"1111111111111111_1111111111111111_1111011100010000_1000110111101000"; -- -0.03490365104942984
	pesos_i(2659) := b"1111111111111111_1111111111111111_1101110010001000_0001010101110000"; -- -0.13854852698034678
	pesos_i(2660) := b"0000000000000000_0000000000000000_0001101011101101_1011110110100111"; -- 0.10519013715168032
	pesos_i(2661) := b"0000000000000000_0000000000000000_0001110111100010_0000010000110101"; -- 0.11672998699633895
	pesos_i(2662) := b"0000000000000000_0000000000000000_0000011010101110_1100011011110100"; -- 0.02610438772344584
	pesos_i(2663) := b"0000000000000000_0000000000000000_0001011110001010_1110001000011110"; -- 0.09196294044330597
	pesos_i(2664) := b"1111111111111111_1111111111111111_1101100111110000_0110011001001110"; -- -0.14867554290195198
	pesos_i(2665) := b"0000000000000000_0000000000000000_0000100001110100_1011110100100100"; -- 0.03303129329528527
	pesos_i(2666) := b"0000000000000000_0000000000000000_0000011000101101_1000100000000100"; -- 0.024132252643955396
	pesos_i(2667) := b"1111111111111111_1111111111111111_1110010100001100_0100000011101111"; -- -0.10528177407898184
	pesos_i(2668) := b"0000000000000000_0000000000000000_0010001111100010_0100101001010111"; -- 0.1401716672158267
	pesos_i(2669) := b"1111111111111111_1111111111111111_1101101010111101_0000001110101010"; -- -0.14555337048630748
	pesos_i(2670) := b"0000000000000000_0000000000000000_0001111001111001_0100110001011100"; -- 0.11903836495150026
	pesos_i(2671) := b"1111111111111111_1111111111111111_1111000001001110_1001111101011010"; -- -0.0613003164597472
	pesos_i(2672) := b"0000000000000000_0000000000000000_0001010111011001_0110101011000101"; -- 0.08534877118050224
	pesos_i(2673) := b"1111111111111111_1111111111111111_1101100100000001_0011011110001100"; -- -0.15232518029011582
	pesos_i(2674) := b"1111111111111111_1111111111111111_1110100000110010_1110111100111110"; -- -0.09297280067011861
	pesos_i(2675) := b"0000000000000000_0000000000000000_0010001011001100_1100010111101011"; -- 0.13593708989338832
	pesos_i(2676) := b"0000000000000000_0000000000000000_0000001110111100_0010111010011011"; -- 0.014590180195445408
	pesos_i(2677) := b"0000000000000000_0000000000000000_0010000101011011_0010010110111100"; -- 0.13029704893040425
	pesos_i(2678) := b"1111111111111111_1111111111111111_1111011011100010_1111011100101000"; -- -0.03559928202271138
	pesos_i(2679) := b"0000000000000000_0000000000000000_0001101100110110_1111110010111000"; -- 0.1063077878142982
	pesos_i(2680) := b"0000000000000000_0000000000000000_0000110000010100_1010011000010000"; -- 0.04719007377498849
	pesos_i(2681) := b"1111111111111111_1111111111111111_1111101000001001_0110000010110101"; -- -0.023294406722722816
	pesos_i(2682) := b"1111111111111111_1111111111111111_1101100111010001_1011000101010001"; -- -0.14914409413896948
	pesos_i(2683) := b"0000000000000000_0000000000000000_0001001001000000_0000111001011010"; -- 0.07128991803124111
	pesos_i(2684) := b"1111111111111111_1111111111111111_1111000011111011_1100011001111011"; -- -0.05865821370065196
	pesos_i(2685) := b"1111111111111111_1111111111111111_1111011000001110_1100101111011111"; -- -0.038836725298765654
	pesos_i(2686) := b"1111111111111111_1111111111111111_1111001100010100_0001110011010111"; -- -0.050474355275918974
	pesos_i(2687) := b"0000000000000000_0000000000000000_0010110110001110_0001001101001100"; -- 0.17794914814654483
	pesos_i(2688) := b"1111111111111111_1111111111111111_1101111111001010_0011000010010000"; -- -0.12582108005768022
	pesos_i(2689) := b"0000000000000000_0000000000000000_0001011001101111_0110001111100000"; -- 0.08763717864504189
	pesos_i(2690) := b"0000000000000000_0000000000000000_0000010010101010_0101101011111111"; -- 0.018224417866278052
	pesos_i(2691) := b"1111111111111111_1111111111111111_1101011111010111_1101101101000100"; -- -0.15686254107318479
	pesos_i(2692) := b"0000000000000000_0000000000000000_0010010010111100_1111101110100010"; -- 0.14350865083715075
	pesos_i(2693) := b"0000000000000000_0000000000000000_0010101101111011_0000011000001111"; -- 0.16984594229000713
	pesos_i(2694) := b"0000000000000000_0000000000000000_0001011000000000_0000000001000101"; -- 0.08593751617902136
	pesos_i(2695) := b"0000000000000000_0000000000000000_0001111011110111_1011010001110101"; -- 0.12096717694257667
	pesos_i(2696) := b"1111111111111111_1111111111111111_1111011111001111_0000001000011001"; -- -0.03199755563395454
	pesos_i(2697) := b"1111111111111111_1111111111111111_1111011011100100_1000101001110010"; -- -0.03557524419530514
	pesos_i(2698) := b"1111111111111111_1111111111111111_1111100001100010_1101010111100101"; -- -0.029741889527337317
	pesos_i(2699) := b"0000000000000000_0000000000000000_0010000111100110_1001100001001111"; -- 0.13242484968855978
	pesos_i(2700) := b"0000000000000000_0000000000000000_0001111001010100_1100011110111101"; -- 0.11848114354606787
	pesos_i(2701) := b"1111111111111111_1111111111111111_1110000111010101_0111110010100001"; -- -0.1178361994055992
	pesos_i(2702) := b"0000000000000000_0000000000000000_0000110011000010_0111001101111001"; -- 0.0498420876878209
	pesos_i(2703) := b"0000000000000000_0000000000000000_0001001111010000_0000110111100110"; -- 0.07739340653764966
	pesos_i(2704) := b"0000000000000000_0000000000000000_0000001001000010_1000110000011111"; -- 0.008827931830264563
	pesos_i(2705) := b"1111111111111111_1111111111111111_1101110100000001_1110111100110110"; -- -0.13668923318740614
	pesos_i(2706) := b"0000000000000000_0000000000000000_0001111101000001_0110101000111111"; -- 0.1220919040739939
	pesos_i(2707) := b"0000000000000000_0000000000000000_0001100100111001_0110100101110000"; -- 0.0985322856341613
	pesos_i(2708) := b"0000000000000000_0000000000000000_0000100111110000_1100001010100110"; -- 0.03882996139893478
	pesos_i(2709) := b"0000000000000000_0000000000000000_0000011100111100_1101110101101011"; -- 0.02827247480613783
	pesos_i(2710) := b"0000000000000000_0000000000000000_0010110111011011_1011110010010110"; -- 0.1791341653454943
	pesos_i(2711) := b"1111111111111111_1111111111111111_1101100111000110_1001010100010100"; -- -0.14931362400596934
	pesos_i(2712) := b"0000000000000000_0000000000000000_0000010111110010_1101100001111000"; -- 0.023236779398642306
	pesos_i(2713) := b"1111111111111111_1111111111111111_1101110001001101_0101011101000110"; -- -0.1394448713056114
	pesos_i(2714) := b"0000000000000000_0000000000000000_0010011100010111_1111000111110001"; -- 0.1527091229505172
	pesos_i(2715) := b"1111111111111111_1111111111111111_1101101011011010_0100101110110001"; -- -0.14510657250578476
	pesos_i(2716) := b"0000000000000000_0000000000000000_0000101101010100_0100000110010001"; -- 0.04425439638183504
	pesos_i(2717) := b"1111111111111111_1111111111111111_1101111110100100_1111001011111110"; -- -0.12638932501595496
	pesos_i(2718) := b"1111111111111111_1111111111111111_1101111110011110_1010110010110100"; -- -0.1264850675313997
	pesos_i(2719) := b"1111111111111111_1111111111111111_1101101101000011_1110110001110101"; -- -0.14349481718007218
	pesos_i(2720) := b"1111111111111111_1111111111111111_1110001101011110_0100111110101110"; -- -0.11184217447688172
	pesos_i(2721) := b"0000000000000000_0000000000000000_0010111101000000_1101011010011101"; -- 0.184583104367053
	pesos_i(2722) := b"1111111111111111_1111111111111111_1101101101001111_1111011110010011"; -- -0.14331104918468476
	pesos_i(2723) := b"0000000000000000_0000000000000000_0000100011111110_1100001000001101"; -- 0.03513729883254692
	pesos_i(2724) := b"0000000000000000_0000000000000000_0000011000011001_0100101000000010"; -- 0.02382338099300436
	pesos_i(2725) := b"1111111111111111_1111111111111111_1101110001011011_0110110001001011"; -- -0.13922999540705866
	pesos_i(2726) := b"0000000000000000_0000000000000000_0001011101101000_0000101110110001"; -- 0.09143136090083889
	pesos_i(2727) := b"1111111111111111_1111111111111111_1101001100011011_1000110111101110"; -- -0.1753608029235476
	pesos_i(2728) := b"1111111111111111_1111111111111111_1110110100000011_1010101011011111"; -- -0.07416278901308355
	pesos_i(2729) := b"0000000000000000_0000000000000000_0000011101101011_1111010110101101"; -- 0.028991083933235753
	pesos_i(2730) := b"0000000000000000_0000000000000000_0001101100000101_1111010010100100"; -- 0.10555962556643571
	pesos_i(2731) := b"1111111111111111_1111111111111111_1101101000010110_0000101001000111"; -- -0.14810119406199432
	pesos_i(2732) := b"0000000000000000_0000000000000000_0000001111111100_0100010000111100"; -- 0.015568031832717402
	pesos_i(2733) := b"1111111111111111_1111111111111111_1111100110110010_1000010100001100"; -- -0.024619755411418916
	pesos_i(2734) := b"0000000000000000_0000000000000000_0010100110000100_0100011001110001"; -- 0.16217460885201038
	pesos_i(2735) := b"0000000000000000_0000000000000000_0010101101100110_0010010000010001"; -- 0.16952729611303047
	pesos_i(2736) := b"1111111111111111_1111111111111111_1111011111111100_0001100010001000"; -- -0.03130957288012867
	pesos_i(2737) := b"0000000000000000_0000000000000000_0000000100100001_1000111010010010"; -- 0.0044182878329211755
	pesos_i(2738) := b"0000000000000000_0000000000000000_0010001100010001_0000110110110110"; -- 0.1369789665532812
	pesos_i(2739) := b"1111111111111111_1111111111111111_1111000101010100_0110010101110011"; -- -0.05730596484016524
	pesos_i(2740) := b"0000000000000000_0000000000000000_0001010001100100_0001101101101110"; -- 0.07965251377916983
	pesos_i(2741) := b"1111111111111111_1111111111111111_1101011001000100_1101101000000111"; -- -0.16301190688316744
	pesos_i(2742) := b"1111111111111111_1111111111111111_1101010010010000_1110110101110100"; -- -0.16966358113186333
	pesos_i(2743) := b"0000000000000000_0000000000000000_0001101111011101_1101010110101111"; -- 0.10885367887126733
	pesos_i(2744) := b"0000000000000000_0000000000000000_0001100101000111_1000011001011011"; -- 0.09874763229787079
	pesos_i(2745) := b"0000000000000000_0000000000000000_0000110001101010_1111101000011010"; -- 0.04850733893551531
	pesos_i(2746) := b"0000000000000000_0000000000000000_0001110111111000_1010010111111010"; -- 0.11707532262901134
	pesos_i(2747) := b"1111111111111111_1111111111111111_1110010101000110_1101001100110111"; -- -0.10438804544867887
	pesos_i(2748) := b"0000000000000000_0000000000000000_0010001111101001_0111011001100100"; -- 0.14028110456011086
	pesos_i(2749) := b"1111111111111111_1111111111111111_1110001111101011_0111001000110100"; -- -0.10968862743537741
	pesos_i(2750) := b"0000000000000000_0000000000000000_0001101111101111_0101010000011100"; -- 0.10912061388565869
	pesos_i(2751) := b"1111111111111111_1111111111111111_1110111101010000_0010001110000101"; -- -0.06518342983176613
	pesos_i(2752) := b"1111111111111111_1111111111111111_1110010001110100_1101100111011011"; -- -0.10759199522847326
	pesos_i(2753) := b"0000000000000000_0000000000000000_0001101001001000_0010000100010000"; -- 0.10266310352383091
	pesos_i(2754) := b"1111111111111111_1111111111111111_1110001111011110_0101111000001101"; -- -0.10988819298415403
	pesos_i(2755) := b"0000000000000000_0000000000000000_0001100010101101_1111101110000100"; -- 0.09640476194628939
	pesos_i(2756) := b"1111111111111111_1111111111111111_1101111011011100_1101010000110011"; -- -0.12944291830419916
	pesos_i(2757) := b"1111111111111111_1111111111111111_1110001101111010_1101100010101011"; -- -0.11140676320619655
	pesos_i(2758) := b"1111111111111111_1111111111111111_1111100111000011_0111100001110011"; -- -0.024361106788904734
	pesos_i(2759) := b"1111111111111111_1111111111111111_1111101101000011_1010100010001101"; -- -0.018498864638202345
	pesos_i(2760) := b"0000000000000000_0000000000000000_0000011011110101_0011001000011000"; -- 0.027178889102435842
	pesos_i(2761) := b"0000000000000000_0000000000000000_0001011100111110_1101111111011101"; -- 0.09080313824261128
	pesos_i(2762) := b"1111111111111111_1111111111111111_1101100111001110_0000110100011100"; -- -0.1491996581015588
	pesos_i(2763) := b"1111111111111111_1111111111111111_1110011000011001_0001100101000010"; -- -0.10117952480590162
	pesos_i(2764) := b"0000000000000000_0000000000000000_0000100001100110_1110110100110101"; -- 0.03282053519886395
	pesos_i(2765) := b"1111111111111111_1111111111111111_1110101110111100_0010100111110100"; -- -0.07916009694606169
	pesos_i(2766) := b"0000000000000000_0000000000000000_0010100101101111_0110001011100000"; -- 0.16185586898389043
	pesos_i(2767) := b"1111111111111111_1111111111111111_1111111001000111_0010000011100010"; -- -0.006727166028297835
	pesos_i(2768) := b"1111111111111111_1111111111111111_1110111010010001_0110111010011101"; -- -0.0680933824333735
	pesos_i(2769) := b"1111111111111111_1111111111111111_1101101000011100_0110100000010100"; -- -0.14800405043834386
	pesos_i(2770) := b"1111111111111111_1111111111111111_1101101010001001_0011010010011110"; -- -0.1463439096373757
	pesos_i(2771) := b"0000000000000000_0000000000000000_0001111111000010_1110100100110001"; -- 0.12406785434422876
	pesos_i(2772) := b"0000000000000000_0000000000000000_0001000001101111_0100010110001101"; -- 0.06419787119694056
	pesos_i(2773) := b"1111111111111111_1111111111111111_1101010011001001_1000011001100110"; -- -0.16879997258253118
	pesos_i(2774) := b"1111111111111111_1111111111111111_1101111110100100_0110011000011110"; -- -0.1263977220064346
	pesos_i(2775) := b"0000000000000000_0000000000000000_0010011011010001_0010011000110010"; -- 0.1516288635395976
	pesos_i(2776) := b"1111111111111111_1111111111111111_1101000011000100_1111001101100111"; -- -0.1844947695434404
	pesos_i(2777) := b"1111111111111111_1111111111111111_1101010100011000_1101011000101101"; -- -0.16758977314918788
	pesos_i(2778) := b"1111111111111111_1111111111111111_1111101110000001_0011010010001011"; -- -0.01755973450255065
	pesos_i(2779) := b"0000000000000000_0000000000000000_0001011000111011_1010110010010111"; -- 0.08684805560350758
	pesos_i(2780) := b"0000000000000000_0000000000000000_0001100110101101_0011110101110010"; -- 0.10029968291254536
	pesos_i(2781) := b"1111111111111111_1111111111111111_1111110010111001_1100101011000000"; -- -0.01279003909186586
	pesos_i(2782) := b"0000000000000000_0000000000000000_0000110011010101_0011100010000001"; -- 0.05012848996919184
	pesos_i(2783) := b"1111111111111111_1111111111111111_1101101000001110_0111111010101000"; -- -0.1482163276646613
	pesos_i(2784) := b"0000000000000000_0000000000000000_0001011011001000_0001111100111000"; -- 0.08899111858298628
	pesos_i(2785) := b"1111111111111111_1111111111111111_1110001110001111_1111000110110100"; -- -0.11108483643729541
	pesos_i(2786) := b"0000000000000000_0000000000000000_0001111111011101_0100101101110111"; -- 0.12447044047188897
	pesos_i(2787) := b"1111111111111111_1111111111111111_1101110100100110_1001000001110000"; -- -0.1361303068513186
	pesos_i(2788) := b"0000000000000000_0000000000000000_0001000000110111_1111101010101111"; -- 0.06335417521033802
	pesos_i(2789) := b"0000000000000000_0000000000000000_0000101001100101_1010100110011010"; -- 0.04061374681321441
	pesos_i(2790) := b"0000000000000000_0000000000000000_0010000011101110_0001011001101110"; -- 0.12863292866117626
	pesos_i(2791) := b"1111111111111111_1111111111111111_1101110011101110_0010111101000101"; -- -0.13699059082281195
	pesos_i(2792) := b"1111111111111111_1111111111111111_1110110100111100_0100101111111100"; -- -0.07329869374207694
	pesos_i(2793) := b"0000000000000000_0000000000000000_0001111001110001_0001001111100001"; -- 0.11891292815362647
	pesos_i(2794) := b"0000000000000000_0000000000000000_0000110111000101_0101010010111110"; -- 0.05379228246573541
	pesos_i(2795) := b"0000000000000000_0000000000000000_0001000100111111_1111100000011100"; -- 0.06738234220199515
	pesos_i(2796) := b"0000000000000000_0000000000000000_0001010000011001_0011010101100001"; -- 0.07850965144288526
	pesos_i(2797) := b"1111111111111111_1111111111111111_1111011110001100_0100111110100010"; -- -0.033015272991348696
	pesos_i(2798) := b"0000000000000000_0000000000000000_0001101001001001_0100011100010111"; -- 0.1026806289644583
	pesos_i(2799) := b"1111111111111111_1111111111111111_1101011011010000_1100010100010101"; -- -0.1608769248919229
	pesos_i(2800) := b"1111111111111111_1111111111111111_1111100010011001_1000100101110101"; -- -0.02890721227701956
	pesos_i(2801) := b"0000000000000000_0000000000000000_0001101000101010_1110100001100110"; -- 0.10221722107403437
	pesos_i(2802) := b"0000000000000000_0000000000000000_0001011100101101_0111100001011010"; -- 0.09053756894267496
	pesos_i(2803) := b"0000000000000000_0000000000000000_0001110100010111_0001101100101101"; -- 0.11363382194772532
	pesos_i(2804) := b"1111111111111111_1111111111111111_1101101110011001_1101010001110011"; -- -0.14218399228736417
	pesos_i(2805) := b"0000000000000000_0000000000000000_0010100110001100_1001011011010001"; -- 0.1623014698204408
	pesos_i(2806) := b"1111111111111111_1111111111111111_1110011011111110_1111000100110010"; -- -0.09767239113767824
	pesos_i(2807) := b"1111111111111111_1111111111111111_1111010011101110_1000001110100001"; -- -0.04323556250500976
	pesos_i(2808) := b"0000000000000000_0000000000000000_0000101001111010_1010111000000111"; -- 0.040934445064492564
	pesos_i(2809) := b"0000000000000000_0000000000000000_0000101111110010_1010010110000110"; -- 0.04667124301709305
	pesos_i(2810) := b"0000000000000000_0000000000000000_0000111111010111_0111001100101010"; -- 0.061881253910440505
	pesos_i(2811) := b"1111111111111111_1111111111111111_1110001111001000_0001111110111111"; -- -0.1102276000870972
	pesos_i(2812) := b"0000000000000000_0000000000000000_0000111100110011_1100100000000010"; -- 0.05938386967288819
	pesos_i(2813) := b"0000000000000000_0000000000000000_0010100010100000_1100111001001111"; -- 0.15870370317655302
	pesos_i(2814) := b"0000000000000000_0000000000000000_0001010110010110_1011010010100001"; -- 0.08433083458884152
	pesos_i(2815) := b"1111111111111111_1111111111111111_1111100001010001_1011101001011110"; -- -0.030002929664706544
	pesos_i(2816) := b"0000000000000000_0000000000000000_0010011000000100_1111100111100011"; -- 0.1485134295973898
	pesos_i(2817) := b"0000000000000000_0000000000000000_0001011010000011_0111011011010011"; -- 0.08794348382797189
	pesos_i(2818) := b"1111111111111111_1111111111111111_1110001001100001_1111111111111100"; -- -0.11569213958903214
	pesos_i(2819) := b"1111111111111111_1111111111111111_1110100101010111_1001010000000010"; -- -0.08850741328490302
	pesos_i(2820) := b"0000000000000000_0000000000000000_0001000100110011_0110100110011100"; -- 0.06719074305234486
	pesos_i(2821) := b"0000000000000000_0000000000000000_0000100101111111_0101111001010010"; -- 0.03709973813203395
	pesos_i(2822) := b"1111111111111111_1111111111111111_1111111101011101_0011110111110001"; -- -0.002483490683945036
	pesos_i(2823) := b"1111111111111111_1111111111111111_1111100100100100_1100100010011010"; -- -0.026782476757964024
	pesos_i(2824) := b"0000000000000000_0000000000000000_0000100110101011_0101010001111100"; -- 0.03777053862842131
	pesos_i(2825) := b"0000000000000000_0000000000000000_0000000101011111_1101010111100111"; -- 0.0053685845390506965
	pesos_i(2826) := b"1111111111111111_1111111111111111_1111101111010101_0000111010110110"; -- -0.01628025113615244
	pesos_i(2827) := b"1111111111111111_1111111111111111_1110110001000111_0111011000010010"; -- -0.07703458847186764
	pesos_i(2828) := b"1111111111111111_1111111111111111_1111100101011110_1000101011100101"; -- -0.025901144981510544
	pesos_i(2829) := b"0000000000000000_0000000000000000_0000010100101110_0001100001001011"; -- 0.020234602213464715
	pesos_i(2830) := b"0000000000000000_0000000000000000_0010011110001110_0101111101011100"; -- 0.15451618191897734
	pesos_i(2831) := b"0000000000000000_0000000000000000_0010100111100001_1010000110111100"; -- 0.16359911765529614
	pesos_i(2832) := b"0000000000000000_0000000000000000_0000010000111101_0010101110011101"; -- 0.01655838569513257
	pesos_i(2833) := b"1111111111111111_1111111111111111_1101010100100010_0001000011000000"; -- -0.16744895280372898
	pesos_i(2834) := b"0000000000000000_0000000000000000_0001010011000010_1110010111100010"; -- 0.08109890720618325
	pesos_i(2835) := b"1111111111111111_1111111111111111_1110001010010011_0100100101001110"; -- -0.11494008873841455
	pesos_i(2836) := b"1111111111111111_1111111111111111_1111000000100111_0011110110101001"; -- -0.06190123201961926
	pesos_i(2837) := b"1111111111111111_1111111111111111_1101010010011010_1001101110100111"; -- -0.16951586896327903
	pesos_i(2838) := b"1111111111111111_1111111111111111_1110001110111001_0010011010000011"; -- -0.11045607846218916
	pesos_i(2839) := b"1111111111111111_1111111111111111_1101110010011111_1101110000111010"; -- -0.13818572592036607
	pesos_i(2840) := b"1111111111111111_1111111111111111_1110011101000001_1000000011101100"; -- -0.09665674430326984
	pesos_i(2841) := b"0000000000000000_0000000000000000_0001110100000111_1110110011101000"; -- 0.11340218218634039
	pesos_i(2842) := b"0000000000000000_0000000000000000_0001010000100000_1010011110011110"; -- 0.0786232720544224
	pesos_i(2843) := b"0000000000000000_0000000000000000_0000011101011101_0101111110110011"; -- 0.02876852155597757
	pesos_i(2844) := b"1111111111111111_1111111111111111_1110001110001101_0001010101001101"; -- -0.11112849102604092
	pesos_i(2845) := b"0000000000000000_0000000000000000_0010101101101011_1011000101101101"; -- 0.16961201574697704
	pesos_i(2846) := b"0000000000000000_0000000000000000_0001101001101110_1111011011000011"; -- 0.10325567502824047
	pesos_i(2847) := b"0000000000000000_0000000000000000_0001110101001111_1111101011101101"; -- 0.11450165075168947
	pesos_i(2848) := b"1111111111111111_1111111111111111_1110000000110010_0001110100010001"; -- -0.12423532800349374
	pesos_i(2849) := b"0000000000000000_0000000000000000_0001101110110011_1001100101000111"; -- 0.10820920924500309
	pesos_i(2850) := b"1111111111111111_1111111111111111_1111100011110011_1000011010110100"; -- -0.027534085271541227
	pesos_i(2851) := b"0000000000000000_0000000000000000_0001110011011000_0010111010101011"; -- 0.11267368011837865
	pesos_i(2852) := b"1111111111111111_1111111111111111_1110000110100010_0111111110110010"; -- -0.1186142148434598
	pesos_i(2853) := b"0000000000000000_0000000000000000_0010010110111110_1010110010110000"; -- 0.1474407128276537
	pesos_i(2854) := b"0000000000000000_0000000000000000_0000000111010001_1110010111111001"; -- 0.007109044448113795
	pesos_i(2855) := b"0000000000000000_0000000000000000_0010101001010001_0011100110001111"; -- 0.16530189266977566
	pesos_i(2856) := b"0000000000000000_0000000000000000_0001011001001101_1100111110111100"; -- 0.08712480877873643
	pesos_i(2857) := b"1111111111111111_1111111111111111_1111110010110010_0000011110001001"; -- -0.012908486382282418
	pesos_i(2858) := b"1111111111111111_1111111111111111_1111101001011110_0011010010100010"; -- -0.022000036693808244
	pesos_i(2859) := b"0000000000000000_0000000000000000_0010110100101110_0110001000100001"; -- 0.1764890031258408
	pesos_i(2860) := b"0000000000000000_0000000000000000_0010010101101101_0001100011110011"; -- 0.14619594507308678
	pesos_i(2861) := b"0000000000000000_0000000000000000_0000110011011101_0110011111000110"; -- 0.05025337784438043
	pesos_i(2862) := b"0000000000000000_0000000000000000_0000000111000111_1110110110000010"; -- 0.0069569055014507076
	pesos_i(2863) := b"1111111111111111_1111111111111111_1111111110011111_1100100001101010"; -- -0.0014681570166245293
	pesos_i(2864) := b"1111111111111111_1111111111111111_1111100000110000_1001111100100101"; -- -0.030508092275816467
	pesos_i(2865) := b"1111111111111111_1111111111111111_1110010001101100_1100101001000101"; -- -0.10771499450680937
	pesos_i(2866) := b"1111111111111111_1111111111111111_1111110101000101_0010101000000010"; -- -0.010663389747991825
	pesos_i(2867) := b"1111111111111111_1111111111111111_1111010100000011_1111001100010010"; -- -0.04290848544742355
	pesos_i(2868) := b"0000000000000000_0000000000000000_0010000111101100_0100101001001111"; -- 0.13251175325460413
	pesos_i(2869) := b"1111111111111111_1111111111111111_1111010111011110_1000100000011100"; -- -0.0395731860100106
	pesos_i(2870) := b"0000000000000000_0000000000000000_0000110000110010_1001100000101100"; -- 0.047647009654011634
	pesos_i(2871) := b"0000000000000000_0000000000000000_0000101110010110_0011100101111001"; -- 0.04526099392274367
	pesos_i(2872) := b"0000000000000000_0000000000000000_0010001011101001_1101100011001010"; -- 0.1363807193803003
	pesos_i(2873) := b"1111111111111111_1111111111111111_1101111101001101_0000001110101010"; -- -0.1277311048813623
	pesos_i(2874) := b"0000000000000000_0000000000000000_0000000110111110_1011011110110100"; -- 0.006816369406453165
	pesos_i(2875) := b"0000000000000000_0000000000000000_0010111001000101_1011001001111111"; -- 0.18075099574114398
	pesos_i(2876) := b"0000000000000000_0000000000000000_0010101000101001_0001000011101111"; -- 0.1646891196618015
	pesos_i(2877) := b"0000000000000000_0000000000000000_0000111101111010_1011110101010110"; -- 0.06046660752210555
	pesos_i(2878) := b"0000000000000000_0000000000000000_0001000100001101_0110000101000111"; -- 0.06661041243577438
	pesos_i(2879) := b"1111111111111111_1111111111111111_1110110000100100_0110111000110000"; -- -0.07756911581179048
	pesos_i(2880) := b"0000000000000000_0000000000000000_0001011100000100_0010001110100110"; -- 0.08990691001403753
	pesos_i(2881) := b"0000000000000000_0000000000000000_0000100111011011_1101111011000101"; -- 0.03851120281708207
	pesos_i(2882) := b"0000000000000000_0000000000000000_0010011011011000_1000111000010000"; -- 0.1517418659194873
	pesos_i(2883) := b"0000000000000000_0000000000000000_0000011110100011_0101000010101110"; -- 0.029835741617455138
	pesos_i(2884) := b"0000000000000000_0000000000000000_0010010000111111_0100101100001110"; -- 0.14159077728579428
	pesos_i(2885) := b"1111111111111111_1111111111111111_1110101001001001_0011110111011100"; -- -0.0848199213209565
	pesos_i(2886) := b"0000000000000000_0000000000000000_0000010010001111_0101010000000110"; -- 0.017812015094166463
	pesos_i(2887) := b"0000000000000000_0000000000000000_0000010010111001_0110001011001111"; -- 0.01845376532986312
	pesos_i(2888) := b"1111111111111111_1111111111111111_1101011000010000_1101110111011100"; -- -0.16380513546481032
	pesos_i(2889) := b"0000000000000000_0000000000000000_0000100011110101_1011101001110110"; -- 0.03499951729971147
	pesos_i(2890) := b"1111111111111111_1111111111111111_1110100100010001_1010100000100110"; -- -0.08957432811952681
	pesos_i(2891) := b"0000000000000000_0000000000000000_0010001101010100_1011010010100111"; -- 0.13801125605787865
	pesos_i(2892) := b"0000000000000000_0000000000000000_0001110111011101_1000010010010011"; -- 0.11666134451733108
	pesos_i(2893) := b"1111111111111111_1111111111111111_1101011000111101_1101101000010100"; -- -0.16311871530113464
	pesos_i(2894) := b"0000000000000000_0000000000000000_0001111000100010_0010110101110011"; -- 0.1177090078485474
	pesos_i(2895) := b"1111111111111111_1111111111111111_1111001011101011_1011101110000101"; -- -0.051090507593565176
	pesos_i(2896) := b"0000000000000000_0000000000000000_0001011000000000_1100110100010001"; -- 0.08594972294936779
	pesos_i(2897) := b"0000000000000000_0000000000000000_0001100110000000_1011111000110011"; -- 0.09962071174927126
	pesos_i(2898) := b"0000000000000000_0000000000000000_0000010001011000_0011110011111001"; -- 0.01697140775960749
	pesos_i(2899) := b"0000000000000000_0000000000000000_0000010001010011_0110000011011001"; -- 0.01689725205005404
	pesos_i(2900) := b"1111111111111111_1111111111111111_1110011000101100_1011001000110101"; -- -0.10088049140925884
	pesos_i(2901) := b"1111111111111111_1111111111111111_1110000010001000_0100000110101111"; -- -0.12292088960411739
	pesos_i(2902) := b"1111111111111111_1111111111111111_1110100001111010_0101000100101001"; -- -0.09188359011803154
	pesos_i(2903) := b"0000000000000000_0000000000000000_0001101011101100_0110110010011101"; -- 0.10517004807769048
	pesos_i(2904) := b"0000000000000000_0000000000000000_0000111101110011_0001001101110101"; -- 0.06034967036952815
	pesos_i(2905) := b"1111111111111111_1111111111111111_1111101011111101_1101011100001100"; -- -0.01956420846295684
	pesos_i(2906) := b"0000000000000000_0000000000000000_0001001100000011_0100100000000010"; -- 0.07426881838626974
	pesos_i(2907) := b"0000000000000000_0000000000000000_0000001101101011_0101010010000001"; -- 0.013356477165206089
	pesos_i(2908) := b"1111111111111111_1111111111111111_1101100010110101_1011000010011100"; -- -0.1534776324197981
	pesos_i(2909) := b"0000000000000000_0000000000000000_0010010100110010_0100000101111000"; -- 0.14529809165383348
	pesos_i(2910) := b"0000000000000000_0000000000000000_0001011000110110_1001110111000110"; -- 0.08677087863045817
	pesos_i(2911) := b"0000000000000000_0000000000000000_0010110000000110_0001011111011011"; -- 0.1719679745910753
	pesos_i(2912) := b"1111111111111111_1111111111111111_1101110011101001_0000101010011010"; -- -0.13706907033976606
	pesos_i(2913) := b"0000000000000000_0000000000000000_0010010011111000_1111000001100010"; -- 0.14442350770409196
	pesos_i(2914) := b"0000000000000000_0000000000000000_0000101000110010_1111001100011111"; -- 0.039839930573285755
	pesos_i(2915) := b"1111111111111111_1111111111111111_1110111001001110_1111111010011100"; -- -0.06910713864218719
	pesos_i(2916) := b"1111111111111111_1111111111111111_1110100100011111_1001001001010111"; -- -0.08936200494012642
	pesos_i(2917) := b"1111111111111111_1111111111111111_1111000001110010_0000000000010011"; -- -0.06076049364510805
	pesos_i(2918) := b"0000000000000000_0000000000000000_0010000011001101_0010001110101111"; -- 0.12813017858726047
	pesos_i(2919) := b"1111111111111111_1111111111111111_1101010000010101_1001111101111001"; -- -0.1715450600628621
	pesos_i(2920) := b"0000000000000000_0000000000000000_0000111100100011_1100101010111011"; -- 0.0591398912487128
	pesos_i(2921) := b"1111111111111111_1111111111111111_1110011000011110_0011001111001000"; -- -0.1011016499116965
	pesos_i(2922) := b"1111111111111111_1111111111111111_1110000110011010_1100100110011110"; -- -0.11873187921742198
	pesos_i(2923) := b"1111111111111111_1111111111111111_1110101100100010_0101110010100011"; -- -0.08150692948009623
	pesos_i(2924) := b"1111111111111111_1111111111111111_1111110000111100_0010010010011010"; -- -0.014707290993187828
	pesos_i(2925) := b"0000000000000000_0000000000000000_0001110101110101_0000000010111110"; -- 0.11506657247061615
	pesos_i(2926) := b"1111111111111111_1111111111111111_1111000101001110_0110101100001101"; -- -0.05739718374554109
	pesos_i(2927) := b"1111111111111111_1111111111111111_1111111010001110_1100011011011101"; -- -0.005633898838290009
	pesos_i(2928) := b"1111111111111111_1111111111111111_1110101010100000_0010000001111110"; -- -0.08349415697995864
	pesos_i(2929) := b"0000000000000000_0000000000000000_0001110001101101_0100001001001010"; -- 0.11104215912419331
	pesos_i(2930) := b"0000000000000000_0000000000000000_0010100111110111_0101111100110011"; -- 0.1639308452311668
	pesos_i(2931) := b"0000000000000000_0000000000000000_0010101100100101_1010000011101100"; -- 0.1685429168144222
	pesos_i(2932) := b"1111111111111111_1111111111111111_1110001110100010_0110111010000110"; -- -0.11080273851697145
	pesos_i(2933) := b"0000000000000000_0000000000000000_0000000100110010_0110000011001101"; -- 0.004674959290530997
	pesos_i(2934) := b"0000000000000000_0000000000000000_0010100111001010_0001101011110110"; -- 0.1632401323338239
	pesos_i(2935) := b"0000000000000000_0000000000000000_0001100111010010_1000001111000011"; -- 0.10086844919777048
	pesos_i(2936) := b"0000000000000000_0000000000000000_0010110000111111_0110010001111010"; -- 0.17284229250058927
	pesos_i(2937) := b"0000000000000000_0000000000000000_0000100010111000_0001011100011101"; -- 0.03405899486528398
	pesos_i(2938) := b"1111111111111111_1111111111111111_1111001111101110_0010100110001100"; -- -0.047147181931456984
	pesos_i(2939) := b"1111111111111111_1111111111111111_1111101101110010_0101011101001111"; -- -0.017786544165477276
	pesos_i(2940) := b"0000000000000000_0000000000000000_0000011100001010_1010110101001110"; -- 0.027506667707215923
	pesos_i(2941) := b"0000000000000000_0000000000000000_0001110100000000_0101010001001101"; -- 0.11328627463853097
	pesos_i(2942) := b"1111111111111111_1111111111111111_1101101010101010_1110111011010110"; -- -0.1458292701185864
	pesos_i(2943) := b"0000000000000000_0000000000000000_0001010110001011_0111010100100011"; -- 0.0841592036203713
	pesos_i(2944) := b"0000000000000000_0000000000000000_0000010101100111_1110101000110111"; -- 0.021116865460270834
	pesos_i(2945) := b"1111111111111111_1111111111111111_1110100111000110_1101011100111111"; -- -0.08680968000982922
	pesos_i(2946) := b"0000000000000000_0000000000000000_0000001011101101_1000010111000000"; -- 0.011436805080461156
	pesos_i(2947) := b"1111111111111111_1111111111111111_1101100001000101_0010011000011011"; -- -0.1551948723795792
	pesos_i(2948) := b"1111111111111111_1111111111111111_1101100010101011_0011001111000010"; -- -0.1536376619910416
	pesos_i(2949) := b"1111111111111111_1111111111111111_1101110110110111_1111011001010001"; -- -0.13391170988841875
	pesos_i(2950) := b"0000000000000000_0000000000000000_0000000111010001_0111101011110001"; -- 0.007102664732728659
	pesos_i(2951) := b"1111111111111111_1111111111111111_1110111110001000_1010000101000010"; -- -0.06432144287739776
	pesos_i(2952) := b"1111111111111111_1111111111111111_1111001011100111_1000011010111100"; -- -0.05115468887620539
	pesos_i(2953) := b"1111111111111111_1111111111111111_1101011100010111_1001000010111110"; -- -0.15979667045601045
	pesos_i(2954) := b"0000000000000000_0000000000000000_0000111011001110_1101011001101100"; -- 0.05784359107291006
	pesos_i(2955) := b"1111111111111111_1111111111111111_1101110000010001_1101001010100100"; -- -0.14035304549830674
	pesos_i(2956) := b"1111111111111111_1111111111111111_1111011100000100_0100100000010010"; -- -0.035090919003668675
	pesos_i(2957) := b"1111111111111111_1111111111111111_1101101010111110_1011101110101001"; -- -0.14552714457424334
	pesos_i(2958) := b"1111111111111111_1111111111111111_1111011111110001_1110010111111111"; -- -0.031465172975507626
	pesos_i(2959) := b"0000000000000000_0000000000000000_0010000101011011_1011011000101011"; -- 0.13030565776497283
	pesos_i(2960) := b"1111111111111111_1111111111111111_1111000100101110_1100111001111000"; -- -0.05787953919755305
	pesos_i(2961) := b"0000000000000000_0000000000000000_0000100011110111_1000101001000110"; -- 0.03502716274736543
	pesos_i(2962) := b"0000000000000000_0000000000000000_0010010000001001_1000000010101111"; -- 0.14076999922422348
	pesos_i(2963) := b"0000000000000000_0000000000000000_0001101101010100_1000010001000111"; -- 0.10675837267637767
	pesos_i(2964) := b"1111111111111111_1111111111111111_1111110101110110_1110110110111110"; -- -0.009904042302942886
	pesos_i(2965) := b"1111111111111111_1111111111111111_1110000000111010_1100111110101100"; -- -0.12410261193787449
	pesos_i(2966) := b"0000000000000000_0000000000000000_0001010100001011_1100101110001111"; -- 0.0822112297212559
	pesos_i(2967) := b"0000000000000000_0000000000000000_0001000010011110_1100111101100000"; -- 0.064923249254029
	pesos_i(2968) := b"0000000000000000_0000000000000000_0000010101100001_1000101011010010"; -- 0.0210196269681001
	pesos_i(2969) := b"1111111111111111_1111111111111111_1110100011000001_0101110000010101"; -- -0.09079956511673733
	pesos_i(2970) := b"1111111111111111_1111111111111111_1110100001111101_1101111101011101"; -- -0.09182933783374729
	pesos_i(2971) := b"0000000000000000_0000000000000000_0001111011101101_1001000111001001"; -- 0.1208125225355319
	pesos_i(2972) := b"0000000000000000_0000000000000000_0010101101011000_0101010101100110"; -- 0.16931661366828546
	pesos_i(2973) := b"0000000000000000_0000000000000000_0000100001001101_0101011001000010"; -- 0.032430068044417476
	pesos_i(2974) := b"1111111111111111_1111111111111111_1111010111000010_0000001101000110"; -- -0.040008349719394556
	pesos_i(2975) := b"0000000000000000_0000000000000000_0001111110100101_1011011101000000"; -- 0.12362237283851549
	pesos_i(2976) := b"1111111111111111_1111111111111111_1111011110110001_1101010110100100"; -- -0.03244271030567772
	pesos_i(2977) := b"0000000000000000_0000000000000000_0001110001011000_1111110010010000"; -- 0.11073282726419685
	pesos_i(2978) := b"1111111111111111_1111111111111111_1101110001011010_1110010010011000"; -- -0.13923808384429578
	pesos_i(2979) := b"1111111111111111_1111111111111111_1110110001111010_1111011101011101"; -- -0.0762486837242792
	pesos_i(2980) := b"1111111111111111_1111111111111111_1111000110101000_1101110110000111"; -- -0.05601706941803956
	pesos_i(2981) := b"1111111111111111_1111111111111111_1111100001100111_1111101011001000"; -- -0.02966339692022852
	pesos_i(2982) := b"0000000000000000_0000000000000000_0000011100110110_1001011010001111"; -- 0.028176698715215772
	pesos_i(2983) := b"1111111111111111_1111111111111111_1110101101001111_1001111010010000"; -- -0.08081635450255989
	pesos_i(2984) := b"1111111111111111_1111111111111111_1111101001001101_1010110001010100"; -- -0.022252301729900115
	pesos_i(2985) := b"0000000000000000_0000000000000000_0010011111100001_1000000101000101"; -- 0.15578468261410802
	pesos_i(2986) := b"0000000000000000_0000000000000000_0000100101001111_0110010001100101"; -- 0.03636767837071499
	pesos_i(2987) := b"1111111111111111_1111111111111111_1110010101001100_1101110100011111"; -- -0.10429590224350656
	pesos_i(2988) := b"1111111111111111_1111111111111111_1110011111100010_0100100110011010"; -- -0.0942033766345803
	pesos_i(2989) := b"0000000000000000_0000000000000000_0000100100010111_0011011110111010"; -- 0.03551052364217394
	pesos_i(2990) := b"0000000000000000_0000000000000000_0001110100000111_1001101100100110"; -- 0.11339730909009396
	pesos_i(2991) := b"1111111111111111_1111111111111111_1110101001010001_0011110100011001"; -- -0.08469789635854565
	pesos_i(2992) := b"1111111111111111_1111111111111111_1110110100101111_1110001110000101"; -- -0.07348802566183436
	pesos_i(2993) := b"1111111111111111_1111111111111111_1111010010100011_1110001111001011"; -- -0.044374239901595905
	pesos_i(2994) := b"0000000000000000_0000000000000000_0000101011011001_1110010110100110"; -- 0.042387345347729595
	pesos_i(2995) := b"0000000000000000_0000000000000000_0000000111011111_0111010010111111"; -- 0.00731591845795657
	pesos_i(2996) := b"1111111111111111_1111111111111111_1111110101011001_1101000001100101"; -- -0.010348296509224988
	pesos_i(2997) := b"0000000000000000_0000000000000000_0010100110010101_0110100111101101"; -- 0.16243612333089852
	pesos_i(2998) := b"0000000000000000_0000000000000000_0010100101100110_0100010000010110"; -- 0.16171670468030477
	pesos_i(2999) := b"0000000000000000_0000000000000000_0001110001100101_1000000110001011"; -- 0.11092385917084682
	pesos_i(3000) := b"0000000000000000_0000000000000000_0001110000000010_0010110000001100"; -- 0.10940814302161492
	pesos_i(3001) := b"1111111111111111_1111111111111111_1101010001010011_1010101001100110"; -- -0.17059836408064738
	pesos_i(3002) := b"1111111111111111_1111111111111111_1101110111000011_0010011101001000"; -- -0.13374094482513685
	pesos_i(3003) := b"1111111111111111_1111111111111111_1110001110010111_1101001001000011"; -- -0.11096464031871499
	pesos_i(3004) := b"0000000000000000_0000000000000000_0001011101010010_0100101100111100"; -- 0.09109945492792242
	pesos_i(3005) := b"0000000000000000_0000000000000000_0000111101011010_0000110001011000"; -- 0.0599677766556016
	pesos_i(3006) := b"1111111111111111_1111111111111111_1110000011001000_0101110111111100"; -- -0.12194264037578151
	pesos_i(3007) := b"0000000000000000_0000000000000000_0000111110001101_0010011110010111"; -- 0.06074759901551824
	pesos_i(3008) := b"0000000000000000_0000000000000000_0010100101101000_1101011011001011"; -- 0.16175596670091827
	pesos_i(3009) := b"1111111111111111_1111111111111111_1111010111001010_1111110010001111"; -- -0.0398714210223332
	pesos_i(3010) := b"1111111111111111_1111111111111111_1110011010101100_0100101001101011"; -- -0.09893355271846956
	pesos_i(3011) := b"1111111111111111_1111111111111111_1110010100000101_1001101111000110"; -- -0.10538317126259537
	pesos_i(3012) := b"0000000000000000_0000000000000000_0000111100000001_1010011110111011"; -- 0.05861900630490102
	pesos_i(3013) := b"0000000000000000_0000000000000000_0000100100001010_0000010110111110"; -- 0.035309180056743154
	pesos_i(3014) := b"0000000000000000_0000000000000000_0000110111011100_1111100000001011"; -- 0.05415296819169083
	pesos_i(3015) := b"1111111111111111_1111111111111111_1110101101010111_1011101111010101"; -- -0.08069253971762638
	pesos_i(3016) := b"0000000000000000_0000000000000000_0010010000111101_0100110000000011"; -- 0.14156031668678118
	pesos_i(3017) := b"0000000000000000_0000000000000000_0000010101001011_0100111111111100"; -- 0.0206804265688376
	pesos_i(3018) := b"1111111111111111_1111111111111111_1111011000101000_1110111100001010"; -- -0.038437900701296504
	pesos_i(3019) := b"0000000000000000_0000000000000000_0001000001100000_0101100101011010"; -- 0.06397016952004858
	pesos_i(3020) := b"0000000000000000_0000000000000000_0001110111000110_1010101111110101"; -- 0.11631273972786133
	pesos_i(3021) := b"0000000000000000_0000000000000000_0001110001000111_1111101110011111"; -- 0.11047337176045613
	pesos_i(3022) := b"1111111111111111_1111111111111111_1101010101001001_0110100000111111"; -- -0.16684864488512247
	pesos_i(3023) := b"0000000000000000_0000000000000000_0001011000111111_1111111101000100"; -- 0.08691401871939203
	pesos_i(3024) := b"0000000000000000_0000000000000000_0000111101110101_0000100101100111"; -- 0.06037958881377459
	pesos_i(3025) := b"1111111111111111_1111111111111111_1101111011001001_0110011101000100"; -- -0.12973932823861092
	pesos_i(3026) := b"0000000000000000_0000000000000000_0010010101101010_0011011101110110"; -- 0.14615198746494404
	pesos_i(3027) := b"1111111111111111_1111111111111111_1111010111111001_1010111110110001"; -- -0.03915883943331468
	pesos_i(3028) := b"0000000000000000_0000000000000000_0010010111001101_0000000011110110"; -- 0.14765935899250007
	pesos_i(3029) := b"1111111111111111_1111111111111111_1111000000111111_0011111001010101"; -- -0.061534980993046384
	pesos_i(3030) := b"0000000000000000_0000000000000000_0000111001011110_1100011001110101"; -- 0.05613365519161838
	pesos_i(3031) := b"0000000000000000_0000000000000000_0001100101101010_0100011101000000"; -- 0.099277928540524
	pesos_i(3032) := b"0000000000000000_0000000000000000_0000010110110001_1110101011111101"; -- 0.022246062159021956
	pesos_i(3033) := b"1111111111111111_1111111111111111_1110100110011001_1100111111100010"; -- -0.0874967644488971
	pesos_i(3034) := b"0000000000000000_0000000000000000_0010100011001110_1001000011000011"; -- 0.15940193897983948
	pesos_i(3035) := b"1111111111111111_1111111111111111_1111100001111011_0110101100110100"; -- -0.029366779073910453
	pesos_i(3036) := b"1111111111111111_1111111111111111_1101100010000010_0000100110010111"; -- -0.1542657857934662
	pesos_i(3037) := b"0000000000000000_0000000000000000_0000110001011001_1010001000010110"; -- 0.048242693265323676
	pesos_i(3038) := b"0000000000000000_0000000000000000_0010011111010101_0100110010100010"; -- 0.15559843982556967
	pesos_i(3039) := b"1111111111111111_1111111111111111_1101100011110001_1110010010001101"; -- -0.15255900913096426
	pesos_i(3040) := b"0000000000000000_0000000000000000_0010101101000100_1111000011001100"; -- 0.1690207003782879
	pesos_i(3041) := b"0000000000000000_0000000000000000_0001000110101111_1100111111000011"; -- 0.06908892153512525
	pesos_i(3042) := b"0000000000000000_0000000000000000_0010001000110010_1000101001001000"; -- 0.13358368161620063
	pesos_i(3043) := b"1111111111111111_1111111111111111_1101101011101001_1101010011010100"; -- -0.14486951669624776
	pesos_i(3044) := b"0000000000000000_0000000000000000_0010101011111011_0110000100011010"; -- 0.16789824385216515
	pesos_i(3045) := b"1111111111111111_1111111111111111_1101011100001100_0001010111101011"; -- -0.15997183803797843
	pesos_i(3046) := b"0000000000000000_0000000000000000_0010011110111101_0011001110011100"; -- 0.1552307373837353
	pesos_i(3047) := b"1111111111111111_1111111111111111_1110011101001110_0000110011011101"; -- -0.09646529772361638
	pesos_i(3048) := b"0000000000000000_0000000000000000_0000111001110010_1000001100101010"; -- 0.056434819998487346
	pesos_i(3049) := b"0000000000000000_0000000000000000_0010011001101000_0100111100111111"; -- 0.15002913751588845
	pesos_i(3050) := b"0000000000000000_0000000000000000_0010100101010000_0000101000101010"; -- 0.16137755900912887
	pesos_i(3051) := b"0000000000000000_0000000000000000_0001000001011111_1111110100010110"; -- 0.0639646701083261
	pesos_i(3052) := b"0000000000000000_0000000000000000_0001110111011111_0010011011101010"; -- 0.11668627937444398
	pesos_i(3053) := b"1111111111111111_1111111111111111_1101101000000000_0000111010011100"; -- -0.14843662912941277
	pesos_i(3054) := b"1111111111111111_1111111111111111_1110011100101111_0101010011101011"; -- -0.09693402536568034
	pesos_i(3055) := b"0000000000000000_0000000000000000_0010100011111001_1101000010000100"; -- 0.16006186696722044
	pesos_i(3056) := b"1111111111111111_1111111111111111_1101010111110101_0111110000110001"; -- -0.16422294431738038
	pesos_i(3057) := b"1111111111111111_1111111111111111_1101110011011001_0001111111100100"; -- -0.13731194199012584
	pesos_i(3058) := b"1111111111111111_1111111111111111_1101011101001111_1110101000010011"; -- -0.15893685378882302
	pesos_i(3059) := b"1111111111111111_1111111111111111_1101011001110011_1101110110101100"; -- -0.16229452660289914
	pesos_i(3060) := b"1111111111111111_1111111111111111_1110101011111010_0000000010110001"; -- -0.0821227614569174
	pesos_i(3061) := b"1111111111111111_1111111111111111_1101101110011110_0000110010100011"; -- -0.14211960802562965
	pesos_i(3062) := b"0000000000000000_0000000000000000_0010001001000000_1010101111101101"; -- 0.1337993100152476
	pesos_i(3063) := b"0000000000000000_0000000000000000_0001011011010101_0011011111010110"; -- 0.0891909500435461
	pesos_i(3064) := b"1111111111111111_1111111111111111_1101010010100101_0100111111011010"; -- -0.16935254031299224
	pesos_i(3065) := b"1111111111111111_1111111111111111_1111010011111010_0000011110010010"; -- -0.04305985146558818
	pesos_i(3066) := b"0000000000000000_0000000000000000_0010001010010101_1100001101001110"; -- 0.1350977007288755
	pesos_i(3067) := b"1111111111111111_1111111111111111_1101111000011100_1011011100010001"; -- -0.13237434222414843
	pesos_i(3068) := b"1111111111111111_1111111111111111_1111011110100110_0001010101011010"; -- -0.03262201832519031
	pesos_i(3069) := b"0000000000000000_0000000000000000_0010010011110001_0101001110010110"; -- 0.14430735030010153
	pesos_i(3070) := b"1111111111111111_1111111111111111_1110001101010000_1101110011001000"; -- -0.11204738726848688
	pesos_i(3071) := b"0000000000000000_0000000000000000_0001000111000010_0010000001100111"; -- 0.06936838639444068
	pesos_i(3072) := b"0000000000000000_0000000000000000_0000111001011110_0011100001110011"; -- 0.05612519075860714
	pesos_i(3073) := b"0000000000000000_0000000000000000_0000111110101010_1011001000010000"; -- 0.06119835739927887
	pesos_i(3074) := b"0000000000000000_0000000000000000_0000011010010101_0111101100100100"; -- 0.025718399308340193
	pesos_i(3075) := b"0000000000000000_0000000000000000_0001101110010010_1010010000101010"; -- 0.1077063180975087
	pesos_i(3076) := b"0000000000000000_0000000000000000_0000110011001001_1101001001000000"; -- 0.049954548491480906
	pesos_i(3077) := b"0000000000000000_0000000000000000_0000010011100100_1010110010010101"; -- 0.019114290511490238
	pesos_i(3078) := b"0000000000000000_0000000000000000_0010010100100011_0001111000001011"; -- 0.14506709831957454
	pesos_i(3079) := b"1111111111111111_1111111111111111_1110101111000100_0000010100000111"; -- -0.07904022778452448
	pesos_i(3080) := b"0000000000000000_0000000000000000_0011110001001100_1000111000100001"; -- 0.2355431393993759
	pesos_i(3081) := b"1111111111111111_1111111111111111_1101111100100111_0111100101111000"; -- -0.12830391704982805
	pesos_i(3082) := b"1111111111111111_1111111111111111_1110110000001011_0001110011001011"; -- -0.07795543715490215
	pesos_i(3083) := b"0000000000000000_0000000000000000_0000111111000100_1000001110111001"; -- 0.06159232395266457
	pesos_i(3084) := b"1111111111111111_1111111111111111_1111110011000000_0011010000100011"; -- -0.012692204894650142
	pesos_i(3085) := b"1111111111111111_1111111111111111_1101011011100001_0111000110110011"; -- -0.16062249553834518
	pesos_i(3086) := b"1111111111111111_1111111111111111_1111010001000110_0110000101111000"; -- -0.04580107510752149
	pesos_i(3087) := b"0000000000000000_0000000000000000_0001000011010001_1011001011001011"; -- 0.06569974383808565
	pesos_i(3088) := b"1111111111111111_1111111111111111_1101011000011000_0000001000100001"; -- -0.16369616225367234
	pesos_i(3089) := b"1111111111111111_1111111111111111_1110110010000111_0011011100010111"; -- -0.07606177993708531
	pesos_i(3090) := b"1111111111111111_1111111111111111_1111110110010011_0000110000110011"; -- -0.0094749809697005
	pesos_i(3091) := b"0000000000000000_0000000000000000_0000110111010111_1100100001101111"; -- 0.054073836499542595
	pesos_i(3092) := b"0000000000000000_0000000000000000_0000111101111111_1110001100010110"; -- 0.06054515165546654
	pesos_i(3093) := b"0000000000000000_0000000000000000_0000011001101111_1111010011101101"; -- 0.025145824283178197
	pesos_i(3094) := b"1111111111111111_1111111111111111_1101100001100100_1011110111110101"; -- -0.15471279880319372
	pesos_i(3095) := b"1111111111111111_1111111111111111_1101000000100100_0011101000100010"; -- -0.18694721861349317
	pesos_i(3096) := b"1111111111111111_1111111111111111_1110000001111000_1000100001111010"; -- -0.12316081063521728
	pesos_i(3097) := b"1111111111111111_1111111111111111_1110001000001101_1011101011001111"; -- -0.11697800101590085
	pesos_i(3098) := b"0000000000000000_0000000000000000_0001110101010100_1110110100111100"; -- 0.11457712862954317
	pesos_i(3099) := b"1111111111111111_1111111111111111_1111010010100101_0111111000010100"; -- -0.044349784928192956
	pesos_i(3100) := b"0000000000000000_0000000000000000_0001000111110111_1011111100110110"; -- 0.070186568036171
	pesos_i(3101) := b"0000000000000000_0000000000000000_0001000000011001_0111111100010111"; -- 0.0628890448929572
	pesos_i(3102) := b"0000000000000000_0000000000000000_0001110001100110_1100111100011001"; -- 0.11094374040002622
	pesos_i(3103) := b"0000000000000000_0000000000000000_0000111100111010_1110001110010001"; -- 0.059492323869966834
	pesos_i(3104) := b"1111111111111111_1111111111111111_1111010010001011_0110101011000000"; -- -0.044747665623801364
	pesos_i(3105) := b"1111111111111111_1111111111111111_1110010000100010_0010010101011100"; -- -0.1088539744579037
	pesos_i(3106) := b"0000000000000000_0000000000000000_0010100010100010_1100000000110000"; -- 0.15873337911489502
	pesos_i(3107) := b"1111111111111111_1111111111111111_1111010011011101_1010000111010000"; -- -0.043493162766431864
	pesos_i(3108) := b"0000000000000000_0000000000000000_0001001110010000_1010000011100000"; -- 0.07642560459365302
	pesos_i(3109) := b"1111111111111111_1111111111111111_1111001001011000_1100101111011101"; -- -0.05333257532481639
	pesos_i(3110) := b"0000000000000000_0000000000000000_0001110100100000_1011111100110001"; -- 0.11378092725530937
	pesos_i(3111) := b"1111111111111111_1111111111111111_1111111111110011_1101110011001001"; -- -0.0001852045180342765
	pesos_i(3112) := b"1111111111111111_1111111111111111_1101110011100111_0001000000101111"; -- -0.13709925508268384
	pesos_i(3113) := b"1111111111111111_1111111111111111_1101110011111011_1010101010011010"; -- -0.136784875335552
	pesos_i(3114) := b"0000000000000000_0000000000000000_0010010001010111_0000000000000000"; -- 0.14195251471609388
	pesos_i(3115) := b"0000000000000000_0000000000000000_0001110011000111_1111001100101111"; -- 0.11242599393961464
	pesos_i(3116) := b"1111111111111111_1111111111111111_1111100010101111_0111010111110000"; -- -0.028572682376060157
	pesos_i(3117) := b"0000000000000000_0000000000000000_0010101010100101_0011101110001001"; -- 0.1665837488100091
	pesos_i(3118) := b"1111111111111111_1111111111111111_1111110101110000_0110110010110101"; -- -0.010003286065906968
	pesos_i(3119) := b"0000000000000000_0000000000000000_0011000111110110_0111011111000110"; -- 0.1951670511694507
	pesos_i(3120) := b"1111111111111111_1111111111111111_1110101111101010_1101101100000101"; -- -0.07844763867151311
	pesos_i(3121) := b"0000000000000000_0000000000000000_0001101101100101_1010011101001111"; -- 0.10701986005424613
	pesos_i(3122) := b"0000000000000000_0000000000000000_0000101000101111_0100110100010101"; -- 0.039784257616024526
	pesos_i(3123) := b"1111111111111111_1111111111111111_1111010001010100_1111101011010000"; -- -0.045578312030366865
	pesos_i(3124) := b"0000000000000000_0000000000000000_0010010111001101_0011111100010001"; -- 0.14766306091901435
	pesos_i(3125) := b"0000000000000000_0000000000000000_0001000100110100_1110001111111101"; -- 0.06721329624055135
	pesos_i(3126) := b"0000000000000000_0000000000000000_0001000010010100_1010000000100011"; -- 0.06476784566655429
	pesos_i(3127) := b"0000000000000000_0000000000000000_0000100011001100_1111111000110101"; -- 0.03437794487487463
	pesos_i(3128) := b"0000000000000000_0000000000000000_0010011001001001_0001101010001110"; -- 0.14955297441860185
	pesos_i(3129) := b"0000000000000000_0000000000000000_0001101100010101_1011111010000111"; -- 0.10580054080005477
	pesos_i(3130) := b"0000000000000000_0000000000000000_0000111111000111_0011011110010111"; -- 0.061633562446320865
	pesos_i(3131) := b"0000000000000000_0000000000000000_0000111111100010_0000101111110101"; -- 0.06204294898147809
	pesos_i(3132) := b"0000000000000000_0000000000000000_0000000000001111_1110011010100101"; -- 0.0002426292767935278
	pesos_i(3133) := b"1111111111111111_1111111111111111_1111001011110010_0001000101111010"; -- -0.05099383125920612
	pesos_i(3134) := b"0000000000000000_0000000000000000_0010001110011110_1000001110110100"; -- 0.13913748874122736
	pesos_i(3135) := b"1111111111111111_1111111111111111_1111011100111001_0111001011110011"; -- -0.03427964755254146
	pesos_i(3136) := b"1111111111111111_1111111111111111_1110101100110011_0011110000100101"; -- -0.08124946691832971
	pesos_i(3137) := b"1111111111111111_1111111111111111_1110011101000011_1000100101010001"; -- -0.09662572636558499
	pesos_i(3138) := b"1111111111111111_1111111111111111_1101101100110001_1010010111111010"; -- -0.14377367638042804
	pesos_i(3139) := b"0000000000000000_0000000000000000_0001001111010000_0001000010011111"; -- 0.07739356893030841
	pesos_i(3140) := b"0000000000000000_0000000000000000_0001100111001000_0001101100000000"; -- 0.10070961717426226
	pesos_i(3141) := b"1111111111111111_1111111111111111_1111110010111100_0000001101110110"; -- -0.012756141286048244
	pesos_i(3142) := b"1111111111111111_1111111111111111_1110101100001001_0001001001101110"; -- -0.08189282243485141
	pesos_i(3143) := b"0000000000000000_0000000000000000_0010001101111110_1100010110110010"; -- 0.1386531408995691
	pesos_i(3144) := b"1111111111111111_1111111111111111_1110000011010100_0010001010000001"; -- -0.12176308007321959
	pesos_i(3145) := b"0000000000000000_0000000000000000_0001101000100100_1010000101000001"; -- 0.10212142780173854
	pesos_i(3146) := b"1111111111111111_1111111111111111_1101110001010100_0000000110001000"; -- -0.13934317056338832
	pesos_i(3147) := b"0000000000000000_0000000000000000_0001111100111110_1101111000010001"; -- 0.12205303117399888
	pesos_i(3148) := b"1111111111111111_1111111111111111_1110111111110011_0100110001010010"; -- -0.06269381528305487
	pesos_i(3149) := b"0000000000000000_0000000000000000_0000101010111000_1011001101010010"; -- 0.04188080550423498
	pesos_i(3150) := b"1111111111111111_1111111111111111_1110001001001011_0111001100111100"; -- -0.11603622234995957
	pesos_i(3151) := b"1111111111111111_1111111111111111_1111101101011100_0010100010010110"; -- -0.01812502238484413
	pesos_i(3152) := b"0000000000000000_0000000000000000_0001111010000000_1011001110000001"; -- 0.1191513242482293
	pesos_i(3153) := b"1111111111111111_1111111111111111_1101110000101100_0000010111111000"; -- -0.13995325755492294
	pesos_i(3154) := b"1111111111111111_1111111111111111_1101110000000100_1001111110010100"; -- -0.14055445332042532
	pesos_i(3155) := b"0000000000000000_0000000000000000_0000000101101100_0001000101000101"; -- 0.005555228589754998
	pesos_i(3156) := b"1111111111111111_1111111111111111_1110011001101111_1111000001000001"; -- -0.0998544541035833
	pesos_i(3157) := b"0000000000000000_0000000000000000_0000100001000100_1011101010001110"; -- 0.032298717114613476
	pesos_i(3158) := b"0000000000000000_0000000000000000_0001001000110001_1000100010101000"; -- 0.07106832610185725
	pesos_i(3159) := b"0000000000000000_0000000000000000_0010001001010010_0111000000001100"; -- 0.1340703993325307
	pesos_i(3160) := b"1111111111111111_1111111111111111_1111001011011101_0011100001000101"; -- -0.05131195359034589
	pesos_i(3161) := b"0000000000000000_0000000000000000_0001001010101011_1011001110011000"; -- 0.07293245761833922
	pesos_i(3162) := b"1111111111111111_1111111111111111_1110001111000011_0000000000001111"; -- -0.11030578273376569
	pesos_i(3163) := b"0000000000000000_0000000000000000_0010101110111000_1011001010111000"; -- 0.1707870196386528
	pesos_i(3164) := b"1111111111111111_1111111111111111_1111100001001010_0100110110000010"; -- -0.030116229674757435
	pesos_i(3165) := b"0000000000000000_0000000000000000_0000011011110011_0110000001001111"; -- 0.027151126186328388
	pesos_i(3166) := b"1111111111111111_1111111111111111_1110100111010111_1001110000011110"; -- -0.0865538050188601
	pesos_i(3167) := b"1111111111111111_1111111111111111_1101011101100010_0010101010100001"; -- -0.15865834790720723
	pesos_i(3168) := b"0000000000000000_0000000000000000_0010101000111110_1101101101001011"; -- 0.1650216158895614
	pesos_i(3169) := b"0000000000000000_0000000000000000_0000100011100111_1011001010000110"; -- 0.03478542102906599
	pesos_i(3170) := b"0000000000000000_0000000000000000_0000001110110001_1011100100111010"; -- 0.01443059612443983
	pesos_i(3171) := b"1111111111111111_1111111111111111_1101110001000111_0000100110010010"; -- -0.13954105542603754
	pesos_i(3172) := b"1111111111111111_1111111111111111_1101110110001111_0000001011100101"; -- -0.13453657068411917
	pesos_i(3173) := b"0000000000000000_0000000000000000_0010100001001011_0111001111000101"; -- 0.15740130964491222
	pesos_i(3174) := b"0000000000000000_0000000000000000_0000100011010011_0001010101011000"; -- 0.03447087678330152
	pesos_i(3175) := b"0000000000000000_0000000000000000_0010100110110010_1011111000101100"; -- 0.16288364963410276
	pesos_i(3176) := b"0000000000000000_0000000000000000_0000010010011100_0001011011010011"; -- 0.018006731536991227
	pesos_i(3177) := b"1111111111111111_1111111111111111_1110110101110110_1010011000100011"; -- -0.07240831038506149
	pesos_i(3178) := b"1111111111111111_1111111111111111_1110110101100011_0111011100100000"; -- -0.07270102947183313
	pesos_i(3179) := b"0000000000000000_0000000000000000_0000011000111001_1111001100011010"; -- 0.02432174107323204
	pesos_i(3180) := b"0000000000000000_0000000000000000_0010101100110011_0000001001000011"; -- 0.16874708304179967
	pesos_i(3181) := b"1111111111111111_1111111111111111_1101010010101010_1101001001001001"; -- -0.1692684719491147
	pesos_i(3182) := b"1111111111111111_1111111111111111_1111110000101110_1010100011110111"; -- -0.014913024541603556
	pesos_i(3183) := b"0000000000000000_0000000000000000_0001110101011100_1111001111001011"; -- 0.11469958988276409
	pesos_i(3184) := b"0000000000000000_0000000000000000_0010010011100010_0011001000011100"; -- 0.14407647310750335
	pesos_i(3185) := b"1111111111111111_1111111111111111_1110101010101010_0011111101001001"; -- -0.08333973385870037
	pesos_i(3186) := b"1111111111111111_1111111111111111_1111110101010000_0011111010011100"; -- -0.010494315042637684
	pesos_i(3187) := b"1111111111111111_1111111111111111_1101101010101100_0011111001001111"; -- -0.1458092744440658
	pesos_i(3188) := b"0000000000000000_0000000000000000_0000001110010001_0100001110111111"; -- 0.013935312432127527
	pesos_i(3189) := b"1111111111111111_1111111111111111_1101100111101001_0011000001100001"; -- -0.1487855685519856
	pesos_i(3190) := b"1111111111111111_1111111111111111_1101011000000110_1000011100101100"; -- -0.16396289043069753
	pesos_i(3191) := b"0000000000000000_0000000000000000_0000001101000000_1010010000011000"; -- 0.012705093207027113
	pesos_i(3192) := b"1111111111111111_1111111111111111_1111110001010111_1000100110100011"; -- -0.01428928147139008
	pesos_i(3193) := b"0000000000000000_0000000000000000_0000000010101000_1110001001010010"; -- 0.0025769664152591886
	pesos_i(3194) := b"0000000000000000_0000000000000000_0001101000000010_0110011011101010"; -- 0.10159915165845873
	pesos_i(3195) := b"1111111111111111_1111111111111111_1110001001100011_1011101101000100"; -- -0.11566571791323198
	pesos_i(3196) := b"1111111111111111_1111111111111111_1110110110010010_0110110110010111"; -- -0.07198443473254883
	pesos_i(3197) := b"0000000000000000_0000000000000000_0000010011110110_0101001111101011"; -- 0.01938366402274786
	pesos_i(3198) := b"1111111111111111_1111111111111111_1101101010111100_0010011000000110"; -- -0.14556658121362784
	pesos_i(3199) := b"1111111111111111_1111111111111111_1101111001000011_0101000010100101"; -- -0.13178535444672054
	pesos_i(3200) := b"0000000000000000_0000000000000000_0001001111000100_1101111110001011"; -- 0.07722279691949083
	pesos_i(3201) := b"0000000000000000_0000000000000000_0010000111001111_1101000000111101"; -- 0.13207723137405875
	pesos_i(3202) := b"1111111111111111_1111111111111111_1101001111010101_1000010110111110"; -- -0.17252315632158124
	pesos_i(3203) := b"0000000000000000_0000000000000000_0001000101011111_0011011001010100"; -- 0.06785907315200944
	pesos_i(3204) := b"0000000000000000_0000000000000000_0001111011000000_1110111011001111"; -- 0.12013142156315491
	pesos_i(3205) := b"1111111111111111_1111111111111111_1110001100000000_1001111000000000"; -- -0.11327183238031356
	pesos_i(3206) := b"0000000000000000_0000000000000000_0000011101100110_0101101110010100"; -- 0.028905605043695614
	pesos_i(3207) := b"0000000000000000_0000000000000000_0001010011100010_0010101000110010"; -- 0.08157600124945777
	pesos_i(3208) := b"1111111111111111_1111111111111111_1110100111110010_1000101110110101"; -- -0.08614279579729725
	pesos_i(3209) := b"0000000000000000_0000000000000000_0010110000111001_0111000111000011"; -- 0.17275153159072115
	pesos_i(3210) := b"1111111111111111_1111111111111111_1111010101111010_1011100111011011"; -- -0.04109610000143696
	pesos_i(3211) := b"1111111111111111_1111111111111111_1111000000111011_0110101110100010"; -- -0.06159331597042873
	pesos_i(3212) := b"0000000000000000_0000000000000000_0000000101011011_0111001001100110"; -- 0.005301618548502354
	pesos_i(3213) := b"0000000000000000_0000000000000000_0010100101110011_0111100101010001"; -- 0.1619182417027679
	pesos_i(3214) := b"1111111111111111_1111111111111111_1111101111010110_0010110111001101"; -- -0.01626313926408424
	pesos_i(3215) := b"1111111111111111_1111111111111111_1110101011000001_1111010100100011"; -- -0.08297794243130721
	pesos_i(3216) := b"0000000000000000_0000000000000000_0000111101010110_0011000011110010"; -- 0.05990892328375788
	pesos_i(3217) := b"1111111111111111_1111111111111111_1110100101000011_1010101011101010"; -- -0.08881122393031467
	pesos_i(3218) := b"0000000000000000_0000000000000000_0000100101111000_1110000111000101"; -- 0.037000761633543204
	pesos_i(3219) := b"0000000000000000_0000000000000000_0001010100100011_0010001111001100"; -- 0.08256744124871163
	pesos_i(3220) := b"0000000000000000_0000000000000000_0001000101100010_0110011111011001"; -- 0.06790780119405969
	pesos_i(3221) := b"0000000000000000_0000000000000000_0001001101010101_0100111101011100"; -- 0.07552047721434636
	pesos_i(3222) := b"0000000000000000_0000000000000000_0000001011000011_0011100000111000"; -- 0.010791314767644349
	pesos_i(3223) := b"1111111111111111_1111111111111111_1111111111000011_1111000111001110"; -- -0.0009163734111400854
	pesos_i(3224) := b"1111111111111111_1111111111111111_1110001000001110_0000111111001000"; -- -0.11697293637331067
	pesos_i(3225) := b"1111111111111111_1111111111111111_1110101100100100_1111010100001011"; -- -0.08146732781075282
	pesos_i(3226) := b"0000000000000000_0000000000000000_0000000011100010_0110011100111001"; -- 0.0034546387902900226
	pesos_i(3227) := b"1111111111111111_1111111111111111_1101100101011000_1010011110110001"; -- -0.15099098131070915
	pesos_i(3228) := b"1111111111111111_1111111111111111_1111001111100101_0100011001100001"; -- -0.04728279228036279
	pesos_i(3229) := b"1111111111111111_1111111111111111_1101101101111100_1110001111100001"; -- -0.14262557756134703
	pesos_i(3230) := b"0000000000000000_0000000000000000_0000000000001011_0100101000110001"; -- 0.00017226887137250716
	pesos_i(3231) := b"0000000000000000_0000000000000000_0010010101101010_1100111001000111"; -- 0.14616097671742798
	pesos_i(3232) := b"1111111111111111_1111111111111111_1101110110001111_1001010001011001"; -- -0.13452790104258228
	pesos_i(3233) := b"1111111111111111_1111111111111111_1101110110111010_1100100101100001"; -- -0.13386861204161274
	pesos_i(3234) := b"1111111111111111_1111111111111111_1110010011001100_0110110110101000"; -- -0.10625567106505797
	pesos_i(3235) := b"0000000000000000_0000000000000000_0010011010001101_1000111101111111"; -- 0.15059754236216186
	pesos_i(3236) := b"1111111111111111_1111111111111111_1101111111111000_0000001000010000"; -- -0.12512194733686607
	pesos_i(3237) := b"1111111111111111_1111111111111111_1110111110000000_0010100000000000"; -- -0.0644507407688704
	pesos_i(3238) := b"1111111111111111_1111111111111111_1110101111010011_1001011100101001"; -- -0.07880263572807304
	pesos_i(3239) := b"1111111111111111_1111111111111111_1111101001101100_1001010111110111"; -- -0.021780612068780514
	pesos_i(3240) := b"0000000000000000_0000000000000000_0010100111000110_0111000000000101"; -- 0.1631841671556669
	pesos_i(3241) := b"1111111111111111_1111111111111111_1101101000010011_1000011100011010"; -- -0.1481395304262995
	pesos_i(3242) := b"0000000000000000_0000000000000000_0000111011011011_1000101011101101"; -- 0.058037455384047365
	pesos_i(3243) := b"1111111111111111_1111111111111111_1111100011100111_1100010010111010"; -- -0.02771349384583129
	pesos_i(3244) := b"0000000000000000_0000000000000000_0010100000001101_1111001111001101"; -- 0.15646289581665881
	pesos_i(3245) := b"1111111111111111_1111111111111111_1111100101011010_1001100001101001"; -- -0.025961374732776394
	pesos_i(3246) := b"0000000000000000_0000000000000000_0000010001101110_0110100001110011"; -- 0.01730969239187655
	pesos_i(3247) := b"1111111111111111_1111111111111111_1110110111010010_1001011011010111"; -- -0.0710054135986585
	pesos_i(3248) := b"1111111111111111_1111111111111111_1110011011000101_1011101111001001"; -- -0.0985453257519628
	pesos_i(3249) := b"1111111111111111_1111111111111111_1111100001011001_0010111001011000"; -- -0.02988920551827337
	pesos_i(3250) := b"0000000000000000_0000000000000000_0001100101011100_0100011000100110"; -- 0.09906423969091967
	pesos_i(3251) := b"0000000000000000_0000000000000000_0000001101111111_1011110001001110"; -- 0.013667839996538157
	pesos_i(3252) := b"0000000000000000_0000000000000000_0001011011000110_1001011001001101"; -- 0.08896769875385525
	pesos_i(3253) := b"1111111111111111_1111111111111111_1110010000100100_1101011000100110"; -- -0.10881291945290056
	pesos_i(3254) := b"0000000000000000_0000000000000000_0000011000001000_0001011111001101"; -- 0.023560988900126617
	pesos_i(3255) := b"0000000000000000_0000000000000000_0000011111011100_1001111010101001"; -- 0.03071014055383223
	pesos_i(3256) := b"1111111111111111_1111111111111111_1111100001111010_0001010101000100"; -- -0.029387160187567873
	pesos_i(3257) := b"0000000000000000_0000000000000000_0010001100100100_1011011011111000"; -- 0.13727897221681393
	pesos_i(3258) := b"0000000000000000_0000000000000000_0010010101111001_1101111001010010"; -- 0.1463908148983424
	pesos_i(3259) := b"1111111111111111_1111111111111111_1111000010001001_0111010010000101"; -- -0.060402600829960205
	pesos_i(3260) := b"0000000000000000_0000000000000000_0001110100000001_1100110110001010"; -- 0.11330875996442802
	pesos_i(3261) := b"0000000000000000_0000000000000000_0001010100011011_1101001110010000"; -- 0.08245584744068207
	pesos_i(3262) := b"1111111111111111_1111111111111111_1111100111011000_0110000011010011"; -- -0.02404208029337651
	pesos_i(3263) := b"1111111111111111_1111111111111111_1111101010001000_0101100111011011"; -- -0.021356948948982178
	pesos_i(3264) := b"0000000000000000_0000000000000000_0001101000100100_0101111011100111"; -- 0.10211747292924686
	pesos_i(3265) := b"0000000000000000_0000000000000000_0010000000000000_1100010111010100"; -- 0.12501179138718269
	pesos_i(3266) := b"0000000000000000_0000000000000000_0001011010111101_0001111101000101"; -- 0.08882327496869795
	pesos_i(3267) := b"0000000000000000_0000000000000000_0010000100010101_0000100100001111"; -- 0.1292272243976547
	pesos_i(3268) := b"0000000000000000_0000000000000000_0001100110000111_0110001011101011"; -- 0.09972208253436983
	pesos_i(3269) := b"1111111111111111_1111111111111111_1111100110011100_0100010101000000"; -- -0.024959251179186622
	pesos_i(3270) := b"0000000000000000_0000000000000000_0000100001100100_0010110010101111"; -- 0.03277854217006012
	pesos_i(3271) := b"0000000000000000_0000000000000000_0010001001010010_1000110100000101"; -- 0.13407212616491115
	pesos_i(3272) := b"1111111111111111_1111111111111111_1101010010110011_0111100111100100"; -- -0.16913641151072628
	pesos_i(3273) := b"0000000000000000_0000000000000000_0001001001111100_1011110011101111"; -- 0.07221585115764484
	pesos_i(3274) := b"0000000000000000_0000000000000000_0000111111000010_0101111001101011"; -- 0.061559582812770096
	pesos_i(3275) := b"0000000000000000_0000000000000000_0001010010100001_0101101111101100"; -- 0.08058714400613391
	pesos_i(3276) := b"1111111111111111_1111111111111111_1111111000111001_1100111110110011"; -- -0.0069303692866310345
	pesos_i(3277) := b"0000000000000000_0000000000000000_0001011010011001_1111000001010101"; -- 0.08828641966453275
	pesos_i(3278) := b"0000000000000000_0000000000000000_0000000101000010_1101000110100101"; -- 0.004925825801091006
	pesos_i(3279) := b"0000000000000000_0000000000000000_0000000000110110_0111110100011000"; -- 0.0008314307641527041
	pesos_i(3280) := b"0000000000000000_0000000000000000_0010010000111101_0100110001111100"; -- 0.141560345020567
	pesos_i(3281) := b"0000000000000000_0000000000000000_0001011100100101_1011001101110010"; -- 0.09041902104875758
	pesos_i(3282) := b"0000000000000000_0000000000000000_0000000001010100_0001001101010101"; -- 0.0012828906571912494
	pesos_i(3283) := b"0000000000000000_0000000000000000_0001100011110001_0111000110101000"; -- 0.0974341425356891
	pesos_i(3284) := b"0000000000000000_0000000000000000_0001000111011110_1000001011100010"; -- 0.06980150251115462
	pesos_i(3285) := b"1111111111111111_1111111111111111_1110010000000110_0111100101111101"; -- -0.10927620605470229
	pesos_i(3286) := b"0000000000000000_0000000000000000_0001010010100110_1000111000111001"; -- 0.08066643610220775
	pesos_i(3287) := b"1111111111111111_1111111111111111_1111110100101000_0101011000110101"; -- -0.011103260126547393
	pesos_i(3288) := b"1111111111111111_1111111111111111_1101101110100100_1111111111001001"; -- -0.1420135625647553
	pesos_i(3289) := b"1111111111111111_1111111111111111_1111001001000111_0111101010110111"; -- -0.053596811494996816
	pesos_i(3290) := b"1111111111111111_1111111111111111_1101101000011110_0111100110100000"; -- -0.1479724868313568
	pesos_i(3291) := b"0000000000000000_0000000000000000_0001001001111010_1011001101011111"; -- 0.07218476356341699
	pesos_i(3292) := b"0000000000000000_0000000000000000_0000010011111111_1010110001101010"; -- 0.01952626794108162
	pesos_i(3293) := b"1111111111111111_1111111111111111_1111110000100010_1000010001100010"; -- -0.015098310454097005
	pesos_i(3294) := b"1111111111111111_1111111111111111_1110010111010000_1010001111100011"; -- -0.10228515356090905
	pesos_i(3295) := b"1111111111111111_1111111111111111_1111001100001001_1011010000100101"; -- -0.05063318338826561
	pesos_i(3296) := b"0000000000000000_0000000000000000_0000111110010011_0110001010010101"; -- 0.060842667993610544
	pesos_i(3297) := b"0000000000000000_0000000000000000_0000001011010011_1010000110100110"; -- 0.011041739407622727
	pesos_i(3298) := b"0000000000000000_0000000000000000_0000111101100001_1101001011011000"; -- 0.06008641984562249
	pesos_i(3299) := b"1111111111111111_1111111111111111_1110011010010010_0111011110110111"; -- -0.09932758116977089
	pesos_i(3300) := b"1111111111111111_1111111111111111_1110111100010011_1110000111000100"; -- -0.06610287641359894
	pesos_i(3301) := b"0000000000000000_0000000000000000_0001111011110101_1111110000010011"; -- 0.12094092822721593
	pesos_i(3302) := b"1111111111111111_1111111111111111_1101011010101100_1010001101010110"; -- -0.1614282527601927
	pesos_i(3303) := b"1111111111111111_1111111111111111_1110011100000001_0100101110111100"; -- -0.09763647710694189
	pesos_i(3304) := b"0000000000000000_0000000000000000_0000100001011110_0000111101101100"; -- 0.03268524545512691
	pesos_i(3305) := b"0000000000000000_0000000000000000_0001010010111100_0011101101100100"; -- 0.08099719221209149
	pesos_i(3306) := b"0000000000000000_0000000000000000_0000111011111111_0110010111111010"; -- 0.05858456951605638
	pesos_i(3307) := b"1111111111111111_1111111111111111_1110001011100101_0100100101111111"; -- -0.11368885648653623
	pesos_i(3308) := b"0000000000000000_0000000000000000_0000011001100010_1011100000100110"; -- 0.024943837478293897
	pesos_i(3309) := b"0000000000000000_0000000000000000_0001001011110111_1000000011011111"; -- 0.07408910232812123
	pesos_i(3310) := b"1111111111111111_1111111111111111_1101111011110100_0110100111010110"; -- -0.12908304724651776
	pesos_i(3311) := b"1111111111111111_1111111111111111_1111111010000111_1110101110000001"; -- -0.005738526276962097
	pesos_i(3312) := b"1111111111111111_1111111111111111_1101110001010011_1110111110000110"; -- -0.1393442438361738
	pesos_i(3313) := b"0000000000000000_0000000000000000_0000011110010110_0110010010001001"; -- 0.029638560639757096
	pesos_i(3314) := b"1111111111111111_1111111111111111_1111111111111101_1111011110110011"; -- -3.101227339270833e-05
	pesos_i(3315) := b"0000000000000000_0000000000000000_0001001100101111_0101101001100101"; -- 0.07494130111197075
	pesos_i(3316) := b"0000000000000000_0000000000000000_0001110110011101_0011111111100010"; -- 0.115680687703165
	pesos_i(3317) := b"1111111111111111_1111111111111111_1111010111111111_0000111111010011"; -- -0.039076815670211464
	pesos_i(3318) := b"1111111111111111_1111111111111111_1111100101011111_0011110100110101"; -- -0.025890516703009375
	pesos_i(3319) := b"0000000000000000_0000000000000000_0001110100101110_1110000110110100"; -- 0.11399660724144912
	pesos_i(3320) := b"0000000000000000_0000000000000000_0000011101010111_1101110001011000"; -- 0.02868439822051519
	pesos_i(3321) := b"1111111111111111_1111111111111111_1101111010100101_0100111001110010"; -- -0.1302901241486645
	pesos_i(3322) := b"0000000000000000_0000000000000000_0010010000000011_1110000011110111"; -- 0.1406841852631843
	pesos_i(3323) := b"1111111111111111_1111111111111111_1101101011100111_1000101111000000"; -- -0.14490439004843017
	pesos_i(3324) := b"1111111111111111_1111111111111111_1110110011101111_1101110101000001"; -- -0.0744649617356373
	pesos_i(3325) := b"0000000000000000_0000000000000000_0001011110110101_1100111111111010"; -- 0.09261798722771113
	pesos_i(3326) := b"1111111111111111_1111111111111111_1111110010011111_0011111011110111"; -- -0.013195099454396382
	pesos_i(3327) := b"1111111111111111_1111111111111111_1100111100010110_1111101010010010"; -- -0.19105562149207164
	pesos_i(3328) := b"1111111111111111_1111111111111111_1110101001111010_1011010000111110"; -- -0.08406518444268375
	pesos_i(3329) := b"1111111111111111_1111111111111111_1110010000010110_0110010100101110"; -- -0.10903327593419103
	pesos_i(3330) := b"0000000000000000_0000000000000000_0010110110001011_1001000111000101"; -- 0.17791091029330952
	pesos_i(3331) := b"1111111111111111_1111111111111111_1110000011010100_1100101101000000"; -- -0.12175302210048133
	pesos_i(3332) := b"0000000000000000_0000000000000000_0001101100111010_0011111111001101"; -- 0.1063575624789638
	pesos_i(3333) := b"0000000000000000_0000000000000000_0001100111011101_0101001100111001"; -- 0.10103340282549894
	pesos_i(3334) := b"0000000000000000_0000000000000000_0000000000101100_1011100101100110"; -- 0.0006824373176688236
	pesos_i(3335) := b"1111111111111111_1111111111111111_1101100010010110_1101011011000011"; -- -0.15394838089356305
	pesos_i(3336) := b"0000000000000000_0000000000000000_0000101100011101_1100000100100110"; -- 0.04342276739889237
	pesos_i(3337) := b"1111111111111111_1111111111111111_1101010100010101_0001101111111011"; -- -0.16764664774782695
	pesos_i(3338) := b"1111111111111111_1111111111111111_1101100011010010_1001010111001010"; -- -0.15303672612626879
	pesos_i(3339) := b"1111111111111111_1111111111111111_1110110010010101_1011011011010011"; -- -0.07584054334263055
	pesos_i(3340) := b"1111111111111111_1111111111111111_1101101111010110_0001010100001110"; -- -0.14126461419301847
	pesos_i(3341) := b"1111111111111111_1111111111111111_1111101100110101_1011010110110011"; -- -0.018711704049220353
	pesos_i(3342) := b"0000000000000000_0000000000000000_0010001000011101_0011100000011010"; -- 0.13325834876183007
	pesos_i(3343) := b"1111111111111111_1111111111111111_1110010011010101_0101001111010001"; -- -0.106119882046755
	pesos_i(3344) := b"1111111111111111_1111111111111111_1111110000010010_0010100010100100"; -- -0.015347919439825192
	pesos_i(3345) := b"0000000000000000_0000000000000000_0001010110001110_0110111100000101"; -- 0.08420461522606631
	pesos_i(3346) := b"1111111111111111_1111111111111111_1111101001011001_1011101011101011"; -- -0.022068326514988763
	pesos_i(3347) := b"1111111111111111_1111111111111111_1111101101100011_1101000100011101"; -- -0.01800816564933713
	pesos_i(3348) := b"1111111111111111_1111111111111111_1101010101110001_0100011100111101"; -- -0.16624026059430572
	pesos_i(3349) := b"0000000000000000_0000000000000000_0000000110000110_1001110001110011"; -- 0.005960252904354857
	pesos_i(3350) := b"1111111111111111_1111111111111111_1101111000100001_0110111011110100"; -- -0.1323023466601318
	pesos_i(3351) := b"1111111111111111_1111111111111111_1111100100011100_1111100110101110"; -- -0.026901621928236766
	pesos_i(3352) := b"0000000000000000_0000000000000000_0000001110010010_1010011010101100"; -- 0.013956467603279402
	pesos_i(3353) := b"0000000000000000_0000000000000000_0010100100111101_1001011000001011"; -- 0.16109597941397819
	pesos_i(3354) := b"1111111111111111_1111111111111111_1101100000011110_0001101001010110"; -- -0.15579066667769828
	pesos_i(3355) := b"0000000000000000_0000000000000000_0010011110011000_1000111000110000"; -- 0.15467156091980333
	pesos_i(3356) := b"0000000000000000_0000000000000000_0010110110111110_1111101011001010"; -- 0.17869536802149139
	pesos_i(3357) := b"1111111111111111_1111111111111111_1110000010100110_1101001001000100"; -- -0.1224545081159491
	pesos_i(3358) := b"0000000000000000_0000000000000000_0001100100000001_0001011000011000"; -- 0.09767282558177554
	pesos_i(3359) := b"0000000000000000_0000000000000000_0010000110101101_0101110101101011"; -- 0.1315515887344277
	pesos_i(3360) := b"1111111111111111_1111111111111111_1111010100011001_0011001111111011"; -- -0.04258418206571954
	pesos_i(3361) := b"0000000000000000_0000000000000000_0000100100110101_1101100110001111"; -- 0.035977933306613634
	pesos_i(3362) := b"0000000000000000_0000000000000000_0010000000001100_0111100000000100"; -- 0.12519025884689333
	pesos_i(3363) := b"1111111111111111_1111111111111111_1110110011101101_1010101001110110"; -- -0.07449850672767135
	pesos_i(3364) := b"1111111111111111_1111111111111111_1110110110100011_0000000011101100"; -- -0.07173151246797285
	pesos_i(3365) := b"1111111111111111_1111111111111111_1110000011000000_0111001110001101"; -- -0.12206342522326116
	pesos_i(3366) := b"0000000000000000_0000000000000000_0010111100110110_1011101111101011"; -- 0.18442892531850325
	pesos_i(3367) := b"1111111111111111_1111111111111111_1110101011111111_0101110011011001"; -- -0.08204097474700735
	pesos_i(3368) := b"0000000000000000_0000000000000000_0010000101110100_1010011111011010"; -- 0.1306862742525439
	pesos_i(3369) := b"0000000000000000_0000000000000000_0000000011010010_1110101010000110"; -- 0.003218324307674721
	pesos_i(3370) := b"1111111111111111_1111111111111111_1110100000100110_0000101100111100"; -- -0.09316949633440261
	pesos_i(3371) := b"1111111111111111_1111111111111111_1110010100100111_1010011101000101"; -- -0.10486368720550686
	pesos_i(3372) := b"0000000000000000_0000000000000000_0000000110101010_1100100101110000"; -- 0.006512250803448396
	pesos_i(3373) := b"1111111111111111_1111111111111111_1111111111110111_0001101110100110"; -- -0.00013568117018921324
	pesos_i(3374) := b"1111111111111111_1111111111111111_1110011000001000_0000011100110101"; -- -0.10144000000294087
	pesos_i(3375) := b"0000000000000000_0000000000000000_0011000001001000_0000111100111100"; -- 0.18859954079257543
	pesos_i(3376) := b"0000000000000000_0000000000000000_0001000011011011_0001001001001010"; -- 0.06584276502687758
	pesos_i(3377) := b"0000000000000000_0000000000000000_0000111000100000_0100000101111001"; -- 0.05517968370129388
	pesos_i(3378) := b"1111111111111111_1111111111111111_1110111110110000_0011110101101110"; -- -0.0637170415894513
	pesos_i(3379) := b"0000000000000000_0000000000000000_0000111111111111_0100000000100101"; -- 0.06248856451859352
	pesos_i(3380) := b"0000000000000000_0000000000000000_0010001000101011_0110000001110000"; -- 0.13347437605584128
	pesos_i(3381) := b"1111111111111111_1111111111111111_1111110111111101_0111110010100110"; -- -0.007850846634422384
	pesos_i(3382) := b"1111111111111111_1111111111111111_1111100001000011_1010110100100100"; -- -0.030217341243105548
	pesos_i(3383) := b"1111111111111111_1111111111111111_1111000111001110_1100011110001111"; -- -0.05543854489709452
	pesos_i(3384) := b"1111111111111111_1111111111111111_1111010100110000_1011010000001110"; -- -0.0422255960707843
	pesos_i(3385) := b"1111111111111111_1111111111111111_1110001011000101_1110111001111011"; -- -0.11416730391692746
	pesos_i(3386) := b"1111111111111111_1111111111111111_1101011111100010_0110010000011000"; -- -0.15670179755272667
	pesos_i(3387) := b"0000000000000000_0000000000000000_0001110010000110_1111101101010010"; -- 0.111434657643619
	pesos_i(3388) := b"1111111111111111_1111111111111111_1110101110100000_0110011000111110"; -- -0.07958374963627621
	pesos_i(3389) := b"0000000000000000_0000000000000000_0000111111001100_1000011000100101"; -- 0.061714538556391384
	pesos_i(3390) := b"1111111111111111_1111111111111111_1110010100010001_1101001000111101"; -- -0.10519681936892526
	pesos_i(3391) := b"0000000000000000_0000000000000000_0001000000111000_0111110001011010"; -- 0.06336190416207753
	pesos_i(3392) := b"1111111111111111_1111111111111111_1101010011000100_1110100111001011"; -- -0.16887034214996485
	pesos_i(3393) := b"1111111111111111_1111111111111111_1110000010100111_0101101000101110"; -- -0.12244640720390705
	pesos_i(3394) := b"1111111111111111_1111111111111111_1110000010010110_0110001100110100"; -- -0.12270526869366342
	pesos_i(3395) := b"0000000000000000_0000000000000000_0001000100011111_0011101011100000"; -- 0.06688278173746741
	pesos_i(3396) := b"0000000000000000_0000000000000000_0001101011000110_1111110101010011"; -- 0.10459883960692208
	pesos_i(3397) := b"0000000000000000_0000000000000000_0000001111110011_0111100100111111"; -- 0.015433862683691043
	pesos_i(3398) := b"1111111111111111_1111111111111111_1111011110010010_0100110111011101"; -- -0.03292382578637889
	pesos_i(3399) := b"1111111111111111_1111111111111111_1101100010110010_1011110010101100"; -- -0.1535226897403319
	pesos_i(3400) := b"0000000000000000_0000000000000000_0010110000101001_1111001010110100"; -- 0.1725150765071307
	pesos_i(3401) := b"1111111111111111_1111111111111111_1110010111010010_0001000011110000"; -- -0.10226339483343425
	pesos_i(3402) := b"1111111111111111_1111111111111111_1101101000011001_0110011001100001"; -- -0.14804992809815454
	pesos_i(3403) := b"0000000000000000_0000000000000000_0001001010111010_1011101111111000"; -- 0.0731618386486771
	pesos_i(3404) := b"1111111111111111_1111111111111111_1110110101101111_0100001000010100"; -- -0.07252108585707501
	pesos_i(3405) := b"0000000000000000_0000000000000000_0001101001110001_0100000011111010"; -- 0.10329061605007522
	pesos_i(3406) := b"1111111111111111_1111111111111111_1111100011100111_0110101101000001"; -- -0.027718826804590768
	pesos_i(3407) := b"1111111111111111_1111111111111111_1111010111101100_0000110101010000"; -- -0.03936688224865134
	pesos_i(3408) := b"0000000000000000_0000000000000000_0000101110010011_0001001001001101"; -- 0.04521288271562654
	pesos_i(3409) := b"1111111111111111_1111111111111111_1100111110100111_0011110000101010"; -- -0.1888544460638442
	pesos_i(3410) := b"1111111111111111_1111111111111111_1111000010010111_1011010100110111"; -- -0.060185121517329514
	pesos_i(3411) := b"1111111111111111_1111111111111111_1111011000111011_0111111100000111"; -- -0.038154660070563645
	pesos_i(3412) := b"0000000000000000_0000000000000000_0010001001110101_0010001000101110"; -- 0.1345998154868282
	pesos_i(3413) := b"0000000000000000_0000000000000000_0010000001100100_1010010001111110"; -- 0.12653568349700267
	pesos_i(3414) := b"0000000000000000_0000000000000000_0001110101110111_0101010010111100"; -- 0.11510209638674936
	pesos_i(3415) := b"0000000000000000_0000000000000000_0010111010101000_1111110101000110"; -- 0.18226607274361148
	pesos_i(3416) := b"0000000000000000_0000000000000000_0000101110110001_0011111100010010"; -- 0.04567331500822143
	pesos_i(3417) := b"1111111111111111_1111111111111111_1110110010010000_0110000101010110"; -- -0.07592193271674569
	pesos_i(3418) := b"0000000000000000_0000000000000000_0000110111110001_1000110110101110"; -- 0.05446706293297478
	pesos_i(3419) := b"0000000000000000_0000000000000000_0000010100010111_0010011100000001"; -- 0.019884526867891505
	pesos_i(3420) := b"1111111111111111_1111111111111111_1101110001000100_1001111010011000"; -- -0.13957794938795054
	pesos_i(3421) := b"1111111111111111_1111111111111111_1110010110011110_1000110101100000"; -- -0.10304943472357672
	pesos_i(3422) := b"0000000000000000_0000000000000000_0001110110101001_0010111000110011"; -- 0.11586273914254636
	pesos_i(3423) := b"1111111111111111_1111111111111111_1101011100110010_1011110010100101"; -- -0.15938206649313405
	pesos_i(3424) := b"0000000000000000_0000000000000000_0001000010100110_1101001100111110"; -- 0.0650455499937336
	pesos_i(3425) := b"1111111111111111_1111111111111111_1110011101110000_1000100101101110"; -- -0.09593907408826821
	pesos_i(3426) := b"1111111111111111_1111111111111111_1110100001111000_0011001000010100"; -- -0.09191596042296717
	pesos_i(3427) := b"1111111111111111_1111111111111111_1110000111110010_0010110011111111"; -- -0.1173984410921906
	pesos_i(3428) := b"1111111111111111_1111111111111111_1111100101111000_1000011001000011"; -- -0.02550469257745176
	pesos_i(3429) := b"1111111111111111_1111111111111111_1111001011111101_0000101011000011"; -- -0.05082638484842887
	pesos_i(3430) := b"0000000000000000_0000000000000000_0010011000000111_0101101000000101"; -- 0.14854967709603265
	pesos_i(3431) := b"0000000000000000_0000000000000000_0000010110100111_1100101011111100"; -- 0.022091566608740232
	pesos_i(3432) := b"1111111111111111_1111111111111111_1111111011100011_0010010011100100"; -- -0.004346555986078554
	pesos_i(3433) := b"1111111111111111_1111111111111111_1111001111110101_0100011011001000"; -- -0.04703862775540842
	pesos_i(3434) := b"1111111111111111_1111111111111111_1101110000001111_0011001111100010"; -- -0.14039302561121259
	pesos_i(3435) := b"1111111111111111_1111111111111111_1101110110010111_1000110111001010"; -- -0.13440622159963894
	pesos_i(3436) := b"1111111111111111_1111111111111111_1110001111101011_0001100111001000"; -- -0.1096938979140691
	pesos_i(3437) := b"0000000000000000_0000000000000000_0000100000110111_0010010000001010"; -- 0.03209138157113814
	pesos_i(3438) := b"1111111111111111_1111111111111111_1110101100111100_0110010101111010"; -- -0.08110967421835079
	pesos_i(3439) := b"0000000000000000_0000000000000000_0010001110010001_0110001000010111"; -- 0.13893712092217514
	pesos_i(3440) := b"0000000000000000_0000000000000000_0000010101001000_1111010100010101"; -- 0.020644490936269938
	pesos_i(3441) := b"1111111111111111_1111111111111111_1111100000101011_0000000011000101"; -- -0.030593826086421444
	pesos_i(3442) := b"1111111111111111_1111111111111111_1110111111010011_1100000110000000"; -- -0.06317511193603782
	pesos_i(3443) := b"1111111111111111_1111111111111111_1111101111010111_1111010001011111"; -- -0.01623604466533643
	pesos_i(3444) := b"1111111111111111_1111111111111111_1111110010010111_1001010110110001"; -- -0.013312000490119463
	pesos_i(3445) := b"1111111111111111_1111111111111111_1111111100101100_1101100101100101"; -- -0.0032219055216389674
	pesos_i(3446) := b"0000000000000000_0000000000000000_0000011111010011_0010001000111011"; -- 0.030565394778568417
	pesos_i(3447) := b"1111111111111111_1111111111111111_1110011011100111_1111001011001001"; -- -0.09802324867509964
	pesos_i(3448) := b"0000000000000000_0000000000000000_0000100000010010_0000101010011011"; -- 0.03152529032556095
	pesos_i(3449) := b"1111111111111111_1111111111111111_1111000111000110_1000011101101001"; -- -0.05556443871650351
	pesos_i(3450) := b"0000000000000000_0000000000000000_0001010101100111_1101000000001001"; -- 0.08361530521895576
	pesos_i(3451) := b"0000000000000000_0000000000000000_0000001111110110_1111010101001000"; -- 0.015487031920900972
	pesos_i(3452) := b"0000000000000000_0000000000000000_0000000000100100_1110010100100000"; -- 0.0005629734105389195
	pesos_i(3453) := b"1111111111111111_1111111111111111_1110111010000010_1011010110111011"; -- -0.06831802539533893
	pesos_i(3454) := b"1111111111111111_1111111111111111_1111010111111101_1000111110011111"; -- -0.03909971581977029
	pesos_i(3455) := b"0000000000000000_0000000000000000_0010001100000000_1010101100110001"; -- 0.13672895379766886
	pesos_i(3456) := b"1111111111111111_1111111111111111_1101101100011010_1011110011101001"; -- -0.14412326156914032
	pesos_i(3457) := b"1111111111111111_1111111111111111_1111001010100011_1010010001110110"; -- -0.0521905147712522
	pesos_i(3458) := b"1111111111111111_1111111111111111_1111110110110000_0101101110011011"; -- -0.009027742999239924
	pesos_i(3459) := b"1111111111111111_1111111111111111_1111000110110011_0010101101111010"; -- -0.05585983535127178
	pesos_i(3460) := b"0000000000000000_0000000000000000_0001111000001110_0101010011111011"; -- 0.11740618827046811
	pesos_i(3461) := b"1111111111111111_1111111111111111_1101010011001100_0001100000010100"; -- -0.16876077192176017
	pesos_i(3462) := b"1111111111111111_1111111111111111_1111111110000010_1010011001010110"; -- -0.0019126931163739795
	pesos_i(3463) := b"1111111111111111_1111111111111111_1111001111000101_1111000010111010"; -- -0.04776092019654824
	pesos_i(3464) := b"1111111111111111_1111111111111111_1111100000101101_0000111010011111"; -- -0.030562483011362718
	pesos_i(3465) := b"1111111111111111_1111111111111111_1110011111100010_0011101110011011"; -- -0.09420421102493332
	pesos_i(3466) := b"0000000000000000_0000000000000000_0001101000111100_1111111011100110"; -- 0.10249322046114281
	pesos_i(3467) := b"1111111111111111_1111111111111111_1111111001000011_1011100100001011"; -- -0.006779131765841929
	pesos_i(3468) := b"0000000000000000_0000000000000000_0000111010011011_0000011101001110"; -- 0.057053047605099994
	pesos_i(3469) := b"1111111111111111_1111111111111111_1111000110110100_1100001111001101"; -- -0.05583549733262341
	pesos_i(3470) := b"1111111111111111_1111111111111111_1111000000010000_1101000101111001"; -- -0.06224337378818155
	pesos_i(3471) := b"0000000000000000_0000000000000000_0011011101010101_0111000011111101"; -- 0.21614748166864461
	pesos_i(3472) := b"0000000000000000_0000000000000000_0001101010101011_1001100110000011"; -- 0.10418090304235614
	pesos_i(3473) := b"0000000000000000_0000000000000000_0001101110010001_1111011001110111"; -- 0.10769596477377433
	pesos_i(3474) := b"0000000000000000_0000000000000000_0001011111010000_0011110110101111"; -- 0.09302125478262853
	pesos_i(3475) := b"0000000000000000_0000000000000000_0001001110101001_0000011110101000"; -- 0.0767979416292289
	pesos_i(3476) := b"1111111111111111_1111111111111111_1111001101001011_0101011101010010"; -- -0.04963163607718664
	pesos_i(3477) := b"0000000000000000_0000000000000000_0010000101110010_1101011100001010"; -- 0.1306585692246183
	pesos_i(3478) := b"0000000000000000_0000000000000000_0010001101111110_0101001011011111"; -- 0.13864629701381104
	pesos_i(3479) := b"1111111111111111_1111111111111111_1101110111001110_1001010000100110"; -- -0.13356660922269115
	pesos_i(3480) := b"0000000000000000_0000000000000000_0010001111111001_0011011011110101"; -- 0.14052146408187885
	pesos_i(3481) := b"1111111111111111_1111111111111111_1111110110110001_1011011110001001"; -- -0.009007004813407075
	pesos_i(3482) := b"0000000000000000_0000000000000000_0001001111101111_1101000011110110"; -- 0.07787805574268993
	pesos_i(3483) := b"1111111111111111_1111111111111111_1110000101110111_0111110010101111"; -- -0.11927052246940832
	pesos_i(3484) := b"1111111111111111_1111111111111111_1111101001111001_0110110010111100"; -- -0.021584705359658254
	pesos_i(3485) := b"1111111111111111_1111111111111111_1111011101110011_1011010100111101"; -- -0.03339068659510885
	pesos_i(3486) := b"0000000000000000_0000000000000000_0000011010110001_0000101111011010"; -- 0.026139012066456357
	pesos_i(3487) := b"0000000000000000_0000000000000000_0001001000100111_1000001010000011"; -- 0.07091537195652661
	pesos_i(3488) := b"1111111111111111_1111111111111111_1101101011101000_0100101010011110"; -- -0.14489301349432995
	pesos_i(3489) := b"1111111111111111_1111111111111111_1111010011111001_1011110101100110"; -- -0.043064272594254674
	pesos_i(3490) := b"1111111111111111_1111111111111111_1110000011001111_0001101100001000"; -- -0.1218398194551171
	pesos_i(3491) := b"1111111111111111_1111111111111111_1110111001101111_1111100100110110"; -- -0.06860392023401482
	pesos_i(3492) := b"0000000000000000_0000000000000000_0000000111010010_0110010010101110"; -- 0.0071165967941143465
	pesos_i(3493) := b"0000000000000000_0000000000000000_0001110000110010_1010110100101100"; -- 0.11014826125197924
	pesos_i(3494) := b"1111111111111111_1111111111111111_1101001100101100_1001001011001000"; -- -0.1751011143280932
	pesos_i(3495) := b"1111111111111111_1111111111111111_1110111101111111_0110100001000001"; -- -0.06446216981001408
	pesos_i(3496) := b"0000000000000000_0000000000000000_0000101011101111_0110011111010011"; -- 0.04271553894820532
	pesos_i(3497) := b"0000000000000000_0000000000000000_0001110011010101_1101001010110011"; -- 0.11263768068460732
	pesos_i(3498) := b"0000000000000000_0000000000000000_0001101011000001_0100100011111010"; -- 0.10451179596037855
	pesos_i(3499) := b"1111111111111111_1111111111111111_1110100110100010_1100110001010110"; -- -0.08735964674025612
	pesos_i(3500) := b"1111111111111111_1111111111111111_1110101110000000_0001100101010100"; -- -0.08007661533437394
	pesos_i(3501) := b"0000000000000000_0000000000000000_0001100010000010_0011001100101011"; -- 0.09573669243620081
	pesos_i(3502) := b"0000000000000000_0000000000000000_0001001110101000_1001110101111001"; -- 0.07679161269513333
	pesos_i(3503) := b"0000000000000000_0000000000000000_0010010101110110_0011111010000100"; -- 0.1463355134158642
	pesos_i(3504) := b"1111111111111111_1111111111111111_1101010101011111_0000000001101000"; -- -0.16651914074544533
	pesos_i(3505) := b"1111111111111111_1111111111111111_1111001101100010_1110111000110100"; -- -0.049271690697331304
	pesos_i(3506) := b"1111111111111111_1111111111111111_1101100101101101_0101010111111110"; -- -0.1506754165722772
	pesos_i(3507) := b"1111111111111111_1111111111111111_1110010010000101_1010100000111000"; -- -0.1073355544061463
	pesos_i(3508) := b"0000000000000000_0000000000000000_0001001110110100_1110110011010110"; -- 0.0769794485796595
	pesos_i(3509) := b"0000000000000000_0000000000000000_0001101111101001_1101001110111011"; -- 0.10903666806174521
	pesos_i(3510) := b"1111111111111111_1111111111111111_1111111111000001_0011100011101001"; -- -0.0009579116879711264
	pesos_i(3511) := b"0000000000000000_0000000000000000_0000000000011100_0111110110001111"; -- 0.00043472995565428625
	pesos_i(3512) := b"1111111111111111_1111111111111111_1101111101111011_1111011100001010"; -- -0.12701469417039596
	pesos_i(3513) := b"0000000000000000_0000000000000000_0011000110101110_1111110000000111"; -- 0.19407630138027446
	pesos_i(3514) := b"1111111111111111_1111111111111111_1110010100100101_1100000000101100"; -- -0.10489272050910771
	pesos_i(3515) := b"1111111111111111_1111111111111111_1111101101101110_1100001100110111"; -- -0.017841147429716802
	pesos_i(3516) := b"1111111111111111_1111111111111111_1111010011010111_1010001000111011"; -- -0.043584690701860516
	pesos_i(3517) := b"0000000000000000_0000000000000000_0000000110101100_0101111001000110"; -- 0.006536380785472263
	pesos_i(3518) := b"1111111111111111_1111111111111111_1110111011111110_1001110000111111"; -- -0.06642745454556163
	pesos_i(3519) := b"1111111111111111_1111111111111111_1111010101001101_0001010110001111"; -- -0.041792538264624264
	pesos_i(3520) := b"1111111111111111_1111111111111111_1111010000110101_0110000001111001"; -- -0.04606053403944446
	pesos_i(3521) := b"1111111111111111_1111111111111111_1101111000010001_0101011101100010"; -- -0.13254789210699366
	pesos_i(3522) := b"1111111111111111_1111111111111111_1110100001011001_0100100010011011"; -- -0.09238764012972754
	pesos_i(3523) := b"0000000000000000_0000000000000000_0001101001000101_0110110000110101"; -- 0.10262180605471813
	pesos_i(3524) := b"1111111111111111_1111111111111111_1110011100001001_1101010010001100"; -- -0.09750625222787022
	pesos_i(3525) := b"0000000000000000_0000000000000000_0000001011111000_0001100000000001"; -- 0.011598110400982234
	pesos_i(3526) := b"1111111111111111_1111111111111111_1111000010101110_1000110100000010"; -- -0.05983656607474344
	pesos_i(3527) := b"0000000000000000_0000000000000000_0010000010111100_1000110100110001"; -- 0.127877068109165
	pesos_i(3528) := b"0000000000000000_0000000000000000_0000011110000010_0101001001111000"; -- 0.029332308131749064
	pesos_i(3529) := b"0000000000000000_0000000000000000_0000100001111001_1010100100101001"; -- 0.03310639620651727
	pesos_i(3530) := b"0000000000000000_0000000000000000_0010000011000101_1001011010100010"; -- 0.12801495993891257
	pesos_i(3531) := b"0000000000000000_0000000000000000_0010001000101000_0110101111001011"; -- 0.13342927642349625
	pesos_i(3532) := b"1111111111111111_1111111111111111_1110000010010111_1100110011111111"; -- -0.12268370416033776
	pesos_i(3533) := b"0000000000000000_0000000000000000_0000000100110100_1000101011000011"; -- 0.004707977901212803
	pesos_i(3534) := b"0000000000000000_0000000000000000_0000111101110100_1010110110001000"; -- 0.0603741128187954
	pesos_i(3535) := b"1111111111111111_1111111111111111_1110111000111010_0010110000001101"; -- -0.06942486463411754
	pesos_i(3536) := b"0000000000000000_0000000000000000_0000100110011001_0110110011001011"; -- 0.03749732927306473
	pesos_i(3537) := b"0000000000000000_0000000000000000_0000111010110010_1100101111110010"; -- 0.05741572062020231
	pesos_i(3538) := b"0000000000000000_0000000000000000_0001110110110000_1100011100111110"; -- 0.11597867258760201
	pesos_i(3539) := b"1111111111111111_1111111111111111_1111000111001011_0000001001001001"; -- -0.055496079651407786
	pesos_i(3540) := b"1111111111111111_1111111111111111_1101111010001010_0000011001100010"; -- -0.13070640659041377
	pesos_i(3541) := b"1111111111111111_1111111111111111_1111101111110100_1110111010010001"; -- -0.015793885706687674
	pesos_i(3542) := b"1111111111111111_1111111111111111_1101101000100100_1000111110001001"; -- -0.14787962818212186
	pesos_i(3543) := b"0000000000000000_0000000000000000_0001001110101000_0101111101000001"; -- 0.07678790413508947
	pesos_i(3544) := b"1111111111111111_1111111111111111_1110111110010111_0001001011001000"; -- -0.06410105342547304
	pesos_i(3545) := b"0000000000000000_0000000000000000_0010011000111101_0101111000111000"; -- 0.14937390196642047
	pesos_i(3546) := b"0000000000000000_0000000000000000_0000001110110100_1101111011010111"; -- 0.01447861436860789
	pesos_i(3547) := b"0000000000000000_0000000000000000_0001011110001100_1010010110101001"; -- 0.09198985446834548
	pesos_i(3548) := b"0000000000000000_0000000000000000_0000000111011011_1000010000000110"; -- 0.007255794069544114
	pesos_i(3549) := b"1111111111111111_1111111111111111_1110111011110100_1001010011100001"; -- -0.06658048152818725
	pesos_i(3550) := b"1111111111111111_1111111111111111_1111000000010010_0010010010100111"; -- -0.06222315724195934
	pesos_i(3551) := b"0000000000000000_0000000000000000_0001110011111100_0110110000111110"; -- 0.11322666655555688
	pesos_i(3552) := b"1111111111111111_1111111111111111_1101011011001010_1101110100100111"; -- -0.1609670429522041
	pesos_i(3553) := b"1111111111111111_1111111111111111_1111010011110100_1001101000000110"; -- -0.043142674997188456
	pesos_i(3554) := b"0000000000000000_0000000000000000_0000001111100000_0011101000001100"; -- 0.015140178502766694
	pesos_i(3555) := b"0000000000000000_0000000000000000_0001010000110010_1011011011110101"; -- 0.07889884450670254
	pesos_i(3556) := b"1111111111111111_1111111111111111_1110010110010011_0111011101001100"; -- -0.10321859737149965
	pesos_i(3557) := b"0000000000000000_0000000000000000_0010101001000010_1010000101010010"; -- 0.1650791956108673
	pesos_i(3558) := b"0000000000000000_0000000000000000_0000001000101010_0100000111101101"; -- 0.008457298544292408
	pesos_i(3559) := b"1111111111111111_1111111111111111_1111100111111100_0000010101111100"; -- -0.023498208204713295
	pesos_i(3560) := b"0000000000000000_0000000000000000_0000100100000010_0101110010110101"; -- 0.035192293246458034
	pesos_i(3561) := b"0000000000000000_0000000000000000_0001110110111001_1111111010110000"; -- 0.11611930650357685
	pesos_i(3562) := b"1111111111111111_1111111111111111_1111001001000100_1111110010010110"; -- -0.05363484712841733
	pesos_i(3563) := b"0000000000000000_0000000000000000_0001100010110001_0101000101110011"; -- 0.09645566050022351
	pesos_i(3564) := b"1111111111111111_1111111111111111_1110011111010001_1101010011000110"; -- -0.0944544807678335
	pesos_i(3565) := b"1111111111111111_1111111111111111_1101010101000110_1101000001001110"; -- -0.1668882188910327
	pesos_i(3566) := b"1111111111111111_1111111111111111_1101011010010001_0111001011010000"; -- -0.16184313211724494
	pesos_i(3567) := b"0000000000000000_0000000000000000_0000001010100100_0010010011110010"; -- 0.010317143409358895
	pesos_i(3568) := b"1111111111111111_1111111111111111_1101001110101010_1101110010011010"; -- -0.17317410691780233
	pesos_i(3569) := b"0000000000000000_0000000000000000_0000010010111101_0001100101110101"; -- 0.018510428440294987
	pesos_i(3570) := b"0000000000000000_0000000000000000_0010011101110111_1001101001010110"; -- 0.15416874500452304
	pesos_i(3571) := b"0000000000000000_0000000000000000_0000010100000101_1110101001101111"; -- 0.019621517168635052
	pesos_i(3572) := b"0000000000000000_0000000000000000_0010000000001111_1001001111001010"; -- 0.12523769083784125
	pesos_i(3573) := b"0000000000000000_0000000000000000_0000001011001000_1010000111111111"; -- 0.01087391358002936
	pesos_i(3574) := b"0000000000000000_0000000000000000_0010000011111011_1101100100010100"; -- 0.1288428950112967
	pesos_i(3575) := b"1111111111111111_1111111111111111_1110101111111011_1001110011010011"; -- -0.0781919465969914
	pesos_i(3576) := b"0000000000000000_0000000000000000_0000100100000010_1000100000010111"; -- 0.03519487924536169
	pesos_i(3577) := b"1111111111111111_1111111111111111_1101101100100101_1010101001111010"; -- -0.1439565137078284
	pesos_i(3578) := b"0000000000000000_0000000000000000_0000001101011100_0011101100100110"; -- 0.013126084016287318
	pesos_i(3579) := b"1111111111111111_1111111111111111_1111001110010100_0000111001101110"; -- -0.04852208915159144
	pesos_i(3580) := b"0000000000000000_0000000000000000_0010000111011011_0011101011100010"; -- 0.13225143454743962
	pesos_i(3581) := b"1111111111111111_1111111111111111_1101111010010001_1110110111000100"; -- -0.13058580369060738
	pesos_i(3582) := b"0000000000000000_0000000000000000_0000011111000110_0100111001010000"; -- 0.030369657937094115
	pesos_i(3583) := b"0000000000000000_0000000000000000_0000110000110010_0010010011011101"; -- 0.047640136789034525
	pesos_i(3584) := b"1111111111111111_1111111111111111_1110110100101011_1110101010010110"; -- -0.07354863959026559
	pesos_i(3585) := b"0000000000000000_0000000000000000_0000110000011001_1001010000001010"; -- 0.04726529348593966
	pesos_i(3586) := b"0000000000000000_0000000000000000_0000111000110000_1101010001100101"; -- 0.055432581542378206
	pesos_i(3587) := b"1111111111111111_1111111111111111_1101111010011101_0101100011100000"; -- -0.1304115727942437
	pesos_i(3588) := b"0000000000000000_0000000000000000_0001000101000001_0010010111100011"; -- 0.06740032958751434
	pesos_i(3589) := b"1111111111111111_1111111111111111_1110000101001100_0100011011100101"; -- -0.11992985645179498
	pesos_i(3590) := b"1111111111111111_1111111111111111_1110000000001000_0111111000011011"; -- -0.12487041327781614
	pesos_i(3591) := b"1111111111111111_1111111111111111_1111011100000111_0100101101011010"; -- -0.035044947134763915
	pesos_i(3592) := b"1111111111111111_1111111111111111_1111111011100010_0100101011001111"; -- -0.004359554780772924
	pesos_i(3593) := b"1111111111111111_1111111111111111_1101110111000010_1000111110101111"; -- -0.13374998063142374
	pesos_i(3594) := b"1111111111111111_1111111111111111_1110010111101000_1011111100111111"; -- -0.10191731169074245
	pesos_i(3595) := b"0000000000000000_0000000000000000_0001101100110000_1000000110100111"; -- 0.10620889968920315
	pesos_i(3596) := b"1111111111111111_1111111111111111_1110011100110100_1111111011001001"; -- -0.0968476065631122
	pesos_i(3597) := b"0000000000000000_0000000000000000_0001001100000111_0110000111101100"; -- 0.07433139817963562
	pesos_i(3598) := b"0000000000000000_0000000000000000_0010001101000100_1011000011100001"; -- 0.13776689042637116
	pesos_i(3599) := b"1111111111111111_1111111111111111_1110010111100100_1100111111101101"; -- -0.10197735270307524
	pesos_i(3600) := b"1111111111111111_1111111111111111_1110100010010010_1111000100011011"; -- -0.09150784570975569
	pesos_i(3601) := b"0000000000000000_0000000000000000_0000110100111111_1010101011010100"; -- 0.0517527358976491
	pesos_i(3602) := b"1111111111111111_1111111111111111_1111010001011010_1101100010100001"; -- -0.04548879688821599
	pesos_i(3603) := b"1111111111111111_1111111111111111_1110100011110110_0101000100100001"; -- -0.08999150212084356
	pesos_i(3604) := b"1111111111111111_1111111111111111_1111000011111111_1111101101101011"; -- -0.05859402319862926
	pesos_i(3605) := b"1111111111111111_1111111111111111_1111011110001111_1101010101000011"; -- -0.03296153168041675
	pesos_i(3606) := b"0000000000000000_0000000000000000_0000111000111111_1110010100001010"; -- 0.055662455478290664
	pesos_i(3607) := b"0000000000000000_0000000000000000_0000110111100010_1110110011110101"; -- 0.0542438600301848
	pesos_i(3608) := b"0000000000000000_0000000000000000_0010100010101001_1001000000111011"; -- 0.1588373321775287
	pesos_i(3609) := b"1111111111111111_1111111111111111_1111001110001110_0101111001100010"; -- -0.048608876277044945
	pesos_i(3610) := b"0000000000000000_0000000000000000_0010010101011001_0001000111011010"; -- 0.14589034617213784
	pesos_i(3611) := b"1111111111111111_1111111111111111_1111010001110001_0001010001101001"; -- -0.045149540309195935
	pesos_i(3612) := b"1111111111111111_1111111111111111_1110000010111010_0100011011110100"; -- -0.12215763605862844
	pesos_i(3613) := b"0000000000000000_0000000000000000_0010101001110010_0000110011101110"; -- 0.16580277259539938
	pesos_i(3614) := b"0000000000000000_0000000000000000_0001011110101011_0011001100100010"; -- 0.09245605076683079
	pesos_i(3615) := b"0000000000000000_0000000000000000_0010100010011100_1100010011100100"; -- 0.15864210668851544
	pesos_i(3616) := b"0000000000000000_0000000000000000_0001111011000011_1010100000000101"; -- 0.12017297853061329
	pesos_i(3617) := b"1111111111111111_1111111111111111_1110010110001110_1111000010100111"; -- -0.10328765800921517
	pesos_i(3618) := b"1111111111111111_1111111111111111_1110100100110001_0011111101000100"; -- -0.08909229851468166
	pesos_i(3619) := b"1111111111111111_1111111111111111_1111011000010001_1100011010001111"; -- -0.03879126549115682
	pesos_i(3620) := b"0000000000000000_0000000000000000_0010011101110000_0010100101011111"; -- 0.15405520028488895
	pesos_i(3621) := b"1111111111111111_1111111111111111_1101100011111110_1010011100000011"; -- -0.15236431283719706
	pesos_i(3622) := b"1111111111111111_1111111111111111_1101010100011011_0101000000100111"; -- -0.16755198533244897
	pesos_i(3623) := b"0000000000000000_0000000000000000_0000100101010101_1010111011101011"; -- 0.03646367289444086
	pesos_i(3624) := b"0000000000000000_0000000000000000_0001100011001110_0001101101010000"; -- 0.09689493852269213
	pesos_i(3625) := b"1111111111111111_1111111111111111_1110001001101100_0111101110100100"; -- -0.11553218131289007
	pesos_i(3626) := b"0000000000000000_0000000000000000_0000011111001010_0001100000010001"; -- 0.03042745982942462
	pesos_i(3627) := b"1111111111111111_1111111111111111_1110100000010010_1010100101010001"; -- -0.09346524970798273
	pesos_i(3628) := b"1111111111111111_1111111111111111_1110111010001000_0111010000000001"; -- -0.06823039028158644
	pesos_i(3629) := b"0000000000000000_0000000000000000_0000100111001000_0011001010001011"; -- 0.038211020323285994
	pesos_i(3630) := b"0000000000000000_0000000000000000_0000100010111010_1011011011101010"; -- 0.034099037350349914
	pesos_i(3631) := b"1111111111111111_1111111111111111_1110101000110110_1110111011001011"; -- -0.08509929212066852
	pesos_i(3632) := b"0000000000000000_0000000000000000_0000010011100110_1011010011101010"; -- 0.019145304910877042
	pesos_i(3633) := b"0000000000000000_0000000000000000_0010010001110001_0001100100111001"; -- 0.14235074652992735
	pesos_i(3634) := b"1111111111111111_1111111111111111_1111000011111000_0001011111011111"; -- -0.05871439754654871
	pesos_i(3635) := b"0000000000000000_0000000000000000_0001011000000110_1000110010110100"; -- 0.0860374393459073
	pesos_i(3636) := b"1111111111111111_1111111111111111_1110100111100101_1011000111100010"; -- -0.08633888474294492
	pesos_i(3637) := b"1111111111111111_1111111111111111_1101100111001101_0111001100010100"; -- -0.14920883914649796
	pesos_i(3638) := b"1111111111111111_1111111111111111_1101011010001000_0100111010000111"; -- -0.1619826240600428
	pesos_i(3639) := b"1111111111111111_1111111111111111_1101101001000111_1010100000100100"; -- -0.14734410406974535
	pesos_i(3640) := b"0000000000000000_0000000000000000_0000001110010100_0011101101001000"; -- 0.013980584291894166
	pesos_i(3641) := b"0000000000000000_0000000000000000_0000111100111011_0111110110011001"; -- 0.05950150484596796
	pesos_i(3642) := b"1111111111111111_1111111111111111_1101100110111001_1101010011010001"; -- -0.1495081891749027
	pesos_i(3643) := b"1111111111111111_1111111111111111_1111101010011101_0010101110101111"; -- -0.021039266410635048
	pesos_i(3644) := b"0000000000000000_0000000000000000_0001010010111110_1001101111101000"; -- 0.08103346270079624
	pesos_i(3645) := b"0000000000000000_0000000000000000_0001100111001100_1001001001000001"; -- 0.10077776046136137
	pesos_i(3646) := b"0000000000000000_0000000000000000_0000010100111101_0111101011001000"; -- 0.02046935435123131
	pesos_i(3647) := b"0000000000000000_0000000000000000_0001110001110110_0101011001001000"; -- 0.11118067995660916
	pesos_i(3648) := b"0000000000000000_0000000000000000_0000101010100100_0010011011000010"; -- 0.04156725143557061
	pesos_i(3649) := b"1111111111111111_1111111111111111_1101100011100010_1100001110011011"; -- -0.15278985468110926
	pesos_i(3650) := b"0000000000000000_0000000000000000_0000101010010100_0001101110000010"; -- 0.04132244048642492
	pesos_i(3651) := b"0000000000000000_0000000000000000_0010010110011111_0111100000100100"; -- 0.14696455846700693
	pesos_i(3652) := b"0000000000000000_0000000000000000_0001110100010000_0100010011110100"; -- 0.11352950049551327
	pesos_i(3653) := b"0000000000000000_0000000000000000_0001011010100100_0100100110100011"; -- 0.08844433054722671
	pesos_i(3654) := b"0000000000000000_0000000000000000_0001100000000110_1100000011101110"; -- 0.0938530521550899
	pesos_i(3655) := b"0000000000000000_0000000000000000_0001101011110100_0100001000101011"; -- 0.10528958849092229
	pesos_i(3656) := b"0000000000000000_0000000000000000_0000001100110001_1010111010110101"; -- 0.012476843952673197
	pesos_i(3657) := b"1111111111111111_1111111111111111_1110101011100011_1000100011011001"; -- -0.0824655981192383
	pesos_i(3658) := b"0000000000000000_0000000000000000_0001010101001101_0010010010001001"; -- 0.08320835442878961
	pesos_i(3659) := b"1111111111111111_1111111111111111_1101010100010010_0001100111001110"; -- -0.16769255376609726
	pesos_i(3660) := b"0000000000000000_0000000000000000_0001101010101101_1000101111100001"; -- 0.10421060785128813
	pesos_i(3661) := b"1111111111111111_1111111111111111_1110001101100011_0110111001001000"; -- -0.11176405657612178
	pesos_i(3662) := b"1111111111111111_1111111111111111_1111110101011101_0000111111001110"; -- -0.010298740599665951
	pesos_i(3663) := b"0000000000000000_0000000000000000_0000000111011100_1000001111011100"; -- 0.007271042929670058
	pesos_i(3664) := b"0000000000000000_0000000000000000_0001100001111110_0110101111001001"; -- 0.09567903195475222
	pesos_i(3665) := b"1111111111111111_1111111111111111_1111100110010110_0011011010111100"; -- -0.025051669243847604
	pesos_i(3666) := b"0000000000000000_0000000000000000_0000011110000110_0011101011100000"; -- 0.02939193690517077
	pesos_i(3667) := b"0000000000000000_0000000000000000_0010010001101101_1000110111110110"; -- 0.14229666958923484
	pesos_i(3668) := b"1111111111111111_1111111111111111_1111000101010011_0001011000011001"; -- -0.057325953403761724
	pesos_i(3669) := b"1111111111111111_1111111111111111_1110110011111011_1111011000001100"; -- -0.07428037833042495
	pesos_i(3670) := b"0000000000000000_0000000000000000_0010001001101001_1001000110100001"; -- 0.13442335310249612
	pesos_i(3671) := b"0000000000000000_0000000000000000_0011000101011111_0000111101010100"; -- 0.19285674858936538
	pesos_i(3672) := b"1111111111111111_1111111111111111_1011110101010000_0010011100110101"; -- -0.2604957099687403
	pesos_i(3673) := b"0000000000000000_0000000000000000_0000111001111001_1000001100000001"; -- 0.05654162197769835
	pesos_i(3674) := b"0000000000000000_0000000000000000_0010000110100001_1110010011100011"; -- 0.1313765577614931
	pesos_i(3675) := b"0000000000000000_0000000000000000_0001111011111110_1001111101101011"; -- 0.12107273453685027
	pesos_i(3676) := b"1111111111111111_1111111111111111_1101010101010001_1001000101000111"; -- -0.16672412889179092
	pesos_i(3677) := b"1111111111111111_1111111111111111_1101110000001100_0000000000100010"; -- -0.14044188664655896
	pesos_i(3678) := b"1111111111111111_1111111111111111_1101111111010000_1011100001101110"; -- -0.1257214291245951
	pesos_i(3679) := b"1111111111111111_1111111111111111_1101111001000101_1011110100000111"; -- -0.1317483766031956
	pesos_i(3680) := b"0000000000000000_0000000000000000_0000000001001010_0100110101101011"; -- 0.0011337648654744514
	pesos_i(3681) := b"0000000000000000_0000000000000000_0000100011011001_1010100001010100"; -- 0.03457119029008145
	pesos_i(3682) := b"1111111111111111_1111111111111111_1110111111110111_0101110011100100"; -- -0.06263179235497841
	pesos_i(3683) := b"1111111111111111_1111111111111111_1111010010010010_1101101100001100"; -- -0.04463416054435546
	pesos_i(3684) := b"0000000000000000_0000000000000000_0010111010101011_0111110110111001"; -- 0.18230424648963484
	pesos_i(3685) := b"1111111111111111_1111111111111111_1111011011100000_1010100111101100"; -- -0.035634403047478516
	pesos_i(3686) := b"1111111111111111_1111111111111111_1110010111111111_0100000100111001"; -- -0.10157387114328878
	pesos_i(3687) := b"0000000000000000_0000000000000000_0001000010110101_1111001000001101"; -- 0.06527626810829132
	pesos_i(3688) := b"0000000000000000_0000000000000000_0000011110111100_0001001101111001"; -- 0.03021356298409214
	pesos_i(3689) := b"0000000000000000_0000000000000000_0000010011010011_1010000101101110"; -- 0.018854226553720044
	pesos_i(3690) := b"1111111111111111_1111111111111111_1110010001110110_1001010010000000"; -- -0.10756561155344123
	pesos_i(3691) := b"1111111111111111_1111111111111111_1111110010100001_0110011011100110"; -- -0.013162201730212266
	pesos_i(3692) := b"0000000000000000_0000000000000000_0000010100011100_1010000010000011"; -- 0.01996806341982909
	pesos_i(3693) := b"1111111111111111_1111111111111111_1111001000111011_1110010110101100"; -- -0.053773541943460526
	pesos_i(3694) := b"0000000000000000_0000000000000000_0000011011001100_1001100001001001"; -- 0.026559369961201916
	pesos_i(3695) := b"0000000000000000_0000000000000000_0010000110000011_1110110100110111"; -- 0.13091929043011719
	pesos_i(3696) := b"1111111111111111_1111111111111111_1110110110111000_0001010110010000"; -- -0.07140984752896073
	pesos_i(3697) := b"0000000000000000_0000000000000000_0000110110110011_0001111100010111"; -- 0.05351442639135098
	pesos_i(3698) := b"1111111111111111_1111111111111111_1110010101001110_0110000100011011"; -- -0.10427277660800438
	pesos_i(3699) := b"1111111111111111_1111111111111111_1101110111000111_0100011101000000"; -- -0.13367800423622753
	pesos_i(3700) := b"1111111111111111_1111111111111111_1110100100101011_1101111000011101"; -- -0.08917438298209988
	pesos_i(3701) := b"1111111111111111_1111111111111111_1110010111011110_1100100110011000"; -- -0.10206928292973198
	pesos_i(3702) := b"0000000000000000_0000000000000000_0001111010010000_0000110000111100"; -- 0.1193854948987775
	pesos_i(3703) := b"1111111111111111_1111111111111111_1110110001100001_0001100100101001"; -- -0.07664339787458108
	pesos_i(3704) := b"1111111111111111_1111111111111111_1101101010000010_1100001100001100"; -- -0.14644223181825733
	pesos_i(3705) := b"1111111111111111_1111111111111111_1110010100110111_0000111100011111"; -- -0.10462861541479618
	pesos_i(3706) := b"0000000000000000_0000000000000000_0000001011101000_1111001010110010"; -- 0.011367004833661432
	pesos_i(3707) := b"0000000000000000_0000000000000000_0000001001001110_0000001100100010"; -- 0.009002872337150516
	pesos_i(3708) := b"1111111111111111_1111111111111111_1111011100110001_1110100110001101"; -- -0.03439464863861418
	pesos_i(3709) := b"1111111111111111_1111111111111111_1110000001110101_0000010100010001"; -- -0.12321441963178566
	pesos_i(3710) := b"0000000000000000_0000000000000000_0000110101110001_1000011110110101"; -- 0.05251358189516998
	pesos_i(3711) := b"0000000000000000_0000000000000000_0000101011000000_0011000011010000"; -- 0.04199509702627502
	pesos_i(3712) := b"0000000000000000_0000000000000000_0010000001110001_1101101111010001"; -- 0.126737345334917
	pesos_i(3713) := b"1111111111111111_1111111111111111_1110110110010010_0100111001110110"; -- -0.07198629017423475
	pesos_i(3714) := b"1111111111111111_1111111111111111_1110010100111011_1010010010011100"; -- -0.10455867005846284
	pesos_i(3715) := b"1111111111111111_1111111111111111_1100110101011001_1110100010111111"; -- -0.19784684508133535
	pesos_i(3716) := b"1111111111111111_1111111111111111_1101010000011101_1110001000101001"; -- -0.1714190149191735
	pesos_i(3717) := b"1111111111111111_1111111111111111_1101001101111111_0001100011110010"; -- -0.17384189687338775
	pesos_i(3718) := b"1111111111111111_1111111111111111_1111000100010011_1000101111011110"; -- -0.05829549629070294
	pesos_i(3719) := b"1111111111111111_1111111111111111_1111001100001011_0101110010111011"; -- -0.05060787611013035
	pesos_i(3720) := b"0000000000000000_0000000000000000_0010010110001110_1101011000001011"; -- 0.14671075589798394
	pesos_i(3721) := b"1111111111111111_1111111111111111_1111001100110010_1100000010101000"; -- -0.050006827261108805
	pesos_i(3722) := b"0000000000000000_0000000000000000_0010101000111101_1001011011100001"; -- 0.16500227917635857
	pesos_i(3723) := b"1111111111111111_1111111111111111_1111111001011100_0100001100001110"; -- -0.006404694590144519
	pesos_i(3724) := b"1111111111111111_1111111111111111_1110010101100101_0100001001111011"; -- -0.10392364974925258
	pesos_i(3725) := b"0000000000000000_0000000000000000_0010001011111010_0000000001110101"; -- 0.13662722456620577
	pesos_i(3726) := b"0000000000000000_0000000000000000_0010101100110101_0000000000110001"; -- 0.16877747718487954
	pesos_i(3727) := b"0000000000000000_0000000000000000_0001111000110100_0100011010100111"; -- 0.11798516819729944
	pesos_i(3728) := b"0000000000000000_0000000000000000_0000101010100001_1011110000001110"; -- 0.04153037388072109
	pesos_i(3729) := b"0000000000000000_0000000000000000_0010101000111111_0010110111011010"; -- 0.16502653663857114
	pesos_i(3730) := b"0000000000000000_0000000000000000_0000100000101010_1101001111101101"; -- 0.031903500945098355
	pesos_i(3731) := b"1111111111111111_1111111111111111_1101111110010001_0010010000001011"; -- -0.12669157714403065
	pesos_i(3732) := b"1111111111111111_1111111111111111_1111011010001111_0001101110001000"; -- -0.03687885226645224
	pesos_i(3733) := b"1111111111111111_1111111111111111_1110100111111010_1011110000011110"; -- -0.08601784002951117
	pesos_i(3734) := b"1111111111111111_1111111111111111_1110100100100110_0011111000111111"; -- -0.08926020574920987
	pesos_i(3735) := b"0000000000000000_0000000000000000_0010101110110100_1000110110100110"; -- 0.17072377494864
	pesos_i(3736) := b"1111111111111111_1111111111111111_1101111010000110_1011101011001010"; -- -0.13075668866865822
	pesos_i(3737) := b"1111111111111111_1111111111111111_1110100011100010_0000000110011110"; -- -0.09030141734655577
	pesos_i(3738) := b"0000000000000000_0000000000000000_0000101110001000_0011011010000101"; -- 0.04504719488891196
	pesos_i(3739) := b"1111111111111111_1111111111111111_1101111000100011_0001101011100111"; -- -0.13227683885957714
	pesos_i(3740) := b"0000000000000000_0000000000000000_0010101010110100_1011010000101101"; -- 0.16681982143473095
	pesos_i(3741) := b"1111111111111111_1111111111111111_1111010001101011_1100111101000011"; -- -0.04522995576596459
	pesos_i(3742) := b"0000000000000000_0000000000000000_0010111111110111_0010010000110110"; -- 0.1873648291671217
	pesos_i(3743) := b"0000000000000000_0000000000000000_0010100111010111_1010100110010000"; -- 0.1634469963835495
	pesos_i(3744) := b"1111111111111111_1111111111111111_1111100001111110_0111100000010001"; -- -0.02932023617166396
	pesos_i(3745) := b"1111111111111111_1111111111111111_1110101111100010_0011001100110011"; -- -0.07857971187131843
	pesos_i(3746) := b"0000000000000000_0000000000000000_0001110100110010_1101100000101000"; -- 0.1140570734703429
	pesos_i(3747) := b"1111111111111111_1111111111111111_1110010101010010_0000110011010111"; -- -0.10421676399213778
	pesos_i(3748) := b"1111111111111111_1111111111111111_1110001110101110_0110111001110000"; -- -0.11061963806661917
	pesos_i(3749) := b"0000000000000000_0000000000000000_0001010110101011_0010000000101001"; -- 0.08464241974368193
	pesos_i(3750) := b"0000000000000000_0000000000000000_0000111100110010_0010101001110111"; -- 0.05935922063664155
	pesos_i(3751) := b"1111111111111111_1111111111111111_1111010110000111_1110111111010100"; -- -0.04089451858794768
	pesos_i(3752) := b"0000000000000000_0000000000000000_0001110000111001_0011101100010110"; -- 0.11024827266394424
	pesos_i(3753) := b"0000000000000000_0000000000000000_0000100101000011_0010000011110100"; -- 0.03618055313433318
	pesos_i(3754) := b"0000000000000000_0000000000000000_0010011001110010_1101001100100010"; -- 0.15018958653094264
	pesos_i(3755) := b"1111111111111111_1111111111111111_1110011011100100_1100001000010111"; -- -0.09807192750305088
	pesos_i(3756) := b"1111111111111111_1111111111111111_1111101011001110_0010010010110101"; -- -0.020292001644344606
	pesos_i(3757) := b"1111111111111111_1111111111111111_1111001000100111_0100111100101000"; -- -0.05408768916497114
	pesos_i(3758) := b"0000000000000000_0000000000000000_0010010110010101_0100111100100000"; -- 0.14680952568424968
	pesos_i(3759) := b"0000000000000000_0000000000000000_0010111010001000_1000011010001110"; -- 0.1817707153219141
	pesos_i(3760) := b"1111111111111111_1111111111111111_1111011100011000_0001010010010001"; -- -0.034788813135589014
	pesos_i(3761) := b"0000000000000000_0000000000000000_0000100110100000_1110110000000001"; -- 0.03761172320328111
	pesos_i(3762) := b"0000000000000000_0000000000000000_0010010110100010_1001000100011110"; -- 0.14701182350934908
	pesos_i(3763) := b"1111111111111111_1111111111111111_1110100011101101_1001110001000001"; -- -0.09012435355549764
	pesos_i(3764) := b"0000000000000000_0000000000000000_0010100111000101_1001011101000101"; -- 0.16317124771741262
	pesos_i(3765) := b"0000000000000000_0000000000000000_0000101010000001_1011001110100011"; -- 0.04104159088943109
	pesos_i(3766) := b"0000000000000000_0000000000000000_0010001100001001_1010110001010011"; -- 0.13686635037584532
	pesos_i(3767) := b"0000000000000000_0000000000000000_0000100010010000_0001010011001001"; -- 0.033448504531733474
	pesos_i(3768) := b"1111111111111111_1111111111111111_1111111001010100_1110000011001001"; -- -0.00651736357983787
	pesos_i(3769) := b"1111111111111111_1111111111111111_1111100011011011_1000100010110101"; -- -0.027900176832661515
	pesos_i(3770) := b"0000000000000000_0000000000000000_0010101101001010_0000011000101001"; -- 0.1690982675208159
	pesos_i(3771) := b"1111111111111111_1111111111111111_1111001000100010_1111111101101001"; -- -0.054153477460644396
	pesos_i(3772) := b"1111111111111111_1111111111111111_1110010101100010_0100101100101010"; -- -0.10396890842909409
	pesos_i(3773) := b"1111111111111111_1111111111111111_1110101111111001_1011110001110010"; -- -0.07822057941514565
	pesos_i(3774) := b"0000000000000000_0000000000000000_0010100000100101_0111110100111001"; -- 0.1568220391332065
	pesos_i(3775) := b"1111111111111111_1111111111111111_1110100000010100_1111000011100011"; -- -0.09343046614762224
	pesos_i(3776) := b"1111111111111111_1111111111111111_1111010111101111_1100001110011000"; -- -0.03931024105327241
	pesos_i(3777) := b"0000000000000000_0000000000000000_0001011101111010_1101100001011100"; -- 0.0917182182785962
	pesos_i(3778) := b"1111111111111111_1111111111111111_1111011111011000_1000011011011110"; -- -0.03185231293831277
	pesos_i(3779) := b"0000000000000000_0000000000000000_0010001010110010_1010111001101110"; -- 0.1355389612717871
	pesos_i(3780) := b"0000000000000000_0000000000000000_0000101000000111_1111100110011100"; -- 0.039184189504192925
	pesos_i(3781) := b"0000000000000000_0000000000000000_0001000011011101_0101001110011100"; -- 0.06587717583945771
	pesos_i(3782) := b"1111111111111111_1111111111111111_1110111011010100_0010001001100100"; -- -0.06707558679021608
	pesos_i(3783) := b"0000000000000000_0000000000000000_0001011010100110_0001000100000010"; -- 0.08847147279564412
	pesos_i(3784) := b"0000000000000000_0000000000000000_0100010100001011_0000001011111100"; -- 0.26969927450488057
	pesos_i(3785) := b"1111111111111111_1111111111111111_1110010010101010_1110101000010001"; -- -0.10676705451572617
	pesos_i(3786) := b"0000000000000000_0000000000000000_0000010110101001_1101011100011111"; -- 0.022122807539207923
	pesos_i(3787) := b"0000000000000000_0000000000000000_0000100100111010_0110001011110101"; -- 0.03604715808656832
	pesos_i(3788) := b"1111111111111111_1111111111111111_1110011010000011_0110011001011001"; -- -0.09955749821596117
	pesos_i(3789) := b"0000000000000000_0000000000000000_0010100010000000_0100011111001010"; -- 0.15820740384931606
	pesos_i(3790) := b"0000000000000000_0000000000000000_0000101101111101_0110110010010101"; -- 0.04488257056625005
	pesos_i(3791) := b"1111111111111111_1111111111111111_1111011011001101_0111100101011110"; -- -0.03592721426364873
	pesos_i(3792) := b"0000000000000000_0000000000000000_0001001011000001_1011101100111110"; -- 0.07326860684462919
	pesos_i(3793) := b"1111111111111111_1111111111111111_1110100110111100_0000111011111001"; -- -0.08697420525474168
	pesos_i(3794) := b"1111111111111111_1111111111111111_1101001110010011_0000010010101001"; -- -0.17353793019189256
	pesos_i(3795) := b"0000000000000000_0000000000000000_0010001000111011_0111101111010100"; -- 0.13372014933093104
	pesos_i(3796) := b"0000000000000000_0000000000000000_0010000001001001_1101100101110110"; -- 0.12612685321237133
	pesos_i(3797) := b"1111111111111111_1111111111111111_1111100000001010_0001010110101111"; -- -0.03109611973675135
	pesos_i(3798) := b"0000000000000000_0000000000000000_0001001100100001_0010001010011101"; -- 0.07472435305306649
	pesos_i(3799) := b"1111111111111111_1111111111111111_1110001000111001_0000110100010101"; -- -0.1163169692392655
	pesos_i(3800) := b"0000000000000000_0000000000000000_0000111000011010_0011011000011100"; -- 0.05508745363335275
	pesos_i(3801) := b"1111111111111111_1111111111111111_1110011000010110_1101010011110010"; -- -0.10121411409424817
	pesos_i(3802) := b"0000000000000000_0000000000000000_0000001000111001_0100010110000000"; -- 0.008686393614317788
	pesos_i(3803) := b"0000000000000000_0000000000000000_0001011011111101_1001000010001010"; -- 0.08980658894818468
	pesos_i(3804) := b"0000000000000000_0000000000000000_0000010111000111_0011101011110110"; -- 0.02257126336317318
	pesos_i(3805) := b"1111111111111111_1111111111111111_1101111100111010_0000001001101101"; -- -0.12802109561263236
	pesos_i(3806) := b"0000000000000000_0000000000000000_0010011000010110_1000100101011111"; -- 0.14878138129816548
	pesos_i(3807) := b"0000000000000000_0000000000000000_0001100011001101_1000101011111001"; -- 0.09688633511440417
	pesos_i(3808) := b"0000000000000000_0000000000000000_0000001110100100_1011000101101011"; -- 0.014231766413060593
	pesos_i(3809) := b"0000000000000000_0000000000000000_0010101100000110_1001100010000000"; -- 0.16806939252084638
	pesos_i(3810) := b"1111111111111111_1111111111111111_1111111011101101_1000010111101000"; -- -0.004188185651442582
	pesos_i(3811) := b"0000000000000000_0000000000000000_0010001101010011_0110110000010011"; -- 0.13799167127439596
	pesos_i(3812) := b"1111111111111111_1111111111111111_1111000101100011_0001001101000111"; -- -0.05708198090522915
	pesos_i(3813) := b"1111111111111111_1111111111111111_1110011010111000_0011000011110101"; -- -0.09875196463625267
	pesos_i(3814) := b"0000000000000000_0000000000000000_0010011111110100_0000100010010001"; -- 0.1560674051342311
	pesos_i(3815) := b"1111111111111111_1111111111111111_1111011000110000_1010110101111111"; -- -0.03831973684885803
	pesos_i(3816) := b"1111111111111111_1111111111111111_1110111000101110_0101011011111101"; -- -0.06960541068273793
	pesos_i(3817) := b"1111111111111111_1111111111111111_1111000111011010_0001100001000111"; -- -0.05526588689162292
	pesos_i(3818) := b"1111111111111111_1111111111111111_1101010010010100_1110010011011110"; -- -0.16960305757827668
	pesos_i(3819) := b"0000000000000000_0000000000000000_0010000111001001_0001110001111000"; -- 0.13197496339832065
	pesos_i(3820) := b"0000000000000000_0000000000000000_0000110100101010_1111000001011111"; -- 0.05143644625833234
	pesos_i(3821) := b"0000000000000000_0000000000000000_0010001001100010_1010000010101011"; -- 0.1343174378100836
	pesos_i(3822) := b"1111111111111111_1111111111111111_1101111010101110_0001111011111000"; -- -0.13015562493177418
	pesos_i(3823) := b"0000000000000000_0000000000000000_0000100001010000_0101011111011001"; -- 0.0324759391726782
	pesos_i(3824) := b"1111111111111111_1111111111111111_1110011101101111_1101111011000001"; -- -0.09594924719391958
	pesos_i(3825) := b"0000000000000000_0000000000000000_0001011001001010_0011010010011001"; -- 0.08706978552002924
	pesos_i(3826) := b"0000000000000000_0000000000000000_0001001100110110_0010101101001010"; -- 0.07504530488975814
	pesos_i(3827) := b"0000000000000000_0000000000000000_0001100111110000_0010000000111110"; -- 0.10132028114193199
	pesos_i(3828) := b"0000000000000000_0000000000000000_0000000011111011_0010110101000000"; -- 0.003832653149023404
	pesos_i(3829) := b"0000000000000000_0000000000000000_0001000100100111_0000110011000111"; -- 0.06700210432983604
	pesos_i(3830) := b"0000000000000000_0000000000000000_0010010100010101_1111100110101110"; -- 0.1448665666314394
	pesos_i(3831) := b"0000000000000000_0000000000000000_0000111011010010_0010001101000010"; -- 0.057893947276674185
	pesos_i(3832) := b"1111111111111111_1111111111111111_1110011101001100_0001100010100100"; -- -0.09649511331970484
	pesos_i(3833) := b"0000000000000000_0000000000000000_0000000010011110_0110101101100011"; -- 0.0024172895182811125
	pesos_i(3834) := b"1111111111111111_1111111111111111_1110010110110011_0001000011001010"; -- -0.10273642613846484
	pesos_i(3835) := b"0000000000000000_0000000000000000_0001001111010100_0110010001101001"; -- 0.07745959811229351
	pesos_i(3836) := b"1111111111111111_1111111111111111_1111011011110001_1001001001000010"; -- -0.035376414122838575
	pesos_i(3837) := b"1111111111111111_1111111111111111_1101101010100101_0111101111000010"; -- -0.1459124232803725
	pesos_i(3838) := b"0000000000000000_0000000000000000_0010011101010011_0001001000100100"; -- 0.15361131067025557
	pesos_i(3839) := b"1111111111111111_1111111111111111_1101101100000100_1101111101011000"; -- -0.1444569025641845
	pesos_i(3840) := b"1111111111111111_1111111111111111_1111000110110000_1011011010100001"; -- -0.05589731748774529
	pesos_i(3841) := b"0000000000000000_0000000000000000_0000011110011010_1101011100010001"; -- 0.0297064225382155
	pesos_i(3842) := b"1111111111111111_1111111111111111_1101100101010111_0010101101101111"; -- -0.15101364654534102
	pesos_i(3843) := b"1111111111111111_1111111111111111_1101100111110110_1101100101100111"; -- -0.1485771296868072
	pesos_i(3844) := b"1111111111111111_1111111111111111_1110011000000011_1001001011100010"; -- -0.10150796865387646
	pesos_i(3845) := b"1111111111111111_1111111111111111_1111110100101110_1100111101011100"; -- -0.011004486137811973
	pesos_i(3846) := b"1111111111111111_1111111111111111_1110101001111000_1100010101101101"; -- -0.0840946778130099
	pesos_i(3847) := b"1111111111111111_1111111111111111_1101110001100110_1111010010100001"; -- -0.13905402239009315
	pesos_i(3848) := b"0000000000000000_0000000000000000_0001110100101000_1101010010001001"; -- 0.11390426970255223
	pesos_i(3849) := b"1111111111111111_1111111111111111_1110101101100000_1110100001001111"; -- -0.08055255949023758
	pesos_i(3850) := b"0000000000000000_0000000000000000_0000101001001000_0100011001000000"; -- 0.04016532005675207
	pesos_i(3851) := b"0000000000000000_0000000000000000_0001110110001011_1101100000001000"; -- 0.11541509803338547
	pesos_i(3852) := b"1111111111111111_1111111111111111_1110100011000001_1100101001000111"; -- -0.09079299701554845
	pesos_i(3853) := b"0000000000000000_0000000000000000_0010100101000110_1101000001111010"; -- 0.16123679147884265
	pesos_i(3854) := b"1111111111111111_1111111111111111_1110111000101010_1010011000011101"; -- -0.06966172972863238
	pesos_i(3855) := b"1111111111111111_1111111111111111_1111001000110101_1000100010110110"; -- -0.05387063546792672
	pesos_i(3856) := b"0000000000000000_0000000000000000_0010010010000111_0110000000111001"; -- 0.14269067181508974
	pesos_i(3857) := b"0000000000000000_0000000000000000_0001010111110100_1000101010111111"; -- 0.08576266451991671
	pesos_i(3858) := b"0000000000000000_0000000000000000_0001011010101001_1011100111010010"; -- 0.0885273111551096
	pesos_i(3859) := b"1111111111111111_1111111111111111_1111100101000110_1110110011110110"; -- -0.02626151082149076
	pesos_i(3860) := b"1111111111111111_1111111111111111_1111011110001011_1101011101100101"; -- -0.0330224397506341
	pesos_i(3861) := b"1111111111111111_1111111111111111_1111010000010011_0001001011011011"; -- -0.04658395903976355
	pesos_i(3862) := b"1111111111111111_1111111111111111_1111101110011101_1000100100000010"; -- -0.01712745372227695
	pesos_i(3863) := b"1111111111111111_1111111111111111_1111101101000011_1010101100011010"; -- -0.018498712578935754
	pesos_i(3864) := b"1111111111111111_1111111111111111_1100111001100101_1110011110010010"; -- -0.19375755960681734
	pesos_i(3865) := b"1111111111111111_1111111111111111_1101111011111010_0101101110000000"; -- -0.12899234884088523
	pesos_i(3866) := b"0000000000000000_0000000000000000_0001110111001110_0101101110101000"; -- 0.11643002380056253
	pesos_i(3867) := b"0000000000000000_0000000000000000_0000011000111110_1000110010110110"; -- 0.024391932026563392
	pesos_i(3868) := b"1111111111111111_1111111111111111_1111001010101111_0100001101001001"; -- -0.05201320148629057
	pesos_i(3869) := b"0000000000000000_0000000000000000_0000111111000100_1001000000111010"; -- 0.06159306913684414
	pesos_i(3870) := b"0000000000000000_0000000000000000_0010010010100101_1011011001101111"; -- 0.14315357404620419
	pesos_i(3871) := b"0000000000000000_0000000000000000_0001011010110011_0011111000011111"; -- 0.08867252605008788
	pesos_i(3872) := b"1111111111111111_1111111111111111_1101011101110011_1100101111101110"; -- -0.1583893341018375
	pesos_i(3873) := b"1111111111111111_1111111111111111_1101101010110011_1000111111001001"; -- -0.1456976064414476
	pesos_i(3874) := b"0000000000000000_0000000000000000_0000101001110000_1011111010100000"; -- 0.04078284649999115
	pesos_i(3875) := b"0000000000000000_0000000000000000_0000100011011111_1110011111100011"; -- 0.0346665315683328
	pesos_i(3876) := b"1111111111111111_1111111111111111_1110011000001111_0010011101001100"; -- -0.1013312759337441
	pesos_i(3877) := b"1111111111111111_1111111111111111_1110100111100101_0110111111001101"; -- -0.0863428234738816
	pesos_i(3878) := b"0000000000000000_0000000000000000_0000111001000110_0011110000001101"; -- 0.05575919447168101
	pesos_i(3879) := b"1111111111111111_1111111111111111_1101010110011011_1011011100110000"; -- -0.165592718872766
	pesos_i(3880) := b"0000000000000000_0000000000000000_0000010011000011_1100110101111011"; -- 0.01861271150137686
	pesos_i(3881) := b"0000000000000000_0000000000000000_0001000111010011_1110000011001010"; -- 0.06963925286761273
	pesos_i(3882) := b"1111111111111111_1111111111111111_1110000111101011_0000001100010100"; -- -0.11750775103956912
	pesos_i(3883) := b"0000000000000000_0000000000000000_0000110100100000_1001101111110111"; -- 0.05127882750974978
	pesos_i(3884) := b"1111111111111111_1111111111111111_1110111110011011_1110011011011110"; -- -0.06402737682693817
	pesos_i(3885) := b"1111111111111111_1111111111111111_1101111000001001_0110100010011100"; -- -0.13266893574022018
	pesos_i(3886) := b"1111111111111111_1111111111111111_1110100111111000_0000100010011110"; -- -0.0860590567851233
	pesos_i(3887) := b"1111111111111111_1111111111111111_1111111000011111_0011111100101101"; -- -0.007335712079079153
	pesos_i(3888) := b"0000000000000000_0000000000000000_0000111101000000_1101111100111110"; -- 0.0595836186796134
	pesos_i(3889) := b"1111111111111111_1111111111111111_1101101110111100_1100011111001011"; -- -0.1416506891691437
	pesos_i(3890) := b"1111111111111111_1111111111111111_1111001001110101_1100101010101110"; -- -0.052890140934913614
	pesos_i(3891) := b"1111111111111111_1111111111111111_1111000011111011_0000001000100001"; -- -0.058669917152042735
	pesos_i(3892) := b"0000000000000000_0000000000000000_0010110011011110_1000010111000011"; -- 0.17527042398847242
	pesos_i(3893) := b"0000000000000000_0000000000000000_0001101111100011_1101101011011010"; -- 0.10894553978269769
	pesos_i(3894) := b"0000000000000000_0000000000000000_0001100001001110_0100111110001111"; -- 0.094944927704567
	pesos_i(3895) := b"0000000000000000_0000000000000000_0010001100010111_0101001001101010"; -- 0.1370746144065574
	pesos_i(3896) := b"0000000000000000_0000000000000000_0000111100010110_1000010101110000"; -- 0.05893739691881708
	pesos_i(3897) := b"0000000000000000_0000000000000000_0001100010001000_0001011011100010"; -- 0.09582655915550149
	pesos_i(3898) := b"1111111111111111_1111111111111111_1110000111100010_0000010011101111"; -- -0.117644969517459
	pesos_i(3899) := b"0000000000000000_0000000000000000_0010100011111001_0100001111010001"; -- 0.16005348072813755
	pesos_i(3900) := b"0000000000000000_0000000000000000_0000110010011001_0011010011111001"; -- 0.04921275219634885
	pesos_i(3901) := b"0000000000000000_0000000000000000_0010001010011100_0111111001011000"; -- 0.13520040171878178
	pesos_i(3902) := b"1111111111111111_1111111111111111_1101010010000001_0000011111110011"; -- -0.16990614245474703
	pesos_i(3903) := b"1111111111111111_1111111111111111_1110111111001110_0010011101100011"; -- -0.06326059178279618
	pesos_i(3904) := b"1111111111111111_1111111111111111_1101111110110111_0110010010010110"; -- -0.12610789623290142
	pesos_i(3905) := b"1111111111111111_1111111111111111_1111001110110101_1110110000000101"; -- -0.04800534128660638
	pesos_i(3906) := b"1111111111111111_1111111111111111_1111110110110000_1111010110000000"; -- -0.009018570152986585
	pesos_i(3907) := b"0000000000000000_0000000000000000_0010010111100001_0011001000101000"; -- 0.14796746699750488
	pesos_i(3908) := b"0000000000000000_0000000000000000_0001110000011111_1111101101001100"; -- 0.10986300083633756
	pesos_i(3909) := b"0000000000000000_0000000000000000_0001010001010010_0010110110111011"; -- 0.07937894656673897
	pesos_i(3910) := b"1111111111111111_1111111111111111_1101101000010001_0100100001100001"; -- -0.14817378649925886
	pesos_i(3911) := b"0000000000000000_0000000000000000_0000110110011001_1001000111111111"; -- 0.0531245466869089
	pesos_i(3912) := b"0000000000000000_0000000000000000_0001110001010000_0011011111111110"; -- 0.11059904057833249
	pesos_i(3913) := b"1111111111111111_1111111111111111_1101011100101100_0000011111110101"; -- -0.15948438899364453
	pesos_i(3914) := b"0000000000000000_0000000000000000_0001101111100010_0000101101010000"; -- 0.10891791068337252
	pesos_i(3915) := b"1111111111111111_1111111111111111_1111100010010111_1101100110110100"; -- -0.028932946794835598
	pesos_i(3916) := b"1111111111111111_1111111111111111_1101010010000111_1000100001010001"; -- -0.16980693836873698
	pesos_i(3917) := b"1111111111111111_1111111111111111_1101001100010011_1001101001110101"; -- -0.1754821266028458
	pesos_i(3918) := b"1111111111111111_1111111111111111_1101110010001111_1111010110011100"; -- -0.13842835377220736
	pesos_i(3919) := b"1111111111111111_1111111111111111_1110011101101011_1011101101100001"; -- -0.09601239085809021
	pesos_i(3920) := b"1111111111111111_1111111111111111_1110010000001110_0111001110101100"; -- -0.10915448243059982
	pesos_i(3921) := b"0000000000000000_0000000000000000_0000001011000100_1001100111110010"; -- 0.010812398491356377
	pesos_i(3922) := b"1111111111111111_1111111111111111_1111010011110110_1101011000011010"; -- -0.04310857644962784
	pesos_i(3923) := b"1111111111111111_1111111111111111_1101100001100011_1010001011011110"; -- -0.15472967226426812
	pesos_i(3924) := b"0000000000000000_0000000000000000_0010010000110001_0011111001100110"; -- 0.14137639982143765
	pesos_i(3925) := b"0000000000000000_0000000000000000_0000010100100101_1111111101010000"; -- 0.020111043108438892
	pesos_i(3926) := b"1111111111111111_1111111111111111_1110011010111111_1010011010001101"; -- -0.09863814413778983
	pesos_i(3927) := b"0000000000000000_0000000000000000_0000110100110110_0011001010110011"; -- 0.05160824659250501
	pesos_i(3928) := b"0000000000000000_0000000000000000_0010011110010010_0111000110111101"; -- 0.15457831256017754
	pesos_i(3929) := b"1111111111111111_1111111111111111_1101111111010100_0111101001010010"; -- -0.12566409597074304
	pesos_i(3930) := b"1111111111111111_1111111111111111_1101100010111000_1111011110110001"; -- -0.15342761928998488
	pesos_i(3931) := b"1111111111111111_1111111111111111_1101101111010111_1111101011110000"; -- -0.14123565338198227
	pesos_i(3932) := b"0000000000000000_0000000000000000_0001000110101010_1100100001111100"; -- 0.06901219384878227
	pesos_i(3933) := b"0000000000000000_0000000000000000_0001100010001100_0101000000011000"; -- 0.09589100444550527
	pesos_i(3934) := b"1111111111111111_1111111111111111_1111001100001010_0011100101010000"; -- -0.050625246048535515
	pesos_i(3935) := b"1111111111111111_1111111111111111_1101110100111001_1101001100110110"; -- -0.13583640983185255
	pesos_i(3936) := b"0000000000000000_0000000000000000_0000101110100010_0001010101110010"; -- 0.04544195214841887
	pesos_i(3937) := b"1111111111111111_1111111111111111_1101101011110011_0111101101110000"; -- -0.14472225688984872
	pesos_i(3938) := b"1111111111111111_1111111111111111_1110100001100001_1001011010011010"; -- -0.09226092096221643
	pesos_i(3939) := b"1111111111111111_1111111111111111_1110111101001001_0110100101110011"; -- -0.06528607304016565
	pesos_i(3940) := b"0000000000000000_0000000000000000_0000110011010001_1000000001100000"; -- 0.05007173865419896
	pesos_i(3941) := b"1111111111111111_1111111111111111_1110111110001011_1110010101110001"; -- -0.06427160250251558
	pesos_i(3942) := b"0000000000000000_0000000000000000_0001010011001001_0001010011000011"; -- 0.08119325402129754
	pesos_i(3943) := b"0000000000000000_0000000000000000_0010000011010100_0011011111110011"; -- 0.12823819803473221
	pesos_i(3944) := b"1111111111111111_1111111111111111_1110110001001101_0000111100001100"; -- -0.07694917642004895
	pesos_i(3945) := b"1111111111111111_1111111111111111_1111011110010010_0010100101000100"; -- -0.03292600711376467
	pesos_i(3946) := b"0000000000000000_0000000000000000_0000111110010001_1000100010010100"; -- 0.060814415092531486
	pesos_i(3947) := b"0000000000000000_0000000000000000_0010101000110101_0010011000011011"; -- 0.16487348706862534
	pesos_i(3948) := b"1111111111111111_1111111111111111_1101110110000010_1000011110001111"; -- -0.13472702751787197
	pesos_i(3949) := b"1111111111111111_1111111111111111_1111100011010000_0000101100010101"; -- -0.028075511410927217
	pesos_i(3950) := b"1111111111111111_1111111111111111_1101110110101111_1011101010111100"; -- -0.134037331608813
	pesos_i(3951) := b"1111111111111111_1111111111111111_1111100100000110_1001111111000010"; -- -0.02724267484284054
	pesos_i(3952) := b"1111111111111111_1111111111111111_1111011000010100_1111100111101001"; -- -0.03874242834592673
	pesos_i(3953) := b"0000000000000000_0000000000000000_0010010101111101_0101001001001000"; -- 0.14644350287158242
	pesos_i(3954) := b"0000000000000000_0000000000000000_0010001010111000_1011011111111011"; -- 0.13563108332257895
	pesos_i(3955) := b"0000000000000000_0000000000000000_0010000000100001_1111101111000011"; -- 0.1255185461898854
	pesos_i(3956) := b"1111111111111111_1111111111111111_1111010101011101_1010101110101100"; -- -0.041539450181484305
	pesos_i(3957) := b"0000000000000000_0000000000000000_0001101000101101_1110111111101001"; -- 0.10226344533725006
	pesos_i(3958) := b"0000000000000000_0000000000000000_0010111010011111_0101011111100011"; -- 0.18211888588767022
	pesos_i(3959) := b"1111111111111111_1111111111111111_1110001000001111_1100001001110001"; -- -0.11694702859127508
	pesos_i(3960) := b"0000000000000000_0000000000000000_0001001100111010_1000001010111001"; -- 0.0751115515072727
	pesos_i(3961) := b"1111111111111111_1111111111111111_1111111111101101_0011001011111011"; -- -0.00028687835763108643
	pesos_i(3962) := b"0000000000000000_0000000000000000_0000110010011101_1101111011110111"; -- 0.049283919600966834
	pesos_i(3963) := b"1111111111111111_1111111111111111_1110010011000110_0001100111100101"; -- -0.106352216300745
	pesos_i(3964) := b"0000000000000000_0000000000000000_0001100101110111_0111010001111100"; -- 0.09947898882764024
	pesos_i(3965) := b"0000000000000000_0000000000000000_0000011010010111_1000101000101000"; -- 0.025749811810395623
	pesos_i(3966) := b"1111111111111111_1111111111111111_1101100000011101_0110110000011100"; -- -0.155801051278229
	pesos_i(3967) := b"0000000000000000_0000000000000000_0001110100011011_1110110010000111"; -- 0.11370733535511084
	pesos_i(3968) := b"0000000000000000_0000000000000000_0000011100111011_1000011010100010"; -- 0.028252043320658365
	pesos_i(3969) := b"0000000000000000_0000000000000000_0001001000011110_0110000000101100"; -- 0.07077599599324118
	pesos_i(3970) := b"1111111111111111_1111111111111111_1101011110010010_1010111011001010"; -- -0.1579180484859241
	pesos_i(3971) := b"1111111111111111_1111111111111111_1111000110111100_0001110001110110"; -- -0.05572340127679386
	pesos_i(3972) := b"0000000000000000_0000000000000000_0000101100000000_0100010010001000"; -- 0.042972834707664984
	pesos_i(3973) := b"0000000000000000_0000000000000000_0000010011110001_1011101101100001"; -- 0.019313536901743575
	pesos_i(3974) := b"1111111111111111_1111111111111111_1101001011101001_1001111111000000"; -- -0.17612268025370545
	pesos_i(3975) := b"0000000000000000_0000000000000000_0010001000011011_1001101101001110"; -- 0.13323374425015075
	pesos_i(3976) := b"0000000000000000_0000000000000000_0001001010011110_0000110110100100"; -- 0.07272420164620359
	pesos_i(3977) := b"0000000000000000_0000000000000000_0000001000001010_0101100011100101"; -- 0.007970386451678222
	pesos_i(3978) := b"1111111111111111_1111111111111111_1110010100001011_1010101101001100"; -- -0.1052906932444959
	pesos_i(3979) := b"0000000000000000_0000000000000000_0001011010100001_1001100011010010"; -- 0.08840327392175845
	pesos_i(3980) := b"0000000000000000_0000000000000000_0010110010101010_1100100110111011"; -- 0.17448101820876336
	pesos_i(3981) := b"1111111111111111_1111111111111111_1110110110000110_0010111011100111"; -- -0.07217127661967884
	pesos_i(3982) := b"0000000000000000_0000000000000000_0010010000000001_0001101000111010"; -- 0.14064182205545409
	pesos_i(3983) := b"0000000000000000_0000000000000000_0001001001101110_0101100101100011"; -- 0.07199629461118648
	pesos_i(3984) := b"1111111111111111_1111111111111111_1111100010001110_1110100100111101"; -- -0.029069349892536844
	pesos_i(3985) := b"0000000000000000_0000000000000000_0001101100010110_0111001100110100"; -- 0.10581131007622396
	pesos_i(3986) := b"0000000000000000_0000000000000000_0001111110010000_0010011000110000"; -- 0.12329329171598498
	pesos_i(3987) := b"0000000000000000_0000000000000000_0000010111100111_0100110101011100"; -- 0.023060641352669716
	pesos_i(3988) := b"0000000000000000_0000000000000000_0000101110101110_0010101000001100"; -- 0.045626285533000875
	pesos_i(3989) := b"1111111111111111_1111111111111111_1111100011011110_0010011010111100"; -- -0.02786024009165144
	pesos_i(3990) := b"0000000000000000_0000000000000000_0010100101010000_0101101011001011"; -- 0.16138236490348828
	pesos_i(3991) := b"1111111111111111_1111111111111111_1111000111001010_1101110111110010"; -- -0.055498245688258424
	pesos_i(3992) := b"0000000000000000_0000000000000000_0000111001110001_0100001101100100"; -- 0.056415760044944814
	pesos_i(3993) := b"1111111111111111_1111111111111111_1101001011101001_0100111111001100"; -- -0.1761274459907886
	pesos_i(3994) := b"0000000000000000_0000000000000000_0001010101001110_0110100010100101"; -- 0.08322767292290563
	pesos_i(3995) := b"1111111111111111_1111111111111111_1110111100001001_1101010100011010"; -- -0.06625621911609748
	pesos_i(3996) := b"0000000000000000_0000000000000000_0000011101001111_1101011100011011"; -- 0.028562015550186923
	pesos_i(3997) := b"1111111111111111_1111111111111111_1101010101110110_1001111001111101"; -- -0.16615876632428964
	pesos_i(3998) := b"0000000000000000_0000000000000000_0001100010101100_0110110111000000"; -- 0.09638105331123582
	pesos_i(3999) := b"0000000000000000_0000000000000000_0000100110010110_1101111111000010"; -- 0.03745840529036851
	pesos_i(4000) := b"1111111111111111_1111111111111111_1111010110010000_0110100110101111"; -- -0.04076518504277504
	pesos_i(4001) := b"0000000000000000_0000000000000000_0010101001011100_0001011000000000"; -- 0.16546762000171028
	pesos_i(4002) := b"0000000000000000_0000000000000000_0010101000000010_0110000001000111"; -- 0.1640987562619658
	pesos_i(4003) := b"0000000000000000_0000000000000000_0001110110111101_0101010100100110"; -- 0.11617023626889864
	pesos_i(4004) := b"0000000000000000_0000000000000000_0010011001110101_0101011010011010"; -- 0.15022794022991814
	pesos_i(4005) := b"0000000000000000_0000000000000000_0001011001111110_1110100100101011"; -- 0.08787400539962112
	pesos_i(4006) := b"1111111111111111_1111111111111111_1101111111101001_0001111011111001"; -- -0.12534910608340696
	pesos_i(4007) := b"0000000000000000_0000000000000000_0000110110000000_0110111100001001"; -- 0.05274099314772179
	pesos_i(4008) := b"1111111111111111_1111111111111111_1101011110010110_0001111010011111"; -- -0.15786560640189565
	pesos_i(4009) := b"0000000000000000_0000000000000000_0000000111010000_1001001101100001"; -- 0.007088862619122554
	pesos_i(4010) := b"0000000000000000_0000000000000000_0000101101101100_1100011110000000"; -- 0.044628590262470964
	pesos_i(4011) := b"0000000000000000_0000000000000000_0010010001101110_0110110010100000"; -- 0.14230994145498777
	pesos_i(4012) := b"0000000000000000_0000000000000000_0001011001101101_1000011101100111"; -- 0.08760877858282644
	pesos_i(4013) := b"1111111111111111_1111111111111111_1111110001001001_1000000110001000"; -- -0.014503387715784228
	pesos_i(4014) := b"1111111111111111_1111111111111111_1110010000101010_1000101101111111"; -- -0.10872581622367151
	pesos_i(4015) := b"0000000000000000_0000000000000000_0010110000000000_1100010100000000"; -- 0.17188674203764595
	pesos_i(4016) := b"1111111111111111_1111111111111111_1111111000011110_0000010000111011"; -- -0.0073544842848466685
	pesos_i(4017) := b"0000000000000000_0000000000000000_0001000110110001_0111001001010111"; -- 0.06911387085716532
	pesos_i(4018) := b"0000000000000000_0000000000000000_0001110001110111_0011001100101010"; -- 0.111193845539978
	pesos_i(4019) := b"1111111111111111_1111111111111111_1101101000000011_0110111001111011"; -- -0.14838513856179336
	pesos_i(4020) := b"0000000000000000_0000000000000000_0000110110001011_0011111000000100"; -- 0.0529059181352795
	pesos_i(4021) := b"1111111111111111_1111111111111111_1111111000010111_0100100100001011"; -- -0.007457194233890458
	pesos_i(4022) := b"1111111111111111_1111111111111111_1101100110110110_1001000001000111"; -- -0.14955805090067026
	pesos_i(4023) := b"1111111111111111_1111111111111111_1110001100111010_0000101101010101"; -- -0.11239556484736273
	pesos_i(4024) := b"1111111111111111_1111111111111111_1101011100110100_0101110011011100"; -- -0.15935725811471763
	pesos_i(4025) := b"0000000000000000_0000000000000000_0000000111000000_0000001110111101"; -- 0.006836160385860021
	pesos_i(4026) := b"0000000000000000_0000000000000000_0000100010111011_1001010011100101"; -- 0.034112268251807465
	pesos_i(4027) := b"0000000000000000_0000000000000000_0001110011100110_1101110111011011"; -- 0.11289774512939094
	pesos_i(4028) := b"1111111111111111_1111111111111111_1101110110011110_1111110011100100"; -- -0.13429278776822695
	pesos_i(4029) := b"1111111111111111_1111111111111111_1111101011110101_1001011000001011"; -- -0.019690153496548877
	pesos_i(4030) := b"1111111111111111_1111111111111111_1101010111011000_0101110100001110"; -- -0.16466730502614785
	pesos_i(4031) := b"0000000000000000_0000000000000000_0000011100011011_1100011110101011"; -- 0.027767638527323273
	pesos_i(4032) := b"0000000000000000_0000000000000000_0000100111000101_1010111110111010"; -- 0.03817270556929481
	pesos_i(4033) := b"1111111111111111_1111111111111111_1111100011011010_1110111110000011"; -- -0.027909307971124044
	pesos_i(4034) := b"1111111111111111_1111111111111111_1111110100100010_1000011010110110"; -- -0.01119192188860912
	pesos_i(4035) := b"1111111111111111_1111111111111111_1111110101101000_0100111111110011"; -- -0.010127070685749955
	pesos_i(4036) := b"1111111111111111_1111111111111111_1111111000011000_0010001000001001"; -- -0.007444260435767958
	pesos_i(4037) := b"0000000000000000_0000000000000000_0001010001100000_0011111110100100"; -- 0.07959363703479248
	pesos_i(4038) := b"1111111111111111_1111111111111111_1111011010101100_1101010010010100"; -- -0.03642531766163946
	pesos_i(4039) := b"1111111111111111_1111111111111111_1110111111111111_0001100110000100"; -- -0.0625137379993646
	pesos_i(4040) := b"1111111111111111_1111111111111111_1101001111100111_0100011011110111"; -- -0.17225223995008837
	pesos_i(4041) := b"0000000000000000_0000000000000000_0000101010010100_1101110000110111"; -- 0.041333926651142223
	pesos_i(4042) := b"1111111111111111_1111111111111111_1110010111101001_0100110001100111"; -- -0.10190889817585576
	pesos_i(4043) := b"0000000000000000_0000000000000000_0010010101001011_0001010001001011"; -- 0.1456768686507179
	pesos_i(4044) := b"1111111111111111_1111111111111111_1111101100110110_0110101100100110"; -- -0.018700888860191296
	pesos_i(4045) := b"0000000000000000_0000000000000000_0001011010100011_0110011111101110"; -- 0.08843087730115926
	pesos_i(4046) := b"1111111111111111_1111111111111111_1101011111011110_0011100110101010"; -- -0.1567653617244356
	pesos_i(4047) := b"1111111111111111_1111111111111111_1101011111010000_1011000011101100"; -- -0.156971876408315
	pesos_i(4048) := b"0000000000000000_0000000000000000_0010001000100111_1010111100101110"; -- 0.13341803436384223
	pesos_i(4049) := b"1111111111111111_1111111111111111_1101100110011010_0010110010110110"; -- -0.14999123158297042
	pesos_i(4050) := b"0000000000000000_0000000000000000_0010001110101100_1000010101100110"; -- 0.13935121288228758
	pesos_i(4051) := b"1111111111111111_1111111111111111_1101110110100111_0110100100001101"; -- -0.13416427067133077
	pesos_i(4052) := b"0000000000000000_0000000000000000_0010001101010111_0001010010010011"; -- 0.13804749100633365
	pesos_i(4053) := b"0000000000000000_0000000000000000_0010010110111100_0101011111011000"; -- 0.14740513817856618
	pesos_i(4054) := b"1111111111111111_1111111111111111_1110101110010010_1110111110110001"; -- -0.07978918000604053
	pesos_i(4055) := b"1111111111111111_1111111111111111_1111011100000000_0100010110010010"; -- -0.03515210321552732
	pesos_i(4056) := b"1111111111111111_1111111111111111_1101111110011101_1000011011011100"; -- -0.12650258177773283
	pesos_i(4057) := b"0000000000000000_0000000000000000_0001011101000101_1101011100100110"; -- 0.09090943030549668
	pesos_i(4058) := b"0000000000000000_0000000000000000_0001011110100111_1110000100010100"; -- 0.09240538343760112
	pesos_i(4059) := b"0000000000000000_0000000000000000_0010101101110111_0001010011111110"; -- 0.1697857971764811
	pesos_i(4060) := b"0000000000000000_0000000000000000_0000000000001111_1001010010000000"; -- 0.00023773302080750327
	pesos_i(4061) := b"0000000000000000_0000000000000000_0000011101111110_1100010000000011"; -- 0.029278040636031656
	pesos_i(4062) := b"0000000000000000_0000000000000000_0001111111101001_1100101010111110"; -- 0.12466113216682188
	pesos_i(4063) := b"1111111111111111_1111111111111111_1110011001000101_1101110011001111"; -- -0.10049648233379198
	pesos_i(4064) := b"1111111111111111_1111111111111111_1101111100111101_1111101100011011"; -- -0.12796049677390509
	pesos_i(4065) := b"1111111111111111_1111111111111111_1111101101100011_0011011100101111"; -- -0.018017340615456026
	pesos_i(4066) := b"1111111111111111_1111111111111111_1111000001001000_0101110001111001"; -- -0.061395855403816695
	pesos_i(4067) := b"0000000000000000_0000000000000000_0001111110001001_0011100110101100"; -- 0.12318764159854745
	pesos_i(4068) := b"0000000000000000_0000000000000000_0001011100000111_0001111111111000"; -- 0.08995246700767992
	pesos_i(4069) := b"0000000000000000_0000000000000000_0001111010111011_0110010110011101"; -- 0.12004695009404641
	pesos_i(4070) := b"0000000000000000_0000000000000000_0001111110111010_1101010100100101"; -- 0.12394458911795679
	pesos_i(4071) := b"1111111111111111_1111111111111111_1111111010110111_0101110010011001"; -- -0.005014622237820482
	pesos_i(4072) := b"1111111111111111_1111111111111111_1110000100001100_1011011111110001"; -- -0.12089968085548833
	pesos_i(4073) := b"0000000000000000_0000000000000000_0001110100100110_1110101010001100"; -- 0.11387506398740177
	pesos_i(4074) := b"0000000000000000_0000000000000000_0010000111101010_0011111100000101"; -- 0.1324805630080751
	pesos_i(4075) := b"0000000000000000_0000000000000000_0000111111110100_1101111110010101"; -- 0.06233022099304452
	pesos_i(4076) := b"1111111111111111_1111111111111111_1110111001000101_1110101101011010"; -- -0.06924561551106226
	pesos_i(4077) := b"0000000000000000_0000000000000000_0001000110100111_0000111101001001"; -- 0.06895537879428752
	pesos_i(4078) := b"0000000000000000_0000000000000000_0001000101001010_0011111100111011"; -- 0.06753916912384353
	pesos_i(4079) := b"0000000000000000_0000000000000000_0011100001000011_0111110011000100"; -- 0.21977977548816716
	pesos_i(4080) := b"0000000000000000_0000000000000000_0001001110000011_1110010110000001"; -- 0.07623133094520748
	pesos_i(4081) := b"0000000000000000_0000000000000000_0001001001110110_0001111100010010"; -- 0.07211488907382649
	pesos_i(4082) := b"1111111111111111_1111111111111111_1110101111010000_1100101111000101"; -- -0.07884527629799572
	pesos_i(4083) := b"0000000000000000_0000000000000000_0010100110010100_1110001011011101"; -- 0.1624280728744495
	pesos_i(4084) := b"1111111111111111_1111111111111111_1101101011000111_0011010111101111"; -- -0.1453977863031806
	pesos_i(4085) := b"0000000000000000_0000000000000000_0001000110010111_1000111000111101"; -- 0.06871880513303057
	pesos_i(4086) := b"1111111111111111_1111111111111111_1101101100101001_1000100011110011"; -- -0.14389747693339855
	pesos_i(4087) := b"0000000000000000_0000000000000000_0010011001101010_1001110100010110"; -- 0.15006429476626243
	pesos_i(4088) := b"1111111111111111_1111111111111111_1111111111100010_0100110100110000"; -- -0.00045316302956813215
	pesos_i(4089) := b"0000000000000000_0000000000000000_0000111000111111_1010011010101110"; -- 0.05565873864972157
	pesos_i(4090) := b"1111111111111111_1111111111111111_1111111010011111_0011010101110010"; -- -0.00538316697935703
	pesos_i(4091) := b"1111111111111111_1111111111111111_1110110010010111_0100001000111100"; -- -0.07581697496373642
	pesos_i(4092) := b"1111111111111111_1111111111111111_1110000010011011_0000101000111111"; -- -0.12263427690133567
	pesos_i(4093) := b"1111111111111111_1111111111111111_1110111100101001_0101000001011111"; -- -0.06577584925612248
	pesos_i(4094) := b"0000000000000000_0000000000000000_0000101010101000_0101001010000000"; -- 0.04163089397195615
	pesos_i(4095) := b"1111111111111111_1111111111111111_1111100000111100_0000111111000011"; -- -0.030333533089360643
	pesos_i(4096) := b"0000000000000000_0000000000000000_0000101000000010_1011110001010010"; -- 0.03910424239805463
	pesos_i(4097) := b"0000000000000000_0000000000000000_0001011000111010_0001100110000011"; -- 0.08682403029023936
	pesos_i(4098) := b"1111111111111111_1111111111111111_1110010111010100_1111101011010010"; -- -0.10221893657169091
	pesos_i(4099) := b"0000000000000000_0000000000000000_0010001001111110_0011110001110101"; -- 0.13473871101505824
	pesos_i(4100) := b"0000000000000000_0000000000000000_0010100011001101_1011111101111000"; -- 0.15938946408803717
	pesos_i(4101) := b"1111111111111111_1111111111111111_1101100000111010_0000000001010110"; -- -0.1553649701763497
	pesos_i(4102) := b"0000000000000000_0000000000000000_0010100000101000_1001010000101111"; -- 0.1568691840983617
	pesos_i(4103) := b"1111111111111111_1111111111111111_1110100100000010_1000101011110111"; -- -0.08980494952445697
	pesos_i(4104) := b"0000000000000000_0000000000000000_0001100001011001_1001001110001000"; -- 0.09511682586170257
	pesos_i(4105) := b"1111111111111111_1111111111111111_1111001110000001_1110111011000011"; -- -0.048798634941239
	pesos_i(4106) := b"1111111111111111_1111111111111111_1111001011011011_1001101011010101"; -- -0.05133659640085577
	pesos_i(4107) := b"0000000000000000_0000000000000000_0010000111101111_1010011110111101"; -- 0.13256309855961756
	pesos_i(4108) := b"1111111111111111_1111111111111111_1111000011110101_0001110101101100"; -- -0.05875984300413465
	pesos_i(4109) := b"0000000000000000_0000000000000000_0001101000111100_0100111011001011"; -- 0.1024827238354471
	pesos_i(4110) := b"0000000000000000_0000000000000000_0001001011101100_0110011111101011"; -- 0.07391976821036068
	pesos_i(4111) := b"0000000000000000_0000000000000000_0000100101011001_1110100011000111"; -- 0.03652815694096329
	pesos_i(4112) := b"1111111111111111_1111111111111111_1110110011011100_0010111000111110"; -- -0.07476531004226844
	pesos_i(4113) := b"1111111111111111_1111111111111111_1110000110001101_1001100110010010"; -- -0.11893310717600383
	pesos_i(4114) := b"1111111111111111_1111111111111111_1101011010110001_0000000111100111"; -- -0.1613615810245976
	pesos_i(4115) := b"1111111111111111_1111111111111111_1101101110011101_0010100000000011"; -- -0.142133235273818
	pesos_i(4116) := b"1111111111111111_1111111111111111_1101100010000100_0100010100011100"; -- -0.15423172052790127
	pesos_i(4117) := b"0000000000000000_0000000000000000_0010011010101000_1000100010101110"; -- 0.15100912330244956
	pesos_i(4118) := b"0000000000000000_0000000000000000_0001111111010101_1111110001001001"; -- 0.12435890938479162
	pesos_i(4119) := b"0000000000000000_0000000000000000_0001011111101111_1101001001001101"; -- 0.09350313537411968
	pesos_i(4120) := b"0000000000000000_0000000000000000_0001000110010010_0001000111111100"; -- 0.06863510520558169
	pesos_i(4121) := b"0000000000000000_0000000000000000_0001010101000110_1000111010111011"; -- 0.08310787264966338
	pesos_i(4122) := b"1111111111111111_1111111111111111_1110010000111010_0010001110010001"; -- -0.10848787029974262
	pesos_i(4123) := b"0000000000000000_0000000000000000_0010000111001111_1101101011101010"; -- 0.13207786771180763
	pesos_i(4124) := b"1111111111111111_1111111111111111_1101101101101101_1000010011001000"; -- -0.14286012760591016
	pesos_i(4125) := b"0000000000000000_0000000000000000_0001011101011110_1100100101100101"; -- 0.09129008027497211
	pesos_i(4126) := b"0000000000000000_0000000000000000_0010100000101110_0100011011110110"; -- 0.15695613386027732
	pesos_i(4127) := b"0000000000000000_0000000000000000_0001010000011011_1010000111101111"; -- 0.07854663937173853
	pesos_i(4128) := b"0000000000000000_0000000000000000_0001101100100011_1011100110101111"; -- 0.10601387526496306
	pesos_i(4129) := b"0000000000000000_0000000000000000_0000110010101110_1101100101110100"; -- 0.049542990489316735
	pesos_i(4130) := b"1111111111111111_1111111111111111_1111101010110011_1000000101100101"; -- -0.020698464299919835
	pesos_i(4131) := b"1111111111111111_1111111111111111_1111101100010110_1111111100001000"; -- -0.019180355518364736
	pesos_i(4132) := b"1111111111111111_1111111111111111_1110111110000101_0110000101011110"; -- -0.06437102748768478
	pesos_i(4133) := b"0000000000000000_0000000000000000_0010000110001011_1000100110000100"; -- 0.1310354181795267
	pesos_i(4134) := b"0000000000000000_0000000000000000_0000010001001001_0111011011101111"; -- 0.016745980540445113
	pesos_i(4135) := b"0000000000000000_0000000000000000_0001011111011001_1111101100110001"; -- 0.09316987941270147
	pesos_i(4136) := b"1111111111111111_1111111111111111_1110001001001110_1000011101000111"; -- -0.11598925128836077
	pesos_i(4137) := b"1111111111111111_1111111111111111_1111100001001100_0100010011010000"; -- -0.030086230413178545
	pesos_i(4138) := b"1111111111111111_1111111111111111_1110111110000101_0011111000100011"; -- -0.0643731274228582
	pesos_i(4139) := b"0000000000000000_0000000000000000_0000001111010001_1111100110000000"; -- 0.014922708250457438
	pesos_i(4140) := b"1111111111111111_1111111111111111_1101010110000001_1000101000100011"; -- -0.16599213255621798
	pesos_i(4141) := b"1111111111111111_1111111111111111_1110011010101110_0110001001110110"; -- -0.09890160199907135
	pesos_i(4142) := b"1111111111111111_1111111111111111_1101010101101011_0111110111001010"; -- -0.1663285618783878
	pesos_i(4143) := b"0000000000000000_0000000000000000_0001100011111000_1111101011100111"; -- 0.0975491347043979
	pesos_i(4144) := b"0000000000000000_0000000000000000_0010010011100101_0111110111011101"; -- 0.1441267647887299
	pesos_i(4145) := b"1111111111111111_1111111111111111_1111010110011011_1011100101011110"; -- -0.040592588878849804
	pesos_i(4146) := b"1111111111111111_1111111111111111_1111011000111000_0011000010000011"; -- -0.038205116376768065
	pesos_i(4147) := b"0000000000000000_0000000000000000_0000011110100111_0011011100101001"; -- 0.02989525546096446
	pesos_i(4148) := b"0000000000000000_0000000000000000_0001011100001100_1011010110101000"; -- 0.09003768311382607
	pesos_i(4149) := b"1111111111111111_1111111111111111_1111011001100011_1000110010110010"; -- -0.03754349367288648
	pesos_i(4150) := b"0000000000000000_0000000000000000_0010101110000100_0011011001010101"; -- 0.169986148686158
	pesos_i(4151) := b"0000000000000000_0000000000000000_0000111010101001_1010001100101010"; -- 0.05727596063582538
	pesos_i(4152) := b"1111111111111111_1111111111111111_1111111100011111_0111000100001101"; -- -0.003426489128217608
	pesos_i(4153) := b"1111111111111111_1111111111111111_1111111100110001_1001110101111001"; -- -0.0031491833053203058
	pesos_i(4154) := b"0000000000000000_0000000000000000_0001001011001010_1111100110101101"; -- 0.0734096573296714
	pesos_i(4155) := b"1111111111111111_1111111111111111_1110110011100111_1000101000001010"; -- -0.07459199201360163
	pesos_i(4156) := b"1111111111111111_1111111111111111_1111010010001000_1010101001111101"; -- -0.044789642773893606
	pesos_i(4157) := b"0000000000000000_0000000000000000_0001011011101111_1101010001000010"; -- 0.08959700222710419
	pesos_i(4158) := b"0000000000000000_0000000000000000_0001101000001001_1001011110110101"; -- 0.10170887149698472
	pesos_i(4159) := b"0000000000000000_0000000000000000_0000100101111101_0101111001001010"; -- 0.0370692187296321
	pesos_i(4160) := b"1111111111111111_1111111111111111_1101101110011011_1110111110100101"; -- -0.14215185372676198
	pesos_i(4161) := b"0000000000000000_0000000000000000_0000100100000011_1111110101000100"; -- 0.03521712211736061
	pesos_i(4162) := b"0000000000000000_0000000000000000_0001110110100001_1100010000100111"; -- 0.11574960670265196
	pesos_i(4163) := b"1111111111111111_1111111111111111_1101110100010100_1100000100011001"; -- -0.13640206479973382
	pesos_i(4164) := b"0000000000000000_0000000000000000_0010000000111001_1011111011111001"; -- 0.12588113394083333
	pesos_i(4165) := b"0000000000000000_0000000000000000_0000001110110011_1010101110101011"; -- 0.014460305386168448
	pesos_i(4166) := b"1111111111111111_1111111111111111_1101110001100101_0100110000111010"; -- -0.13907931884047692
	pesos_i(4167) := b"0000000000000000_0000000000000000_0000010100111011_1011101010110000"; -- 0.020442645975508808
	pesos_i(4168) := b"0000000000000000_0000000000000000_0001101011110101_1011000111001100"; -- 0.10531150077509045
	pesos_i(4169) := b"1111111111111111_1111111111111111_1111111110010001_0010101100011001"; -- -0.001691156720377756
	pesos_i(4170) := b"0000000000000000_0000000000000000_0000001111010011_0101000000101001"; -- 0.014943132370749887
	pesos_i(4171) := b"1111111111111111_1111111111111111_1101110111011001_1110100011000000"; -- -0.13339371975788486
	pesos_i(4172) := b"1111111111111111_1111111111111111_1111001101010111_1001100101010011"; -- -0.04944459640790155
	pesos_i(4173) := b"1111111111111111_1111111111111111_1101110100111111_1110110110010110"; -- -0.1357432849622969
	pesos_i(4174) := b"1111111111111111_1111111111111111_1111110011111000_0010000110101000"; -- -0.011838814176185477
	pesos_i(4175) := b"1111111111111111_1111111111111111_1111111110100000_1111010001111100"; -- -0.0014502713844460119
	pesos_i(4176) := b"0000000000000000_0000000000000000_0001011111110101_0110110010110000"; -- 0.09358863163971307
	pesos_i(4177) := b"0000000000000000_0000000000000000_0001000111000110_0100011001001101"; -- 0.0694316805704778
	pesos_i(4178) := b"1111111111111111_1111111111111111_1101011010110000_0101101010010011"; -- -0.1613715544217255
	pesos_i(4179) := b"0000000000000000_0000000000000000_0010000111001000_1000001000011001"; -- 0.13196576223217693
	pesos_i(4180) := b"1111111111111111_1111111111111111_1101111000011011_0011110000101100"; -- -0.13239692618067672
	pesos_i(4181) := b"1111111111111111_1111111111111111_1101010110101000_1110011010011100"; -- -0.1653915280519862
	pesos_i(4182) := b"0000000000000000_0000000000000000_0010111110111000_1011101100011011"; -- 0.18641251965472735
	pesos_i(4183) := b"0000000000000000_0000000000000000_0010110010100010_0011010100110111"; -- 0.17435009570904453
	pesos_i(4184) := b"1111111111111111_1111111111111111_1111000100100110_0010110010010010"; -- -0.05801125934016683
	pesos_i(4185) := b"0000000000000000_0000000000000000_0001000100100110_0001111010101010"; -- 0.06698791159734967
	pesos_i(4186) := b"0000000000000000_0000000000000000_0010101111101110_1100000101011010"; -- 0.17161186643855275
	pesos_i(4187) := b"1111111111111111_1111111111111111_1111100101110111_0111110101111101"; -- -0.025520474365765808
	pesos_i(4188) := b"0000000000000000_0000000000000000_0000001001000010_1011110010110010"; -- 0.008830827302656026
	pesos_i(4189) := b"1111111111111111_1111111111111111_1110100101100101_1000001010110011"; -- -0.08829482201836111
	pesos_i(4190) := b"0000000000000000_0000000000000000_0001110001010000_0010010110001011"; -- 0.110597940880021
	pesos_i(4191) := b"1111111111111111_1111111111111111_1110110001111100_1000111011101110"; -- -0.07622439099720506
	pesos_i(4192) := b"1111111111111111_1111111111111111_1101010011000100_1001101111111110"; -- -0.1688749793752347
	pesos_i(4193) := b"1111111111111111_1111111111111111_1101010110010110_1100011000000010"; -- -0.16566812934937805
	pesos_i(4194) := b"0000000000000000_0000000000000000_0001000000010111_1010001100001010"; -- 0.06286066992255379
	pesos_i(4195) := b"1111111111111111_1111111111111111_1110011001011001_1000110001000011"; -- -0.10019610754406841
	pesos_i(4196) := b"1111111111111111_1111111111111111_1111010000000001_0101010101100011"; -- -0.046854651716846545
	pesos_i(4197) := b"0000000000000000_0000000000000000_0010011101101111_1011111010011001"; -- 0.1540488360846076
	pesos_i(4198) := b"0000000000000000_0000000000000000_0010001001101000_1011001011100010"; -- 0.13441007628134508
	pesos_i(4199) := b"1111111111111111_1111111111111111_1111001010000010_1000101010111111"; -- -0.05269558757230053
	pesos_i(4200) := b"0000000000000000_0000000000000000_0001000010010110_1011001101110011"; -- 0.06479951425599087
	pesos_i(4201) := b"1111111111111111_1111111111111111_1110100100110010_0101100100010001"; -- -0.08907550181153574
	pesos_i(4202) := b"0000000000000000_0000000000000000_0001100001010000_0000110010100101"; -- 0.09497145681698983
	pesos_i(4203) := b"0000000000000000_0000000000000000_0000111100000111_0111010000110100"; -- 0.058707487774395876
	pesos_i(4204) := b"0000000000000000_0000000000000000_0001100100011100_0010100011001000"; -- 0.09808592695613909
	pesos_i(4205) := b"1111111111111111_1111111111111111_1110000110110111_1110011111011101"; -- -0.1182875715552376
	pesos_i(4206) := b"1111111111111111_1111111111111111_1110111011010111_1100110111010100"; -- -0.06701959211801664
	pesos_i(4207) := b"0000000000000000_0000000000000000_0001101110110000_0011000001110001"; -- 0.10815718413933083
	pesos_i(4208) := b"0000000000000000_0000000000000000_0010011110101000_1011011110111110"; -- 0.15491817846544717
	pesos_i(4209) := b"1111111111111111_1111111111111111_1111001101001110_0110111001010001"; -- -0.04958448918036921
	pesos_i(4210) := b"1111111111111111_1111111111111111_1110000100111000_0101111011101100"; -- -0.12023360011044953
	pesos_i(4211) := b"0000000000000000_0000000000000000_0010000001000000_0100001010001111"; -- 0.1259805296870197
	pesos_i(4212) := b"1111111111111111_1111111111111111_1110001001111001_1001101100011011"; -- -0.11533194141292741
	pesos_i(4213) := b"0000000000000000_0000000000000000_0000000011101001_1010000101011100"; -- 0.0035649156760938962
	pesos_i(4214) := b"1111111111111111_1111111111111111_1101001111111011_0111110000111110"; -- -0.17194388850688921
	pesos_i(4215) := b"0000000000000000_0000000000000000_0000010000001110_1011011100010101"; -- 0.01584953555570208
	pesos_i(4216) := b"1111111111111111_1111111111111111_1111110100010001_0101101001011010"; -- -0.011453965117524861
	pesos_i(4217) := b"1111111111111111_1111111111111111_1101111000001111_1111010101111001"; -- -0.1325689869043223
	pesos_i(4218) := b"1111111111111111_1111111111111111_1111011111011000_1101110101000001"; -- -0.03184716369118145
	pesos_i(4219) := b"1111111111111111_1111111111111111_1111101111000101_1101000111110110"; -- -0.01651275398647466
	pesos_i(4220) := b"1111111111111111_1111111111111111_1101101101000000_1110101111100010"; -- -0.1435406278023961
	pesos_i(4221) := b"0000000000000000_0000000000000000_0000000001100011_0110011001010101"; -- 0.0015167196075503648
	pesos_i(4222) := b"0000000000000000_0000000000000000_0001001011100100_0001011111110111"; -- 0.0737929324031568
	pesos_i(4223) := b"0000000000000000_0000000000000000_0001001011000011_0000100010000110"; -- 0.07328847180610722
	pesos_i(4224) := b"0000000000000000_0000000000000000_0001100100001011_0111110010011111"; -- 0.09783152474352477
	pesos_i(4225) := b"0000000000000000_0000000000000000_0000011110010101_0101010011011001"; -- 0.029622366946106825
	pesos_i(4226) := b"1111111111111111_1111111111111111_1101111100010011_1011001111111110"; -- -0.12860560452970762
	pesos_i(4227) := b"1111111111111111_1111111111111111_1111111001010010_0101000000000110"; -- -0.006556509594702516
	pesos_i(4228) := b"0000000000000000_0000000000000000_0010100001111110_1011111111000011"; -- 0.15818403727071179
	pesos_i(4229) := b"1111111111111111_1111111111111111_1111001010101010_0101000011011100"; -- -0.052088686362924
	pesos_i(4230) := b"1111111111111111_1111111111111111_1101101110110000_0010001111000101"; -- -0.14184357116581417
	pesos_i(4231) := b"0000000000000000_0000000000000000_0001001110111110_1000111000101000"; -- 0.0771263930354168
	pesos_i(4232) := b"0000000000000000_0000000000000000_0000000010110100_1011110111110101"; -- 0.0027579043444387434
	pesos_i(4233) := b"0000000000000000_0000000000000000_0010011101110110_0101011000000001"; -- 0.1541494133443268
	pesos_i(4234) := b"0000000000000000_0000000000000000_0000111111100010_0010110011011100"; -- 0.062044910205388284
	pesos_i(4235) := b"0000000000000000_0000000000000000_0001110010110101_0001101101100010"; -- 0.11213847288084448
	pesos_i(4236) := b"1111111111111111_1111111111111111_1111010011110001_0101001001011111"; -- -0.043192722137925924
	pesos_i(4237) := b"1111111111111111_1111111111111111_1101011110110001_0001111011011101"; -- -0.1574536048255472
	pesos_i(4238) := b"0000000000000000_0000000000000000_0000110100110101_0011110001010010"; -- 0.051593561252255
	pesos_i(4239) := b"0000000000000000_0000000000000000_0000000100100101_0001101111110011"; -- 0.004472491051746189
	pesos_i(4240) := b"1111111111111111_1111111111111111_1101011010011010_1111101110101001"; -- -0.16169764638195638
	pesos_i(4241) := b"0000000000000000_0000000000000000_0000010000001100_1000001001100101"; -- 0.015815877686822306
	pesos_i(4242) := b"1111111111111111_1111111111111111_1111100110100011_0100000101001111"; -- -0.02485267468303782
	pesos_i(4243) := b"1111111111111111_1111111111111111_1111001000110101_0011000111010100"; -- -0.05387581425494147
	pesos_i(4244) := b"1111111111111111_1111111111111111_1101100111000101_1100001000011011"; -- -0.14932619890691237
	pesos_i(4245) := b"1111111111111111_1111111111111111_1101111101010000_0010111111010011"; -- -0.12768269635764332
	pesos_i(4246) := b"0000000000000000_0000000000000000_0001100000111110_0001111100011001"; -- 0.0946978984306325
	pesos_i(4247) := b"0000000000000000_0000000000000000_0000101011010000_0101100001100010"; -- 0.04224159614797522
	pesos_i(4248) := b"0000000000000000_0000000000000000_0001111111100001_0110010110100010"; -- 0.12453303526683647
	pesos_i(4249) := b"0000000000000000_0000000000000000_0010000000001000_0111001011100001"; -- 0.12512891765268436
	pesos_i(4250) := b"0000000000000000_0000000000000000_0001010100110001_1001000111100111"; -- 0.08278762702309456
	pesos_i(4251) := b"1111111111111111_1111111111111111_1110000001010001_0000101101001111"; -- -0.12376336393463322
	pesos_i(4252) := b"1111111111111111_1111111111111111_1110010110110011_1101111111101110"; -- -0.10272407957843745
	pesos_i(4253) := b"0000000000000000_0000000000000000_0001111100001100_1101011100001111"; -- 0.121289673939645
	pesos_i(4254) := b"1111111111111111_1111111111111111_1110100111110100_1010100000100101"; -- -0.08611058329447417
	pesos_i(4255) := b"1111111111111111_1111111111111111_1111100011101011_1011001101110011"; -- -0.027653488456851144
	pesos_i(4256) := b"0000000000000000_0000000000000000_0001000011000000_1001011001000110"; -- 0.06543864443334182
	pesos_i(4257) := b"1111111111111111_1111111111111111_1110010010010001_0111101010011001"; -- -0.10715516827298587
	pesos_i(4258) := b"0000000000000000_0000000000000000_0001110110010100_1100010110000000"; -- 0.11555132269129542
	pesos_i(4259) := b"1111111111111111_1111111111111111_1110100001111001_0010101000110011"; -- -0.09190117116138852
	pesos_i(4260) := b"1111111111111111_1111111111111111_1110101111000000_0010100110010011"; -- -0.07909908457076154
	pesos_i(4261) := b"1111111111111111_1111111111111111_1101100000111011_1101000011000110"; -- -0.15533728757413096
	pesos_i(4262) := b"1111111111111111_1111111111111111_1111101011011110_1000000101100001"; -- -0.02004233715947736
	pesos_i(4263) := b"0000000000000000_0000000000000000_0010000011100000_0110010010000100"; -- 0.1284239600433776
	pesos_i(4264) := b"0000000000000000_0000000000000000_0001000011100000_0110100110101101"; -- 0.06592426746824187
	pesos_i(4265) := b"1111111111111111_1111111111111111_1111100111110100_0101110000000011"; -- -0.023615121208810916
	pesos_i(4266) := b"1111111111111111_1111111111111111_1101110000010011_0000100011000010"; -- -0.14033456100195982
	pesos_i(4267) := b"0000000000000000_0000000000000000_0000100111000010_0110000000100010"; -- 0.03812218510524642
	pesos_i(4268) := b"1111111111111111_1111111111111111_1101110001100110_1101100011000011"; -- -0.13905568359311354
	pesos_i(4269) := b"0000000000000000_0000000000000000_0010000000100110_0000100000000111"; -- 0.12558031243985998
	pesos_i(4270) := b"1111111111111111_1111111111111111_1110010000000110_0101101010101000"; -- -0.10927804383699428
	pesos_i(4271) := b"1111111111111111_1111111111111111_1110011110011000_0100001000001010"; -- -0.09533297780243992
	pesos_i(4272) := b"1111111111111111_1111111111111111_1111100111000010_0111110010100001"; -- -0.024376116479734755
	pesos_i(4273) := b"1111111111111111_1111111111111111_1110111001010001_0001101000000000"; -- -0.0690749883144314
	pesos_i(4274) := b"0000000000000000_0000000000000000_0001010110101101_0011000000000101"; -- 0.08467388270496368
	pesos_i(4275) := b"1111111111111111_1111111111111111_1101111000111101_0000001001110000"; -- -0.13188156865728834
	pesos_i(4276) := b"0000000000000000_0000000000000000_0001100010001110_1100011111010001"; -- 0.09592865814630186
	pesos_i(4277) := b"1111111111111111_1111111111111111_1111110011000110_0000110000110101"; -- -0.012603032059511006
	pesos_i(4278) := b"0000000000000000_0000000000000000_0010101011001100_0101111011100000"; -- 0.16718094806949352
	pesos_i(4279) := b"1111111111111111_1111111111111111_1110100110100110_1001001001011101"; -- -0.08730206714591955
	pesos_i(4280) := b"0000000000000000_0000000000000000_0010100110110010_0101010010101001"; -- 0.1628773605585794
	pesos_i(4281) := b"1111111111111111_1111111111111111_1110011101000001_0010010100011010"; -- -0.09666221739515296
	pesos_i(4282) := b"0000000000000000_0000000000000000_0010100111010110_0011000000101100"; -- 0.16342450207260548
	pesos_i(4283) := b"0000000000000000_0000000000000000_0000001100010011_1110100101000000"; -- 0.012022569821711087
	pesos_i(4284) := b"1111111111111111_1111111111111111_1110011101000111_1000000111011000"; -- -0.0965651366325623
	pesos_i(4285) := b"0000000000000000_0000000000000000_0001000110011101_0111110011111000"; -- 0.06880932853455647
	pesos_i(4286) := b"1111111111111111_1111111111111111_1101101000010111_1110000110011000"; -- -0.1480731014748874
	pesos_i(4287) := b"0000000000000000_0000000000000000_0001101011110111_1101101001101101"; -- 0.10534444004958077
	pesos_i(4288) := b"1111111111111111_1111111111111111_1110101010110010_0111111011110010"; -- -0.08321386902484176
	pesos_i(4289) := b"1111111111111111_1111111111111111_1111101101111111_0100101001110001"; -- -0.017588946743478277
	pesos_i(4290) := b"0000000000000000_0000000000000000_0000011111110110_0011011101001111"; -- 0.031100708736451814
	pesos_i(4291) := b"0000000000000000_0000000000000000_0000111110100100_1111011000100100"; -- 0.06111086247886095
	pesos_i(4292) := b"1111111111111111_1111111111111111_1101011010000001_0100101001000011"; -- -0.16208968980125948
	pesos_i(4293) := b"1111111111111111_1111111111111111_1110110101111010_1101011110010100"; -- -0.07234432834423504
	pesos_i(4294) := b"0000000000000000_0000000000000000_0010011101010100_0111001100100001"; -- 0.15363235042000944
	pesos_i(4295) := b"1111111111111111_1111111111111111_1110101001010100_0000001100011001"; -- -0.08465557707651196
	pesos_i(4296) := b"0000000000000000_0000000000000000_0011101100100010_0001001101010011"; -- 0.2309887006916392
	pesos_i(4297) := b"0000000000000000_0000000000000000_0000101101010111_1011101101000000"; -- 0.04430742569022793
	pesos_i(4298) := b"1111111111111111_1111111111111111_1101101000100100_1111110011110001"; -- -0.14787310717047297
	pesos_i(4299) := b"0000000000000000_0000000000000000_0010000010111111_1001011100000111"; -- 0.12792343059630326
	pesos_i(4300) := b"0000000000000000_0000000000000000_0000100010110000_0100100101110111"; -- 0.033939925703436125
	pesos_i(4301) := b"0000000000000000_0000000000000000_0001101011110011_0101001101100110"; -- 0.10527535670366805
	pesos_i(4302) := b"0000000000000000_0000000000000000_0001010100110100_0001111111100000"; -- 0.0828266069396084
	pesos_i(4303) := b"0000000000000000_0000000000000000_0001100101110101_0101101110110111"; -- 0.09944699485274336
	pesos_i(4304) := b"0000000000000000_0000000000000000_0001000011101001_1101001110101111"; -- 0.06606791525687042
	pesos_i(4305) := b"1111111111111111_1111111111111111_1101111100011110_1010011101111001"; -- -0.128438504096028
	pesos_i(4306) := b"1111111111111111_1111111111111111_1110111010111000_0000001110011100"; -- -0.06750466772606578
	pesos_i(4307) := b"1111111111111111_1111111111111111_1110110000010101_1010000111111111"; -- -0.07779490961214176
	pesos_i(4308) := b"1111111111111111_1111111111111111_1111011101100011_0000110010111110"; -- -0.033644870335184346
	pesos_i(4309) := b"0000000000000000_0000000000000000_0010011001110000_1000110101001110"; -- 0.1501549067375712
	pesos_i(4310) := b"1111111111111111_1111111111111111_1111000000010100_0101100101011110"; -- -0.062189497416389336
	pesos_i(4311) := b"0000000000000000_0000000000000000_0001111011101011_0101000010010001"; -- 0.12077811754365379
	pesos_i(4312) := b"0000000000000000_0000000000000000_0010100110000110_1110110001100110"; -- 0.16221501823136777
	pesos_i(4313) := b"1111111111111111_1111111111111111_1101111110011000_1001110101011011"; -- -0.12657753491881985
	pesos_i(4314) := b"1111111111111111_1111111111111111_1110011111111111_0100101110110000"; -- -0.09376074737696237
	pesos_i(4315) := b"1111111111111111_1111111111111111_1111010011010010_1001110001111110"; -- -0.04366132674062566
	pesos_i(4316) := b"0000000000000000_0000000000000000_0010010010101011_1100001100100000"; -- 0.1432458831896586
	pesos_i(4317) := b"0000000000000000_0000000000000000_0010000111111000_1011000100110000"; -- 0.13270099092885032
	pesos_i(4318) := b"0000000000000000_0000000000000000_0001110010000110_1110111111001011"; -- 0.11143397045213675
	pesos_i(4319) := b"0000000000000000_0000000000000000_0000111000011111_1000111010010110"; -- 0.055169021305017524
	pesos_i(4320) := b"0000000000000000_0000000000000000_0010000010001100_0100110110010001"; -- 0.12714085374540032
	pesos_i(4321) := b"0000000000000000_0000000000000000_0001101111010000_1011000101100011"; -- 0.10865315125893249
	pesos_i(4322) := b"0000000000000000_0000000000000000_0010011111010100_0001101010100010"; -- 0.15558020077008233
	pesos_i(4323) := b"0000000000000000_0000000000000000_0001000000110010_0011111011100010"; -- 0.0632666876017102
	pesos_i(4324) := b"0000000000000000_0000000000000000_0000100100001101_1101010100110000"; -- 0.03536732119347782
	pesos_i(4325) := b"0000000000000000_0000000000000000_0000101101000010_1101011010000010"; -- 0.04398861564670951
	pesos_i(4326) := b"1111111111111111_1111111111111111_1101100001101110_1001010111010010"; -- -0.15456260318103482
	pesos_i(4327) := b"0000000000000000_0000000000000000_0010101000100110_0001111011101111"; -- 0.16464417788584787
	pesos_i(4328) := b"0000000000000000_0000000000000000_0000111000100101_1110110101111011"; -- 0.0552662302297329
	pesos_i(4329) := b"0000000000000000_0000000000000000_0000000010001101_0010010000000010"; -- 0.0021536354399051116
	pesos_i(4330) := b"1111111111111111_1111111111111111_1101010001010010_1101110110000000"; -- -0.17061057686621586
	pesos_i(4331) := b"1111111111111111_1111111111111111_1110010111111111_1101111111000000"; -- -0.10156442217082515
	pesos_i(4332) := b"0000000000000000_0000000000000000_0010100010001000_0010001110100111"; -- 0.1583273202942278
	pesos_i(4333) := b"1111111111111111_1111111111111111_1111010001111001_1000111111011111"; -- -0.045020111252791005
	pesos_i(4334) := b"1111111111111111_1111111111111111_1101011101011110_1101100010000111"; -- -0.15870901778978092
	pesos_i(4335) := b"1111111111111111_1111111111111111_1101101111111110_1110101100101101"; -- -0.1406415001138053
	pesos_i(4336) := b"1111111111111111_1111111111111111_1101011011001001_0101000110100010"; -- -0.16099061763611963
	pesos_i(4337) := b"1111111111111111_1111111111111111_1101111111111111_0000101110110000"; -- -0.12501456218317544
	pesos_i(4338) := b"1111111111111111_1111111111111111_1111100001000110_0111001010000000"; -- -0.03017506014608607
	pesos_i(4339) := b"1111111111111111_1111111111111111_1101001110100111_1101010010010011"; -- -0.17322036190977058
	pesos_i(4340) := b"0000000000000000_0000000000000000_0001101000010000_0110001000111101"; -- 0.10181249602753473
	pesos_i(4341) := b"1111111111111111_1111111111111111_1111001001011101_0100000001111110"; -- -0.05326458861400679
	pesos_i(4342) := b"1111111111111111_1111111111111111_1110111011100001_1000010100001000"; -- -0.06687134309490748
	pesos_i(4343) := b"1111111111111111_1111111111111111_1101000101110011_1111001100010001"; -- -0.1818245013029572
	pesos_i(4344) := b"1111111111111111_1111111111111111_1111010101001110_1010111101010011"; -- -0.04176811421959856
	pesos_i(4345) := b"1111111111111111_1111111111111111_1110111101100000_0110111010100010"; -- -0.0649348120600893
	pesos_i(4346) := b"1111111111111111_1111111111111111_1110111111100001_1001101111111000"; -- -0.0629637259777984
	pesos_i(4347) := b"0000000000000000_0000000000000000_0000010100111010_1010010110100110"; -- 0.020426133100627866
	pesos_i(4348) := b"0000000000000000_0000000000000000_0000011011010011_0111001010000100"; -- 0.026663930103715077
	pesos_i(4349) := b"1111111111111111_1111111111111111_1110011000111011_0110001010011110"; -- -0.10065635346378957
	pesos_i(4350) := b"0000000000000000_0000000000000000_0001100011010101_0100110001000010"; -- 0.09700466750063219
	pesos_i(4351) := b"1111111111111111_1111111111111111_1111001010100000_1111000100110101"; -- -0.05223171658708871
	pesos_i(4352) := b"1111111111111111_1111111111111111_1110101110000101_0000110001010011"; -- -0.08000109656558532
	pesos_i(4353) := b"0000000000000000_0000000000000000_0001110100110011_1010011111101010"; -- 0.11406945675086849
	pesos_i(4354) := b"1111111111111111_1111111111111111_1111000101000101_0101011000011001"; -- -0.05753576169429388
	pesos_i(4355) := b"0000000000000000_0000000000000000_0010101110111010_0101100010101111"; -- 0.170812170811528
	pesos_i(4356) := b"0000000000000000_0000000000000000_0000101001100101_0010011000011111"; -- 0.040605909787296675
	pesos_i(4357) := b"0000000000000000_0000000000000000_0010000010010001_1111100000110110"; -- 0.127227319022834
	pesos_i(4358) := b"1111111111111111_1111111111111111_1111110101100010_0010111110001000"; -- -0.010220555472809967
	pesos_i(4359) := b"0000000000000000_0000000000000000_0001011101011101_0101110100111100"; -- 0.09126837453519206
	pesos_i(4360) := b"0000000000000000_0000000000000000_0000110100011000_1000101001101010"; -- 0.05115571104773546
	pesos_i(4361) := b"0000000000000000_0000000000000000_0000001101110101_1110100111001001"; -- 0.0135179630037753
	pesos_i(4362) := b"1111111111111111_1111111111111111_1110001010111000_1100001110111110"; -- -0.1143682155547708
	pesos_i(4363) := b"1111111111111111_1111111111111111_1110011000110110_0100000000101001"; -- -0.10073470124944184
	pesos_i(4364) := b"0000000000000000_0000000000000000_0000111011011110_0001111010101110"; -- 0.05807677984557293
	pesos_i(4365) := b"0000000000000000_0000000000000000_0001100011010001_1001001010111101"; -- 0.09694783319333371
	pesos_i(4366) := b"1111111111111111_1111111111111111_1101110010011011_1011001001000000"; -- -0.13824926319585104
	pesos_i(4367) := b"1111111111111111_1111111111111111_1111001000011101_1011011001000111"; -- -0.054234130651542645
	pesos_i(4368) := b"0000000000000000_0000000000000000_0010100010001010_1011011001111100"; -- 0.15836658971503778
	pesos_i(4369) := b"1111111111111111_1111111111111111_1111100101001101_0011110111111010"; -- -0.026165129254247743
	pesos_i(4370) := b"1111111111111111_1111111111111111_1111011101110001_0101010101010110"; -- -0.033426920328391126
	pesos_i(4371) := b"1111111111111111_1111111111111111_1111111010010100_0100000111111101"; -- -0.0055502660549806735
	pesos_i(4372) := b"0000000000000000_0000000000000000_0000000110111011_1110100100111110"; -- 0.006773545908259159
	pesos_i(4373) := b"0000000000000000_0000000000000000_0001101011010000_1000111101011001"; -- 0.10474487241248782
	pesos_i(4374) := b"1111111111111111_1111111111111111_1111001100101000_1110111110011111"; -- -0.05015661599545416
	pesos_i(4375) := b"1111111111111111_1111111111111111_1111101100101011_0100011110111011"; -- -0.018870846487435658
	pesos_i(4376) := b"0000000000000000_0000000000000000_0001001011010111_0110110100110001"; -- 0.07359964804643938
	pesos_i(4377) := b"1111111111111111_1111111111111111_1110100001011110_0011010101111100"; -- -0.0923124859868806
	pesos_i(4378) := b"1111111111111111_1111111111111111_1111001101101010_1111100110110011"; -- -0.04914893509684047
	pesos_i(4379) := b"0000000000000000_0000000000000000_0000001011101101_1001110011101111"; -- 0.01143818699450293
	pesos_i(4380) := b"1111111111111111_1111111111111111_1111011110111010_1101100000110101"; -- -0.03230522834702052
	pesos_i(4381) := b"0000000000000000_0000000000000000_0001001011000110_0000000110011110"; -- 0.07333383657387436
	pesos_i(4382) := b"0000000000000000_0000000000000000_0001111110101000_1000000110101001"; -- 0.12366495495165142
	pesos_i(4383) := b"1111111111111111_1111111111111111_1111111000101010_0101011111000111"; -- -0.007166399001276136
	pesos_i(4384) := b"1111111111111111_1111111111111111_1110010111000010_0101110101001101"; -- -0.10250298369021091
	pesos_i(4385) := b"0000000000000000_0000000000000000_0000000001101011_1110010110010110"; -- 0.0016463749153689334
	pesos_i(4386) := b"0000000000000000_0000000000000000_0010011001101101_0101010100101110"; -- 0.15010578522199072
	pesos_i(4387) := b"1111111111111111_1111111111111111_1111000101100111_0110010000011010"; -- -0.05701612820474538
	pesos_i(4388) := b"1111111111111111_1111111111111111_1111111111110100_1101111101010010"; -- -0.00016979442921710684
	pesos_i(4389) := b"1111111111111111_1111111111111111_1111101100010010_0000101000101101"; -- -0.019255985306109592
	pesos_i(4390) := b"0000000000000000_0000000000000000_0001011101000110_1000101110111101"; -- 0.0909201942903363
	pesos_i(4391) := b"0000000000000000_0000000000000000_0010001100000111_0010000111010111"; -- 0.13682757844397855
	pesos_i(4392) := b"1111111111111111_1111111111111111_1110101110010001_1010100001010101"; -- -0.07980869225077172
	pesos_i(4393) := b"0000000000000000_0000000000000000_0010010100001011_1110101110100010"; -- 0.14471314149389153
	pesos_i(4394) := b"1111111111111111_1111111111111111_1111000000110110_0001101100010000"; -- -0.06167441243052004
	pesos_i(4395) := b"0000000000000000_0000000000000000_0010100010011111_0000100111100000"; -- 0.1586767360401631
	pesos_i(4396) := b"1111111111111111_1111111111111111_1110100111110001_0011011110001001"; -- -0.0861630715751664
	pesos_i(4397) := b"0000000000000000_0000000000000000_0001000101110110_1101000001110110"; -- 0.0682192123438233
	pesos_i(4398) := b"0000000000000000_0000000000000000_0010010000011110_1011001111111000"; -- 0.14109349065674795
	pesos_i(4399) := b"0000000000000000_0000000000000000_0010001001100001_0110110010001001"; -- 0.1342990717622932
	pesos_i(4400) := b"1111111111111111_1111111111111111_1111100111000001_1011101001111000"; -- -0.02438768941721986
	pesos_i(4401) := b"1111111111111111_1111111111111111_1110101101010001_0000010110100011"; -- -0.08079495210124053
	pesos_i(4402) := b"0000000000000000_0000000000000000_0001101111010000_0101010011001111"; -- 0.10864763304602973
	pesos_i(4403) := b"0000000000000000_0000000000000000_0000101101100101_1101010011100010"; -- 0.04452257651474128
	pesos_i(4404) := b"0000000000000000_0000000000000000_0001010011101110_0011100100101110"; -- 0.08175999987955056
	pesos_i(4405) := b"0000000000000000_0000000000000000_0000001011110110_1010110100001010"; -- 0.011576476146151872
	pesos_i(4406) := b"1111111111111111_1111111111111111_1101100000111100_1010110011011111"; -- -0.15532416883111144
	pesos_i(4407) := b"1111111111111111_1111111111111111_1110101000010010_1110110101000111"; -- -0.08564869899849135
	pesos_i(4408) := b"0000000000000000_0000000000000000_0010001011000100_0110001100001111"; -- 0.13580912710694962
	pesos_i(4409) := b"0000000000000000_0000000000000000_0001001000111000_0101000100111001"; -- 0.07117183332495036
	pesos_i(4410) := b"0000000000000000_0000000000000000_0001100011110101_1111100001111111"; -- 0.09750321493288451
	pesos_i(4411) := b"1111111111111111_1111111111111111_1111000000111101_0111001001110011"; -- -0.06156239213843668
	pesos_i(4412) := b"1111111111111111_1111111111111111_1110110000111111_1110100100110010"; -- -0.07714979666562585
	pesos_i(4413) := b"0000000000000000_0000000000000000_0001111011101010_1000000011001000"; -- 0.12076573261662112
	pesos_i(4414) := b"1111111111111111_1111111111111111_1110111101000011_1001110011101110"; -- -0.0653745573487203
	pesos_i(4415) := b"0000000000000000_0000000000000000_0001110010100110_1010010001101010"; -- 0.1119177588638116
	pesos_i(4416) := b"0000000000000000_0000000000000000_0000000010011010_0101011000101010"; -- 0.0023549892530469185
	pesos_i(4417) := b"0000000000000000_0000000000000000_0000000111011110_1110100110000000"; -- 0.007307618887662182
	pesos_i(4418) := b"0000000000000000_0000000000000000_0001111010011001_1101110110101011"; -- 0.11953530718068371
	pesos_i(4419) := b"0000000000000000_0000000000000000_0001011111111001_1111001101000100"; -- 0.09365768814924096
	pesos_i(4420) := b"0000000000000000_0000000000000000_0001100111010000_0001111001101011"; -- 0.10083189113815139
	pesos_i(4421) := b"1111111111111111_1111111111111111_1110010101001111_1001100110010100"; -- -0.10425415162271605
	pesos_i(4422) := b"1111111111111111_1111111111111111_1110110100101110_1111111010100101"; -- -0.07350166765039352
	pesos_i(4423) := b"0000000000000000_0000000000000000_0000110110000100_1110111111111001"; -- 0.052809713624771645
	pesos_i(4424) := b"1111111111111111_1111111111111111_1111110001011011_0110110110110110"; -- -0.014229910971426393
	pesos_i(4425) := b"0000000000000000_0000000000000000_0000101010011110_1011100000101110"; -- 0.041484366749581315
	pesos_i(4426) := b"1111111111111111_1111111111111111_1101111101001001_0010010111111101"; -- -0.1277900941996216
	pesos_i(4427) := b"1111111111111111_1111111111111111_1101010100110000_1011111001111101"; -- -0.16722497403724593
	pesos_i(4428) := b"1111111111111111_1111111111111111_1101100001000110_0001000011010001"; -- -0.1551808824086396
	pesos_i(4429) := b"1111111111111111_1111111111111111_1111011010110011_0010010011100111"; -- -0.03632897728115387
	pesos_i(4430) := b"0000000000000000_0000000000000000_0001001111001011_0000101001110000"; -- 0.07731690620493968
	pesos_i(4431) := b"0000000000000000_0000000000000000_0001001101110101_1011010000000100"; -- 0.07601475806337761
	pesos_i(4432) := b"1111111111111111_1111111111111111_1111111111001110_1110110000010001"; -- -0.0007488688469599603
	pesos_i(4433) := b"0000000000000000_0000000000000000_0000110111110111_0110110010110010"; -- 0.05455664975123794
	pesos_i(4434) := b"0000000000000000_0000000000000000_0010100101001010_0111110110010011"; -- 0.1612928852497523
	pesos_i(4435) := b"1111111111111111_1111111111111111_1101010011111111_1101110011101010"; -- -0.1679708412702787
	pesos_i(4436) := b"1111111111111111_1111111111111111_1101111011110101_0110110001010001"; -- -0.12906764062319007
	pesos_i(4437) := b"0000000000000000_0000000000000000_0001100010000111_0000000001011101"; -- 0.0958099582431835
	pesos_i(4438) := b"0000000000000000_0000000000000000_0001111110100110_0011111001111000"; -- 0.12363043244802815
	pesos_i(4439) := b"1111111111111111_1111111111111111_1111101110011101_1011101111001100"; -- -0.017124426546042872
	pesos_i(4440) := b"1111111111111111_1111111111111111_1111010011000000_1100000111110011"; -- -0.043933752250800276
	pesos_i(4441) := b"0000000000000000_0000000000000000_0001111011110111_1001100100001001"; -- 0.12096554241378825
	pesos_i(4442) := b"0000000000000000_0000000000000000_0001101110000011_0010100001000010"; -- 0.10747005099390045
	pesos_i(4443) := b"0000000000000000_0000000000000000_0000111111001001_1001111100010010"; -- 0.061670247990685746
	pesos_i(4444) := b"0000000000000000_0000000000000000_0010011101011010_1011101010000100"; -- 0.15372815820149457
	pesos_i(4445) := b"1111111111111111_1111111111111111_1110001001000000_1111010111111111"; -- -0.11619627498296904
	pesos_i(4446) := b"0000000000000000_0000000000000000_0001001100011000_0010101000100110"; -- 0.07458747322943174
	pesos_i(4447) := b"0000000000000000_0000000000000000_0010110100001110_1011001010010111"; -- 0.17600551777342419
	pesos_i(4448) := b"0000000000000000_0000000000000000_0000111001111000_0101101110101001"; -- 0.056524017968823476
	pesos_i(4449) := b"1111111111111111_1111111111111111_1110110101100101_1101101001110101"; -- -0.07266459121050653
	pesos_i(4450) := b"1111111111111111_1111111111111111_1111101101110101_0101110011101000"; -- -0.01774043393543691
	pesos_i(4451) := b"1111111111111111_1111111111111111_1111111111110011_1011001011001100"; -- -0.0001877072018783723
	pesos_i(4452) := b"0000000000000000_0000000000000000_0001000100010101_1011010010111011"; -- 0.06673745686034097
	pesos_i(4453) := b"0000000000000000_0000000000000000_0010010000000111_1110100000011010"; -- 0.14074564575634477
	pesos_i(4454) := b"0000000000000000_0000000000000000_0000110000010100_0001010100100000"; -- 0.04718143486962942
	pesos_i(4455) := b"0000000000000000_0000000000000000_0010110100000010_1001110110001000"; -- 0.17582115707492066
	pesos_i(4456) := b"1111111111111111_1111111111111111_1101100110001011_1000111011110110"; -- -0.15021425707974104
	pesos_i(4457) := b"1111111111111111_1111111111111111_1111100100101100_0000101110100001"; -- -0.02667167003064068
	pesos_i(4458) := b"0000000000000000_0000000000000000_0000101011001111_1101101000101101"; -- 0.0422340737179678
	pesos_i(4459) := b"0000000000000000_0000000000000000_0000001001111010_1110011101110110"; -- 0.009687868346954356
	pesos_i(4460) := b"1111111111111111_1111111111111111_1101101101011100_0101010110001000"; -- -0.14312234325545212
	pesos_i(4461) := b"1111111111111111_1111111111111111_1101100111101111_0101101011001010"; -- -0.14869148805560817
	pesos_i(4462) := b"0000000000000000_0000000000000000_0000011110001000_1111010011110101"; -- 0.029433545965641326
	pesos_i(4463) := b"0000000000000000_0000000000000000_0000111100000110_1100001100101010"; -- 0.058696935420166366
	pesos_i(4464) := b"0000000000000000_0000000000000000_0000101101010010_1000011111101101"; -- 0.04422807259188924
	pesos_i(4465) := b"0000000000000000_0000000000000000_0010111000100101_0110101110100001"; -- 0.1802584904484337
	pesos_i(4466) := b"0000000000000000_0000000000000000_0001010011001011_0010001011101010"; -- 0.08122461517023258
	pesos_i(4467) := b"1111111111111111_1111111111111111_1101011110101010_1100100111011001"; -- -0.157550224882073
	pesos_i(4468) := b"1111111111111111_1111111111111111_1111111010110101_1000110111101001"; -- -0.005042200727243448
	pesos_i(4469) := b"1111111111111111_1111111111111111_1101010111010001_1111100010110010"; -- -0.164764839760625
	pesos_i(4470) := b"1111111111111111_1111111111111111_1110001001111000_0110000000110010"; -- -0.11535071163204906
	pesos_i(4471) := b"0000000000000000_0000000000000000_0010001010010011_1000010101111001"; -- 0.1350634974661903
	pesos_i(4472) := b"0000000000000000_0000000000000000_0010000010000110_1101000110110000"; -- 0.12705717602803032
	pesos_i(4473) := b"0000000000000000_0000000000000000_0010100110110111_1111011001110011"; -- 0.16296329784777944
	pesos_i(4474) := b"1111111111111111_1111111111111111_1110100000000101_1010010010011101"; -- -0.09366389438116256
	pesos_i(4475) := b"1111111111111111_1111111111111111_1110111110111111_0001100111101001"; -- -0.06349027689904768
	pesos_i(4476) := b"1111111111111111_1111111111111111_1101011000110100_0101001001000011"; -- -0.1632641398615169
	pesos_i(4477) := b"1111111111111111_1111111111111111_1111000001101010_1001111101001010"; -- -0.060873073909096055
	pesos_i(4478) := b"0000000000000000_0000000000000000_0001100111001010_0111101110101101"; -- 0.10074589710346003
	pesos_i(4479) := b"0000000000000000_0000000000000000_0000101011110101_1101010111001010"; -- 0.042813646079320575
	pesos_i(4480) := b"1111111111111111_1111111111111111_1110110100111100_0110100100110011"; -- -0.07329695230337445
	pesos_i(4481) := b"0000000000000000_0000000000000000_0001001011011011_0111001001101101"; -- 0.07366099512106418
	pesos_i(4482) := b"1111111111111111_1111111111111111_1110110100100011_1010110100111101"; -- -0.07367436649150821
	pesos_i(4483) := b"1111111111111111_1111111111111111_1111000001110100_1111100000101001"; -- -0.060715188936702295
	pesos_i(4484) := b"0000000000000000_0000000000000000_0000100100011011_0011110110000101"; -- 0.0355719040718644
	pesos_i(4485) := b"0000000000000000_0000000000000000_0010000000110010_0010000000111111"; -- 0.12576486137824106
	pesos_i(4486) := b"1111111111111111_1111111111111111_1111101111001011_0101100001110111"; -- -0.016428442868129525
	pesos_i(4487) := b"1111111111111111_1111111111111111_1111101111101001_1000000010010111"; -- -0.015968287509471112
	pesos_i(4488) := b"1111111111111111_1111111111111111_1110110111101110_1100111110010001"; -- -0.07057478639489838
	pesos_i(4489) := b"1111111111111111_1111111111111111_1110110111011111_0001000110001110"; -- -0.07081499369465774
	pesos_i(4490) := b"0000000000000000_0000000000000000_0000000011001011_0110101011001000"; -- 0.0031038989031164925
	pesos_i(4491) := b"0000000000000000_0000000000000000_0010100010101111_1010111110101011"; -- 0.15893075867233222
	pesos_i(4492) := b"1111111111111111_1111111111111111_1101011101111100_1110110111100011"; -- -0.15824998090726344
	pesos_i(4493) := b"1111111111111111_1111111111111111_1111110000010011_0101010011100001"; -- -0.015330023787412208
	pesos_i(4494) := b"0000000000000000_0000000000000000_0010000001100011_1000101011011111"; -- 0.12651889739651537
	pesos_i(4495) := b"0000000000000000_0000000000000000_0010011110110110_0101010000110011"; -- 0.15512586819569335
	pesos_i(4496) := b"0000000000000000_0000000000000000_0010110001001101_1110110110110011"; -- 0.17306409462562153
	pesos_i(4497) := b"0000000000000000_0000000000000000_0010101111000001_0110001111000100"; -- 0.1709196427097292
	pesos_i(4498) := b"0000000000000000_0000000000000000_0010000110111111_0111000100010000"; -- 0.1318274178155626
	pesos_i(4499) := b"1111111111111111_1111111111111111_1111001011111001_0110010001100000"; -- -0.050882078648679156
	pesos_i(4500) := b"1111111111111111_1111111111111111_1111110001010001_1100001111011111"; -- -0.014377363315025793
	pesos_i(4501) := b"1111111111111111_1111111111111111_1110111111110000_0001010110001110"; -- -0.0627428557593498
	pesos_i(4502) := b"1111111111111111_1111111111111111_1110110011000111_0000000110101010"; -- -0.07508840175822706
	pesos_i(4503) := b"1111111111111111_1111111111111111_1101110011110001_1010101001111110"; -- -0.1369374698004475
	pesos_i(4504) := b"1111111111111111_1111111111111111_1100010111000000_1000001001010001"; -- -0.2275312949620147
	pesos_i(4505) := b"1111111111111111_1111111111111111_1110000111111101_1001011010001110"; -- -0.11722430265392261
	pesos_i(4506) := b"1111111111111111_1111111111111111_1110101001010000_0100010001111000"; -- -0.08471271576844253
	pesos_i(4507) := b"0000000000000000_0000000000000000_0001111001011101_1111001001101000"; -- 0.11862101586647397
	pesos_i(4508) := b"0000000000000000_0000000000000000_0010001001100010_0010001100011001"; -- 0.13430995335370213
	pesos_i(4509) := b"1111111111111111_1111111111111111_1111000010101101_0001001110110011"; -- -0.059859055371247555
	pesos_i(4510) := b"0000000000000000_0000000000000000_0000101100100000_1111100010111000"; -- 0.04347185606139222
	pesos_i(4511) := b"1111111111111111_1111111111111111_1110001110100011_1011111100001010"; -- -0.11078268048896438
	pesos_i(4512) := b"1111111111111111_1111111111111111_1111111111001100_1011010111101111"; -- -0.0007826128540905641
	pesos_i(4513) := b"1111111111111111_1111111111111111_1110100111110111_0111001111010010"; -- -0.08606792561204107
	pesos_i(4514) := b"0000000000000000_0000000000000000_0001111010001101_0010101101000101"; -- 0.11934156839683784
	pesos_i(4515) := b"1111111111111111_1111111111111111_1101001001111010_1101111011001101"; -- -0.17781264786263798
	pesos_i(4516) := b"0000000000000000_0000000000000000_0001010111111101_0010100001001010"; -- 0.08589412493901755
	pesos_i(4517) := b"1111111111111111_1111111111111111_1110011101110111_1100100101101100"; -- -0.09582844846415033
	pesos_i(4518) := b"0000000000000000_0000000000000000_0001001100010001_0000100011100001"; -- 0.07447867854591227
	pesos_i(4519) := b"1111111111111111_1111111111111111_1110110001111001_0111001101110010"; -- -0.0762718053540697
	pesos_i(4520) := b"0000000000000000_0000000000000000_0001010110101100_1010010001111011"; -- 0.08466556559937014
	pesos_i(4521) := b"1111111111111111_1111111111111111_1111010011010101_1011011110011101"; -- -0.043613933787106825
	pesos_i(4522) := b"0000000000000000_0000000000000000_0000111010110111_0011100010110101"; -- 0.05748323843954688
	pesos_i(4523) := b"1111111111111111_1111111111111111_1111011111111100_0100101110000010"; -- -0.03130653443789537
	pesos_i(4524) := b"0000000000000000_0000000000000000_0001010110101101_0010100011010011"; -- 0.08467345373631165
	pesos_i(4525) := b"1111111111111111_1111111111111111_1101100010000001_1100001101001101"; -- -0.15426997526651115
	pesos_i(4526) := b"1111111111111111_1111111111111111_1111111110001111_1110001100010011"; -- -0.0017107084984541996
	pesos_i(4527) := b"0000000000000000_0000000000000000_0010111000011110_0111110011100001"; -- 0.18015270699919095
	pesos_i(4528) := b"0000000000000000_0000000000000000_0001110101010000_0100100001101110"; -- 0.1145062703475184
	pesos_i(4529) := b"0000000000000000_0000000000000000_0000110000000001_0011111001001010"; -- 0.04689397156371669
	pesos_i(4530) := b"0000000000000000_0000000000000000_0000011000011001_0000001000001111"; -- 0.023819092451234886
	pesos_i(4531) := b"0000000000000000_0000000000000000_0010001001010110_1000111010101010"; -- 0.1341332591969672
	pesos_i(4532) := b"1111111111111111_1111111111111111_1101001111100101_0101011100111100"; -- -0.17228178763512125
	pesos_i(4533) := b"0000000000000000_0000000000000000_0000001111000101_1110011011111001"; -- 0.014738498509458022
	pesos_i(4534) := b"1111111111111111_1111111111111111_1101011010111101_1100011111000111"; -- -0.16116668129868028
	pesos_i(4535) := b"1111111111111111_1111111111111111_1101010101000110_1010010000011100"; -- -0.16689085307036675
	pesos_i(4536) := b"0000000000000000_0000000000000000_0000011011100111_1101100011100111"; -- 0.026975208616438817
	pesos_i(4537) := b"0000000000000000_0000000000000000_0000011111011001_0101011001101011"; -- 0.030660058186163318
	pesos_i(4538) := b"0000000000000000_0000000000000000_0001111011101100_1101001010111100"; -- 0.12080113499694174
	pesos_i(4539) := b"1111111111111111_1111111111111111_1101100001101110_0000011101101111"; -- -0.15457109012451398
	pesos_i(4540) := b"0000000000000000_0000000000000000_0000111100011110_0010110110000000"; -- 0.05905422557877627
	pesos_i(4541) := b"0000000000000000_0000000000000000_0000111001111111_0011001011010111"; -- 0.056628396440297366
	pesos_i(4542) := b"0000000000000000_0000000000000000_0010110000110011_0111101000101001"; -- 0.1726604795354355
	pesos_i(4543) := b"0000000000000000_0000000000000000_0001110001100010_1010010000000000"; -- 0.1108801364196602
	pesos_i(4544) := b"0000000000000000_0000000000000000_0000100110110100_0100011100011010"; -- 0.037907069927828746
	pesos_i(4545) := b"0000000000000000_0000000000000000_0001011101001101_1100111011110110"; -- 0.09103101260752183
	pesos_i(4546) := b"0000000000000000_0000000000000000_0001000101001101_1000110101011011"; -- 0.06758960214585485
	pesos_i(4547) := b"1111111111111111_1111111111111111_1111110111000100_0110010110101101"; -- -0.008721967083844267
	pesos_i(4548) := b"0000000000000000_0000000000000000_0010100001010001_0001000100101001"; -- 0.15748698467360786
	pesos_i(4549) := b"1111111111111111_1111111111111111_1101011000011001_0110100110000111"; -- -0.16367474040084665
	pesos_i(4550) := b"0000000000000000_0000000000000000_0000011110010011_0011011111101001"; -- 0.029590124421583344
	pesos_i(4551) := b"1111111111111111_1111111111111111_1111000101010011_0001010010110101"; -- -0.057326036185245004
	pesos_i(4552) := b"1111111111111111_1111111111111111_1111001000001001_1111001111000000"; -- -0.054535642201832664
	pesos_i(4553) := b"0000000000000000_0000000000000000_0000010000100001_0000110011000111"; -- 0.016129301582396744
	pesos_i(4554) := b"1111111111111111_1111111111111111_1101011100010000_0001101111110110"; -- -0.15991044274566016
	pesos_i(4555) := b"0000000000000000_0000000000000000_0000001001101001_0111000111000100"; -- 0.00942145386692915
	pesos_i(4556) := b"1111111111111111_1111111111111111_1111011010000101_0010010000010100"; -- -0.037030930569169285
	pesos_i(4557) := b"0000000000000000_0000000000000000_0000010000000100_1010100000001000"; -- 0.01569605064256775
	pesos_i(4558) := b"0000000000000000_0000000000000000_0000001100100110_0111011101001000"; -- 0.012305693614797875
	pesos_i(4559) := b"1111111111111111_1111111111111111_1110011110001101_0001010101001001"; -- -0.09550349211863272
	pesos_i(4560) := b"1111111111111111_1111111111111111_1110110001001000_0001101100101101"; -- -0.07702474749899467
	pesos_i(4561) := b"0000000000000000_0000000000000000_0000100001011111_0101000110001000"; -- 0.03270444454899072
	pesos_i(4562) := b"1111111111111111_1111111111111111_1110110001000100_1101101011101011"; -- -0.07707435382325913
	pesos_i(4563) := b"0000000000000000_0000000000000000_0010100000001111_0001011000110110"; -- 0.1564802057664504
	pesos_i(4564) := b"1111111111111111_1111111111111111_1110001011101110_1101111000001101"; -- -0.11354267284446092
	pesos_i(4565) := b"1111111111111111_1111111111111111_1101001101110111_0001101100110110"; -- -0.17396383227481368
	pesos_i(4566) := b"0000000000000000_0000000000000000_0001110000010011_1111110101110000"; -- 0.10968002304103285
	pesos_i(4567) := b"0000000000000000_0000000000000000_0010101010100010_0010010100001011"; -- 0.16653663170734506
	pesos_i(4568) := b"1111111111111111_1111111111111111_1100111000010101_1101100000010010"; -- -0.19497918660662852
	pesos_i(4569) := b"0000000000000000_0000000000000000_0010101111101001_1110011111011011"; -- 0.1715378676018828
	pesos_i(4570) := b"0000000000000000_0000000000000000_0000011111001100_0110001100111011"; -- 0.030462457554210398
	pesos_i(4571) := b"1111111111111111_1111111111111111_1110110101000110_1010000100010000"; -- -0.07314103470036024
	pesos_i(4572) := b"1111111111111111_1111111111111111_1111110010101110_1001010010111000"; -- -0.012961106458862563
	pesos_i(4573) := b"0000000000000000_0000000000000000_0010100110110001_0011101100111001"; -- 0.16286058565499992
	pesos_i(4574) := b"0000000000000000_0000000000000000_0010010111101110_0001010000011110"; -- 0.14816404078704198
	pesos_i(4575) := b"1111111111111111_1111111111111111_1110011010110100_1001111100011011"; -- -0.09880643445276924
	pesos_i(4576) := b"1111111111111111_1111111111111111_1101011101111100_0001000110100101"; -- -0.1582631084331233
	pesos_i(4577) := b"1111111111111111_1111111111111111_1111111100010110_0010001110110111"; -- -0.00356842797411525
	pesos_i(4578) := b"0000000000000000_0000000000000000_0010001011000010_1111101110100110"; -- 0.1357877045874871
	pesos_i(4579) := b"0000000000000000_0000000000000000_0010101011101110_0111111010011010"; -- 0.16770163773465016
	pesos_i(4580) := b"1111111111111111_1111111111111111_1101011101110010_0010101010110001"; -- -0.15841420344023352
	pesos_i(4581) := b"0000000000000000_0000000000000000_0000000101000010_1101000000000010"; -- 0.004925728314159748
	pesos_i(4582) := b"1111111111111111_1111111111111111_1110011101111001_0100110010101010"; -- -0.09580536687884914
	pesos_i(4583) := b"0000000000000000_0000000000000000_0010001111010100_0100111100010001"; -- 0.13995832590116006
	pesos_i(4584) := b"1111111111111111_1111111111111111_1111100000110101_0111000110010011"; -- -0.030434514708137878
	pesos_i(4585) := b"1111111111111111_1111111111111111_1101010101101011_0011001011101111"; -- -0.16633302378510567
	pesos_i(4586) := b"1111111111111111_1111111111111111_1110000010000000_0001001101110111"; -- -0.12304571473876932
	pesos_i(4587) := b"1111111111111111_1111111111111111_1101011101001111_0011101000110010"; -- -0.15894733696128033
	pesos_i(4588) := b"1111111111111111_1111111111111111_1111001010110001_1000010100010101"; -- -0.05197876196342739
	pesos_i(4589) := b"1111111111111111_1111111111111111_1111010101011001_1000111100110000"; -- -0.04160218309245488
	pesos_i(4590) := b"1111111111111111_1111111111111111_1110101011110001_0110100010000011"; -- -0.08225390240857837
	pesos_i(4591) := b"1111111111111111_1111111111111111_1101111110010100_1100110101110010"; -- -0.12663570381031164
	pesos_i(4592) := b"1111111111111111_1111111111111111_1111111110011101_0001011111010100"; -- -0.001509199738192163
	pesos_i(4593) := b"1111111111111111_1111111111111111_1111011111001000_0100100000100010"; -- -0.032100192798617595
	pesos_i(4594) := b"1111111111111111_1111111111111111_1111010101111000_0100100100000000"; -- -0.04113334427614189
	pesos_i(4595) := b"1111111111111111_1111111111111111_1110100001101011_1011000100111011"; -- -0.09210674575217659
	pesos_i(4596) := b"1111111111111111_1111111111111111_1111011111010010_0000101000011001"; -- -0.031951302345768595
	pesos_i(4597) := b"0000000000000000_0000000000000000_0000011110000110_1011001100001110"; -- 0.029399100183542946
	pesos_i(4598) := b"1111111111111111_1111111111111111_1101010001010111_1010100000000001"; -- -0.17053747146835793
	pesos_i(4599) := b"0000000000000000_0000000000000000_0010011100000010_1101010110110111"; -- 0.1523870059690891
	pesos_i(4600) := b"0000000000000000_0000000000000000_0000001111011001_0000001101001010"; -- 0.015030103378000564
	pesos_i(4601) := b"1111111111111111_1111111111111111_1101011100100001_0010110000110011"; -- -0.1596500754402337
	pesos_i(4602) := b"1111111111111111_1111111111111111_1111110110010000_0011011000110110"; -- -0.009518253053841285
	pesos_i(4603) := b"0000000000000000_0000000000000000_0001111100100010_1011100100011100"; -- 0.12162358213811138
	pesos_i(4604) := b"1111111111111111_1111111111111111_1101101111111111_1101100101111111"; -- -0.1406272950232077
	pesos_i(4605) := b"0000000000000000_0000000000000000_0000000100110111_0011111110110010"; -- 0.004749279824929783
	pesos_i(4606) := b"0000000000000000_0000000000000000_0000010001001110_0110000000111111"; -- 0.016820922210933155
	pesos_i(4607) := b"0000000000000000_0000000000000000_0000001110000001_1000001101101011"; -- 0.01369496684955152
	pesos_i(4608) := b"0000000000000000_0000000000000000_0000111011011101_0110101101010011"; -- 0.05806608941410299
	pesos_i(4609) := b"1111111111111111_1111111111111111_1110110111100100_1100010101010100"; -- -0.07072798444399896
	pesos_i(4610) := b"1111111111111111_1111111111111111_1111001110101000_1110100011101110"; -- -0.048203889710105544
	pesos_i(4611) := b"0000000000000000_0000000000000000_0001000001010100_1001010010011101"; -- 0.06379059621930831
	pesos_i(4612) := b"0000000000000000_0000000000000000_0000000101000110_0111000100100000"; -- 0.004981107953528099
	pesos_i(4613) := b"1111111111111111_1111111111111111_1110000100011010_1011100111111110"; -- -0.12068593550367884
	pesos_i(4614) := b"1111111111111111_1111111111111111_1111001010111110_0000000000000111"; -- -0.051788328345338766
	pesos_i(4615) := b"0000000000000000_0000000000000000_0000101001100110_0000011111001000"; -- 0.04061936023291038
	pesos_i(4616) := b"0000000000000000_0000000000000000_0000000101110110_0101110011011000"; -- 0.005712321022712013
	pesos_i(4617) := b"1111111111111111_1111111111111111_1110100101011010_0111100011101000"; -- -0.08846325245954245
	pesos_i(4618) := b"1111111111111111_1111111111111111_1111010011101011_0011000101101010"; -- -0.04328623916368553
	pesos_i(4619) := b"0000000000000000_0000000000000000_0000100110110011_0000110000010111"; -- 0.037888293919466534
	pesos_i(4620) := b"1111111111111111_1111111111111111_1110010001101010_1000000000111000"; -- -0.10774992587218644
	pesos_i(4621) := b"1111111111111111_1111111111111111_1111111100111000_1011111011010110"; -- -0.0030403831882706406
	pesos_i(4622) := b"1111111111111111_1111111111111111_1110000110101110_0010101110010101"; -- -0.11843612298064495
	pesos_i(4623) := b"0000000000000000_0000000000000000_0001101110011100_1001111001111000"; -- 0.1078585664517998
	pesos_i(4624) := b"0000000000000000_0000000000000000_0010000011101001_1100011011000010"; -- 0.1285671447887747
	pesos_i(4625) := b"0000000000000000_0000000000000000_0001010111110101_0101001100010101"; -- 0.08577460544669019
	pesos_i(4626) := b"0000000000000000_0000000000000000_0001000111001100_0111110101100010"; -- 0.06952651637140206
	pesos_i(4627) := b"0000000000000000_0000000000000000_0000001110101110_0111110101011000"; -- 0.014381250283011297
	pesos_i(4628) := b"1111111111111111_1111111111111111_1110110011101111_0101000100001111"; -- -0.0744733180371166
	pesos_i(4629) := b"1111111111111111_1111111111111111_1101001101100001_0100101110011000"; -- -0.174296641728738
	pesos_i(4630) := b"0000000000000000_0000000000000000_0000011111010111_1100000010000011"; -- 0.030635864178432858
	pesos_i(4631) := b"1111111111111111_1111111111111111_1110011000010011_0100001011100101"; -- -0.1012685957503537
	pesos_i(4632) := b"1111111111111111_1111111111111111_1111010011101001_1000101000110001"; -- -0.04331146528488037
	pesos_i(4633) := b"1111111111111111_1111111111111111_1110001101110100_1111111110101011"; -- -0.11149599152957919
	pesos_i(4634) := b"0000000000000000_0000000000000000_0010010110001101_1000100100100001"; -- 0.14669091276815752
	pesos_i(4635) := b"0000000000000000_0000000000000000_0001000111001101_0010001101110011"; -- 0.0695364146398613
	pesos_i(4636) := b"1111111111111111_1111111111111111_1101010011100011_1101110001000101"; -- -0.16839812581505703
	pesos_i(4637) := b"0000000000000000_0000000000000000_0001100010010110_0010111101010011"; -- 0.09604163902894058
	pesos_i(4638) := b"0000000000000000_0000000000000000_0001101110110100_1000011100011110"; -- 0.10822338562579258
	pesos_i(4639) := b"1111111111111111_1111111111111111_1101010110111111_1000111101110010"; -- -0.16504577131388146
	pesos_i(4640) := b"1111111111111111_1111111111111111_1110101000110101_0100101010111011"; -- -0.08512432989433215
	pesos_i(4641) := b"1111111111111111_1111111111111111_1111001110000101_0100001010101010"; -- -0.048747857570827176
	pesos_i(4642) := b"1111111111111111_1111111111111111_1101110110001111_1010000100111100"; -- -0.13452713291059024
	pesos_i(4643) := b"0000000000000000_0000000000000000_0001010010010010_0010100111101000"; -- 0.08035528107789232
	pesos_i(4644) := b"1111111111111111_1111111111111111_1111011011111111_1010000000000111"; -- -0.03516197047290228
	pesos_i(4645) := b"1111111111111111_1111111111111111_1101111110110101_0011110100100110"; -- -0.12614076437079733
	pesos_i(4646) := b"1111111111111111_1111111111111111_1101111110001010_1010100110011101"; -- -0.1267904274708542
	pesos_i(4647) := b"1111111111111111_1111111111111111_1110111000000000_0110010011011001"; -- -0.07030648892124097
	pesos_i(4648) := b"0000000000000000_0000000000000000_0000111000110001_0111001111011101"; -- 0.055442086583939926
	pesos_i(4649) := b"1111111111111111_1111111111111111_1101010011101101_0011011001010110"; -- -0.1682554282050287
	pesos_i(4650) := b"0000000000000000_0000000000000000_0000011001110011_1100101000111100"; -- 0.025204314913328935
	pesos_i(4651) := b"1111111111111111_1111111111111111_1111100100000000_1111000001011100"; -- -0.027329423452954322
	pesos_i(4652) := b"0000000000000000_0000000000000000_0001101100111101_1010110101110101"; -- 0.10640987490327282
	pesos_i(4653) := b"0000000000000000_0000000000000000_0001011011101011_1010100111000011"; -- 0.08953343411639464
	pesos_i(4654) := b"1111111111111111_1111111111111111_1110111110111101_0101101001001000"; -- -0.06351695765282797
	pesos_i(4655) := b"0000000000000000_0000000000000000_0000100110000111_0000100011100110"; -- 0.03721671697982224
	pesos_i(4656) := b"1111111111111111_1111111111111111_1101011011101111_0111100011101000"; -- -0.16040844280826705
	pesos_i(4657) := b"1111111111111111_1111111111111111_1110011010111110_1101110111011110"; -- -0.09865010569436528
	pesos_i(4658) := b"0000000000000000_0000000000000000_0010011001101010_1110001111001011"; -- 0.15006850914667982
	pesos_i(4659) := b"0000000000000000_0000000000000000_0001111101100100_1100111100110100"; -- 0.12263197923581416
	pesos_i(4660) := b"1111111111111111_1111111111111111_1101100011100010_1010010101101011"; -- -0.15279165395398356
	pesos_i(4661) := b"1111111111111111_1111111111111111_1111001001101011_1011101110100011"; -- -0.05304362554121513
	pesos_i(4662) := b"0000000000000000_0000000000000000_0010111011011011_0010110110111000"; -- 0.18303189991960697
	pesos_i(4663) := b"0000000000000000_0000000000000000_0001101110100101_1011000100110001"; -- 0.1079970117151719
	pesos_i(4664) := b"0000000000000000_0000000000000000_0001111001000101_0000110010110100"; -- 0.11824111369954274
	pesos_i(4665) := b"0000000000000000_0000000000000000_0001101011001100_1110011010000000"; -- 0.10468903177380658
	pesos_i(4666) := b"1111111111111111_1111111111111111_1101011001011101_1101010001011111"; -- -0.16263077433202922
	pesos_i(4667) := b"0000000000000000_0000000000000000_0010100010111110_0101011010001101"; -- 0.15915432878652275
	pesos_i(4668) := b"1111111111111111_1111111111111111_1110111100111111_1001001011011111"; -- -0.06543619215109205
	pesos_i(4669) := b"1111111111111111_1111111111111111_1110111010011010_0010100011011101"; -- -0.06796021085393643
	pesos_i(4670) := b"1111111111111111_1111111111111111_1101101101101000_0110011111111011"; -- -0.14293813811089554
	pesos_i(4671) := b"0000000000000000_0000000000000000_0001111011101011_1110010010110010"; -- 0.12078694677175687
	pesos_i(4672) := b"1111111111111111_1111111111111111_1111000011010011_1011111001001011"; -- -0.059269053099164706
	pesos_i(4673) := b"0000000000000000_0000000000000000_0000001100101001_0111110001000000"; -- 0.01235176627817739
	pesos_i(4674) := b"1111111111111111_1111111111111111_1110010000111000_1110000000010000"; -- -0.10850715256858025
	pesos_i(4675) := b"0000000000000000_0000000000000000_0000000011100101_0110110011011000"; -- 0.003500750365713368
	pesos_i(4676) := b"0000000000000000_0000000000000000_0001010001111111_0100101111001110"; -- 0.08006738441550083
	pesos_i(4677) := b"1111111111111111_1111111111111111_1101100011100110_0111011001011110"; -- -0.15273342325676245
	pesos_i(4678) := b"1111111111111111_1111111111111111_1101100010100010_1101001101111000"; -- -0.15376547158095805
	pesos_i(4679) := b"1111111111111111_1111111111111111_1111111001101101_0010010010000110"; -- -0.006147115071783819
	pesos_i(4680) := b"1111111111111111_1111111111111111_1101011101101110_1100000110101001"; -- -0.15846624024484363
	pesos_i(4681) := b"0000000000000000_0000000000000000_0010000110000000_0101010110111011"; -- 0.13086448489896316
	pesos_i(4682) := b"1111111111111111_1111111111111111_1111010000101110_1111010011101001"; -- -0.046158497942720686
	pesos_i(4683) := b"0000000000000000_0000000000000000_0010011100011010_1001101100010000"; -- 0.15274972099642614
	pesos_i(4684) := b"1111111111111111_1111111111111111_1101110100001000_1100100111010001"; -- -0.13658465046768012
	pesos_i(4685) := b"1111111111111111_1111111111111111_1111101101011001_0110010110000011"; -- -0.018167167143095263
	pesos_i(4686) := b"0000000000000000_0000000000000000_0010000110001010_0001001111011010"; -- 0.13101314608426057
	pesos_i(4687) := b"1111111111111111_1111111111111111_1101111000001011_1101111110001111"; -- -0.13263132823281434
	pesos_i(4688) := b"0000000000000000_0000000000000000_0001101110011001_1000110010010000"; -- 0.1078117227926226
	pesos_i(4689) := b"0000000000000000_0000000000000000_0000010100110010_1110001110010001"; -- 0.020307753570917218
	pesos_i(4690) := b"1111111111111111_1111111111111111_1110000001100111_0110011111001011"; -- -0.12342215828060023
	pesos_i(4691) := b"0000000000000000_0000000000000000_0001111110011100_0000111100011111"; -- 0.12347502231847356
	pesos_i(4692) := b"0000000000000000_0000000000000000_0010010110110000_1011000110001110"; -- 0.14722737998498617
	pesos_i(4693) := b"1111111111111111_1111111111111111_1110110000100000_0100100101101101"; -- -0.0776323423290359
	pesos_i(4694) := b"0000000000000000_0000000000000000_0001110100011010_1110000110001111"; -- 0.11369142292858711
	pesos_i(4695) := b"1111111111111111_1111111111111111_1111000011110001_1110100110111111"; -- -0.05880869952861545
	pesos_i(4696) := b"1111111111111111_1111111111111111_1110101110010011_1001101001100010"; -- -0.07977900604078421
	pesos_i(4697) := b"1111111111111111_1111111111111111_1111110100001111_1110001110001000"; -- -0.011476306207207373
	pesos_i(4698) := b"1111111111111111_1111111111111111_1111000011010110_1011111110101100"; -- -0.05922319452401951
	pesos_i(4699) := b"0000000000000000_0000000000000000_0010010110001000_1110111001111100"; -- 0.1466206602030736
	pesos_i(4700) := b"1111111111111111_1111111111111111_1110001010000011_0011011110010110"; -- -0.11518528556711644
	pesos_i(4701) := b"1111111111111111_1111111111111111_1111111011001110_1000001100101111"; -- -0.004661370417456707
	pesos_i(4702) := b"0000000000000000_0000000000000000_0010100100001001_0001000000001100"; -- 0.1602945356206471
	pesos_i(4703) := b"0000000000000000_0000000000000000_0000101100100000_0010010011111010"; -- 0.043459235291440634
	pesos_i(4704) := b"1111111111111111_1111111111111111_1111000011010110_0111111101110001"; -- -0.05922702312351173
	pesos_i(4705) := b"0000000000000000_0000000000000000_0010010111101101_0001111110010110"; -- 0.1481494655930587
	pesos_i(4706) := b"1111111111111111_1111111111111111_1110110101000110_1000100011110011"; -- -0.07314247197389932
	pesos_i(4707) := b"1111111111111111_1111111111111111_1111100110010001_0111010101010111"; -- -0.025124231478230594
	pesos_i(4708) := b"0000000000000000_0000000000000000_0000001010010101_1011010110010011"; -- 0.010096882135280396
	pesos_i(4709) := b"0000000000000000_0000000000000000_0010001101001111_0001101000111001"; -- 0.1379257573619971
	pesos_i(4710) := b"1111111111111111_1111111111111111_1111000011000100_0001110110001111"; -- -0.05950751544818111
	pesos_i(4711) := b"0000000000000000_0000000000000000_0000011011110111_1110011001111101"; -- 0.027220158984711695
	pesos_i(4712) := b"1111111111111111_1111111111111111_1111010101001110_0101001011010101"; -- -0.04177362727419481
	pesos_i(4713) := b"0000000000000000_0000000000000000_0000011111011011_0110010110111001"; -- 0.030691487901824036
	pesos_i(4714) := b"1111111111111111_1111111111111111_1111111001100110_1001100000110011"; -- -0.006247031653390864
	pesos_i(4715) := b"1111111111111111_1111111111111111_1110101011000111_1011011001110010"; -- -0.08289012630296529
	pesos_i(4716) := b"0000000000000000_0000000000000000_0010001001101100_1101101001001100"; -- 0.13447346064683088
	pesos_i(4717) := b"0000000000000000_0000000000000000_0000000010100100_0011100100001111"; -- 0.002505842272651705
	pesos_i(4718) := b"1111111111111111_1111111111111111_1111111111110111_1111011000111011"; -- -0.00012265271444765236
	pesos_i(4719) := b"1111111111111111_1111111111111111_1101011001001010_0001010101100111"; -- -0.1629320739002599
	pesos_i(4720) := b"1111111111111111_1111111111111111_1111010000111101_0100100010000010"; -- -0.045939892123580545
	pesos_i(4721) := b"1111111111111111_1111111111111111_1101111010000010_0101010111100111"; -- -0.13082373726672372
	pesos_i(4722) := b"1111111111111111_1111111111111111_1111010010100111_1000101010111110"; -- -0.04431851254706503
	pesos_i(4723) := b"1111111111111111_1111111111111111_1111001101101010_1001000101111111"; -- -0.049155146122495774
	pesos_i(4724) := b"1111111111111111_1111111111111111_1111101110111100_1110101010110101"; -- -0.016648608082412735
	pesos_i(4725) := b"1111111111111111_1111111111111111_1110110011101100_0011010111001110"; -- -0.07452071872346451
	pesos_i(4726) := b"0000000000000000_0000000000000000_0001010101011010_0011000010100100"; -- 0.08340744013570006
	pesos_i(4727) := b"0000000000000000_0000000000000000_0001001100000010_0111001011001001"; -- 0.0742561092353636
	pesos_i(4728) := b"1111111111111111_1111111111111111_1101111110110000_0000011110111101"; -- -0.12622024198486093
	pesos_i(4729) := b"0000000000000000_0000000000000000_0010010111011000_1100000101111100"; -- 0.14783868107917453
	pesos_i(4730) := b"0000000000000000_0000000000000000_0010100100000111_0001001100000100"; -- 0.16026419502023231
	pesos_i(4731) := b"1111111111111111_1111111111111111_1101111010010011_1111101010001011"; -- -0.13055452459560368
	pesos_i(4732) := b"0000000000000000_0000000000000000_0001000110111101_1110001100101010"; -- 0.0693037010908189
	pesos_i(4733) := b"0000000000000000_0000000000000000_0001011010111101_0110100111011110"; -- 0.0888277213683485
	pesos_i(4734) := b"0000000000000000_0000000000000000_0001011011100000_0010010000101101"; -- 0.08935762495179318
	pesos_i(4735) := b"0000000000000000_0000000000000000_0010011100111111_1001001000100001"; -- 0.153313763614922
	pesos_i(4736) := b"0000000000000000_0000000000000000_0001101010001011_1000111000010011"; -- 0.10369193995209738
	pesos_i(4737) := b"0000000000000000_0000000000000000_0001001010111000_1010100101010110"; -- 0.07313021041826905
	pesos_i(4738) := b"1111111111111111_1111111111111111_1101011011000000_0110101111011001"; -- -0.16112638427210596
	pesos_i(4739) := b"1111111111111111_1111111111111111_1110001000101010_1011100000101001"; -- -0.11653565417157272
	pesos_i(4740) := b"1111111111111111_1111111111111111_1111000011011110_1001011011000101"; -- -0.05910356228413672
	pesos_i(4741) := b"0000000000000000_0000000000000000_0001101111000010_1001011110001101"; -- 0.10843798816878003
	pesos_i(4742) := b"1111111111111111_1111111111111111_1101010000111011_0110000101001001"; -- -0.17096893290531262
	pesos_i(4743) := b"0000000000000000_0000000000000000_0000011000011101_1011101000100100"; -- 0.02389109962714439
	pesos_i(4744) := b"0000000000000000_0000000000000000_0001101001101010_1111011011011001"; -- 0.10319464500799819
	pesos_i(4745) := b"1111111111111111_1111111111111111_1101110111010000_0111000010010111"; -- -0.1335382110119215
	pesos_i(4746) := b"0000000000000000_0000000000000000_0001000111001111_0100110010110111"; -- 0.06956939189855227
	pesos_i(4747) := b"0000000000000000_0000000000000000_0001001010111001_1011001111010001"; -- 0.07314609377621437
	pesos_i(4748) := b"0000000000000000_0000000000000000_0010011010111111_1010011110100010"; -- 0.15136192030242626
	pesos_i(4749) := b"1111111111111111_1111111111111111_1111001111011101_1011000000011011"; -- -0.047398560814489704
	pesos_i(4750) := b"1111111111111111_1111111111111111_1101101010110111_1010111001011101"; -- -0.14563474866024467
	pesos_i(4751) := b"0000000000000000_0000000000000000_0010101110100111_0100010110101110"; -- 0.17052112107437972
	pesos_i(4752) := b"0000000000000000_0000000000000000_0000001011010010_0111101010001110"; -- 0.01102415043342303
	pesos_i(4753) := b"0000000000000000_0000000000000000_0001100111101110_0011010111111011"; -- 0.10129105932662703
	pesos_i(4754) := b"0000000000000000_0000000000000000_0000011111100110_0110001111110110"; -- 0.030859229652982798
	pesos_i(4755) := b"0000000000000000_0000000000000000_0010000011010001_1011111110000000"; -- 0.1282005011660334
	pesos_i(4756) := b"1111111111111111_1111111111111111_1110001101100000_1101100011101101"; -- -0.11180347655329465
	pesos_i(4757) := b"0000000000000000_0000000000000000_0001111101011001_1001110011001111"; -- 0.12246112874402015
	pesos_i(4758) := b"1111111111111111_1111111111111111_1110111110000010_1011001011100111"; -- -0.0644119440933795
	pesos_i(4759) := b"1111111111111111_1111111111111111_1111000011011110_1110101100110001"; -- -0.059098530227122026
	pesos_i(4760) := b"0000000000000000_0000000000000000_0000110001111111_0100101111010000"; -- 0.048817384943807024
	pesos_i(4761) := b"1111111111111111_1111111111111111_1111101101100011_0101010001101001"; -- -0.018015598564769766
	pesos_i(4762) := b"0000000000000000_0000000000000000_0000010100100110_0011101110111100"; -- 0.020114644396489977
	pesos_i(4763) := b"1111111111111111_1111111111111111_1101100110110010_0101001110101010"; -- -0.1496226987974507
	pesos_i(4764) := b"0000000000000000_0000000000000000_0010011100000100_0101001101101001"; -- 0.1524097568338936
	pesos_i(4765) := b"0000000000000000_0000000000000000_0010101000111101_0011100101011010"; -- 0.16499670462945074
	pesos_i(4766) := b"1111111111111111_1111111111111111_1110011111010001_1111010100111010"; -- -0.09445254655210586
	pesos_i(4767) := b"0000000000000000_0000000000000000_0001100110011100_1010000111100111"; -- 0.10004627117160939
	pesos_i(4768) := b"0000000000000000_0000000000000000_0000100110111101_0101101110010111"; -- 0.03804562025148722
	pesos_i(4769) := b"0000000000000000_0000000000000000_0010011011001000_0100111110111111"; -- 0.15149401104262067
	pesos_i(4770) := b"0000000000000000_0000000000000000_0000110100011101_1010001011100110"; -- 0.05123346444174915
	pesos_i(4771) := b"0000000000000000_0000000000000000_0000110000000001_0000110010110010"; -- 0.04689101541069431
	pesos_i(4772) := b"0000000000000000_0000000000000000_0010000111011111_0000100101000010"; -- 0.1323095117652005
	pesos_i(4773) := b"1111111111111111_1111111111111111_1101011001111101_0001101011101000"; -- -0.16215354763678239
	pesos_i(4774) := b"1111111111111111_1111111111111111_1101100001101111_1000010110100001"; -- -0.1545483094645186
	pesos_i(4775) := b"1111111111111111_1111111111111111_1111000111001111_1100010111010110"; -- -0.05542338873069837
	pesos_i(4776) := b"0000000000000000_0000000000000000_0000010010000011_1001111101101110"; -- 0.01763340403582514
	pesos_i(4777) := b"1111111111111111_1111111111111111_1111111111010110_0110010110000001"; -- -0.0006348190077011131
	pesos_i(4778) := b"1111111111111111_1111111111111111_1110011000011011_0110001001001000"; -- -0.10114465458715055
	pesos_i(4779) := b"0000000000000000_0000000000000000_0000010010010011_1101100010000110"; -- 0.017880947787396972
	pesos_i(4780) := b"1111111111111111_1111111111111111_1101000101011110_0111000100111110"; -- -0.1821526739601104
	pesos_i(4781) := b"1111111111111111_1111111111111111_1111011011100100_1010100010101101"; -- -0.035573442225053466
	pesos_i(4782) := b"1111111111111111_1111111111111111_1110001000101101_1111010001010111"; -- -0.116486290599747
	pesos_i(4783) := b"1111111111111111_1111111111111111_1110100010111110_1010001100111000"; -- -0.09084110144054137
	pesos_i(4784) := b"0000000000000000_0000000000000000_0000100111101101_1111101101101111"; -- 0.038787569645316794
	pesos_i(4785) := b"0000000000000000_0000000000000000_0001011111110010_0001110001011111"; -- 0.09353806799753132
	pesos_i(4786) := b"0000000000000000_0000000000000000_0010110110010110_1001110010010100"; -- 0.17807940119419385
	pesos_i(4787) := b"1111111111111111_1111111111111111_1110100000001010_1000011111001101"; -- -0.09358931773707835
	pesos_i(4788) := b"0000000000000000_0000000000000000_0000000011000100_0010010101110100"; -- 0.0029929550275626417
	pesos_i(4789) := b"1111111111111111_1111111111111111_1111100110001000_1100010010001011"; -- -0.02525683973364433
	pesos_i(4790) := b"1111111111111111_1111111111111111_1110011100011111_0100111010010111"; -- -0.09717854321274175
	pesos_i(4791) := b"1111111111111111_1111111111111111_1110000101111111_1010010101111001"; -- -0.11914602079807309
	pesos_i(4792) := b"0000000000000000_0000000000000000_0010101101101001_0101010001100110"; -- 0.16957595333303457
	pesos_i(4793) := b"0000000000000000_0000000000000000_0001001000110101_0110110011101001"; -- 0.07112770741994266
	pesos_i(4794) := b"1111111111111111_1111111111111111_1111101010101101_0100101001101110"; -- -0.020793293212514524
	pesos_i(4795) := b"0000000000000000_0000000000000000_0001000101010010_0110010001010001"; -- 0.06766345011415284
	pesos_i(4796) := b"1111111111111111_1111111111111111_1110000101011101_1010101110000010"; -- -0.1196644600495377
	pesos_i(4797) := b"1111111111111111_1111111111111111_1111110001100000_0011111000001001"; -- -0.014156458580349566
	pesos_i(4798) := b"1111111111111111_1111111111111111_1111101111000001_1100000010101011"; -- -0.016574819882211843
	pesos_i(4799) := b"0000000000000000_0000000000000000_0000101111100000_0110011010100100"; -- 0.04639283670706281
	pesos_i(4800) := b"0000000000000000_0000000000000000_0010101110011110_0110101010000011"; -- 0.17038598718171624
	pesos_i(4801) := b"0000000000000000_0000000000000000_0000000101101100_0000000010000110"; -- 0.005554230436224093
	pesos_i(4802) := b"0000000000000000_0000000000000000_0010110000000011_1011001011011101"; -- 0.1719314374733949
	pesos_i(4803) := b"0000000000000000_0000000000000000_0001001110001000_1100111010111110"; -- 0.0763062680209154
	pesos_i(4804) := b"1111111111111111_1111111111111111_1111101010110000_1100111000010101"; -- -0.02073966967012034
	pesos_i(4805) := b"1111111111111111_1111111111111111_1111101000101110_1100011011111010"; -- -0.02272373582304722
	pesos_i(4806) := b"1111111111111111_1111111111111111_1111001110101000_0110010110011011"; -- -0.04821171735263344
	pesos_i(4807) := b"1111111111111111_1111111111111111_1101110100110011_0111110000101010"; -- -0.13593315091064812
	pesos_i(4808) := b"0000000000000000_0000000000000000_0001001101000000_0101000100011000"; -- 0.07520014617359176
	pesos_i(4809) := b"0000000000000000_0000000000000000_0010101100010111_1101111111011011"; -- 0.16833304485955203
	pesos_i(4810) := b"0000000000000000_0000000000000000_0001101010011000_0101010000000011"; -- 0.10388684336618584
	pesos_i(4811) := b"1111111111111111_1111111111111111_1111001111000011_1100111001100110"; -- -0.04779348380062409
	pesos_i(4812) := b"0000000000000000_0000000000000000_0010101011101010_1110110100011111"; -- 0.16764719008760107
	pesos_i(4813) := b"1111111111111111_1111111111111111_1110110110011010_0101010111111111"; -- -0.07186377083353675
	pesos_i(4814) := b"1111111111111111_1111111111111111_1101011000011101_0001111101001011"; -- -0.16361812985288388
	pesos_i(4815) := b"0000000000000000_0000000000000000_0010100110000001_0111111101101010"; -- 0.1621322282417315
	pesos_i(4816) := b"1111111111111111_1111111111111111_1110111001110011_1101110111101001"; -- -0.06854451241308307
	pesos_i(4817) := b"1111111111111111_1111111111111111_1111001101010110_0010100101100010"; -- -0.04946652745988495
	pesos_i(4818) := b"1111111111111111_1111111111111111_1111100111110101_1000010011101110"; -- -0.023597423554968796
	pesos_i(4819) := b"1111111111111111_1111111111111111_1110101011010111_0110000011101010"; -- -0.08265108382598656
	pesos_i(4820) := b"1111111111111111_1111111111111111_1110100001111001_0111001101000000"; -- -0.0918968170095226
	pesos_i(4821) := b"1111111111111111_1111111111111111_1111000001100101_0111111100101100"; -- -0.06095128219376178
	pesos_i(4822) := b"1111111111111111_1111111111111111_1110001110110111_0110100011101100"; -- -0.11048263788027164
	pesos_i(4823) := b"0000000000000000_0000000000000000_0010010100101111_0001101001001111"; -- 0.1452499810915257
	pesos_i(4824) := b"0000000000000000_0000000000000000_0001100101001000_1001000100000010"; -- 0.09876352600001877
	pesos_i(4825) := b"0000000000000000_0000000000000000_0010110011100111_0100000010010111"; -- 0.17540363003021656
	pesos_i(4826) := b"0000000000000000_0000000000000000_0001110101011001_1101001111110101"; -- 0.11465191579452307
	pesos_i(4827) := b"1111111111111111_1111111111111111_1110010011010010_0010011001010001"; -- -0.10616837039134862
	pesos_i(4828) := b"0000000000000000_0000000000000000_0000100000001111_1001110000101010"; -- 0.031488190040705126
	pesos_i(4829) := b"1111111111111111_1111111111111111_1111101111000001_1111000100111101"; -- -0.016571924807332963
	pesos_i(4830) := b"0000000000000000_0000000000000000_0010011100101010_0101011001000110"; -- 0.15298976143695164
	pesos_i(4831) := b"0000000000000000_0000000000000000_0010010010100101_0110000000000001"; -- 0.14314842238631972
	pesos_i(4832) := b"1111111111111111_1111111111111111_1110000000111111_0111011000001011"; -- -0.12403166032996892
	pesos_i(4833) := b"0000000000000000_0000000000000000_0000100010001101_0001011110001000"; -- 0.03340289189097419
	pesos_i(4834) := b"0000000000000000_0000000000000000_0010000001010100_0111001011010110"; -- 0.12628858304393675
	pesos_i(4835) := b"0000000000000000_0000000000000000_0000110011101101_0111111000111101"; -- 0.05049885751136128
	pesos_i(4836) := b"1111111111111111_1111111111111111_1110110100010000_1010011001100100"; -- -0.07396469172121402
	pesos_i(4837) := b"0000000000000000_0000000000000000_0000000000001111_1001101001110011"; -- 0.00023808776222236156
	pesos_i(4838) := b"0000000000000000_0000000000000000_0001000000110111_1000101111110101"; -- 0.06334757538048373
	pesos_i(4839) := b"0000000000000000_0000000000000000_0001111011110100_0011110001110010"; -- 0.12091424725067132
	pesos_i(4840) := b"1111111111111111_1111111111111111_1111101000000001_0110110001000001"; -- -0.02341578882729703
	pesos_i(4841) := b"1111111111111111_1111111111111111_1101100101111000_1110110000011110"; -- -0.15049862174235393
	pesos_i(4842) := b"1111111111111111_1111111111111111_1111110011101000_1010101111110010"; -- -0.012074712130352978
	pesos_i(4843) := b"1111111111111111_1111111111111111_1101111111011100_1100011011100110"; -- -0.1255374610542629
	pesos_i(4844) := b"1111111111111111_1111111111111111_1101011111000011_1010000011001001"; -- -0.15717120253482095
	pesos_i(4845) := b"1111111111111111_1111111111111111_1111101010010011_1101110001010100"; -- -0.021181325539553493
	pesos_i(4846) := b"0000000000000000_0000000000000000_0010000101010101_0111110101000000"; -- 0.1302107125001603
	pesos_i(4847) := b"0000000000000000_0000000000000000_0000010111000101_0000111010111010"; -- 0.02253810923317359
	pesos_i(4848) := b"0000000000000000_0000000000000000_0000110101010110_1010001100010100"; -- 0.05210322605077497
	pesos_i(4849) := b"1111111111111111_1111111111111111_1110000111110001_1010101000110011"; -- -0.11740623712843568
	pesos_i(4850) := b"1111111111111111_1111111111111111_1110110100110111_0100101101000110"; -- -0.07337502993251947
	pesos_i(4851) := b"0000000000000000_0000000000000000_0000110110111001_1000100011101001"; -- 0.05361228640819476
	pesos_i(4852) := b"1111111111111111_1111111111111111_1111111111011110_1111000000100010"; -- -0.0005044858211329536
	pesos_i(4853) := b"1111111111111111_1111111111111111_1111111000100000_1111101010010110"; -- -0.00730928269046603
	pesos_i(4854) := b"0000000000000000_0000000000000000_0010000100110010_0010101010011101"; -- 0.1296717293102685
	pesos_i(4855) := b"1111111111111111_1111111111111111_1110101100100010_0101100001101100"; -- -0.08150718083148985
	pesos_i(4856) := b"0000000000000000_0000000000000000_0010000111010101_0000000011111111"; -- 0.1321564313480932
	pesos_i(4857) := b"1111111111111111_1111111111111111_1111100110110011_1010111110100001"; -- -0.024601958571167037
	pesos_i(4858) := b"0000000000000000_0000000000000000_0010000010000111_1111110011110000"; -- 0.12707501273426092
	pesos_i(4859) := b"0000000000000000_0000000000000000_0000111101001101_0101111101110011"; -- 0.05977436605073263
	pesos_i(4860) := b"0000000000000000_0000000000000000_0010001111111001_1000011100101111"; -- 0.14052624605134345
	pesos_i(4861) := b"0000000000000000_0000000000000000_0000101111000110_1001010011100001"; -- 0.04599886407161355
	pesos_i(4862) := b"1111111111111111_1111111111111111_1110011111011000_0001011100001101"; -- -0.09435897768200263
	pesos_i(4863) := b"0000000000000000_0000000000000000_0000101100011010_1000101110000100"; -- 0.04337379432344289
	pesos_i(4864) := b"1111111111111111_1111111111111111_1111001010100010_1000111110111011"; -- -0.052207009212793365
	pesos_i(4865) := b"1111111111111111_1111111111111111_1111000111010010_0010001110011100"; -- -0.055387281777132695
	pesos_i(4866) := b"0000000000000000_0000000000000000_0000011001101000_0110100001000011"; -- 0.02503062856528387
	pesos_i(4867) := b"1111111111111111_1111111111111111_1111000101100001_1011001111110011"; -- -0.05710292165092649
	pesos_i(4868) := b"0000000000000000_0000000000000000_0000111001101011_0010011100011001"; -- 0.05632252092649035
	pesos_i(4869) := b"1111111111111111_1111111111111111_1110001100001011_1010000100011100"; -- -0.1131038004909764
	pesos_i(4870) := b"0000000000000000_0000000000000000_0010110010001110_0110111100111011"; -- 0.17404837786879582
	pesos_i(4871) := b"1111111111111111_1111111111111111_1110001011110111_1000000001111010"; -- -0.11341092125351555
	pesos_i(4872) := b"1111111111111111_1111111111111111_1110010100100011_1111101110001011"; -- -0.10491969927970589
	pesos_i(4873) := b"0000000000000000_0000000000000000_0010111100000010_1000000101000100"; -- 0.18363197239253476
	pesos_i(4874) := b"1111111111111111_1111111111111111_1111010010010000_1011101100110001"; -- -0.04466657694769629
	pesos_i(4875) := b"0000000000000000_0000000000000000_0000110010010000_0101100011111011"; -- 0.04907756915935853
	pesos_i(4876) := b"1111111111111111_1111111111111111_1111111101111101_1101111000100101"; -- -0.0019856605675408357
	pesos_i(4877) := b"1111111111111111_1111111111111111_1101101110011111_1000111110101110"; -- -0.14209653861057647
	pesos_i(4878) := b"0000000000000000_0000000000000000_0000011000101000_1001111101111001"; -- 0.02405735696714598
	pesos_i(4879) := b"1111111111111111_1111111111111111_1101100010011111_1011001110011001"; -- -0.15381314778397684
	pesos_i(4880) := b"0000000000000000_0000000000000000_0000101001110110_1010111110111000"; -- 0.040873510732053475
	pesos_i(4881) := b"1111111111111111_1111111111111111_1110011111111110_1001000011101101"; -- -0.09377187934772863
	pesos_i(4882) := b"1111111111111111_1111111111111111_1110010111001010_1001100110110110"; -- -0.10237731279851713
	pesos_i(4883) := b"0000000000000000_0000000000000000_0010001010100101_0010111100000110"; -- 0.13533300312243865
	pesos_i(4884) := b"0000000000000000_0000000000000000_0001110100111101_1101110010001110"; -- 0.11422518221468551
	pesos_i(4885) := b"0000000000000000_0000000000000000_0001011010111110_0010100100000010"; -- 0.08883911421923237
	pesos_i(4886) := b"0000000000000000_0000000000000000_0010100010111111_1000110000011011"; -- 0.15917277960857054
	pesos_i(4887) := b"0000000000000000_0000000000000000_0010010110010110_0110110000010111"; -- 0.14682651110176909
	pesos_i(4888) := b"1111111111111111_1111111111111111_1110000000110000_1111011111100010"; -- -0.1242528031131609
	pesos_i(4889) := b"1111111111111111_1111111111111111_1101011001101001_0001111010001100"; -- -0.16245850645214183
	pesos_i(4890) := b"1111111111111111_1111111111111111_1111011010001101_1011011110100100"; -- -0.036900064919060345
	pesos_i(4891) := b"0000000000000000_0000000000000000_0001000100001101_1110010101100010"; -- 0.06661828655912479
	pesos_i(4892) := b"0000000000000000_0000000000000000_0000110010101100_0100100000000010"; -- 0.04950380377855025
	pesos_i(4893) := b"0000000000000000_0000000000000000_0000100101100101_1110100101110001"; -- 0.036711301915032114
	pesos_i(4894) := b"1111111111111111_1111111111111111_1101010010010100_1011010000111001"; -- -0.16960595716489307
	pesos_i(4895) := b"1111111111111111_1111111111111111_1110111111110111_1000000000001011"; -- -0.06262969706696823
	pesos_i(4896) := b"0000000000000000_0000000000000000_0010011110011001_0001001010011110"; -- 0.15467945437518946
	pesos_i(4897) := b"0000000000000000_0000000000000000_0010010001011001_1110101000011000"; -- 0.1419969852662957
	pesos_i(4898) := b"0000000000000000_0000000000000000_0001010101000011_0000001010010010"; -- 0.08305374202932307
	pesos_i(4899) := b"0000000000000000_0000000000000000_0010100100110001_1100010010011111"; -- 0.16091565019565643
	pesos_i(4900) := b"1111111111111111_1111111111111111_1111000110110011_0001010111010010"; -- -0.05586112610116741
	pesos_i(4901) := b"0000000000000000_0000000000000000_0001100100000000_1000010111001011"; -- 0.097664224617844
	pesos_i(4902) := b"1111111111111111_1111111111111111_1110111011111000_0101101101011000"; -- -0.06652287590786803
	pesos_i(4903) := b"0000000000000000_0000000000000000_0010000101111010_1000001000110011"; -- 0.13077558283291205
	pesos_i(4904) := b"1111111111111111_1111111111111111_1101011001111001_1100101111111111"; -- -0.16220402749075816
	pesos_i(4905) := b"0000000000000000_0000000000000000_0001101100001101_0001001001110001"; -- 0.10566821353709284
	pesos_i(4906) := b"1111111111111111_1111111111111111_1111100101011001_1101111100111010"; -- -0.025972412412567706
	pesos_i(4907) := b"0000000000000000_0000000000000000_0000110110000001_0010100111010001"; -- 0.05275212618185921
	pesos_i(4908) := b"1111111111111111_1111111111111111_1110111001100000_0000000110111101"; -- -0.06884755270571111
	pesos_i(4909) := b"0000000000000000_0000000000000000_0000110011001000_0001010000000000"; -- 0.04992794995748827
	pesos_i(4910) := b"0000000000000000_0000000000000000_0010011111101101_1001000000001011"; -- 0.15596866864285555
	pesos_i(4911) := b"0000000000000000_0000000000000000_0000000111001101_0001001101111101"; -- 0.007035463239782469
	pesos_i(4912) := b"0000000000000000_0000000000000000_0000100010110011_1001011110111110"; -- 0.03399036779494333
	pesos_i(4913) := b"0000000000000000_0000000000000000_0010010000001111_1100111100110001"; -- 0.14086623149235666
	pesos_i(4914) := b"1111111111111111_1111111111111111_1101010000111000_0110011100001010"; -- -0.17101436615950344
	pesos_i(4915) := b"1111111111111111_1111111111111111_1110111111100010_0111100111111100"; -- -0.0629504929443593
	pesos_i(4916) := b"0000000000000000_0000000000000000_0001100001111110_0011011101001111"; -- 0.09567590404188639
	pesos_i(4917) := b"0000000000000000_0000000000000000_0000111010001110_1111000010011011"; -- 0.05686858935480701
	pesos_i(4918) := b"1111111111111111_1111111111111111_1101110101100010_1100001010111110"; -- -0.135211781248916
	pesos_i(4919) := b"1111111111111111_1111111111111111_1110101001110100_1111000001110010"; -- -0.08415314882488484
	pesos_i(4920) := b"0000000000000000_0000000000000000_0001011111000011_1011001110111000"; -- 0.09282992598819792
	pesos_i(4921) := b"1111111111111111_1111111111111111_1101100011110001_1111111010100001"; -- -0.15255745471843446
	pesos_i(4922) := b"0000000000000000_0000000000000000_0000100011001110_1101011010101101"; -- 0.03440610612980664
	pesos_i(4923) := b"1111111111111111_1111111111111111_1111110011010010_1111101111000101"; -- -0.012405647701613948
	pesos_i(4924) := b"0000000000000000_0000000000000000_0001100011111110_1001010010010000"; -- 0.0976345873912723
	pesos_i(4925) := b"1111111111111111_1111111111111111_1101010110011001_0110011011010011"; -- -0.16562802646336894
	pesos_i(4926) := b"1111111111111111_1111111111111111_1101110101001111_1110100010001000"; -- -0.13549944568338507
	pesos_i(4927) := b"0000000000000000_0000000000000000_0001010001001100_1101110100011000"; -- 0.07929784624099703
	pesos_i(4928) := b"0000000000000000_0000000000000000_0010100001000011_0100111010101100"; -- 0.15727702816748265
	pesos_i(4929) := b"1111111111111111_1111111111111111_1111101100101010_1110101100011100"; -- -0.01887636726346662
	pesos_i(4930) := b"0000000000000000_0000000000000000_0010110101100010_0111111100110100"; -- 0.17728419329254894
	pesos_i(4931) := b"0000000000000000_0000000000000000_0000101010110111_0001010101111001"; -- 0.041856138260843584
	pesos_i(4932) := b"0000000000000000_0000000000000000_0010000100100101_0111100111100100"; -- 0.1294780903439662
	pesos_i(4933) := b"1111111111111111_1111111111111111_1101011010001010_0110010001011110"; -- -0.16195080482776444
	pesos_i(4934) := b"0000000000000000_0000000000000000_0010000011000111_1010000011110101"; -- 0.12804609271421621
	pesos_i(4935) := b"0000000000000000_0000000000000000_0000100001011001_1101101011101100"; -- 0.03262108096357263
	pesos_i(4936) := b"1111111111111111_1111111111111111_1110000111111001_0001010111000111"; -- -0.11729301341509063
	pesos_i(4937) := b"0000000000000000_0000000000000000_0001000010011110_0001010111101001"; -- 0.06491219471282592
	pesos_i(4938) := b"1111111111111111_1111111111111111_1110100111010111_1110110001000000"; -- -0.08654902867166615
	pesos_i(4939) := b"0000000000000000_0000000000000000_0000110111011011_1001111001010011"; -- 0.0541323617424051
	pesos_i(4940) := b"0000000000000000_0000000000000000_0001101101000000_1011110101110001"; -- 0.10645660412983796
	pesos_i(4941) := b"0000000000000000_0000000000000000_0001101001110000_0111011011011111"; -- 0.10327856960528342
	pesos_i(4942) := b"0000000000000000_0000000000000000_0000001101000101_1110010000110110"; -- 0.012785208990393386
	pesos_i(4943) := b"1111111111111111_1111111111111111_1110100110010100_1011110001001100"; -- -0.0875742259032342
	pesos_i(4944) := b"0000000000000000_0000000000000000_0001011001010111_0010100010001100"; -- 0.08726743140974433
	pesos_i(4945) := b"0000000000000000_0000000000000000_0010100110101101_0010100010100000"; -- 0.16279844191171536
	pesos_i(4946) := b"0000000000000000_0000000000000000_0000001101001000_0000010111001010"; -- 0.012817727868423378
	pesos_i(4947) := b"0000000000000000_0000000000000000_0001010110110101_0110001001100101"; -- 0.0847989555619561
	pesos_i(4948) := b"1111111111111111_1111111111111111_1101010110100001_1111101000101001"; -- -0.16549717424173233
	pesos_i(4949) := b"0000000000000000_0000000000000000_0001101001101000_1101110101000110"; -- 0.10316260301491234
	pesos_i(4950) := b"1111111111111111_1111111111111111_1101010101000001_0101100011010111"; -- -0.16697163345036312
	pesos_i(4951) := b"1111111111111111_1111111111111111_1111011011000011_0110010110010100"; -- -0.03608098165255631
	pesos_i(4952) := b"0000000000000000_0000000000000000_0001010111000110_1011110111101001"; -- 0.08506380964743784
	pesos_i(4953) := b"1111111111111111_1111111111111111_1101101000111001_1001010010010000"; -- -0.14755889408081171
	pesos_i(4954) := b"0000000000000000_0000000000000000_0001100000011010_1000101011001011"; -- 0.09415500127635523
	pesos_i(4955) := b"0000000000000000_0000000000000000_0001100100111001_0001111110010101"; -- 0.09852788329828506
	pesos_i(4956) := b"1111111111111111_1111111111111111_1110000010000100_1010101110011110"; -- -0.12297561065785106
	pesos_i(4957) := b"1111111111111111_1111111111111111_1110010110000111_1000001010010001"; -- -0.103401031043868
	pesos_i(4958) := b"0000000000000000_0000000000000000_0001011001100100_0100110110110010"; -- 0.08746800990070322
	pesos_i(4959) := b"1111111111111111_1111111111111111_1101110010110111_0111111111011111"; -- -0.1378250198131307
	pesos_i(4960) := b"1111111111111111_1111111111111111_1110001011101001_1011100100101001"; -- -0.11362116574810259
	pesos_i(4961) := b"1111111111111111_1111111111111111_1111110100110111_0100110011110111"; -- -0.010874929246739792
	pesos_i(4962) := b"0000000000000000_0000000000000000_0001111100101010_1000101101101011"; -- 0.12174292913904661
	pesos_i(4963) := b"0000000000000000_0000000000000000_0001000110001101_1110100110001111"; -- 0.06857166034367851
	pesos_i(4964) := b"1111111111111111_1111111111111111_1111011110010011_0010010101001001"; -- -0.03291098566693913
	pesos_i(4965) := b"1111111111111111_1111111111111111_1110010011011001_1101000111101101"; -- -0.10605133019691403
	pesos_i(4966) := b"1111111111111111_1111111111111111_1111101010110101_0001001001101001"; -- -0.020674561867523915
	pesos_i(4967) := b"1111111111111111_1111111111111111_1111101111110110_0111110110001100"; -- -0.01577010475398455
	pesos_i(4968) := b"1111111111111111_1111111111111111_1110010100011111_0100111010000110"; -- -0.10499104712604554
	pesos_i(4969) := b"0000000000000000_0000000000000000_0010101101100111_0110101011111100"; -- 0.16954678206519355
	pesos_i(4970) := b"1111111111111111_1111111111111111_1101111001001100_1001111011110011"; -- -0.13164335802775948
	pesos_i(4971) := b"0000000000000000_0000000000000000_0001000011111100_1101010110100000"; -- 0.06635794798685278
	pesos_i(4972) := b"1111111111111111_1111111111111111_1111000000111001_0110110011111100"; -- -0.06162375306524189
	pesos_i(4973) := b"0000000000000000_0000000000000000_0000001000010101_0110000111110101"; -- 0.008138773353748114
	pesos_i(4974) := b"0000000000000000_0000000000000000_0001111000100110_1011110000001101"; -- 0.11777854275289
	pesos_i(4975) := b"1111111111111111_1111111111111111_1111010001000000_1110010010000010"; -- -0.04588481747451422
	pesos_i(4976) := b"1111111111111111_1111111111111111_1111000000001110_1000111100100101"; -- -0.06227784485515225
	pesos_i(4977) := b"0000000000000000_0000000000000000_0000011010011101_1110011100010000"; -- 0.025846902314723797
	pesos_i(4978) := b"1111111111111111_1111111111111111_1110111010101011_0011110101001101"; -- -0.06769959317357824
	pesos_i(4979) := b"1111111111111111_1111111111111111_1111010011110101_0010011111110001"; -- -0.04313421600886076
	pesos_i(4980) := b"0000000000000000_0000000000000000_0001110100001001_0011111100001000"; -- 0.11342233596486377
	pesos_i(4981) := b"1111111111111111_1111111111111111_1111111011110000_0011111100111001"; -- -0.004146622287984943
	pesos_i(4982) := b"1111111111111111_1111111111111111_1111110001011010_1000010101011000"; -- -0.014243760973585791
	pesos_i(4983) := b"0000000000000000_0000000000000000_0001100110100110_0000100000011111"; -- 0.10018969299140416
	pesos_i(4984) := b"0000000000000000_0000000000000000_0010000100010101_1100101111110110"; -- 0.1292388415158768
	pesos_i(4985) := b"0000000000000000_0000000000000000_0010001111110010_1101100110100111"; -- 0.14042435014717128
	pesos_i(4986) := b"1111111111111111_1111111111111111_1111111010001110_0110000001100000"; -- -0.005640007630663361
	pesos_i(4987) := b"1111111111111111_1111111111111111_1111111011000110_0100011100001010"; -- -0.004787025408053466
	pesos_i(4988) := b"1111111111111111_1111111111111111_1111101011110100_1110110000111010"; -- -0.019700275348237928
	pesos_i(4989) := b"1111111111111111_1111111111111111_1110010111101110_0001001010101100"; -- -0.10183604515808095
	pesos_i(4990) := b"0000000000000000_0000000000000000_0010100010111001_1010111101011111"; -- 0.15908332895427393
	pesos_i(4991) := b"0000000000000000_0000000000000000_0010011101100110_0000110010101110"; -- 0.15390090236332846
	pesos_i(4992) := b"1111111111111111_1111111111111111_1110101111100100_1000110101101011"; -- -0.07854381684150107
	pesos_i(4993) := b"0000000000000000_0000000000000000_0010101000111100_0100110001101001"; -- 0.1649825818244183
	pesos_i(4994) := b"0000000000000000_0000000000000000_0000011101100011_1110000001111011"; -- 0.028867750100279917
	pesos_i(4995) := b"1111111111111111_1111111111111111_1101111011011101_0111111000111000"; -- -0.1294327844199733
	pesos_i(4996) := b"1111111111111111_1111111111111111_1111001000100001_1111101101111110"; -- -0.054168969946948954
	pesos_i(4997) := b"0000000000000000_0000000000000000_0010011000010011_0100111011111110"; -- 0.14873212535649238
	pesos_i(4998) := b"1111111111111111_1111111111111111_1110011100000101_1001100000010010"; -- -0.09757089197450179
	pesos_i(4999) := b"0000000000000000_0000000000000000_0010100111110111_0010010111100011"; -- 0.16392742903991056
	pesos_i(5000) := b"1111111111111111_1111111111111111_1111111100110011_1100100111010011"; -- -0.0031160221618879947
	pesos_i(5001) := b"0000000000000000_0000000000000000_0000101001000111_0011000111000011"; -- 0.04014883994876891
	pesos_i(5002) := b"0000000000000000_0000000000000000_0010110110101010_0000011111000000"; -- 0.1783757061608523
	pesos_i(5003) := b"1111111111111111_1111111111111111_1111000111000110_0001000111110111"; -- -0.05557143886665335
	pesos_i(5004) := b"0000000000000000_0000000000000000_0010100011000000_1101110001101011"; -- 0.15919282539559396
	pesos_i(5005) := b"1111111111111111_1111111111111111_1101010101011010_1000101001101010"; -- -0.16658720886328562
	pesos_i(5006) := b"1111111111111111_1111111111111111_1111111100011001_0011100011001011"; -- -0.003521395062459097
	pesos_i(5007) := b"1111111111111111_1111111111111111_1111010010100011_1011110111111100"; -- -0.044376493393213375
	pesos_i(5008) := b"1111111111111111_1111111111111111_1111011000111001_1110000100010111"; -- -0.03817933271404075
	pesos_i(5009) := b"1111111111111111_1111111111111111_1111101011000000_1001111101111111"; -- -0.02049830580059281
	pesos_i(5010) := b"0000000000000000_0000000000000000_0010010111111000_0011010011000110"; -- 0.14831857532315337
	pesos_i(5011) := b"0000000000000000_0000000000000000_0010100010111101_0110000111110101"; -- 0.15913974988068413
	pesos_i(5012) := b"1111111111111111_1111111111111111_1111100110110010_1001100101110100"; -- -0.024618538990561982
	pesos_i(5013) := b"1111111111111111_1111111111111111_1110011010110101_0101111000100111"; -- -0.09879504724332656
	pesos_i(5014) := b"0000000000000000_0000000000000000_0010000000100111_1010010001010001"; -- 0.12560488672912892
	pesos_i(5015) := b"1111111111111111_1111111111111111_1101001000111110_0110101010101101"; -- -0.17873509677252258
	pesos_i(5016) := b"1111111111111111_1111111111111111_1111001001001011_1101111100001111"; -- -0.05352979547541874
	pesos_i(5017) := b"1111111111111111_1111111111111111_1111111011011101_1100110111100111"; -- -0.004428034846450735
	pesos_i(5018) := b"1111111111111111_1111111111111111_1101011101010111_1100001110011111"; -- -0.1588170754617178
	pesos_i(5019) := b"1111111111111111_1111111111111111_1101111010001000_1100100110110111"; -- -0.13072528154222487
	pesos_i(5020) := b"1111111111111111_1111111111111111_1111011100101011_1001100111111110"; -- -0.0344909433329775
	pesos_i(5021) := b"0000000000000000_0000000000000000_0010110010000101_0010111101110100"; -- 0.17390724731061227
	pesos_i(5022) := b"1111111111111111_1111111111111111_1101111111111001_0101000101110010"; -- -0.1251019569527699
	pesos_i(5023) := b"0000000000000000_0000000000000000_0000001010100001_1001110011010101"; -- 0.010278512929069283
	pesos_i(5024) := b"0000000000000000_0000000000000000_0000111111010011_1100000111101101"; -- 0.06182491336213325
	pesos_i(5025) := b"0000000000000000_0000000000000000_0001000010010101_1011001010110001"; -- 0.06478421033162751
	pesos_i(5026) := b"0000000000000000_0000000000000000_0010000000001001_1001010110011010"; -- 0.12514624615295658
	pesos_i(5027) := b"1111111111111111_1111111111111111_1110110100010100_0010110010110101"; -- -0.07391090950969711
	pesos_i(5028) := b"0000000000000000_0000000000000000_0000001111110100_0000011110100010"; -- 0.015442349550070277
	pesos_i(5029) := b"0000000000000000_0000000000000000_0000100110101001_0110011111100001"; -- 0.037741176968435514
	pesos_i(5030) := b"0000000000000000_0000000000000000_0001010111011011_1100010001110010"; -- 0.08538463374455181
	pesos_i(5031) := b"1111111111111111_1111111111111111_1101010001011000_0111111100100000"; -- -0.17052464926926061
	pesos_i(5032) := b"1111111111111111_1111111111111111_1101101100111010_1101100011000011"; -- -0.14363332025465797
	pesos_i(5033) := b"1111111111111111_1111111111111111_1111111111000011_1110010011001110"; -- -0.0009171482883337425
	pesos_i(5034) := b"1111111111111111_1111111111111111_1110111011101001_1100010011010110"; -- -0.06674546974448335
	pesos_i(5035) := b"1111111111111111_1111111111111111_1110101001000001_0011110111101101"; -- -0.08494198766863487
	pesos_i(5036) := b"1111111111111111_1111111111111111_1111001011110111_1011100111010111"; -- -0.05090750207510146
	pesos_i(5037) := b"1111111111111111_1111111111111111_1101110110001010_0011110001101101"; -- -0.13460943535410294
	pesos_i(5038) := b"1111111111111111_1111111111111111_1111010011000101_0000010010110101"; -- -0.0438687380640973
	pesos_i(5039) := b"1111111111111111_1111111111111111_1111011010101110_1101101010000101"; -- -0.036394445890872804
	pesos_i(5040) := b"1111111111111111_1111111111111111_1101001111011100_0010000110000111"; -- -0.17242231804401523
	pesos_i(5041) := b"1111111111111111_1111111111111111_1101101000101100_0001110010110000"; -- -0.1477644033131161
	pesos_i(5042) := b"0000000000000000_0000000000000000_0010011010100011_1000000011000011"; -- 0.15093235735475383
	pesos_i(5043) := b"1111111111111111_1111111111111111_1101111101010001_1001010101000000"; -- -0.1276613921430701
	pesos_i(5044) := b"1111111111111111_1111111111111111_1101010110110110_1000111101011100"; -- -0.1651831054379505
	pesos_i(5045) := b"1111111111111111_1111111111111111_1110001110011001_0101001011100110"; -- -0.11094171420642619
	pesos_i(5046) := b"0000000000000000_0000000000000000_0010100010100001_0110001101100100"; -- 0.15871258929288398
	pesos_i(5047) := b"1111111111111111_1111111111111111_1111100011100011_0011111000011000"; -- -0.027782553880411537
	pesos_i(5048) := b"0000000000000000_0000000000000000_0010010000001101_1110001000110001"; -- 0.14083684634628688
	pesos_i(5049) := b"0000000000000000_0000000000000000_0001111001111110_0001010010101010"; -- 0.1191113391747216
	pesos_i(5050) := b"1111111111111111_1111111111111111_1110101110111010_0110111010010100"; -- -0.07918652430095394
	pesos_i(5051) := b"0000000000000000_0000000000000000_0001100110100010_1100110110110000"; -- 0.10014043377998641
	pesos_i(5052) := b"1111111111111111_1111111111111111_1101101100110100_0000111010111011"; -- -0.14373691506297145
	pesos_i(5053) := b"1111111111111111_1111111111111111_1111001110100010_0100110011111111"; -- -0.04830473688307712
	pesos_i(5054) := b"0000000000000000_0000000000000000_0000000101110111_0100100011011010"; -- 0.005726388150478499
	pesos_i(5055) := b"0000000000000000_0000000000000000_0000111101110000_1111010111010110"; -- 0.060317387281415
	pesos_i(5056) := b"0000000000000000_0000000000000000_0001001010110100_0000110000010010"; -- 0.07305980136458406
	pesos_i(5057) := b"1111111111111111_1111111111111111_1111101101001100_0010111000110111"; -- -0.018368827396561364
	pesos_i(5058) := b"1111111111111111_1111111111111111_1101111100100111_0000100000110111"; -- -0.1283106676109502
	pesos_i(5059) := b"1111111111111111_1111111111111111_1111000101101111_1001110100100110"; -- -0.05689065764292823
	pesos_i(5060) := b"0000000000000000_0000000000000000_0000010100010011_1010110011111111"; -- 0.01983147830871874
	pesos_i(5061) := b"1111111111111111_1111111111111111_1110010100001110_1010111000000111"; -- -0.1052447541434525
	pesos_i(5062) := b"1111111111111111_1111111111111111_1110011111000000_0010001111010101"; -- -0.09472442683197513
	pesos_i(5063) := b"1111111111111111_1111111111111111_1111001011110110_1110111101101010"; -- -0.05091956779478847
	pesos_i(5064) := b"1111111111111111_1111111111111111_1111010100110101_1110001001000111"; -- -0.04214654706326958
	pesos_i(5065) := b"0000000000000000_0000000000000000_0010001111110010_0011111010001110"; -- 0.14041510552347983
	pesos_i(5066) := b"0000000000000000_0000000000000000_0001110110110000_0001010011110111"; -- 0.11596804650790336
	pesos_i(5067) := b"1111111111111111_1111111111111111_1110110100001100_1001011110000001"; -- -0.07402661416886379
	pesos_i(5068) := b"0000000000000000_0000000000000000_0010000010001010_1010110001110110"; -- 0.12711599232096688
	pesos_i(5069) := b"0000000000000000_0000000000000000_0010001110000110_0000110100100101"; -- 0.13876421113483803
	pesos_i(5070) := b"0000000000000000_0000000000000000_0001100111001011_0001000110101011"; -- 0.10075483716474969
	pesos_i(5071) := b"1111111111111111_1111111111111111_1110001100100000_1101001011010111"; -- -0.11278040172161746
	pesos_i(5072) := b"1111111111111111_1111111111111111_1110010010000010_1101101000111010"; -- -0.10737835014808461
	pesos_i(5073) := b"1111111111111111_1111111111111111_1110110011110100_1000001100110111"; -- -0.07439403442356944
	pesos_i(5074) := b"0000000000000000_0000000000000000_0001000111001011_1001001000000001"; -- 0.06951248669031981
	pesos_i(5075) := b"1111111111111111_1111111111111111_1101011011011001_1110000100111000"; -- -0.1607379186147032
	pesos_i(5076) := b"1111111111111111_1111111111111111_1111110110011100_0101100011001001"; -- -0.009333086915755719
	pesos_i(5077) := b"0000000000000000_0000000000000000_0001101100010000_0010101010100101"; -- 0.10571543255153937
	pesos_i(5078) := b"1111111111111111_1111111111111111_1111101111111010_0010101010110011"; -- -0.015714007691348526
	pesos_i(5079) := b"0000000000000000_0000000000000000_0001101101011110_0001100100110001"; -- 0.10690457776420918
	pesos_i(5080) := b"0000000000000000_0000000000000000_0000101011100101_1110000111011101"; -- 0.04257022521910518
	pesos_i(5081) := b"1111111111111111_1111111111111111_1111110100110000_1110110111110111"; -- -0.010972144408659883
	pesos_i(5082) := b"1111111111111111_1111111111111111_1111011001000000_1011100001010001"; -- -0.038074951271257665
	pesos_i(5083) := b"1111111111111111_1111111111111111_1111111011100101_1010010100110001"; -- -0.004308391017556714
	pesos_i(5084) := b"1111111111111111_1111111111111111_1101101000000001_0010110001011011"; -- -0.14841959752796655
	pesos_i(5085) := b"0000000000000000_0000000000000000_0001101011101101_0100000110011010"; -- 0.10518274318828301
	pesos_i(5086) := b"0000000000000000_0000000000000000_0001100011010100_0100010100101100"; -- 0.09698898621264916
	pesos_i(5087) := b"0000000000000000_0000000000000000_0001011011000001_1011011000010110"; -- 0.08889329934120796
	pesos_i(5088) := b"0000000000000000_0000000000000000_0010011100010000_0110100010111101"; -- 0.1525941334278739
	pesos_i(5089) := b"0000000000000000_0000000000000000_0000110010010010_1010011010100110"; -- 0.049112716248702074
	pesos_i(5090) := b"1111111111111111_1111111111111111_1111100001111000_1001001001110011"; -- -0.02941021624188384
	pesos_i(5091) := b"1111111111111111_1111111111111111_1110110100011010_1100101100001110"; -- -0.07380991839542762
	pesos_i(5092) := b"0000000000000000_0000000000000000_0000000101000000_1110010100111010"; -- 0.00489647541111574
	pesos_i(5093) := b"0000000000000000_0000000000000000_0001110111001011_0111011101011010"; -- 0.11638589808236156
	pesos_i(5094) := b"1111111111111111_1111111111111111_1101011110100111_1110011100111110"; -- -0.1575942492247595
	pesos_i(5095) := b"0000000000000000_0000000000000000_0001001111100011_0010100110001110"; -- 0.0776849718827923
	pesos_i(5096) := b"1111111111111111_1111111111111111_1101101110101000_1101001000001100"; -- -0.1419552536652972
	pesos_i(5097) := b"1111111111111111_1111111111111111_1110011110010101_1110000000010001"; -- -0.0953693350284625
	pesos_i(5098) := b"0000000000000000_0000000000000000_0001111101100100_0010110010100001"; -- 0.12262228893548513
	pesos_i(5099) := b"1111111111111111_1111111111111111_1111111101000001_0001001101101111"; -- -0.002913270458714409
	pesos_i(5100) := b"0000000000000000_0000000000000000_0010001110010101_1010110001110111"; -- 0.13900258937130255
	pesos_i(5101) := b"0000000000000000_0000000000000000_0010001101011111_0100010011001110"; -- 0.13817243607729188
	pesos_i(5102) := b"0000000000000000_0000000000000000_0000111000101010_1101010100000000"; -- 0.05534106498138552
	pesos_i(5103) := b"1111111111111111_1111111111111111_1100111011001111_1100101000011100"; -- -0.1921418839251084
	pesos_i(5104) := b"1111111111111111_1111111111111111_1110101010110001_1110110010111010"; -- -0.08322258431103845
	pesos_i(5105) := b"0000000000000000_0000000000000000_0000101011011001_1000000101010111"; -- 0.04238136657237432
	pesos_i(5106) := b"0000000000000000_0000000000000000_0000110101001000_1101010011110101"; -- 0.05189257614559039
	pesos_i(5107) := b"1111111111111111_1111111111111111_1110110001110101_0001100111010110"; -- -0.0763381818423866
	pesos_i(5108) := b"0000000000000000_0000000000000000_0001110100111001_1111100110100011"; -- 0.11416588045573596
	pesos_i(5109) := b"0000000000000000_0000000000000000_0001110101101001_1001101110100100"; -- 0.11489269970210432
	pesos_i(5110) := b"0000000000000000_0000000000000000_0001111001000000_1000010100000001"; -- 0.11817199015739888
	pesos_i(5111) := b"0000000000000000_0000000000000000_0001100001000011_0001000001001100"; -- 0.09477331030396825
	pesos_i(5112) := b"1111111111111111_1111111111111111_1111100001001100_1010010010000101"; -- -0.030080525913506823
	pesos_i(5113) := b"1111111111111111_1111111111111111_1101011101001010_0110000100111001"; -- -0.15902130465870382
	pesos_i(5114) := b"1111111111111111_1111111111111111_1101011011011111_1111001111001010"; -- -0.16064525910788138
	pesos_i(5115) := b"0000000000000000_0000000000000000_0010110010001011_1100100001100001"; -- 0.17400791518912564
	pesos_i(5116) := b"1111111111111111_1111111111111111_1110011000110110_0110110011100100"; -- -0.10073203492523031
	pesos_i(5117) := b"1111111111111111_1111111111111111_1111110111110100_1010100111110011"; -- -0.007985475683331102
	pesos_i(5118) := b"1111111111111111_1111111111111111_1101100101010100_1110101010100011"; -- -0.15104802638520526
	pesos_i(5119) := b"0000000000000000_0000000000000000_0000100001001100_1100100111010000"; -- 0.03242169699194519
	pesos_i(5120) := b"0000000000000000_0000000000000000_0001010010101101_1000100000101011"; -- 0.08077288684857623
	pesos_i(5121) := b"0000000000000000_0000000000000000_0000101001000000_1011000110111001"; -- 0.040049655632300354
	pesos_i(5122) := b"1111111111111111_1111111111111111_1111100100001001_0100000000110000"; -- -0.027202595011281885
	pesos_i(5123) := b"1111111111111111_1111111111111111_1110010000010101_1100111001111011"; -- -0.10904225814231158
	pesos_i(5124) := b"1111111111111111_1111111111111111_1111111111010101_0010010101011101"; -- -0.0006539009962801701
	pesos_i(5125) := b"1111111111111111_1111111111111111_1110010100010101_1101101111000010"; -- -0.10513521686939337
	pesos_i(5126) := b"0000000000000000_0000000000000000_0000001101010010_1011111001001000"; -- 0.012981312333715293
	pesos_i(5127) := b"1111111111111111_1111111111111111_1111111100111110_1110011111110110"; -- -0.0029463791102462547
	pesos_i(5128) := b"1111111111111111_1111111111111111_1101001100000110_1010000110011011"; -- -0.1756800647397925
	pesos_i(5129) := b"0000000000000000_0000000000000000_0010000111001011_1100010101101100"; -- 0.13201555138581353
	pesos_i(5130) := b"1111111111111111_1111111111111111_1101110111100101_0111111101000100"; -- -0.13321690161550337
	pesos_i(5131) := b"1111111111111111_1111111111111111_1110110011110011_0011000111010101"; -- -0.07441414409863206
	pesos_i(5132) := b"1111111111111111_1111111111111111_1111001011011101_1111100010111010"; -- -0.05130048233749264
	pesos_i(5133) := b"1111111111111111_1111111111111111_1101111110110100_1001000101010100"; -- -0.1261510056753362
	pesos_i(5134) := b"0000000000000000_0000000000000000_0001010111000001_1100010110000101"; -- 0.08498796930555516
	pesos_i(5135) := b"0000000000000000_0000000000000000_0000010101000111_0010101010001011"; -- 0.020617159816004534
	pesos_i(5136) := b"0000000000000000_0000000000000000_0000001100110111_1011010100101100"; -- 0.012568781987887717
	pesos_i(5137) := b"1111111111111111_1111111111111111_1110000101101100_0110100110100111"; -- -0.1194395032967081
	pesos_i(5138) := b"0000000000000000_0000000000000000_0010010001100110_0000001110011111"; -- 0.1421816123262145
	pesos_i(5139) := b"0000000000000000_0000000000000000_0000100011011001_0011011011010110"; -- 0.03456442581766376
	pesos_i(5140) := b"1111111111111111_1111111111111111_1111100010100011_0011000010101010"; -- -0.02875991685553509
	pesos_i(5141) := b"0000000000000000_0000000000000000_0001100000011011_1001110001100010"; -- 0.09417130843284101
	pesos_i(5142) := b"0000000000000000_0000000000000000_0010101001000001_0001010010011110"; -- 0.16505555022606438
	pesos_i(5143) := b"0000000000000000_0000000000000000_0000100100010100_0011110011010001"; -- 0.035465050690946756
	pesos_i(5144) := b"1111111111111111_1111111111111111_1111000001100101_1001110000011101"; -- -0.06094955734419297
	pesos_i(5145) := b"0000000000000000_0000000000000000_0000101011111111_0101001101101100"; -- 0.04295846348361302
	pesos_i(5146) := b"0000000000000000_0000000000000000_0011010010001000_0110100001011011"; -- 0.20520641546696988
	pesos_i(5147) := b"0000000000000000_0000000000000000_0000100110110101_1011111101100100"; -- 0.03792949864600733
	pesos_i(5148) := b"0000000000000000_0000000000000000_0000110110011110_1101011001001101"; -- 0.053204912016276446
	pesos_i(5149) := b"0000000000000000_0000000000000000_0000001011100001_1000100101111010"; -- 0.011253921666751742
	pesos_i(5150) := b"1111111111111111_1111111111111111_1101101011000000_1110010001100101"; -- -0.145494199105468
	pesos_i(5151) := b"1111111111111111_1111111111111111_1101011101000011_1010011010010100"; -- -0.15912398223475985
	pesos_i(5152) := b"1111111111111111_1111111111111111_1110111111101101_1011100110010011"; -- -0.06277885601722794
	pesos_i(5153) := b"1111111111111111_1111111111111111_1100111101011001_1001011000110101"; -- -0.19003926469004342
	pesos_i(5154) := b"1111111111111111_1111111111111111_1101010000010010_0001000100001010"; -- -0.17159932608131817
	pesos_i(5155) := b"0000000000000000_0000000000000000_0010110011011000_0111100000011001"; -- 0.1751780567566982
	pesos_i(5156) := b"0000000000000000_0000000000000000_0001101001001010_1001001111011111"; -- 0.10270046417276603
	pesos_i(5157) := b"0000000000000000_0000000000000000_0001110000111100_1001000010011010"; -- 0.11029914625619396
	pesos_i(5158) := b"0000000000000000_0000000000000000_0010010101001101_0011110111001100"; -- 0.1457098602404448
	pesos_i(5159) := b"0000000000000000_0000000000000000_0001101001011001_0111000011110111"; -- 0.1029272653613931
	pesos_i(5160) := b"0000000000000000_0000000000000000_0000111011101010_0111110010110000"; -- 0.05826548862770878
	pesos_i(5161) := b"1111111111111111_1111111111111111_1111101010100110_0000110101000111"; -- -0.020903749628107662
	pesos_i(5162) := b"1111111111111111_1111111111111111_1101110000100010_1111100110011010"; -- -0.14009132384473724
	pesos_i(5163) := b"1111111111111111_1111111111111111_1110100111011111_1001101101101111"; -- -0.08643177553211542
	pesos_i(5164) := b"0000000000000000_0000000000000000_0010010110011011_0101010110101100"; -- 0.14690146881164526
	pesos_i(5165) := b"0000000000000000_0000000000000000_0001010000001011_1100011001100101"; -- 0.07830467197168985
	pesos_i(5166) := b"0000000000000000_0000000000000000_0011001010011100_1111101101100111"; -- 0.19770785592488704
	pesos_i(5167) := b"0000000000000000_0000000000000000_0001010000011111_0110110111001110"; -- 0.07860456737490076
	pesos_i(5168) := b"0000000000000000_0000000000000000_0010011110010101_0111010000101111"; -- 0.15462423454413957
	pesos_i(5169) := b"0000000000000000_0000000000000000_0001111111110011_0000011011111100"; -- 0.12480205215427519
	pesos_i(5170) := b"0000000000000000_0000000000000000_0000110101011000_1111000101101001"; -- 0.05213841271649888
	pesos_i(5171) := b"1111111111111111_1111111111111111_1111010010011101_1000000001010001"; -- -0.04447172185403575
	pesos_i(5172) := b"1111111111111111_1111111111111111_1111000111101100_0110111010101111"; -- -0.054986078592957094
	pesos_i(5173) := b"1111111111111111_1111111111111111_1110000011011110_1010111100011111"; -- -0.12160211083500085
	pesos_i(5174) := b"1111111111111111_1111111111111111_1110101110011101_0110011100111100"; -- -0.07962946683816054
	pesos_i(5175) := b"1111111111111111_1111111111111111_1110001100011110_0111101001111000"; -- -0.11281618664538527
	pesos_i(5176) := b"0000000000000000_0000000000000000_0010011100000011_0001110101101111"; -- 0.15239128078961703
	pesos_i(5177) := b"0000000000000000_0000000000000000_0010100110101010_0110010001010110"; -- 0.16275622460268682
	pesos_i(5178) := b"1111111111111111_1111111111111111_1110010111000000_0101100000111101"; -- -0.10253380305404919
	pesos_i(5179) := b"1111111111111111_1111111111111111_1110101011001110_1000011000010000"; -- -0.08278619882039819
	pesos_i(5180) := b"0000000000000000_0000000000000000_0001000111001000_1001010111010111"; -- 0.0694669390401413
	pesos_i(5181) := b"1111111111111111_1111111111111111_1111111111100111_1000100001100001"; -- -0.0003733409992687861
	pesos_i(5182) := b"0000000000000000_0000000000000000_0000101100000011_0110100111000000"; -- 0.04302082949181574
	pesos_i(5183) := b"1111111111111111_1111111111111111_1111000001100000_1111100101011001"; -- -0.06102029403045712
	pesos_i(5184) := b"1111111111111111_1111111111111111_1111000101001001_0100101101010000"; -- -0.05747536937172093
	pesos_i(5185) := b"1111111111111111_1111111111111111_1111110001001111_0100100010001011"; -- -0.014415231684832197
	pesos_i(5186) := b"0000000000000000_0000000000000000_0001000011010000_0000110011100000"; -- 0.06567459558613321
	pesos_i(5187) := b"1111111111111111_1111111111111111_1101110001101100_0011110010001000"; -- -0.13897344276250487
	pesos_i(5188) := b"1111111111111111_1111111111111111_1111001011110010_0001110010111100"; -- -0.0509931603526488
	pesos_i(5189) := b"1111111111111111_1111111111111111_1110101111110100_1101110101011011"; -- -0.07829491162869445
	pesos_i(5190) := b"1111111111111111_1111111111111111_1110010000101111_0111111100111101"; -- -0.10865025287552876
	pesos_i(5191) := b"0000000000000000_0000000000000000_0010000101001001_1111110101111001"; -- 0.1300352498374114
	pesos_i(5192) := b"1111111111111111_1111111111111111_1110011110011111_1001011101011011"; -- -0.09522108106848134
	pesos_i(5193) := b"1111111111111111_1111111111111111_1101111011011100_0111110111110111"; -- -0.12944805827562184
	pesos_i(5194) := b"0000000000000000_0000000000000000_0010001000111010_0010110000011010"; -- 0.13370013850355164
	pesos_i(5195) := b"1111111111111111_1111111111111111_1111101000111010_1110011100100000"; -- -0.022538714177224698
	pesos_i(5196) := b"0000000000000000_0000000000000000_0001010101111010_1001011110111001"; -- 0.08390186565797295
	pesos_i(5197) := b"1111111111111111_1111111111111111_1110010000010100_1101100110100110"; -- -0.10905685124983316
	pesos_i(5198) := b"1111111111111111_1111111111111111_1101101010100000_0110100001010010"; -- -0.14598987587249293
	pesos_i(5199) := b"0000000000000000_0000000000000000_0000101111101010_0000011010000101"; -- 0.04653969526418922
	pesos_i(5200) := b"0000000000000000_0000000000000000_0000001011111111_0111111000011001"; -- 0.011711007233398157
	pesos_i(5201) := b"0000000000000000_0000000000000000_0001101111011011_0110001000001100"; -- 0.10881626874170731
	pesos_i(5202) := b"0000000000000000_0000000000000000_0010101100011101_1100111111100111"; -- 0.16842364684631472
	pesos_i(5203) := b"1111111111111111_1111111111111111_1111011110001111_0111100110101101"; -- -0.03296699071846933
	pesos_i(5204) := b"0000000000000000_0000000000000000_0000110101001111_1010000101010001"; -- 0.051996309636721035
	pesos_i(5205) := b"0000000000000000_0000000000000000_0010100000011010_0000001110010010"; -- 0.15664694142751326
	pesos_i(5206) := b"0000000000000000_0000000000000000_0000111100000110_0100001010100101"; -- 0.058689275139408754
	pesos_i(5207) := b"1111111111111111_1111111111111111_1111010110010011_1111000010100011"; -- -0.04071136494777167
	pesos_i(5208) := b"1111111111111111_1111111111111111_1111111000110000_0011001110111101"; -- -0.00707699434335926
	pesos_i(5209) := b"1111111111111111_1111111111111111_1101011100001001_0011100110000111"; -- -0.1600154920690275
	pesos_i(5210) := b"0000000000000000_0000000000000000_0010100010100000_1111011111010000"; -- 0.15870617707887277
	pesos_i(5211) := b"0000000000000000_0000000000000000_0000110111111101_0010101000000000"; -- 0.054644227053740696
	pesos_i(5212) := b"0000000000000000_0000000000000000_0000111001010110_0100000000101010"; -- 0.05600358039270852
	pesos_i(5213) := b"1111111111111111_1111111111111111_1111000001100111_1110000101010100"; -- -0.06091491403115696
	pesos_i(5214) := b"1111111111111111_1111111111111111_1111010101111110_0111011000010011"; -- -0.041039104870575584
	pesos_i(5215) := b"0000000000000000_0000000000000000_0000110001011001_0100101011101011"; -- 0.04823749764520682
	pesos_i(5216) := b"1111111111111111_1111111111111111_1110001011101111_0111111010110111"; -- -0.11353309662312451
	pesos_i(5217) := b"1111111111111111_1111111111111111_1111100000110001_0000011100101001"; -- -0.030501892623065335
	pesos_i(5218) := b"1111111111111111_1111111111111111_1111110101001110_1111011000001101"; -- -0.010513898584723206
	pesos_i(5219) := b"1111111111111111_1111111111111111_1101111111110100_0000011110010100"; -- -0.12518265370898582
	pesos_i(5220) := b"0000000000000000_0000000000000000_0001000111101010_0111011000110100"; -- 0.06998385200019686
	pesos_i(5221) := b"0000000000000000_0000000000000000_0001101101011110_1011111101010001"; -- 0.1069144794122919
	pesos_i(5222) := b"1111111111111111_1111111111111111_1110000100011100_1100111000101011"; -- -0.12065421541984911
	pesos_i(5223) := b"1111111111111111_1111111111111111_1111001111001000_0000011110100011"; -- -0.04772903692813571
	pesos_i(5224) := b"0000000000000000_0000000000000000_0000100010101001_1110010000011001"; -- 0.033842331034672934
	pesos_i(5225) := b"0000000000000000_0000000000000000_0001011001000010_1011011101111011"; -- 0.0869555162553818
	pesos_i(5226) := b"1111111111111111_1111111111111111_1111000001101111_1101111011111110"; -- -0.0607929829401561
	pesos_i(5227) := b"1111111111111111_1111111111111111_1110001010101100_1101111000100100"; -- -0.11454974776230102
	pesos_i(5228) := b"0000000000000000_0000000000000000_0000000110001010_1000000101100001"; -- 0.006019674494696084
	pesos_i(5229) := b"0000000000000000_0000000000000000_0000010111110100_0101111000010010"; -- 0.023260001532837925
	pesos_i(5230) := b"0000000000000000_0000000000000000_0000110100011001_0101101001101011"; -- 0.05116810914556432
	pesos_i(5231) := b"0000000000000000_0000000000000000_0001111100001001_1000010110101000"; -- 0.12123904566079029
	pesos_i(5232) := b"0000000000000000_0000000000000000_0000010100000110_0010001001000011"; -- 0.019624844919616136
	pesos_i(5233) := b"0000000000000000_0000000000000000_0010000100000011_1111110011111100"; -- 0.12896710537407477
	pesos_i(5234) := b"0000000000000000_0000000000000000_0001101101111011_0101101000100111"; -- 0.1073509546432023
	pesos_i(5235) := b"0000000000000000_0000000000000000_0010110000111110_1000101010100110"; -- 0.1728293089268391
	pesos_i(5236) := b"1111111111111111_1111111111111111_1110100010101001_0110000000010000"; -- -0.09116553879593556
	pesos_i(5237) := b"0000000000000000_0000000000000000_0000101101100110_1011001000000111"; -- 0.044535757635114456
	pesos_i(5238) := b"0000000000000000_0000000000000000_0010011001100011_1001011001111111"; -- 0.1499570903032573
	pesos_i(5239) := b"0000000000000000_0000000000000000_0000111101101110_1101101000010011"; -- 0.06028521499318453
	pesos_i(5240) := b"0000000000000000_0000000000000000_0000111100111100_1001001001111110"; -- 0.059518008993833554
	pesos_i(5241) := b"0000000000000000_0000000000000000_0001100111001010_0010100100101111"; -- 0.10074098013756931
	pesos_i(5242) := b"0000000000000000_0000000000000000_0010100010001111_0111000101010101"; -- 0.15843876198125273
	pesos_i(5243) := b"1111111111111111_1111111111111111_1111001110110111_0000110000100111"; -- -0.047988167344124255
	pesos_i(5244) := b"1111111111111111_1111111111111111_1101001110101011_0100001000001000"; -- -0.17316806135670185
	pesos_i(5245) := b"0000000000000000_0000000000000000_0001010000101001_0101000000000111"; -- 0.07875538036071891
	pesos_i(5246) := b"1111111111111111_1111111111111111_1111010010001010_1101000011011001"; -- -0.044756838865527615
	pesos_i(5247) := b"0000000000000000_0000000000000000_0000100111111011_1101110101011101"; -- 0.03899940030675665
	pesos_i(5248) := b"0000000000000000_0000000000000000_0001001100101000_0000110010101110"; -- 0.07482985725092758
	pesos_i(5249) := b"0000000000000000_0000000000000000_0010011101010100_0010000010101111"; -- 0.1536274363672157
	pesos_i(5250) := b"1111111111111111_1111111111111111_1111011010100111_1101010110010100"; -- -0.03650155208382587
	pesos_i(5251) := b"0000000000000000_0000000000000000_0001010100010101_0010101000101000"; -- 0.0823541973622123
	pesos_i(5252) := b"0000000000000000_0000000000000000_0000001010110110_1100101111110000"; -- 0.010601755268356536
	pesos_i(5253) := b"0000000000000000_0000000000000000_0001100111001010_0010111101011110"; -- 0.10074134873382479
	pesos_i(5254) := b"0000000000000000_0000000000000000_0000000110110001_1000001000110111"; -- 0.006614817036806728
	pesos_i(5255) := b"0000000000000000_0000000000000000_0000001001000001_1000011110111001"; -- 0.00881241108893624
	pesos_i(5256) := b"1111111111111111_1111111111111111_1111011100100100_0010101000000010"; -- -0.03460442975040793
	pesos_i(5257) := b"1111111111111111_1111111111111111_1101001001111100_0001011010111011"; -- -0.17779405539877866
	pesos_i(5258) := b"0000000000000000_0000000000000000_0001110011001010_0110011000010010"; -- 0.11246335917090748
	pesos_i(5259) := b"0000000000000000_0000000000000000_0010100101000101_0100000111000001"; -- 0.16121302569625093
	pesos_i(5260) := b"0000000000000000_0000000000000000_0000001101110001_0110000010000111"; -- 0.013448746589639748
	pesos_i(5261) := b"0000000000000000_0000000000000000_0001111010110000_1111101011111000"; -- 0.11988800569377167
	pesos_i(5262) := b"1111111111111111_1111111111111111_1110000010000111_1001100111100001"; -- -0.12293089152645406
	pesos_i(5263) := b"1111111111111111_1111111111111111_1111011011101111_1110100011111101"; -- -0.035401762338191256
	pesos_i(5264) := b"1111111111111111_1111111111111111_1110000001110110_0100111010000001"; -- -0.12319478372466383
	pesos_i(5265) := b"1111111111111111_1111111111111111_1101010010010110_0110101111111100"; -- -0.16957974532631193
	pesos_i(5266) := b"0000000000000000_0000000000000000_0000011100111010_1001100101100000"; -- 0.028237901740637332
	pesos_i(5267) := b"0000000000000000_0000000000000000_0001101000110000_1011111011010011"; -- 0.10230629594347239
	pesos_i(5268) := b"1111111111111111_1111111111111111_1111001000011111_1111011001101111"; -- -0.05419978887055589
	pesos_i(5269) := b"0000000000000000_0000000000000000_0000110001000011_0000001001001111"; -- 0.04789747654166372
	pesos_i(5270) := b"1111111111111111_1111111111111111_1110011100000110_0000100100110100"; -- -0.09756414872621043
	pesos_i(5271) := b"1111111111111111_1111111111111111_1111111000101111_1100011001010000"; -- -0.007083516503837838
	pesos_i(5272) := b"0000000000000000_0000000000000000_0001001111101110_0110001100101111"; -- 0.07785625366985847
	pesos_i(5273) := b"1111111111111111_1111111111111111_1110100110001001_0001001001001010"; -- -0.08775220569935425
	pesos_i(5274) := b"1111111111111111_1111111111111111_1101110010100100_1101010100000111"; -- -0.1381098611078783
	pesos_i(5275) := b"0000000000000000_0000000000000000_0000001000011100_1010101001101110"; -- 0.008249904462912178
	pesos_i(5276) := b"0000000000000000_0000000000000000_0001101111101001_1011011001111101"; -- 0.10903492493922341
	pesos_i(5277) := b"0000000000000000_0000000000000000_0001010001000011_0011000101000101"; -- 0.07915027544376207
	pesos_i(5278) := b"0000000000000000_0000000000000000_0001000010010001_1101101000000001"; -- 0.06472551838298224
	pesos_i(5279) := b"0000000000000000_0000000000000000_0001000010111010_0100101010000000"; -- 0.06534257527326187
	pesos_i(5280) := b"0000000000000000_0000000000000000_0001001101101111_1011001011101010"; -- 0.07592313970854905
	pesos_i(5281) := b"1111111111111111_1111111111111111_1110111000111110_0001000101101110"; -- -0.06936541622763065
	pesos_i(5282) := b"0000000000000000_0000000000000000_0010011001110100_0111110001111010"; -- 0.15021493888374926
	pesos_i(5283) := b"1111111111111111_1111111111111111_1101101011110111_0000111000010000"; -- -0.14466774081843645
	pesos_i(5284) := b"1111111111111111_1111111111111111_1110110101110011_0011111111100010"; -- -0.07246018162506619
	pesos_i(5285) := b"1111111111111111_1111111111111111_1111101110001100_1101111110011001"; -- -0.017381692050495525
	pesos_i(5286) := b"0000000000000000_0000000000000000_0001101100010100_0101110100111000"; -- 0.10577948202368585
	pesos_i(5287) := b"1111111111111111_1111111111111111_1111111101010111_1101100011001011"; -- -0.0025658135111493174
	pesos_i(5288) := b"0000000000000000_0000000000000000_0001110110001011_0101001001101111"; -- 0.11540713513316272
	pesos_i(5289) := b"0000000000000000_0000000000000000_0010010100010010_1110110000110110"; -- 0.14481998746375918
	pesos_i(5290) := b"0000000000000000_0000000000000000_0010100101111001_0010011101101110"; -- 0.16200491361720484
	pesos_i(5291) := b"1111111111111111_1111111111111111_1110111101010100_1001100010111111"; -- -0.06511540727347156
	pesos_i(5292) := b"0000000000000000_0000000000000000_0000101010110010_1010011111010010"; -- 0.04178856739421659
	pesos_i(5293) := b"0000000000000000_0000000000000000_0010100011011110_1000000010101000"; -- 0.15964511959895833
	pesos_i(5294) := b"0000000000000000_0000000000000000_0010100100010110_0110100011110010"; -- 0.16049819856834122
	pesos_i(5295) := b"1111111111111111_1111111111111111_1101011000000110_1100010010110001"; -- -0.16395922353444498
	pesos_i(5296) := b"1111111111111111_1111111111111111_1111010010010101_1101110100010100"; -- -0.044588263071336454
	pesos_i(5297) := b"1111111111111111_1111111111111111_1110111100110101_1000101101010100"; -- -0.06558922952126815
	pesos_i(5298) := b"0000000000000000_0000000000000000_0000000100011011_0101110110101101"; -- 0.0043238207072276045
	pesos_i(5299) := b"1111111111111111_1111111111111111_1101001110000001_0111001010111011"; -- -0.1738060276830632
	pesos_i(5300) := b"0000000000000000_0000000000000000_0010000101000001_1110000000010000"; -- 0.12991142634578773
	pesos_i(5301) := b"1111111111111111_1111111111111111_1111110101110111_0000011010010011"; -- -0.009902562149287811
	pesos_i(5302) := b"0000000000000000_0000000000000000_0000111001100101_1000000011110110"; -- 0.05623632437101854
	pesos_i(5303) := b"0000000000000000_0000000000000000_0010010111001010_1001110100100010"; -- 0.1476228912821513
	pesos_i(5304) := b"0000000000000000_0000000000000000_0010110001000010_0000010101110010"; -- 0.1728824045760148
	pesos_i(5305) := b"0000000000000000_0000000000000000_0000101101111011_1100101110100011"; -- 0.04485771876827072
	pesos_i(5306) := b"0000000000000000_0000000000000000_0010001010110000_1011111110110101"; -- 0.1355094734121756
	pesos_i(5307) := b"0000000000000000_0000000000000000_0000011100010000_1011101101100000"; -- 0.027599059077750777
	pesos_i(5308) := b"1111111111111111_1111111111111111_1101011010111110_0100010011110001"; -- -0.16115922085543238
	pesos_i(5309) := b"1111111111111111_1111111111111111_1111110000111001_1100010001011110"; -- -0.014743544735140916
	pesos_i(5310) := b"0000000000000000_0000000000000000_0001001101000010_0001010101001000"; -- 0.0752270985756302
	pesos_i(5311) := b"1111111111111111_1111111111111111_1101001010101110_0001000010110011"; -- -0.17703147530762514
	pesos_i(5312) := b"1111111111111111_1111111111111111_1111001011111111_1000100111111001"; -- -0.05078828506691932
	pesos_i(5313) := b"1111111111111111_1111111111111111_1111011110001110_1101110110010000"; -- -0.03297629576551657
	pesos_i(5314) := b"0000000000000000_0000000000000000_0000001111111101_1001010000010010"; -- 0.015588049237383867
	pesos_i(5315) := b"0000000000000000_0000000000000000_0000101000100110_0011110001111010"; -- 0.0396459386745397
	pesos_i(5316) := b"0000000000000000_0000000000000000_0001111000010100_0001111000011011"; -- 0.11749447010422855
	pesos_i(5317) := b"0000000000000000_0000000000000000_0001011000110011_0110011110101100"; -- 0.08672187752064885
	pesos_i(5318) := b"0000000000000000_0000000000000000_0000010000101101_1011011101010001"; -- 0.016322571974189893
	pesos_i(5319) := b"1111111111111111_1111111111111111_1101101011101110_1110111101000001"; -- -0.1447916475603359
	pesos_i(5320) := b"0000000000000000_0000000000000000_0010000000011111_1101011011111011"; -- 0.12548583621470694
	pesos_i(5321) := b"0000000000000000_0000000000000000_0001001000110001_0100100101100111"; -- 0.07106455587817234
	pesos_i(5322) := b"0000000000000000_0000000000000000_0001010111111110_1110010100010100"; -- 0.08592063642985238
	pesos_i(5323) := b"1111111111111111_1111111111111111_1110011111011110_0111000100100011"; -- -0.09426205535894383
	pesos_i(5324) := b"0000000000000000_0000000000000000_0001110010010001_1100000000101011"; -- 0.11159897851774692
	pesos_i(5325) := b"1111111111111111_1111111111111111_1101110100001011_1100010100111001"; -- -0.13653914792330052
	pesos_i(5326) := b"1111111111111111_1111111111111111_1101011111011011_0100101101010100"; -- -0.1568100852766493
	pesos_i(5327) := b"0000000000000000_0000000000000000_0000100010111101_0000101001000010"; -- 0.034134522484262506
	pesos_i(5328) := b"1111111111111111_1111111111111111_1101010110111001_1011010000001000"; -- -0.16513514336005614
	pesos_i(5329) := b"0000000000000000_0000000000000000_0001010100101011_0111000101000100"; -- 0.08269412919338932
	pesos_i(5330) := b"0000000000000000_0000000000000000_0000110101110101_1001001010001011"; -- 0.052575262925163166
	pesos_i(5331) := b"1111111111111111_1111111111111111_1111100100110110_0110000011110000"; -- -0.026513997543252024
	pesos_i(5332) := b"0000000000000000_0000000000000000_0001000101101000_0001011001101001"; -- 0.06799449979969449
	pesos_i(5333) := b"1111111111111111_1111111111111111_1101011111100000_1001101001000011"; -- -0.15672908657832757
	pesos_i(5334) := b"1111111111111111_1111111111111111_1111110110010011_1001010111010110"; -- -0.009466777096246918
	pesos_i(5335) := b"1111111111111111_1111111111111111_1101110100100001_0011000110011000"; -- -0.13621225403381418
	pesos_i(5336) := b"1111111111111111_1111111111111111_1111111111100111_1110100101100001"; -- -0.00036755919832653255
	pesos_i(5337) := b"1111111111111111_1111111111111111_1111011001001110_1101111100110001"; -- -0.03785901124579387
	pesos_i(5338) := b"1111111111111111_1111111111111111_1111111010111010_1011000101110111"; -- -0.0049637875108803926
	pesos_i(5339) := b"0000000000000000_0000000000000000_0000011110101111_1011101101000111"; -- 0.030025200574892785
	pesos_i(5340) := b"1111111111111111_1111111111111111_1101110101111000_0000101111000101"; -- -0.13488699375413551
	pesos_i(5341) := b"1111111111111111_1111111111111111_1110110010000001_0101101111101000"; -- -0.07615113824343683
	pesos_i(5342) := b"1111111111111111_1111111111111111_1110111000001010_1001110010001000"; -- -0.07015058210442214
	pesos_i(5343) := b"0000000000000000_0000000000000000_0010000111001010_0110011101100100"; -- 0.13199468791006833
	pesos_i(5344) := b"0000000000000000_0000000000000000_0010110011011100_1111000110110000"; -- 0.1752463391918023
	pesos_i(5345) := b"1111111111111111_1111111111111111_1111110000011000_0000001010100100"; -- -0.015258631776193845
	pesos_i(5346) := b"1111111111111111_1111111111111111_1101010100100111_0010011010000001"; -- -0.16737136229932964
	pesos_i(5347) := b"0000000000000000_0000000000000000_0010000100001011_0000010110100101"; -- 0.12907443303881408
	pesos_i(5348) := b"0000000000000000_0000000000000000_0001111010111000_1110001001001010"; -- 0.12000860515992658
	pesos_i(5349) := b"0000000000000000_0000000000000000_0001100110110110_0000001010101010"; -- 0.100433508353626
	pesos_i(5350) := b"1111111111111111_1111111111111111_1111100001101000_1100011110101101"; -- -0.029651184268501874
	pesos_i(5351) := b"1111111111111111_1111111111111111_1110001101101011_0110110010010011"; -- -0.11164208813285025
	pesos_i(5352) := b"0000000000000000_0000000000000000_0000100111011110_0011001110100100"; -- 0.03854677926870617
	pesos_i(5353) := b"0000000000000000_0000000000000000_0000101101001101_0000100110100000"; -- 0.04414425049378233
	pesos_i(5354) := b"0000000000000000_0000000000000000_0000100110010001_1111101100000010"; -- 0.037383735582669005
	pesos_i(5355) := b"1111111111111111_1111111111111111_1111000101001100_1110011011001001"; -- -0.05742032625627022
	pesos_i(5356) := b"0000000000000000_0000000000000000_0001100010101110_0100010101010011"; -- 0.09640916138206872
	pesos_i(5357) := b"1111111111111111_1111111111111111_1110101101110010_1010010110100111"; -- -0.08028187434508183
	pesos_i(5358) := b"0000000000000000_0000000000000000_0010000110010000_1101010100010000"; -- 0.1311162151333743
	pesos_i(5359) := b"1111111111111111_1111111111111111_1111101101000100_0010011111111100"; -- -0.01849126906728857
	pesos_i(5360) := b"1111111111111111_1111111111111111_1111101000011001_1100110001011101"; -- -0.023043849289285295
	pesos_i(5361) := b"1111111111111111_1111111111111111_1110101111001110_1001010010000000"; -- -0.07887908825191614
	pesos_i(5362) := b"1111111111111111_1111111111111111_1101110001011101_0110111110010111"; -- -0.1391992812802512
	pesos_i(5363) := b"0000000000000000_0000000000000000_0001110010101100_0100101101001001"; -- 0.11200399901747109
	pesos_i(5364) := b"1111111111111111_1111111111111111_1111101100001101_1110011111010110"; -- -0.01931906716217659
	pesos_i(5365) := b"1111111111111111_1111111111111111_1111000010000000_0100100110100001"; -- -0.06054248639877549
	pesos_i(5366) := b"1111111111111111_1111111111111111_1101110011000001_1001101001101010"; -- -0.13767085000850943
	pesos_i(5367) := b"1111111111111111_1111111111111111_1110010100111001_1110010111111001"; -- -0.10458529158734836
	pesos_i(5368) := b"0000000000000000_0000000000000000_0010100110000111_0011001001001001"; -- 0.16221918383037678
	pesos_i(5369) := b"0000000000000000_0000000000000000_0010001100110010_1010000010011011"; -- 0.1374912622361084
	pesos_i(5370) := b"1111111111111111_1111111111111111_1101100110100011_1110100110110101"; -- -0.1498426373015185
	pesos_i(5371) := b"1111111111111111_1111111111111111_1110100000010000_1010001100111101"; -- -0.0934961296846106
	pesos_i(5372) := b"1111111111111111_1111111111111111_1111100011110100_1111010111111110"; -- -0.02751219311186297
	pesos_i(5373) := b"0000000000000000_0000000000000000_0010110100100111_1010111011110110"; -- 0.17638677118948304
	pesos_i(5374) := b"1111111111111111_1111111111111111_1111101010000110_1000100000011111"; -- -0.0213847088567057
	pesos_i(5375) := b"0000000000000000_0000000000000000_0001001101010101_1001010110011000"; -- 0.07552466361593774
	pesos_i(5376) := b"1111111111111111_1111111111111111_1101101110011101_1011011001010010"; -- -0.14212475290227525
	pesos_i(5377) := b"1111111111111111_1111111111111111_1101100001111111_1011000000000101"; -- -0.15430164224535894
	pesos_i(5378) := b"1111111111111111_1111111111111111_1110000001011001_1001011111101101"; -- -0.12363291217677781
	pesos_i(5379) := b"1111111111111111_1111111111111111_1111001001011000_0001111110111010"; -- -0.05334283558621949
	pesos_i(5380) := b"0000000000000000_0000000000000000_0000101001110110_0011001111001001"; -- 0.040866123694904916
	pesos_i(5381) := b"1111111111111111_1111111111111111_1110100110000100_1111001111101011"; -- -0.08781505126486905
	pesos_i(5382) := b"1111111111111111_1111111111111111_1110000001101110_0101111100001111"; -- -0.12331586717433318
	pesos_i(5383) := b"1111111111111111_1111111111111111_1110110111110001_0000010000110001"; -- -0.0705411319892405
	pesos_i(5384) := b"1111111111111111_1111111111111111_1101110000100110_1011111010010111"; -- -0.1400338060142844
	pesos_i(5385) := b"0000000000000000_0000000000000000_0001001110101000_0000011000000101"; -- 0.07678258541280991
	pesos_i(5386) := b"1111111111111111_1111111111111111_1111100101000100_0101010101100111"; -- -0.026301061934373964
	pesos_i(5387) := b"1111111111111111_1111111111111111_1111101010001101_0100111111011110"; -- -0.02128125033085966
	pesos_i(5388) := b"0000000000000000_0000000000000000_0001011111010111_0001110100100001"; -- 0.09312612595041725
	pesos_i(5389) := b"0000000000000000_0000000000000000_0010101011111000_1001010010000110"; -- 0.16785553229613345
	pesos_i(5390) := b"0000000000000000_0000000000000000_0000101011111010_0100010111111111"; -- 0.04288136930342641
	pesos_i(5391) := b"1111111111111111_1111111111111111_1111101111001110_0100010010010110"; -- -0.016383851461953272
	pesos_i(5392) := b"1111111111111111_1111111111111111_1111101101100000_1010011001011101"; -- -0.018056490212173565
	pesos_i(5393) := b"1111111111111111_1111111111111111_1101111010101110_1101011101010010"; -- -0.1301446366647452
	pesos_i(5394) := b"0000000000000000_0000000000000000_0010101101001011_1011100100001110"; -- 0.1691241894119039
	pesos_i(5395) := b"1111111111111111_1111111111111111_1111111101001000_0110111100101111"; -- -0.002800990084991315
	pesos_i(5396) := b"0000000000000000_0000000000000000_0001011000101111_1110100100000101"; -- 0.08666855209824254
	pesos_i(5397) := b"1111111111111111_1111111111111111_1111011110110001_0101100100101010"; -- -0.03245012982232895
	pesos_i(5398) := b"1111111111111111_1111111111111111_1101111100010010_1101101110000101"; -- -0.12861850738370229
	pesos_i(5399) := b"1111111111111111_1111111111111111_1110111110110111_0001110101110110"; -- -0.06361213563993125
	pesos_i(5400) := b"0000000000000000_0000000000000000_0010100111010100_1101010011011100"; -- 0.16340380066505505
	pesos_i(5401) := b"0000000000000000_0000000000000000_0001000000110101_0010100001101010"; -- 0.06331112461507098
	pesos_i(5402) := b"0000000000000000_0000000000000000_0001001101001010_0111100101010111"; -- 0.07535513277024782
	pesos_i(5403) := b"1111111111111111_1111111111111111_1111111101000001_1011001101100011"; -- -0.002903736511472447
	pesos_i(5404) := b"1111111111111111_1111111111111111_1110010100100101_1110111011100001"; -- -0.1048899364333486
	pesos_i(5405) := b"0000000000000000_0000000000000000_0001010001101011_1111011101011110"; -- 0.07977243477423318
	pesos_i(5406) := b"1111111111111111_1111111111111111_1110010101010000_1111101110001010"; -- -0.10423305404031183
	pesos_i(5407) := b"1111111111111111_1111111111111111_1110110010110011_1011000110011001"; -- -0.07538309116978753
	pesos_i(5408) := b"0000000000000000_0000000000000000_0000011100011010_1101101000001000"; -- 0.027753474276929258
	pesos_i(5409) := b"1111111111111111_1111111111111111_1101010010010011_1010111100111001"; -- -0.16962151385613938
	pesos_i(5410) := b"0000000000000000_0000000000000000_0001010010011101_1111000111001001"; -- 0.08053504144252308
	pesos_i(5411) := b"0000000000000000_0000000000000000_0010100000111010_1111010111011111"; -- 0.1571496648455394
	pesos_i(5412) := b"1111111111111111_1111111111111111_1110101111010010_1010100000101011"; -- -0.07881688064843685
	pesos_i(5413) := b"0000000000000000_0000000000000000_0010101100100011_0100011101010011"; -- 0.1685070589111863
	pesos_i(5414) := b"0000000000000000_0000000000000000_0000110111011001_0001101000100101"; -- 0.05409396552630052
	pesos_i(5415) := b"1111111111111111_1111111111111111_1111010110101000_0100011011011110"; -- -0.040401049322970256
	pesos_i(5416) := b"1111111111111111_1111111111111111_1101110010111111_1001010011110001"; -- -0.13770169360256806
	pesos_i(5417) := b"1111111111111111_1111111111111111_1111110001011111_0010011000000011"; -- -0.01417314940175917
	pesos_i(5418) := b"1111111111111111_1111111111111111_1101101111100001_1101011001101000"; -- -0.1410852428484733
	pesos_i(5419) := b"1111111111111111_1111111111111111_1101011011110011_0110100011010110"; -- -0.1603483655443281
	pesos_i(5420) := b"1111111111111111_1111111111111111_1110011011111000_0000011000000101"; -- -0.09777796149890401
	pesos_i(5421) := b"1111111111111111_1111111111111111_1101110010010011_1001010111010000"; -- -0.13837302844150745
	pesos_i(5422) := b"0000000000000000_0000000000000000_0001010010001000_0001110101001110"; -- 0.08020194201020245
	pesos_i(5423) := b"1111111111111111_1111111111111111_1110101000110011_0110010100111110"; -- -0.08515326728232915
	pesos_i(5424) := b"0000000000000000_0000000000000000_0001001001000010_0100001110101001"; -- 0.07132361296051679
	pesos_i(5425) := b"0000000000000000_0000000000000000_0000011011001000_0101101001111001"; -- 0.02649465034073532
	pesos_i(5426) := b"1111111111111111_1111111111111111_1101110000000101_0001000110000100"; -- -0.14054766214452202
	pesos_i(5427) := b"1111111111111111_1111111111111111_1111111011110010_1000000011111101"; -- -0.004112184829743318
	pesos_i(5428) := b"0000000000000000_0000000000000000_0010011011001111_0011101100010101"; -- 0.15159959086941813
	pesos_i(5429) := b"1111111111111111_1111111111111111_1111001111010011_0110000011100100"; -- -0.04755587044152751
	pesos_i(5430) := b"0000000000000000_0000000000000000_0010000000001011_1010100101011010"; -- 0.12517794076330369
	pesos_i(5431) := b"0000000000000000_0000000000000000_0010100011110001_0101011011001101"; -- 0.15993254195072837
	pesos_i(5432) := b"0000000000000000_0000000000000000_0000111111010011_0000111010001000"; -- 0.06181422061154351
	pesos_i(5433) := b"0000000000000000_0000000000000000_0001110000011010_1110110010011000"; -- 0.10978583059011617
	pesos_i(5434) := b"0000000000000000_0000000000000000_0001000000111101_1110010011000011"; -- 0.06344442139797056
	pesos_i(5435) := b"1111111111111111_1111111111111111_1110111100101100_0010000100110001"; -- -0.06573288483084808
	pesos_i(5436) := b"1111111111111111_1111111111111111_1110010101000000_0010000000111111"; -- -0.10449026558453771
	pesos_i(5437) := b"1111111111111111_1111111111111111_1111111111100001_0101100010101000"; -- -0.000467738178279136
	pesos_i(5438) := b"0000000000000000_0000000000000000_0000010111111110_1000010101001011"; -- 0.02341492730669369
	pesos_i(5439) := b"1111111111111111_1111111111111111_1110100011011011_0000100100100000"; -- -0.09040778139454672
	pesos_i(5440) := b"1111111111111111_1111111111111111_1110101101100001_0011000110011101"; -- -0.08054819037826869
	pesos_i(5441) := b"1111111111111111_1111111111111111_1100110111000001_1110111010101001"; -- -0.19625957852618692
	pesos_i(5442) := b"0000000000000000_0000000000000000_0001100000011100_1010010000111011"; -- 0.09418703497424546
	pesos_i(5443) := b"1111111111111111_1111111111111111_1111001011101110_0110111001001010"; -- -0.05104933450666112
	pesos_i(5444) := b"0000000000000000_0000000000000000_0010000101011000_0110110011010110"; -- 0.1302555104840577
	pesos_i(5445) := b"1111111111111111_1111111111111111_1111001011001100_1110001111100111"; -- -0.051561123046291624
	pesos_i(5446) := b"0000000000000000_0000000000000000_0000011001110101_0101000110011111"; -- 0.025227643396417296
	pesos_i(5447) := b"0000000000000000_0000000000000000_0001001000100001_1001001011010111"; -- 0.07082479241776768
	pesos_i(5448) := b"1111111111111111_1111111111111111_1111011111000111_1101011101011101"; -- -0.03210691421220922
	pesos_i(5449) := b"1111111111111111_1111111111111111_1101001110110111_0100000101111010"; -- -0.17298498894628303
	pesos_i(5450) := b"0000000000000000_0000000000000000_0000111011110000_1111111111011100"; -- 0.058364859688673804
	pesos_i(5451) := b"0000000000000000_0000000000000000_0000010000101101_1110100100101111"; -- 0.016325544383922672
	pesos_i(5452) := b"0000000000000000_0000000000000000_0000000010010101_0010111111011000"; -- 0.002276411215765351
	pesos_i(5453) := b"1111111111111111_1111111111111111_1101010000001001_0010101011010100"; -- -0.17173511824144666
	pesos_i(5454) := b"0000000000000000_0000000000000000_0001001010101001_1011001001000100"; -- 0.0729018607201038
	pesos_i(5455) := b"1111111111111111_1111111111111111_1110011000010100_1100110101010001"; -- -0.10124508629913063
	pesos_i(5456) := b"0000000000000000_0000000000000000_0010100110011110_1100000001000000"; -- 0.16257859763173108
	pesos_i(5457) := b"0000000000000000_0000000000000000_0001111101100111_0100001100100011"; -- 0.1226694068257736
	pesos_i(5458) := b"1111111111111111_1111111111111111_1110101011110010_1111011001001000"; -- -0.08223019361494734
	pesos_i(5459) := b"1111111111111111_1111111111111111_1110011000011101_1011111100000010"; -- -0.10110861005266708
	pesos_i(5460) := b"0000000000000000_0000000000000000_0000010101110110_0101010100101111"; -- 0.021336864394555243
	pesos_i(5461) := b"1111111111111111_1111111111111111_1110010101101011_1111001001000000"; -- -0.10382162045602662
	pesos_i(5462) := b"1111111111111111_1111111111111111_1101100011110101_1011011000110100"; -- -0.15250073650941337
	pesos_i(5463) := b"1111111111111111_1111111111111111_1110000101000000_1011101110011111"; -- -0.12010600439758623
	pesos_i(5464) := b"1111111111111111_1111111111111111_1111000100100000_1001000111000111"; -- -0.05809677968246934
	pesos_i(5465) := b"0000000000000000_0000000000000000_0010010110011000_1101110111011011"; -- 0.14686380962752288
	pesos_i(5466) := b"0000000000000000_0000000000000000_0010001110000011_1100010101011011"; -- 0.13872941457169408
	pesos_i(5467) := b"0000000000000000_0000000000000000_0000101101111110_1111000110010101"; -- 0.04490575692395343
	pesos_i(5468) := b"0000000000000000_0000000000000000_0000000101101100_1101001100101100"; -- 0.005566786092894556
	pesos_i(5469) := b"1111111111111111_1111111111111111_1111100110101110_1100011011010001"; -- -0.02467687023651174
	pesos_i(5470) := b"1111111111111111_1111111111111111_1111110001111111_1000011111001110"; -- -0.013679039246133312
	pesos_i(5471) := b"1111111111111111_1111111111111111_1101100100001001_1110000110111100"; -- -0.15219296612695699
	pesos_i(5472) := b"0000000000000000_0000000000000000_0010010001011000_1001011100000110"; -- 0.14197677513090376
	pesos_i(5473) := b"1111111111111111_1111111111111111_1111000010010111_0010100000110000"; -- -0.06019352749533084
	pesos_i(5474) := b"1111111111111111_1111111111111111_1101001110110100_1100101101010100"; -- -0.17302254867023384
	pesos_i(5475) := b"0000000000000000_0000000000000000_0001000100101001_0101101000001111"; -- 0.06703722822757702
	pesos_i(5476) := b"0000000000000000_0000000000000000_0001111101100010_1100100000100111"; -- 0.12260104140118977
	pesos_i(5477) := b"0000000000000000_0000000000000000_0000111011001111_0000100000111111"; -- 0.057846560906943574
	pesos_i(5478) := b"0000000000000000_0000000000000000_0011010100010001_0111010010000101"; -- 0.20729759461476321
	pesos_i(5479) := b"0000000000000000_0000000000000000_0001010000010011_1001100111011000"; -- 0.07842408682847876
	pesos_i(5480) := b"0000000000000000_0000000000000000_0000101010110001_0011000110101000"; -- 0.04176626531538752
	pesos_i(5481) := b"1111111111111111_1111111111111111_1110110110100000_1010010110010001"; -- -0.07176747525299407
	pesos_i(5482) := b"1111111111111111_1111111111111111_1110010010110001_0110000101001000"; -- -0.10666839584237385
	pesos_i(5483) := b"1111111111111111_1111111111111111_1110100000101101_1000011010111001"; -- -0.09305532440789246
	pesos_i(5484) := b"0000000000000000_0000000000000000_0001000100000010_1011101100000100"; -- 0.06644791461596462
	pesos_i(5485) := b"1111111111111111_1111111111111111_1110111110101011_1100011101011100"; -- -0.0637851142195256
	pesos_i(5486) := b"0000000000000000_0000000000000000_0001101000000101_0111110100001001"; -- 0.10164624666005552
	pesos_i(5487) := b"0000000000000000_0000000000000000_0001010000100111_0010100110111111"; -- 0.07872258098728857
	pesos_i(5488) := b"1111111111111111_1111111111111111_1101110011001101_0111001100011010"; -- -0.13749008776031862
	pesos_i(5489) := b"1111111111111111_1111111111111111_1110110100100010_0011001110000011"; -- -0.07369688079451522
	pesos_i(5490) := b"0000000000000000_0000000000000000_0001111001110011_0011011000001100"; -- 0.11894548212564958
	pesos_i(5491) := b"0000000000000000_0000000000000000_0001100110001111_1011100001101010"; -- 0.09984924867528046
	pesos_i(5492) := b"1111111111111111_1111111111111111_1111110100101011_1001010111001110"; -- -0.011053693068793282
	pesos_i(5493) := b"0000000000000000_0000000000000000_0001001000011110_0110001001001110"; -- 0.07077612319946447
	pesos_i(5494) := b"1111111111111111_1111111111111111_1110011110101011_1010110100111011"; -- -0.09503667168892788
	pesos_i(5495) := b"0000000000000000_0000000000000000_0010010010011111_1001110010101110"; -- 0.1430604863818862
	pesos_i(5496) := b"0000000000000000_0000000000000000_0010001110010100_1010010001000101"; -- 0.13898684197842673
	pesos_i(5497) := b"1111111111111111_1111111111111111_1101011111010001_0010110000110000"; -- -0.15696452919486428
	pesos_i(5498) := b"1111111111111111_1111111111111111_1111110001011111_0100011100011101"; -- -0.014171176241711422
	pesos_i(5499) := b"1111111111111111_1111111111111111_1101100100000101_1100010111011110"; -- -0.15225566215427
	pesos_i(5500) := b"0000000000000000_0000000000000000_0010101001010011_1110010001001101"; -- 0.1653425873816388
	pesos_i(5501) := b"1111111111111111_1111111111111111_1111000101110111_1100001000010111"; -- -0.056766385394898165
	pesos_i(5502) := b"0000000000000000_0000000000000000_0000100010000010_1000010110010011"; -- 0.03324160429481185
	pesos_i(5503) := b"1111111111111111_1111111111111111_1110110011100110_1110001100111000"; -- -0.07460193531619227
	pesos_i(5504) := b"0000000000000000_0000000000000000_0010000011100100_0110100100100110"; -- 0.12848527115437322
	pesos_i(5505) := b"1111111111111111_1111111111111111_1111100011100100_0000001110110011"; -- -0.027770775683809527
	pesos_i(5506) := b"0000000000000000_0000000000000000_0000000011100001_0110001101000110"; -- 0.003439144657185732
	pesos_i(5507) := b"0000000000000000_0000000000000000_0000000110110011_1001000100010101"; -- 0.0066462207938799344
	pesos_i(5508) := b"0000000000000000_0000000000000000_0000000011000110_1011101011001001"; -- 0.0030323735745094844
	pesos_i(5509) := b"1111111111111111_1111111111111111_1101111111101000_0001011010111011"; -- -0.12536485612957024
	pesos_i(5510) := b"0000000000000000_0000000000000000_0000101100100101_1101111111111010"; -- 0.043546675232373294
	pesos_i(5511) := b"1111111111111111_1111111111111111_1110100010111111_1010101100001001"; -- -0.0908253767425241
	pesos_i(5512) := b"0000000000000000_0000000000000000_0010101001110011_0010011101001110"; -- 0.1658196034947194
	pesos_i(5513) := b"0000000000000000_0000000000000000_0000101011110101_0100110101110101"; -- 0.04280552019214016
	pesos_i(5514) := b"1111111111111111_1111111111111111_1101111011100001_0000101010010111"; -- -0.12937864123601714
	pesos_i(5515) := b"1111111111111111_1111111111111111_1111111011000001_1001001011101101"; -- -0.004858796193634968
	pesos_i(5516) := b"1111111111111111_1111111111111111_1110000100101101_0011100001011101"; -- -0.12040374492139828
	pesos_i(5517) := b"1111111111111111_1111111111111111_1110011111101101_1001110101100001"; -- -0.09403053641256552
	pesos_i(5518) := b"1111111111111111_1111111111111111_1111010101100001_0100110101010110"; -- -0.04148403799191816
	pesos_i(5519) := b"1111111111111111_1111111111111111_1110110101000010_1010001101001001"; -- -0.07320193745263964
	pesos_i(5520) := b"1111111111111111_1111111111111111_1110101101001111_1100000100100111"; -- -0.0808142928987536
	pesos_i(5521) := b"0000000000000000_0000000000000000_0000111000110100_1101010100111110"; -- 0.0554936673032758
	pesos_i(5522) := b"1111111111111111_1111111111111111_1111010011001010_0000011000001111"; -- -0.04379236357461334
	pesos_i(5523) := b"1111111111111111_1111111111111111_1101100101101101_0001101000000110"; -- -0.15067899087977585
	pesos_i(5524) := b"0000000000000000_0000000000000000_0001000111010011_1101101111101001"; -- 0.06963896206426257
	pesos_i(5525) := b"1111111111111111_1111111111111111_1111000011010111_0110011011110110"; -- -0.05921322347167913
	pesos_i(5526) := b"0000000000000000_0000000000000000_0000001011101111_0111110010000010"; -- 0.01146677188870039
	pesos_i(5527) := b"1111111111111111_1111111111111111_1111111011110100_1011110001001001"; -- -0.004078132823795441
	pesos_i(5528) := b"0000000000000000_0000000000000000_0000110110101011_0010010010000110"; -- 0.053392679877922275
	pesos_i(5529) := b"1111111111111111_1111111111111111_1110110111101111_1100111001110100"; -- -0.07055959380141044
	pesos_i(5530) := b"1111111111111111_1111111111111111_1111101101011010_0001011100111011"; -- -0.018156574377723236
	pesos_i(5531) := b"0000000000000000_0000000000000000_0010100011000001_0100010100010101"; -- 0.15919906399461442
	pesos_i(5532) := b"0000000000000000_0000000000000000_0010111100011011_1010101010010101"; -- 0.18401590478299346
	pesos_i(5533) := b"1111111111111111_1111111111111111_1111011100010101_1111100011101100"; -- -0.03482097848040615
	pesos_i(5534) := b"0000000000000000_0000000000000000_0010110100110001_1101001000100110"; -- 0.17654145657850867
	pesos_i(5535) := b"1111111111111111_1111111111111111_1110101001100111_0001011110011111"; -- -0.08436443689146207
	pesos_i(5536) := b"1111111111111111_1111111111111111_1111000011011010_0111100111000110"; -- -0.05916632577561269
	pesos_i(5537) := b"1111111111111111_1111111111111111_1110010011111111_0010110101100000"; -- -0.1054813043174051
	pesos_i(5538) := b"1111111111111111_1111111111111111_1110001010011001_0010001011000000"; -- -0.1148508340153533
	pesos_i(5539) := b"1111111111111111_1111111111111111_1110100111000110_1001110110000110"; -- -0.08681312073852514
	pesos_i(5540) := b"0000000000000000_0000000000000000_0000111000010010_1001010011110001"; -- 0.05497103591813975
	pesos_i(5541) := b"1111111111111111_1111111111111111_1101011000001110_0111111101100100"; -- -0.16384128377597634
	pesos_i(5542) := b"0000000000000000_0000000000000000_0010111000110100_1010011000111111"; -- 0.18049086598072347
	pesos_i(5543) := b"1111111111111111_1111111111111111_1101010100001000_1001001100000011"; -- -0.16783791714483196
	pesos_i(5544) := b"0000000000000000_0000000000000000_0000111110111011_1010011010101001"; -- 0.061457077389603515
	pesos_i(5545) := b"0000000000000000_0000000000000000_0000001010011011_0011111100001001"; -- 0.010181369518718017
	pesos_i(5546) := b"1111111111111111_1111111111111111_1101110100010000_1001011100001000"; -- -0.13646560709556496
	pesos_i(5547) := b"0000000000000000_0000000000000000_0001001010101111_1000001100010101"; -- 0.07299060110077914
	pesos_i(5548) := b"1111111111111111_1111111111111111_1101101101100010_1101110111100110"; -- -0.14302266242988218
	pesos_i(5549) := b"0000000000000000_0000000000000000_0010001011000100_1110101010110011"; -- 0.13581721172689082
	pesos_i(5550) := b"0000000000000000_0000000000000000_0001010010001001_1011011000100000"; -- 0.08022630969362356
	pesos_i(5551) := b"1111111111111111_1111111111111111_1111010111001100_1100001011100111"; -- -0.0398443398709681
	pesos_i(5552) := b"1111111111111111_1111111111111111_1101101001001011_1111011011110100"; -- -0.14727837137137956
	pesos_i(5553) := b"0000000000000000_0000000000000000_0000100101101101_0111111011100010"; -- 0.03682702085795843
	pesos_i(5554) := b"1111111111111111_1111111111111111_1111011101011111_1110011101000010"; -- -0.033692880885154326
	pesos_i(5555) := b"0000000000000000_0000000000000000_0000010110001111_0101000001011010"; -- 0.021718046243650195
	pesos_i(5556) := b"1111111111111111_1111111111111111_1110110011010100_0011101100100111"; -- -0.07488661089164979
	pesos_i(5557) := b"1111111111111111_1111111111111111_1110101100100110_0011100000011110"; -- -0.08144807108557783
	pesos_i(5558) := b"0000000000000000_0000000000000000_0010000110010011_0110100010011111"; -- 0.1311555279925623
	pesos_i(5559) := b"1111111111111111_1111111111111111_1110110000011111_0110110000010011"; -- -0.07764553592946077
	pesos_i(5560) := b"0000000000000000_0000000000000000_0001011011110110_0001101011100110"; -- 0.08969276531604234
	pesos_i(5561) := b"0000000000000000_0000000000000000_0001100100001000_0010100110111110"; -- 0.09778080829758605
	pesos_i(5562) := b"0000000000000000_0000000000000000_0000111000111111_1001001100101010"; -- 0.05565757526417412
	pesos_i(5563) := b"1111111111111111_1111111111111111_1111011101011110_0011010000110111"; -- -0.03371881156303326
	pesos_i(5564) := b"0000000000000000_0000000000000000_0010001100110001_0100100101000001"; -- 0.1374707969596922
	pesos_i(5565) := b"0000000000000000_0000000000000000_0010101010010101_0010000011111110"; -- 0.16633802598331018
	pesos_i(5566) := b"0000000000000000_0000000000000000_0010100100110111_0000101000001001"; -- 0.16099608151246975
	pesos_i(5567) := b"1111111111111111_1111111111111111_1111001101110001_0001111111100111"; -- -0.04905510521950557
	pesos_i(5568) := b"0000000000000000_0000000000000000_0000110111010111_0100001011001100"; -- 0.054065871023511375
	pesos_i(5569) := b"1111111111111111_1111111111111111_1110100111011000_0100001111010011"; -- -0.08654380903497771
	pesos_i(5570) := b"1111111111111111_1111111111111111_1111111010101111_1010000100000010"; -- -0.005132615173229338
	pesos_i(5571) := b"1111111111111111_1111111111111111_1110000110110001_1010000111010000"; -- -0.11838329952387994
	pesos_i(5572) := b"0000000000000000_0000000000000000_0001011101010110_1111100110100001"; -- 0.09117088501321113
	pesos_i(5573) := b"0000000000000000_0000000000000000_0010011010101000_1100000100000001"; -- 0.15101248052044364
	pesos_i(5574) := b"0000000000000000_0000000000000000_0001011010000110_1010011111010010"; -- 0.08799218059209415
	pesos_i(5575) := b"0000000000000000_0000000000000000_0001111000100000_1100101000000111"; -- 0.11768782300252055
	pesos_i(5576) := b"0000000000000000_0000000000000000_0010111101110011_0000111000101111"; -- 0.18534935606195374
	pesos_i(5577) := b"0000000000000000_0000000000000000_0000011100001111_0011100101010101"; -- 0.02757604898805175
	pesos_i(5578) := b"0000000000000000_0000000000000000_0010001100001001_1010000011001011"; -- 0.13686566301938233
	pesos_i(5579) := b"0000000000000000_0000000000000000_0001110111111000_1010101110111010"; -- 0.11707566540481101
	pesos_i(5580) := b"0000000000000000_0000000000000000_0010011111101111_1000101111101011"; -- 0.1559989403024691
	pesos_i(5581) := b"0000000000000000_0000000000000000_0000001000111011_1111101111101010"; -- 0.008727783802371821
	pesos_i(5582) := b"1111111111111111_1111111111111111_1110010010110100_0011000111101010"; -- -0.1066254429642209
	pesos_i(5583) := b"0000000000000000_0000000000000000_0001000001011111_1010010110000110"; -- 0.06395945086676333
	pesos_i(5584) := b"0000000000000000_0000000000000000_0000011110111001_0100110010110111"; -- 0.030171198651513714
	pesos_i(5585) := b"1111111111111111_1111111111111111_1101100100101111_1000110111010011"; -- -0.1516181336460616
	pesos_i(5586) := b"0000000000000000_0000000000000000_0000011111110110_0110001111011000"; -- 0.03110336333717084
	pesos_i(5587) := b"0000000000000000_0000000000000000_0001001111001001_1110101101011001"; -- 0.07729979437755936
	pesos_i(5588) := b"0000000000000000_0000000000000000_0001000000111011_0101011011001011"; -- 0.06340544178509067
	pesos_i(5589) := b"1111111111111111_1111111111111111_1101011000000000_1000001110010010"; -- -0.16405465775623929
	pesos_i(5590) := b"1111111111111111_1111111111111111_1110001001000101_1111101000001001"; -- -0.11611974018396218
	pesos_i(5591) := b"1111111111111111_1111111111111111_1110000000101001_1111010100110111"; -- -0.12435977376462728
	pesos_i(5592) := b"0000000000000000_0000000000000000_0010010000000000_1110010001010111"; -- 0.14063861011048892
	pesos_i(5593) := b"0000000000000000_0000000000000000_0001001111011011_1000100100110111"; -- 0.07756860351716525
	pesos_i(5594) := b"0000000000000000_0000000000000000_0010110000111011_0001010010100110"; -- 0.17277649923504923
	pesos_i(5595) := b"0000000000000000_0000000000000000_0010011101010000_0010110101001000"; -- 0.153567152091078
	pesos_i(5596) := b"1111111111111111_1111111111111111_1111001100111110_1101000010011100"; -- -0.04982277103898262
	pesos_i(5597) := b"1111111111111111_1111111111111111_1101000100110101_0101100011010001"; -- -0.182779740295539
	pesos_i(5598) := b"0000000000000000_0000000000000000_0001001010111110_0110010001111111"; -- 0.07321765989858241
	pesos_i(5599) := b"1111111111111111_1111111111111111_1110011101010000_1101111100011111"; -- -0.09642224780133926
	pesos_i(5600) := b"1111111111111111_1111111111111111_1110111000001001_1001110101011111"; -- -0.07016579075881409
	pesos_i(5601) := b"1111111111111111_1111111111111111_1110001001100101_1110000100101010"; -- -0.1156329415925203
	pesos_i(5602) := b"1111111111111111_1111111111111111_1110010011001110_0011101110010000"; -- -0.10622813914732494
	pesos_i(5603) := b"1111111111111111_1111111111111111_1111100110111100_1010010100100111"; -- -0.024465253893624243
	pesos_i(5604) := b"0000000000000000_0000000000000000_0010011100010010_0111100011111100"; -- 0.15262561950194906
	pesos_i(5605) := b"1111111111111111_1111111111111111_1111010001001011_0101000110001010"; -- -0.045725730741415956
	pesos_i(5606) := b"0000000000000000_0000000000000000_0010001111111100_1001010011001001"; -- 0.1405728331211281
	pesos_i(5607) := b"0000000000000000_0000000000000000_0000100010011010_1011100011001111"; -- 0.0336108689552822
	pesos_i(5608) := b"0000000000000000_0000000000000000_0001010010101110_0110000000011111"; -- 0.08078575856597223
	pesos_i(5609) := b"1111111111111111_1111111111111111_1111111101001111_1011110001110000"; -- -0.002689573972327317
	pesos_i(5610) := b"0000000000000000_0000000000000000_0000010100101101_1000010001000101"; -- 0.020225779343710833
	pesos_i(5611) := b"0000000000000000_0000000000000000_0010001100010111_1011011100110111"; -- 0.13708062253732906
	pesos_i(5612) := b"1111111111111111_1111111111111111_1110111110110000_1011100100111100"; -- -0.06370966233516823
	pesos_i(5613) := b"1111111111111111_1111111111111111_1111110000001010_1111010000010101"; -- -0.015457863778073375
	pesos_i(5614) := b"0000000000000000_0000000000000000_0000000010100011_0000100111001011"; -- 0.0024877664345725387
	pesos_i(5615) := b"1111111111111111_1111111111111111_1110000011111100_0011111011101111"; -- -0.12115103410640803
	pesos_i(5616) := b"0000000000000000_0000000000000000_0010110001010000_0010011110000101"; -- 0.17309805857608548
	pesos_i(5617) := b"1111111111111111_1111111111111111_1110010000111011_1100101000010011"; -- -0.1084626868984472
	pesos_i(5618) := b"0000000000000000_0000000000000000_0001011011100010_0110110110110111"; -- 0.08939252583362237
	pesos_i(5619) := b"1111111111111111_1111111111111111_1101010010011010_1000110011100101"; -- -0.16951674851231344
	pesos_i(5620) := b"0000000000000000_0000000000000000_0010100001101111_1001101000110011"; -- 0.15795291659376
	pesos_i(5621) := b"0000000000000000_0000000000000000_0010010111100001_0011101100001000"; -- 0.1479679960492954
	pesos_i(5622) := b"0000000000000000_0000000000000000_0010010011111100_1001000010110011"; -- 0.1444788395479073
	pesos_i(5623) := b"1111111111111111_1111111111111111_1111110010110110_0011011001000011"; -- -0.012844666088604099
	pesos_i(5624) := b"1111111111111111_1111111111111111_1110001101100000_1011101011111000"; -- -0.1118052621324998
	pesos_i(5625) := b"1111111111111111_1111111111111111_1110011110101000_0101110000100100"; -- -0.09508728141626582
	pesos_i(5626) := b"1111111111111111_1111111111111111_1110110110100001_1110010101111000"; -- -0.07174840767242927
	pesos_i(5627) := b"0000000000000000_0000000000000000_0001011111001111_0101000001111010"; -- 0.09300711605594346
	pesos_i(5628) := b"0000000000000000_0000000000000000_0000000000000010_1001010111110100"; -- 3.945546903848899e-05
	pesos_i(5629) := b"1111111111111111_1111111111111111_1111000001110011_1000000100011011"; -- -0.060737543882861005
	pesos_i(5630) := b"0000000000000000_0000000000000000_0000011000110000_0011110111000111"; -- 0.024173604107983755
	pesos_i(5631) := b"1111111111111111_1111111111111111_1110010011111110_0110011011011001"; -- -0.10549313729131893
	pesos_i(5632) := b"1111111111111111_1111111111111111_1111001011110101_0010100100001110"; -- -0.050946649521174225
	pesos_i(5633) := b"1111111111111111_1111111111111111_1110001010011010_1001001010100001"; -- -0.11482890666803762
	pesos_i(5634) := b"0000000000000000_0000000000000000_0001001101100110_1011010000001000"; -- 0.0757858771689014
	pesos_i(5635) := b"1111111111111111_1111111111111111_1111011110001000_0011101011001000"; -- -0.03307755101195456
	pesos_i(5636) := b"0000000000000000_0000000000000000_0000111100000001_0010010010001011"; -- 0.058611186999586014
	pesos_i(5637) := b"0000000000000000_0000000000000000_0001001010001011_0111011011000000"; -- 0.07244054977635174
	pesos_i(5638) := b"1111111111111111_1111111111111111_1110000101000111_1100100001011111"; -- -0.11999843297525703
	pesos_i(5639) := b"0000000000000000_0000000000000000_0000110110011010_1110010110001110"; -- 0.053144786063522964
	pesos_i(5640) := b"0000000000000000_0000000000000000_0000100001000000_0111101010101110"; -- 0.032233874892186834
	pesos_i(5641) := b"0000000000000000_0000000000000000_0000001111010001_0111000011111011"; -- 0.01491457114494258
	pesos_i(5642) := b"1111111111111111_1111111111111111_1110010101100001_1001001100001110"; -- -0.10397988225635581
	pesos_i(5643) := b"0000000000000000_0000000000000000_0000101011110101_0011101010110100"; -- 0.04280440240250833
	pesos_i(5644) := b"0000000000000000_0000000000000000_0010000010000100_1101100001100010"; -- 0.12702705747088947
	pesos_i(5645) := b"1111111111111111_1111111111111111_1101010110101000_0001110101111101"; -- -0.16540351581410032
	pesos_i(5646) := b"1111111111111111_1111111111111111_1110100100101100_0010110100000111"; -- -0.0891696795464329
	pesos_i(5647) := b"0000000000000000_0000000000000000_0001010100111111_0111001001011111"; -- 0.08299937071589604
	pesos_i(5648) := b"1111111111111111_1111111111111111_1110010110010010_0101001111110011"; -- -0.10323596308541237
	pesos_i(5649) := b"0000000000000000_0000000000000000_0010001010011110_1111000111111100"; -- 0.13523781201424728
	pesos_i(5650) := b"1111111111111111_1111111111111111_1111111101111100_1011011011001001"; -- -0.0020032653779124875
	pesos_i(5651) := b"1111111111111111_1111111111111111_1101001111000111_0110100011111001"; -- -0.17273849418705278
	pesos_i(5652) := b"0000000000000000_0000000000000000_0000110101110100_1001010010011111"; -- 0.05256012811190706
	pesos_i(5653) := b"0000000000000000_0000000000000000_0010100111100010_1000100001101010"; -- 0.1636128672973416
	pesos_i(5654) := b"1111111111111111_1111111111111111_1101001110100001_0110101100001010"; -- -0.17331820495910766
	pesos_i(5655) := b"1111111111111111_1111111111111111_1111001010011101_1001111100111000"; -- -0.052282379972713997
	pesos_i(5656) := b"0000000000000000_0000000000000000_0010011001101111_1100100011101010"; -- 0.15014320101826323
	pesos_i(5657) := b"1111111111111111_1111111111111111_1110000010010101_0111001001100101"; -- -0.12271962194691895
	pesos_i(5658) := b"1111111111111111_1111111111111111_1110111010101010_1101100011101010"; -- -0.06770557677125538
	pesos_i(5659) := b"0000000000000000_0000000000000000_0000011100111001_0100011101101111"; -- 0.028217758790365033
	pesos_i(5660) := b"1111111111111111_1111111111111111_1111100111010100_1101011001000000"; -- -0.024096116405184113
	pesos_i(5661) := b"1111111111111111_1111111111111111_1110000100100101_0101010000100000"; -- -0.12052416046772003
	pesos_i(5662) := b"0000000000000000_0000000000000000_0000111111101101_1101011000011100"; -- 0.06222284495876643
	pesos_i(5663) := b"0000000000000000_0000000000000000_0010001000100000_0011110100001111"; -- 0.13330442072818013
	pesos_i(5664) := b"1111111111111111_1111111111111111_1101001111101010_0001000101101101"; -- -0.17220965459986737
	pesos_i(5665) := b"1111111111111111_1111111111111111_1111110110001111_1001001010110100"; -- -0.009527998947994222
	pesos_i(5666) := b"0000000000000000_0000000000000000_0000111000011000_1101010100001111"; -- 0.055066410259439515
	pesos_i(5667) := b"1111111111111111_1111111111111111_1101111011100100_0101011011111001"; -- -0.12932831220758453
	pesos_i(5668) := b"0000000000000000_0000000000000000_0000000000110110_0110010001000010"; -- 0.0008299503361966685
	pesos_i(5669) := b"1111111111111111_1111111111111111_1111100001110000_1111111010111001"; -- -0.02952583302179016
	pesos_i(5670) := b"1111111111111111_1111111111111111_1110011011101111_1010010000100011"; -- -0.09790586609145728
	pesos_i(5671) := b"1111111111111111_1111111111111111_1101101110101000_0010001011001010"; -- -0.1419656999640192
	pesos_i(5672) := b"0000000000000000_0000000000000000_0000000111011000_0010011110111100"; -- 0.007204516821328444
	pesos_i(5673) := b"1111111111111111_1111111111111111_1110100011001101_1011000010010100"; -- -0.09061142345722671
	pesos_i(5674) := b"1111111111111111_1111111111111111_1110000001110010_0100011110111100"; -- -0.12325622236643434
	pesos_i(5675) := b"0000000000000000_0000000000000000_0001101011100000_0010010101011111"; -- 0.10498269628348791
	pesos_i(5676) := b"0000000000000000_0000000000000000_0000111000101111_1000011000111111"; -- 0.055412664793898905
	pesos_i(5677) := b"0000000000000000_0000000000000000_0000000110010101_1000010110010011"; -- 0.0061877712423187925
	pesos_i(5678) := b"0000000000000000_0000000000000000_0001101001101001_0110110000011101"; -- 0.10317111680279208
	pesos_i(5679) := b"0000000000000000_0000000000000000_0010011000011000_1011000011011001"; -- 0.14881425197954729
	pesos_i(5680) := b"0000000000000000_0000000000000000_0001111011101011_1101111000010101"; -- 0.12078655243543393
	pesos_i(5681) := b"1111111111111111_1111111111111111_1110111011110110_0011010001101101"; -- -0.06655571308044184
	pesos_i(5682) := b"0000000000000000_0000000000000000_0010100001000001_0110111001011011"; -- 0.1572483990804516
	pesos_i(5683) := b"0000000000000000_0000000000000000_0010001100100101_1110101110001101"; -- 0.13729736504417994
	pesos_i(5684) := b"1111111111111111_1111111111111111_1111010011010101_0011011110110000"; -- -0.04362155868245974
	pesos_i(5685) := b"0000000000000000_0000000000000000_0001001001111010_1001001010000010"; -- 0.07218280475298744
	pesos_i(5686) := b"0000000000000000_0000000000000000_0000000010101101_0010100110111011"; -- 0.0026422577383732556
	pesos_i(5687) := b"0000000000000000_0000000000000000_0000010011110011_0101001110001011"; -- 0.019337865215201592
	pesos_i(5688) := b"0000000000000000_0000000000000000_0010001001110001_0100011101010011"; -- 0.13454099449868143
	pesos_i(5689) := b"0000000000000000_0000000000000000_0000011001111000_0100101100000110"; -- 0.025273026519623477
	pesos_i(5690) := b"1111111111111111_1111111111111111_1111001101101101_1101000000111000"; -- -0.049105631154997255
	pesos_i(5691) := b"1111111111111111_1111111111111111_1110010001010000_0110111100100100"; -- -0.10814767232955647
	pesos_i(5692) := b"0000000000000000_0000000000000000_0000011011100000_1111101001110111"; -- 0.02687039752669366
	pesos_i(5693) := b"0000000000000000_0000000000000000_0000111111000010_1111101111011100"; -- 0.0615689669602575
	pesos_i(5694) := b"1111111111111111_1111111111111111_1101111000110000_1101001100010001"; -- -0.13206749756956349
	pesos_i(5695) := b"0000000000000000_0000000000000000_0001100101111110_1110001111011110"; -- 0.09959243932388176
	pesos_i(5696) := b"0000000000000000_0000000000000000_0000011100001010_1000001100001101"; -- 0.027504149163825375
	pesos_i(5697) := b"1111111111111111_1111111111111111_1111011000110100_0101101100101111"; -- -0.03826360790983085
	pesos_i(5698) := b"1111111111111111_1111111111111111_1110100101110110_1111010101000100"; -- -0.08802859386692366
	pesos_i(5699) := b"1111111111111111_1111111111111111_1110011100100101_0001010011000011"; -- -0.09709043741323595
	pesos_i(5700) := b"1111111111111111_1111111111111111_1110111001100001_0001111111111000"; -- -0.06883049207147277
	pesos_i(5701) := b"0000000000000000_0000000000000000_0000000000011100_0000010001000011"; -- 0.000427500172597912
	pesos_i(5702) := b"0000000000000000_0000000000000000_0010010101111101_1001000010001010"; -- 0.1464472137536381
	pesos_i(5703) := b"0000000000000000_0000000000000000_0001000101011010_1100001100101001"; -- 0.06779117348113413
	pesos_i(5704) := b"1111111111111111_1111111111111111_1111110100110011_0111101011111110"; -- -0.010933220902222214
	pesos_i(5705) := b"0000000000000000_0000000000000000_0010000111110001_1111000100011111"; -- 0.13259799019093005
	pesos_i(5706) := b"0000000000000000_0000000000000000_0000010101110110_0011111011001111"; -- 0.021335530854371752
	pesos_i(5707) := b"0000000000000000_0000000000000000_0010000011111110_0101010000010101"; -- 0.12888074418473955
	pesos_i(5708) := b"0000000000000000_0000000000000000_0000111001111010_1000111010110100"; -- 0.05655757802386507
	pesos_i(5709) := b"0000000000000000_0000000000000000_0010001011101010_0010000111010110"; -- 0.13638507333506447
	pesos_i(5710) := b"0000000000000000_0000000000000000_0000001011011110_0011011110010011"; -- 0.011203263761290987
	pesos_i(5711) := b"1111111111111111_1111111111111111_1101001000110010_1111101110000100"; -- -0.17890956910244216
	pesos_i(5712) := b"1111111111111111_1111111111111111_1101101000010011_0011001000001000"; -- -0.14814460097476373
	pesos_i(5713) := b"0000000000000000_0000000000000000_0001001001100111_1000111011101101"; -- 0.0718926744053359
	pesos_i(5714) := b"1111111111111111_1111111111111111_1101011101111110_1011111110101011"; -- -0.15822221824564775
	pesos_i(5715) := b"1111111111111111_1111111111111111_1111111101111110_1100101100100010"; -- -0.001971534812513662
	pesos_i(5716) := b"0000000000000000_0000000000000000_0010100111000001_0101011010110110"; -- 0.1631063645756336
	pesos_i(5717) := b"1111111111111111_1111111111111111_1101010111111111_1000001101000000"; -- -0.16406993573601647
	pesos_i(5718) := b"0000000000000000_0000000000000000_0010100100011000_1100001011111000"; -- 0.16053408202547104
	pesos_i(5719) := b"0000000000000000_0000000000000000_0000100101000011_0101001010101101"; -- 0.03618351684350345
	pesos_i(5720) := b"0000000000000000_0000000000000000_0010000010101011_0011110001010101"; -- 0.12761284906368597
	pesos_i(5721) := b"0000000000000000_0000000000000000_0010001110110110_1111000011110011"; -- 0.13951021121637197
	pesos_i(5722) := b"1111111111111111_1111111111111111_1110110011001100_0110010111101101"; -- -0.07500613181270337
	pesos_i(5723) := b"1111111111111111_1111111111111111_1111011100011001_0011000111110000"; -- -0.03477180374782252
	pesos_i(5724) := b"1111111111111111_1111111111111111_1111110011000001_0010000110000100"; -- -0.012678056028164868
	pesos_i(5725) := b"1111111111111111_1111111111111111_1101100000110010_1011011111100110"; -- -0.15547609940734064
	pesos_i(5726) := b"0000000000000000_0000000000000000_0001011001011110_1101100010101110"; -- 0.08738474119129794
	pesos_i(5727) := b"1111111111111111_1111111111111111_1111000010001101_0011100001101010"; -- -0.06034514825356248
	pesos_i(5728) := b"1111111111111111_1111111111111111_1110101010111110_1110000110101001"; -- -0.08302487974876278
	pesos_i(5729) := b"1111111111111111_1111111111111111_1110101111001110_0100011110101000"; -- -0.07888366832756509
	pesos_i(5730) := b"1111111111111111_1111111111111111_1110110011011101_0110100101111111"; -- -0.07474651952272403
	pesos_i(5731) := b"0000000000000000_0000000000000000_0000111101100101_0110001111011010"; -- 0.06014083932057257
	pesos_i(5732) := b"1111111111111111_1111111111111111_1101010100011001_1010111100111101"; -- -0.16757683517312502
	pesos_i(5733) := b"1111111111111111_1111111111111111_1101011110010010_0111001011100011"; -- -0.1579216190272023
	pesos_i(5734) := b"1111111111111111_1111111111111111_1110001000011111_1110101000000110"; -- -0.11670052864837648
	pesos_i(5735) := b"0000000000000000_0000000000000000_0000010100111110_0110111111110100"; -- 0.020483967783676615
	pesos_i(5736) := b"1111111111111111_1111111111111111_1111000111011000_1110110001011101"; -- -0.05528376330954064
	pesos_i(5737) := b"1111111111111111_1111111111111111_1111011001010011_0000101001010000"; -- -0.03779540575105175
	pesos_i(5738) := b"0000000000000000_0000000000000000_0010100010001101_1111110101011010"; -- 0.15841659019366955
	pesos_i(5739) := b"1111111111111111_1111111111111111_1110111111001111_1001001100100110"; -- -0.0632389099727242
	pesos_i(5740) := b"1111111111111111_1111111111111111_1111010001000101_1111111001110000"; -- -0.04580697790455779
	pesos_i(5741) := b"0000000000000000_0000000000000000_0010011110110101_1100101010010100"; -- 0.15511766535583263
	pesos_i(5742) := b"0000000000000000_0000000000000000_0000011101011110_0001011010011010"; -- 0.028779423356076368
	pesos_i(5743) := b"1111111111111111_1111111111111111_1111110010010011_1010000000001111"; -- -0.013372417841966909
	pesos_i(5744) := b"0000000000000000_0000000000000000_0001000110111001_0111101010010110"; -- 0.06923643265849938
	pesos_i(5745) := b"0000000000000000_0000000000000000_0011001010010000_0001011011100001"; -- 0.1975111293501715
	pesos_i(5746) := b"1111111111111111_1111111111111111_1101011101001001_0111001010100100"; -- -0.1590355253687197
	pesos_i(5747) := b"0000000000000000_0000000000000000_0001101001101101_0110110000111000"; -- 0.10323215830869543
	pesos_i(5748) := b"1111111111111111_1111111111111111_1111011011110110_0110001010011001"; -- -0.035302960971624504
	pesos_i(5749) := b"0000000000000000_0000000000000000_0001001001000101_0101000010010000"; -- 0.07137015834561647
	pesos_i(5750) := b"0000000000000000_0000000000000000_0001001000001100_0111100000111001"; -- 0.07050277125550133
	pesos_i(5751) := b"0000000000000000_0000000000000000_0000100100101001_1100110001110100"; -- 0.035794046758680594
	pesos_i(5752) := b"1111111111111111_1111111111111111_1110000010111000_0110001111001101"; -- -0.12218643422923556
	pesos_i(5753) := b"1111111111111111_1111111111111111_1111100101011111_1101111011001110"; -- -0.025880884905983066
	pesos_i(5754) := b"0000000000000000_0000000000000000_0010011111000010_1011110100011111"; -- 0.1553152275512912
	pesos_i(5755) := b"0000000000000000_0000000000000000_0000111111101100_0011000111111110"; -- 0.06219780397991557
	pesos_i(5756) := b"0000000000000000_0000000000000000_0001110111001110_1101010001000010"; -- 0.11643721208509988
	pesos_i(5757) := b"1111111111111111_1111111111111111_1110100101010111_1010100111011011"; -- -0.08850611111832997
	pesos_i(5758) := b"0000000000000000_0000000000000000_0001101100010110_1101100001011110"; -- 0.10581733990245674
	pesos_i(5759) := b"1111111111111111_1111111111111111_1110101000110101_1110001111011010"; -- -0.08511520314307655
	pesos_i(5760) := b"0000000000000000_0000000000000000_0000110011101010_0010000011101000"; -- 0.05044751802202754
	pesos_i(5761) := b"0000000000000000_0000000000000000_0000010010100001_1111000101011100"; -- 0.01809605118378354
	pesos_i(5762) := b"0000000000000000_0000000000000000_0010100101011101_0010001011100011"; -- 0.16157739684463884
	pesos_i(5763) := b"0000000000000000_0000000000000000_0000011110001110_0000000000111011"; -- 0.029510511702350747
	pesos_i(5764) := b"1111111111111111_1111111111111111_1101110110001101_0100101011110001"; -- -0.13456279400095855
	pesos_i(5765) := b"0000000000000000_0000000000000000_0010010001000011_1101101000111110"; -- 0.14166034713512543
	pesos_i(5766) := b"1111111111111111_1111111111111111_1110101010000010_0110101101100111"; -- -0.08394745574335406
	pesos_i(5767) := b"1111111111111111_1111111111111111_1111000001110100_1000100111111110"; -- -0.060721755596631066
	pesos_i(5768) := b"0000000000000000_0000000000000000_0001100011100110_0000100101010100"; -- 0.09726007741267068
	pesos_i(5769) := b"1111111111111111_1111111111111111_1111110100101101_0111111110001001"; -- -0.01102450283625693
	pesos_i(5770) := b"1111111111111111_1111111111111111_1110110100010111_0110100001101011"; -- -0.07386157405009795
	pesos_i(5771) := b"0000000000000000_0000000000000000_0001100010111001_0010111111111111"; -- 0.09657573676363859
	pesos_i(5772) := b"0000000000000000_0000000000000000_0001010100011101_1011010111101001"; -- 0.08248459756818921
	pesos_i(5773) := b"0000000000000000_0000000000000000_0000010111011010_0001011100111010"; -- 0.022859050438333285
	pesos_i(5774) := b"0000000000000000_0000000000000000_0001010100011000_0011011000001101"; -- 0.08240068271153522
	pesos_i(5775) := b"0000000000000000_0000000000000000_0000111100111101_1000001001100011"; -- 0.059532307770173515
	pesos_i(5776) := b"0000000000000000_0000000000000000_0001111111100001_1011101111101101"; -- 0.12453817880188248
	pesos_i(5777) := b"0000000000000000_0000000000000000_0000000100111101_0010111111110000"; -- 0.004839893455071817
	pesos_i(5778) := b"0000000000000000_0000000000000000_0001111101000001_1010000110010010"; -- 0.12209520151754111
	pesos_i(5779) := b"1111111111111111_1111111111111111_1111100101001101_0110100011101110"; -- -0.026162568829751463
	pesos_i(5780) := b"1111111111111111_1111111111111111_1111111110010011_1011100001001010"; -- -0.0016522236202448407
	pesos_i(5781) := b"1111111111111111_1111111111111111_1111110111001001_1011111110111000"; -- -0.008640306021559421
	pesos_i(5782) := b"1111111111111111_1111111111111111_1110100001101111_0001000000100011"; -- -0.09205531265006292
	pesos_i(5783) := b"0000000000000000_0000000000000000_0000011101100001_1111110111101000"; -- 0.02883898646065522
	pesos_i(5784) := b"0000000000000000_0000000000000000_0000001010111011_1111011110101000"; -- 0.01068065499988717
	pesos_i(5785) := b"1111111111111111_1111111111111111_1101011011000101_0110010100000011"; -- -0.16105049781599792
	pesos_i(5786) := b"0000000000000000_0000000000000000_0000001010111010_0111001101010101"; -- 0.010657509026651274
	pesos_i(5787) := b"1111111111111111_1111111111111111_1111010111001011_1110001011111111"; -- -0.03985768590191691
	pesos_i(5788) := b"0000000000000000_0000000000000000_0001001011111011_1100110101001001"; -- 0.07415469207126181
	pesos_i(5789) := b"0000000000000000_0000000000000000_0001010010111110_1110011001111000"; -- 0.08103790698123867
	pesos_i(5790) := b"0000000000000000_0000000000000000_0001101110001010_1011011101011010"; -- 0.10758539137913707
	pesos_i(5791) := b"1111111111111111_1111111111111111_1110100010010000_0011000111110001"; -- -0.09154975763963195
	pesos_i(5792) := b"0000000000000000_0000000000000000_0000110001111101_1010010100111101"; -- 0.048792197521832364
	pesos_i(5793) := b"0000000000000000_0000000000000000_0000110011111111_1110011111111011"; -- 0.05077981843482696
	pesos_i(5794) := b"0000000000000000_0000000000000000_0000111100010101_0101100111100010"; -- 0.05891954210112757
	pesos_i(5795) := b"1111111111111111_1111111111111111_1111000011100100_0110000110010111"; -- -0.05901517929532898
	pesos_i(5796) := b"1111111111111111_1111111111111111_1110110100101110_1110110111100010"; -- -0.07350266667717828
	pesos_i(5797) := b"1111111111111111_1111111111111111_1110101011010100_0110110111011101"; -- -0.08269608846505978
	pesos_i(5798) := b"1111111111111111_1111111111111111_1110110101001110_1000100000011000"; -- -0.07302045263298623
	pesos_i(5799) := b"1111111111111111_1111111111111111_1110110000110101_0100000011000001"; -- -0.07731242445512142
	pesos_i(5800) := b"0000000000000000_0000000000000000_0010011000110001_0110000011111101"; -- 0.14919096154097475
	pesos_i(5801) := b"0000000000000000_0000000000000000_0000100100000001_0110001100001011"; -- 0.03517741215541457
	pesos_i(5802) := b"1111111111111111_1111111111111111_1101001111001011_0101100110011101"; -- -0.1726783744018599
	pesos_i(5803) := b"0000000000000000_0000000000000000_0000110111111001_0001001000100010"; -- 0.054581769222220966
	pesos_i(5804) := b"0000000000000000_0000000000000000_0001100010000011_0100011110011111"; -- 0.09575317033697121
	pesos_i(5805) := b"1111111111111111_1111111111111111_1110111001101010_0000110000000001"; -- -0.06869435276131511
	pesos_i(5806) := b"1111111111111111_1111111111111111_1101000000110001_0100101001110110"; -- -0.18674788117201793
	pesos_i(5807) := b"1111111111111111_1111111111111111_1110000011010110_0010011101111011"; -- -0.12173226597322213
	pesos_i(5808) := b"1111111111111111_1111111111111111_1101001110011011_1001010000000001"; -- -0.17340731593332742
	pesos_i(5809) := b"0000000000000000_0000000000000000_0000011011100000_0010100101100011"; -- 0.02685793570463557
	pesos_i(5810) := b"1111111111111111_1111111111111111_1101110011011001_1110011110100011"; -- -0.13730003619393813
	pesos_i(5811) := b"0000000000000000_0000000000000000_0010101011111010_1000111001000111"; -- 0.1678856776696603
	pesos_i(5812) := b"1111111111111111_1111111111111111_1101111110110100_1001111000010100"; -- -0.1261502458072093
	pesos_i(5813) := b"1111111111111111_1111111111111111_1111010000011111_0001111010100100"; -- -0.04640015118885613
	pesos_i(5814) := b"0000000000000000_0000000000000000_0000011101010100_1111010100111011"; -- 0.02864010518067844
	pesos_i(5815) := b"0000000000000000_0000000000000000_0010010100100111_0001100011011100"; -- 0.14512782458862492
	pesos_i(5816) := b"0000000000000000_0000000000000000_0000111111000001_0010100101100100"; -- 0.06154116335310825
	pesos_i(5817) := b"0000000000000000_0000000000000000_0000111001001001_0001100010001001"; -- 0.05580285396203319
	pesos_i(5818) := b"0000000000000000_0000000000000000_0000110000100101_1111010011100010"; -- 0.047454171454390966
	pesos_i(5819) := b"0000000000000000_0000000000000000_0000011111010010_0011111010111101"; -- 0.030551835281979505
	pesos_i(5820) := b"1111111111111111_1111111111111111_1110011100000101_0011010010011011"; -- -0.09757682045883652
	pesos_i(5821) := b"0000000000000000_0000000000000000_0010010111001001_1100000001001101"; -- 0.14760972854174312
	pesos_i(5822) := b"0000000000000000_0000000000000000_0000010101011101_0101000101110100"; -- 0.020955172291101044
	pesos_i(5823) := b"1111111111111111_1111111111111111_1111000011001000_1111000101011000"; -- -0.05943385707006472
	pesos_i(5824) := b"1111111111111111_1111111111111111_1110100010001001_1110110110001001"; -- -0.09164538776874943
	pesos_i(5825) := b"0000000000000000_0000000000000000_0001001110011111_0100101110001011"; -- 0.0766494001990652
	pesos_i(5826) := b"1111111111111111_1111111111111111_1110110010110001_0001111010100001"; -- -0.07542236859464234
	pesos_i(5827) := b"1111111111111111_1111111111111111_1110100011010011_1000000011100111"; -- -0.09052271243373071
	pesos_i(5828) := b"0000000000000000_0000000000000000_0000101101110111_0011000010011110"; -- 0.04478744364147946
	pesos_i(5829) := b"1111111111111111_1111111111111111_1111001111101101_0011111101100111"; -- -0.0471611378962285
	pesos_i(5830) := b"1111111111111111_1111111111111111_1110001111110101_1111111100101001"; -- -0.10952763784043543
	pesos_i(5831) := b"0000000000000000_0000000000000000_0010001010000001_1111001111100111"; -- 0.13479542144387552
	pesos_i(5832) := b"0000000000000000_0000000000000000_0000000000010100_0010000100001001"; -- 0.00030714487253742
	pesos_i(5833) := b"1111111111111111_1111111111111111_1110101111001001_0001011010000100"; -- -0.07896289143675922
	pesos_i(5834) := b"0000000000000000_0000000000000000_0000100111111101_0100111001100110"; -- 0.03902139659915326
	pesos_i(5835) := b"0000000000000000_0000000000000000_0001011010000110_0101001010111111"; -- 0.08798710983393976
	pesos_i(5836) := b"1111111111111111_1111111111111111_1111011101110010_0111111100010000"; -- -0.03340917446127807
	pesos_i(5837) := b"1111111111111111_1111111111111111_1111100011100001_1011001101101111"; -- -0.0278060773062531
	pesos_i(5838) := b"1111111111111111_1111111111111111_1110011000011101_1110110011101100"; -- -0.10110587358022376
	pesos_i(5839) := b"0000000000000000_0000000000000000_0010011001001011_0110011011011001"; -- 0.14958803936691056
	pesos_i(5840) := b"0000000000000000_0000000000000000_0010011101100000_0001010010110101"; -- 0.15380982807550123
	pesos_i(5841) := b"1111111111111111_1111111111111111_1101110110100011_0100111110100001"; -- -0.1342268210899333
	pesos_i(5842) := b"0000000000000000_0000000000000000_0010011110110110_1110000001101101"; -- 0.15513422637293448
	pesos_i(5843) := b"0000000000000000_0000000000000000_0010100011100110_0100100100111001"; -- 0.15976388589978097
	pesos_i(5844) := b"1111111111111111_1111111111111111_1110111010111011_1101001011110011"; -- -0.06744653288669625
	pesos_i(5845) := b"0000000000000000_0000000000000000_0001110101010011_0011011001101011"; -- 0.11455097315428298
	pesos_i(5846) := b"0000000000000000_0000000000000000_0000100100111110_1001101011100010"; -- 0.03611152657662886
	pesos_i(5847) := b"0000000000000000_0000000000000000_0001010001010110_1100111001110000"; -- 0.0794495604902559
	pesos_i(5848) := b"1111111111111111_1111111111111111_1111100001110111_1011110101000000"; -- -0.02942292380797312
	pesos_i(5849) := b"1111111111111111_1111111111111111_1111101111110101_1100111010010011"; -- -0.01578053387824855
	pesos_i(5850) := b"0000000000000000_0000000000000000_0000000110111101_1000110000111100"; -- 0.0067985198368540915
	pesos_i(5851) := b"1111111111111111_1111111111111111_1101111011101111_1010011111110010"; -- -0.12915563915631434
	pesos_i(5852) := b"0000000000000000_0000000000000000_0000110110001101_0010000100100100"; -- 0.05293471455220912
	pesos_i(5853) := b"0000000000000000_0000000000000000_0000111111100000_0110101001000110"; -- 0.062018053157264406
	pesos_i(5854) := b"1111111111111111_1111111111111111_1110001100000011_1111010010000001"; -- -0.11322090017455477
	pesos_i(5855) := b"1111111111111111_1111111111111111_1111001111010011_1101110110001001"; -- -0.04754844108038245
	pesos_i(5856) := b"0000000000000000_0000000000000000_0000001000101101_0100011011100000"; -- 0.00850336992205783
	pesos_i(5857) := b"0000000000000000_0000000000000000_0000100011111111_0101110110000101"; -- 0.035146565382523684
	pesos_i(5858) := b"1111111111111111_1111111111111111_1111110111111000_1010101101011111"; -- -0.0079243558957514
	pesos_i(5859) := b"0000000000000000_0000000000000000_0000010010011101_0101011101100100"; -- 0.018025838828507137
	pesos_i(5860) := b"0000000000000000_0000000000000000_0001010010000101_0000001101010110"; -- 0.08015461783810963
	pesos_i(5861) := b"0000000000000000_0000000000000000_0010000110111101_0000011111110110"; -- 0.13179063567026725
	pesos_i(5862) := b"1111111111111111_1111111111111111_1111011001010101_0001000001000001"; -- -0.03776453410280076
	pesos_i(5863) := b"0000000000000000_0000000000000000_0010010000010000_0000101110011111"; -- 0.14086983332243377
	pesos_i(5864) := b"0000000000000000_0000000000000000_0001101001010000_1011011001001100"; -- 0.10279406888471729
	pesos_i(5865) := b"0000000000000000_0000000000000000_0001011011010011_1011110100010101"; -- 0.08916837472004778
	pesos_i(5866) := b"0000000000000000_0000000000000000_0001100101010111_0000100101001001"; -- 0.09898431801628338
	pesos_i(5867) := b"0000000000000000_0000000000000000_0000110010100001_1010111110010101"; -- 0.04934213059114658
	pesos_i(5868) := b"1111111111111111_1111111111111111_1111101111100001_0010111111111000"; -- -0.01609516319451149
	pesos_i(5869) := b"1111111111111111_1111111111111111_1101001000100101_0100100101001010"; -- -0.17911855632462906
	pesos_i(5870) := b"0000000000000000_0000000000000000_0000101000110010_1111111010101000"; -- 0.039840618259938544
	pesos_i(5871) := b"1111111111111111_1111111111111111_1101100001100001_0010000011111001"; -- -0.15476793217851417
	pesos_i(5872) := b"0000000000000000_0000000000000000_0000100101101101_1011000101010011"; -- 0.03683002735033955
	pesos_i(5873) := b"1111111111111111_1111111111111111_1101111010011100_0110110010111100"; -- -0.13042564785712246
	pesos_i(5874) := b"0000000000000000_0000000000000000_0010110000101011_1110110101011111"; -- 0.17254527626029867
	pesos_i(5875) := b"1111111111111111_1111111111111111_1110010111111000_0010011110110001"; -- -0.1016822044314656
	pesos_i(5876) := b"0000000000000000_0000000000000000_0010001001110110_1011100110110110"; -- 0.13462410641283745
	pesos_i(5877) := b"1111111111111111_1111111111111111_1101101110010101_0010011101001011"; -- -0.1422553483835253
	pesos_i(5878) := b"1111111111111111_1111111111111111_1101110001111100_1100101001010001"; -- -0.1387208512745801
	pesos_i(5879) := b"0000000000000000_0000000000000000_0001100000101000_1001100110111111"; -- 0.09436951555036018
	pesos_i(5880) := b"0000000000000000_0000000000000000_0000111011010001_0001111100011100"; -- 0.05787844110851734
	pesos_i(5881) := b"1111111111111111_1111111111111111_1110001100111111_0000110000011111"; -- -0.11231922377298416
	pesos_i(5882) := b"0000000000000000_0000000000000000_0000000010101101_0100010001101000"; -- 0.002643847777461059
	pesos_i(5883) := b"1111111111111111_1111111111111111_1101011110000010_1100001011011110"; -- -0.15816099245253626
	pesos_i(5884) := b"1111111111111111_1111111111111111_1110100000000000_1011000001010110"; -- -0.09373948964285138
	pesos_i(5885) := b"0000000000000000_0000000000000000_0000001100001110_1111101011110100"; -- 0.011947331007580803
	pesos_i(5886) := b"1111111111111111_1111111111111111_1101111011000000_0101111000011000"; -- -0.1298772039731116
	pesos_i(5887) := b"0000000000000000_0000000000000000_0010100111100110_0000110011000111"; -- 0.16366653307065462
	pesos_i(5888) := b"0000000000000000_0000000000000000_0010101000111010_1000100111111001"; -- 0.16495573348835288
	pesos_i(5889) := b"1111111111111111_1111111111111111_1110010000100011_0010101100000100"; -- -0.10883837839674754
	pesos_i(5890) := b"0000000000000000_0000000000000000_0001110111010101_0001010000110011"; -- 0.11653257596112697
	pesos_i(5891) := b"0000000000000000_0000000000000000_0010110011010001_1000100001100110"; -- 0.17507221681418406
	pesos_i(5892) := b"0000000000000000_0000000000000000_0000001001010001_1010101101100011"; -- 0.009058677464792993
	pesos_i(5893) := b"0000000000000000_0000000000000000_0000101110011101_0011111000011011"; -- 0.045368081661732305
	pesos_i(5894) := b"0000000000000000_0000000000000000_0000110001101001_1101011111001010"; -- 0.04849003496089757
	pesos_i(5895) := b"1111111111111111_1111111111111111_1111100101010011_1110101001000111"; -- -0.026063306531454212
	pesos_i(5896) := b"0000000000000000_0000000000000000_0000110010000111_1001100110001000"; -- 0.04894408763533161
	pesos_i(5897) := b"0000000000000000_0000000000000000_0001110000110100_0100111001011110"; -- 0.11017312819432519
	pesos_i(5898) := b"1111111111111111_1111111111111111_1101101010001111_1001110110011011"; -- -0.1462460991336574
	pesos_i(5899) := b"1111111111111111_1111111111111111_1101001110111111_0000001010010111"; -- -0.1728666669128501
	pesos_i(5900) := b"1111111111111111_1111111111111111_1110001010010110_1100101101001011"; -- -0.11488656449127563
	pesos_i(5901) := b"0000000000000000_0000000000000000_0001001010000000_0011001010010111"; -- 0.07226864039203142
	pesos_i(5902) := b"0000000000000000_0000000000000000_0000111101010011_1000101011001101"; -- 0.05986850262603399
	pesos_i(5903) := b"1111111111111111_1111111111111111_1111100000100011_1001101100001000"; -- -0.030706701911917978
	pesos_i(5904) := b"0000000000000000_0000000000000000_0010011000110111_0110010011111110"; -- 0.14928275310650332
	pesos_i(5905) := b"1111111111111111_1111111111111111_1110100110001001_1011011111010000"; -- -0.08774233991455015
	pesos_i(5906) := b"1111111111111111_1111111111111111_1101111001000110_1111000010111010"; -- -0.13173003628979638
	pesos_i(5907) := b"1111111111111111_1111111111111111_1101111110101000_1000010110101011"; -- -0.12633480615812784
	pesos_i(5908) := b"0000000000000000_0000000000000000_0000010111111101_1010010001001111"; -- 0.023401517129626976
	pesos_i(5909) := b"1111111111111111_1111111111111111_1101011000100010_0000100011000100"; -- -0.16354317866354146
	pesos_i(5910) := b"0000000000000000_0000000000000000_0001101101101100_0110110000111111"; -- 0.10712315120327393
	pesos_i(5911) := b"1111111111111111_1111111111111111_1101111010111100_0010000010010000"; -- -0.1299419066728223
	pesos_i(5912) := b"0000000000000000_0000000000000000_0010010101000100_0111100110000001"; -- 0.1455760898253589
	pesos_i(5913) := b"0000000000000000_0000000000000000_0000101110100000_0001110001110011"; -- 0.045411852030555394
	pesos_i(5914) := b"1111111111111111_1111111111111111_1101100001001111_0101100101000100"; -- -0.15503923497439046
	pesos_i(5915) := b"1111111111111111_1111111111111111_1111111110111010_1001010011001100"; -- -0.0010592461572608584
	pesos_i(5916) := b"1111111111111111_1111111111111111_1111101011101111_0110111110110100"; -- -0.019783991462127712
	pesos_i(5917) := b"1111111111111111_1111111111111111_1101010101110011_0010010011010111"; -- -0.16621179353660423
	pesos_i(5918) := b"1111111111111111_1111111111111111_1110010010111000_0111011000101010"; -- -0.10656033974589417
	pesos_i(5919) := b"1111111111111111_1111111111111111_1101101000010101_0001101010011100"; -- -0.14811547943910147
	pesos_i(5920) := b"0000000000000000_0000000000000000_0000111011101101_1011001111100110"; -- 0.05831455574140204
	pesos_i(5921) := b"1111111111111111_1111111111111111_1110101000011001_1111010011000110"; -- -0.08554144062378409
	pesos_i(5922) := b"0000000000000000_0000000000000000_0010010101010100_1010100101001100"; -- 0.14582307919724274
	pesos_i(5923) := b"0000000000000000_0000000000000000_0000111101001010_1001001100010101"; -- 0.059731667261401125
	pesos_i(5924) := b"1111111111111111_1111111111111111_1110010010011110_0010011100011101"; -- -0.10696178008709699
	pesos_i(5925) := b"0000000000000000_0000000000000000_0010111010001110_1111001001111000"; -- 0.1818687003067532
	pesos_i(5926) := b"1111111111111111_1111111111111111_1111010111101000_0110011000000001"; -- -0.039422631136506826
	pesos_i(5927) := b"1111111111111111_1111111111111111_1111000001101111_1010010110000100"; -- -0.06079640890927772
	pesos_i(5928) := b"1111111111111111_1111111111111111_1101011010100010_0001101100100111"; -- -0.16158895776718105
	pesos_i(5929) := b"1111111111111111_1111111111111111_1110101000100110_0110000100001110"; -- -0.08535188109039603
	pesos_i(5930) := b"0000000000000000_0000000000000000_0010000010110100_0111011001100011"; -- 0.12775363849460286
	pesos_i(5931) := b"1111111111111111_1111111111111111_1110010011011111_0111000010111111"; -- -0.10596556985959929
	pesos_i(5932) := b"1111111111111111_1111111111111111_1101100001101100_1100111001001000"; -- -0.1545897554752674
	pesos_i(5933) := b"1111111111111111_1111111111111111_1111011010011100_0111100001110100"; -- -0.03667494923530157
	pesos_i(5934) := b"1111111111111111_1111111111111111_1111110001001110_0000011101010110"; -- -0.014434377082209167
	pesos_i(5935) := b"1111111111111111_1111111111111111_1110010010100001_0000111101100101"; -- -0.10691741729456795
	pesos_i(5936) := b"0000000000000000_0000000000000000_0000001000011100_0010110010111000"; -- 0.008242411625930063
	pesos_i(5937) := b"0000000000000000_0000000000000000_0001110100000000_1111111110010100"; -- 0.11329648361999589
	pesos_i(5938) := b"1111111111111111_1111111111111111_1110011111011011_0001011111110011"; -- -0.09431314760471217
	pesos_i(5939) := b"1111111111111111_1111111111111111_1111101010100011_1110111010101101"; -- -0.02093609113480617
	pesos_i(5940) := b"0000000000000000_0000000000000000_0010010011110110_1101100100101100"; -- 0.144391606487223
	pesos_i(5941) := b"0000000000000000_0000000000000000_0010111010101111_0011010010110101"; -- 0.18236092964663084
	pesos_i(5942) := b"0000000000000000_0000000000000000_0010000011011011_0100101100100011"; -- 0.12834615329363824
	pesos_i(5943) := b"0000000000000000_0000000000000000_0010110000000010_0001110000011110"; -- 0.17190719355950837
	pesos_i(5944) := b"1111111111111111_1111111111111111_1111000101101110_1010100000101111"; -- -0.05690525875529834
	pesos_i(5945) := b"1111111111111111_1111111111111111_1111101011100110_0110110100110010"; -- -0.019921470052483355
	pesos_i(5946) := b"1111111111111111_1111111111111111_1110101100110111_0100000101000101"; -- -0.08118812627389828
	pesos_i(5947) := b"1111111111111111_1111111111111111_1110000111110111_0001110011011001"; -- -0.11732310975565374
	pesos_i(5948) := b"0000000000000000_0000000000000000_0000100101010100_1101101100110111"; -- 0.03645105445776251
	pesos_i(5949) := b"0000000000000000_0000000000000000_0010001001110101_0010011110110011"; -- 0.13460014451171165
	pesos_i(5950) := b"0000000000000000_0000000000000000_0000010110001010_1000000011110001"; -- 0.021644648465953036
	pesos_i(5951) := b"0000000000000000_0000000000000000_0000010101011101_0100101100110110"; -- 0.020954800223243267
	pesos_i(5952) := b"0000000000000000_0000000000000000_0001111011010111_1010111101111111"; -- 0.12047859992496726
	pesos_i(5953) := b"0000000000000000_0000000000000000_0000101101010110_0110010111010101"; -- 0.04428707542760742
	pesos_i(5954) := b"1111111111111111_1111111111111111_1111101010111111_0111011011110001"; -- -0.02051598187324959
	pesos_i(5955) := b"1111111111111111_1111111111111111_1101011111101001_1010000111010101"; -- -0.15659130629643006
	pesos_i(5956) := b"0000000000000000_0000000000000000_0010000101010011_1101000100110011"; -- 0.13018519882321924
	pesos_i(5957) := b"1111111111111111_1111111111111111_1110100111110011_1100100001100100"; -- -0.08612391999217645
	pesos_i(5958) := b"0000000000000000_0000000000000000_0010011010101010_1110011001011111"; -- 0.15104522524294497
	pesos_i(5959) := b"1111111111111111_1111111111111111_1101111011001010_0101000110110100"; -- -0.129725354749366
	pesos_i(5960) := b"1111111111111111_1111111111111111_1110111000011101_1011101001110011"; -- -0.06985888198731362
	pesos_i(5961) := b"1111111111111111_1111111111111111_1101100111010110_1001011100011111"; -- -0.14906936161717696
	pesos_i(5962) := b"0000000000000000_0000000000000000_0001101100010101_0000001110101100"; -- 0.10578940350857466
	pesos_i(5963) := b"0000000000000000_0000000000000000_0010101000001011_1110000001111100"; -- 0.16424372696518874
	pesos_i(5964) := b"0000000000000000_0000000000000000_0001001100101110_0010000011100111"; -- 0.07492261540574689
	pesos_i(5965) := b"0000000000000000_0000000000000000_0001010000101111_1010010010001000"; -- 0.07885196999240746
	pesos_i(5966) := b"0000000000000000_0000000000000000_0010001111000100_0001001110110000"; -- 0.1397106462255437
	pesos_i(5967) := b"0000000000000000_0000000000000000_0000100110001111_1011001010110100"; -- 0.03734890827329139
	pesos_i(5968) := b"0000000000000000_0000000000000000_0010101001010111_1101001110011100"; -- 0.16540262766445277
	pesos_i(5969) := b"1111111111111111_1111111111111111_1101001101011100_0010100111010111"; -- -0.17437494766519873
	pesos_i(5970) := b"0000000000000000_0000000000000000_0010011010001011_1001001000010010"; -- 0.15056717826447147
	pesos_i(5971) := b"1111111111111111_1111111111111111_1111011010100110_1010111001011100"; -- -0.03651914828394455
	pesos_i(5972) := b"0000000000000000_0000000000000000_0000001000111101_1001000000000111"; -- 0.008751870807920996
	pesos_i(5973) := b"1111111111111111_1111111111111111_1101100101110111_1101110101111100"; -- -0.15051475257319002
	pesos_i(5974) := b"1111111111111111_1111111111111111_1110101100101000_0111110011011110"; -- -0.08141345574193863
	pesos_i(5975) := b"1111111111111111_1111111111111111_1110111110001110_0110110010010101"; -- -0.06423302995535754
	pesos_i(5976) := b"0000000000000000_0000000000000000_0001010001001101_1110010110111101"; -- 0.07931362029381113
	pesos_i(5977) := b"0000000000000000_0000000000000000_0000000100001000_1110101000101101"; -- 0.004042278368047588
	pesos_i(5978) := b"1111111111111111_1111111111111111_1111000101101101_0010011001001110"; -- -0.05692825887079684
	pesos_i(5979) := b"1111111111111111_1111111111111111_1110001011001001_1000100000011101"; -- -0.11411237030424462
	pesos_i(5980) := b"0000000000000000_0000000000000000_0001000000100010_0000001101011000"; -- 0.06301899819589817
	pesos_i(5981) := b"1111111111111111_1111111111111111_1101101011011000_0101011011010101"; -- -0.1451364259664962
	pesos_i(5982) := b"1111111111111111_1111111111111111_1111101101000110_1010000011010110"; -- -0.018453548147221072
	pesos_i(5983) := b"1111111111111111_1111111111111111_1101100100101010_1110010101100001"; -- -0.15168920887191834
	pesos_i(5984) := b"0000000000000000_0000000000000000_0000001001011111_0111111110000000"; -- 0.009269684612445067
	pesos_i(5985) := b"1111111111111111_1111111111111111_1110110111000001_1110011001000001"; -- -0.07126007953783177
	pesos_i(5986) := b"1111111111111111_1111111111111111_1111101100001110_1111100111101000"; -- -0.019302731483779433
	pesos_i(5987) := b"0000000000000000_0000000000000000_0010010110100011_0000010101001001"; -- 0.1470187477387802
	pesos_i(5988) := b"1111111111111111_1111111111111111_1111011000011100_1100111111001011"; -- -0.03862286858159987
	pesos_i(5989) := b"0000000000000000_0000000000000000_0001010000000011_0001101101101001"; -- 0.07817241012048211
	pesos_i(5990) := b"1111111111111111_1111111111111111_1111100001100101_1010001000001110"; -- -0.029699203202973142
	pesos_i(5991) := b"1111111111111111_1111111111111111_1111100000101011_0010100101011000"; -- -0.03059140790287901
	pesos_i(5992) := b"1111111111111111_1111111111111111_1110101001100000_1101110001111000"; -- -0.08445951523531839
	pesos_i(5993) := b"1111111111111111_1111111111111111_1111100010101111_0110000011011100"; -- -0.02857393874851584
	pesos_i(5994) := b"1111111111111111_1111111111111111_1101101001101101_1000001010001000"; -- -0.1467665116184749
	pesos_i(5995) := b"0000000000000000_0000000000000000_0010010101010001_0111010000101000"; -- 0.14577413529938732
	pesos_i(5996) := b"1111111111111111_1111111111111111_1110010001101010_0101111011001001"; -- -0.10775191874299835
	pesos_i(5997) := b"1111111111111111_1111111111111111_1111011110101111_0010101101110100"; -- -0.03248337179826919
	pesos_i(5998) := b"1111111111111111_1111111111111111_1110000011111101_0010000111011111"; -- -0.12113750738365714
	pesos_i(5999) := b"1111111111111111_1111111111111111_1111011011011001_1111110000000101"; -- -0.03573632121053829
	pesos_i(6000) := b"1111111111111111_1111111111111111_1110110001100000_0011110001011101"; -- -0.0766565583199771
	pesos_i(6001) := b"1111111111111111_1111111111111111_1101011011100011_1101001001100001"; -- -0.16058621532806602
	pesos_i(6002) := b"1111111111111111_1111111111111111_1111010110111000_0100101000101101"; -- -0.040156711572479735
	pesos_i(6003) := b"1111111111111111_1111111111111111_1111100001110101_0001000110000001"; -- -0.029463678385414697
	pesos_i(6004) := b"0000000000000000_0000000000000000_0000110111001100_1010111011110100"; -- 0.0539044709124216
	pesos_i(6005) := b"0000000000000000_0000000000000000_0000010100000010_0000111100101110"; -- 0.0195626722719775
	pesos_i(6006) := b"0000000000000000_0000000000000000_0010010011000100_0101100100100110"; -- 0.14362103632158313
	pesos_i(6007) := b"0000000000000000_0000000000000000_0001101110010110_0010111000100011"; -- 0.1077603183528127
	pesos_i(6008) := b"0000000000000000_0000000000000000_0001001100100111_1010101010010011"; -- 0.07482400968669525
	pesos_i(6009) := b"0000000000000000_0000000000000000_0000001011000101_1010001011011001"; -- 0.010828187861646642
	pesos_i(6010) := b"0000000000000000_0000000000000000_0000010100011011_0101010000101100"; -- 0.019948254325551914
	pesos_i(6011) := b"1111111111111111_1111111111111111_1111110001111001_1010101100101001"; -- -0.013768484645514932
	pesos_i(6012) := b"1111111111111111_1111111111111111_1111100000100000_1010100011110110"; -- -0.03075164795837516
	pesos_i(6013) := b"0000000000000000_0000000000000000_0000000100110101_0011100110101000"; -- 0.004718402450184799
	pesos_i(6014) := b"1111111111111111_1111111111111111_1111000110110110_1000111101100001"; -- -0.055808104339127515
	pesos_i(6015) := b"1111111111111111_1111111111111111_1101110110001111_1111111110010011"; -- -0.13452150967361282
	pesos_i(6016) := b"0000000000000000_0000000000000000_0000111001100010_0001000111111110"; -- 0.05618393377109221
	pesos_i(6017) := b"0000000000000000_0000000000000000_0000001101111101_1110001101001000"; -- 0.013639645610559045
	pesos_i(6018) := b"0000000000000000_0000000000000000_0000111111110111_0100101001001110"; -- 0.06236709988565833
	pesos_i(6019) := b"0000000000000000_0000000000000000_0001010111001001_0111100111010001"; -- 0.08510552752579625
	pesos_i(6020) := b"0000000000000000_0000000000000000_0010011011111101_1101010100011001"; -- 0.15231067524363107
	pesos_i(6021) := b"0000000000000000_0000000000000000_0000010010001001_0000000101110001"; -- 0.017715540004575824
	pesos_i(6022) := b"1111111111111111_1111111111111111_1110000111101001_1001000110000100"; -- -0.11752977883888595
	pesos_i(6023) := b"0000000000000000_0000000000000000_0000100001110101_0010111011111000"; -- 0.03303807792627811
	pesos_i(6024) := b"0000000000000000_0000000000000000_0000010010010000_0111001100100000"; -- 0.01782912749593471
	pesos_i(6025) := b"0000000000000000_0000000000000000_0010101011110100_1010110110101001"; -- 0.16779599546029722
	pesos_i(6026) := b"1111111111111111_1111111111111111_1111011011011011_1011001010000110"; -- -0.03571018443096179
	pesos_i(6027) := b"0000000000000000_0000000000000000_0010100000000011_1100011110111001"; -- 0.15630768071127737
	pesos_i(6028) := b"0000000000000000_0000000000000000_0000001100010100_1111101101101110"; -- 0.012038912170873805
	pesos_i(6029) := b"1111111111111111_1111111111111111_1111010111101010_1111110111010000"; -- -0.039383064895909446
	pesos_i(6030) := b"1111111111111111_1111111111111111_1111100011100100_1111011011010100"; -- -0.027756284066751017
	pesos_i(6031) := b"0000000000000000_0000000000000000_0000011110110101_1001101101110010"; -- 0.030114856066287027
	pesos_i(6032) := b"1111111111111111_1111111111111111_1101110100010000_0101000001101101"; -- -0.13646981565569583
	pesos_i(6033) := b"1111111111111111_1111111111111111_1111011110011000_0110000011011111"; -- -0.032831140210613285
	pesos_i(6034) := b"1111111111111111_1111111111111111_1101100010101111_0101001101111101"; -- -0.15357473553508205
	pesos_i(6035) := b"1111111111111111_1111111111111111_1111100001000000_1101010010101010"; -- -0.030260761822606383
	pesos_i(6036) := b"0000000000000000_0000000000000000_0001010011101100_1010011111110011"; -- 0.08173608484290563
	pesos_i(6037) := b"1111111111111111_1111111111111111_1101100101101001_1000001111111100"; -- -0.1507337101770803
	pesos_i(6038) := b"1111111111111111_1111111111111111_1111000001110011_0111100010101111"; -- -0.0607380459094077
	pesos_i(6039) := b"0000000000000000_0000000000000000_0010000101110000_1100110101101101"; -- 0.1306274788082527
	pesos_i(6040) := b"1111111111111111_1111111111111111_1101110101000110_1110110010110100"; -- -0.13563652605272697
	pesos_i(6041) := b"1111111111111111_1111111111111111_1101101010100011_1011011110010000"; -- -0.14593937609791588
	pesos_i(6042) := b"1111111111111111_1111111111111111_1111110100011110_1011001000001010"; -- -0.011250374327806857
	pesos_i(6043) := b"1111111111111111_1111111111111111_1111100111110101_0000110000000001"; -- -0.02360463111899888
	pesos_i(6044) := b"1111111111111111_1111111111111111_1101100011010011_1110010010110100"; -- -0.15301676385403376
	pesos_i(6045) := b"1111111111111111_1111111111111111_1110101011010101_1010111010110001"; -- -0.082676965486313
	pesos_i(6046) := b"0000000000000000_0000000000000000_0001000010000000_0001100000000100"; -- 0.0644545565478016
	pesos_i(6047) := b"0000000000000000_0000000000000000_0010001001110010_0010011001100011"; -- 0.13455428999362776
	pesos_i(6048) := b"1111111111111111_1111111111111111_1111100110000010_1000111101101100"; -- -0.02535155886766996
	pesos_i(6049) := b"0000000000000000_0000000000000000_0000011111000111_1001100001011110"; -- 0.0303893308454741
	pesos_i(6050) := b"1111111111111111_1111111111111111_1110100101001011_1111110000000011"; -- -0.0886843198228017
	pesos_i(6051) := b"1111111111111111_1111111111111111_1111000111111000_0010010011110000"; -- -0.05480736877160341
	pesos_i(6052) := b"1111111111111111_1111111111111111_1110010000101110_0111101111000101"; -- -0.10866571836867912
	pesos_i(6053) := b"0000000000000000_0000000000000000_0001100110001011_1011011100011101"; -- 0.09978813607133849
	pesos_i(6054) := b"0000000000000000_0000000000000000_0001101100000000_1100010010010111"; -- 0.1054804676190948
	pesos_i(6055) := b"1111111111111111_1111111111111111_1111111000110001_1011110111010011"; -- -0.007053504983959874
	pesos_i(6056) := b"1111111111111111_1111111111111111_1101111111001110_0110010101001001"; -- -0.1257569023676965
	pesos_i(6057) := b"0000000000000000_0000000000000000_0000001101000011_1111101110010110"; -- 0.012756084642533127
	pesos_i(6058) := b"0000000000000000_0000000000000000_0010010100010101_0101001110001001"; -- 0.14485666371793107
	pesos_i(6059) := b"0000000000000000_0000000000000000_0000010010101000_1100110100101011"; -- 0.018200705633937005
	pesos_i(6060) := b"1111111111111111_1111111111111111_1111100000000001_1000110110000110"; -- -0.03122630572460927
	pesos_i(6061) := b"0000000000000000_0000000000000000_0000101101111001_1110000010101010"; -- 0.04482845452207149
	pesos_i(6062) := b"1111111111111111_1111111111111111_1110101010011111_0100111011100111"; -- -0.08350664954157007
	pesos_i(6063) := b"1111111111111111_1111111111111111_1111001011110110_1101001000111110"; -- -0.05092130659131073
	pesos_i(6064) := b"1111111111111111_1111111111111111_1111001110011100_0000010101010011"; -- -0.04840056164813025
	pesos_i(6065) := b"1111111111111111_1111111111111111_1111100111100011_1101001000011000"; -- -0.023867482288880377
	pesos_i(6066) := b"0000000000000000_0000000000000000_0000101100101010_0000011000110000"; -- 0.0436099880153342
	pesos_i(6067) := b"0000000000000000_0000000000000000_0001000000110000_1000100110000000"; -- 0.06324061754755213
	pesos_i(6068) := b"1111111111111111_1111111111111111_1110100100100010_0110111101010101"; -- -0.08931831520801743
	pesos_i(6069) := b"1111111111111111_1111111111111111_1110101001000010_1101111010101000"; -- -0.08491714848231306
	pesos_i(6070) := b"1111111111111111_1111111111111111_1101111110110001_1001110010101001"; -- -0.12619610670918407
	pesos_i(6071) := b"1111111111111111_1111111111111111_1100101011111000_1010110000010000"; -- -0.20714306447716668
	pesos_i(6072) := b"1111111111111111_1111111111111111_1111100111000110_1111111100000000"; -- -0.02430731066189526
	pesos_i(6073) := b"1111111111111111_1111111111111111_1110001000011100_1101110000111100"; -- -0.11674712699369157
	pesos_i(6074) := b"1111111111111111_1111111111111111_1110010100000010_0110000111110101"; -- -0.10543239367463027
	pesos_i(6075) := b"0000000000000000_0000000000000000_0010000010111110_1100010111101011"; -- 0.12791096671393717
	pesos_i(6076) := b"0000000000000000_0000000000000000_0000110110110110_0100110111000101"; -- 0.05356298507429992
	pesos_i(6077) := b"1111111111111111_1111111111111111_1111101101011001_0110010011111100"; -- -0.018167198598561307
	pesos_i(6078) := b"0000000000000000_0000000000000000_0010010111101011_0100010101011001"; -- 0.1481211987604521
	pesos_i(6079) := b"1111111111111111_1111111111111111_1110010100100001_1111011001010000"; -- -0.10495052868348405
	pesos_i(6080) := b"0000000000000000_0000000000000000_0010000110010010_0000001010010001"; -- 0.13113418610121744
	pesos_i(6081) := b"1111111111111111_1111111111111111_1110000101000100_0010010000100110"; -- -0.12005399775895685
	pesos_i(6082) := b"0000000000000000_0000000000000000_0010000100001111_1000110111111101"; -- 0.12914359509840037
	pesos_i(6083) := b"1111111111111111_1111111111111111_1111100001101100_0001100110010011"; -- -0.029600526482984182
	pesos_i(6084) := b"0000000000000000_0000000000000000_0001000000110010_1111010111101011"; -- 0.06327759724700081
	pesos_i(6085) := b"1111111111111111_1111111111111111_1110010001110100_1111000110001110"; -- -0.10759058273064782
	pesos_i(6086) := b"1111111111111111_1111111111111111_1110001101111101_1001000000101100"; -- -0.11136530796327343
	pesos_i(6087) := b"0000000000000000_0000000000000000_0000101011101000_0001111100110111"; -- 0.04260439951602607
	pesos_i(6088) := b"0000000000000000_0000000000000000_0000110001111000_1100101100001101"; -- 0.0487181573541636
	pesos_i(6089) := b"1111111111111111_1111111111111111_1110110010100100_1001011011011111"; -- -0.07561356605967186
	pesos_i(6090) := b"1111111111111111_1111111111111111_1110100110101111_1110000000001011"; -- -0.0871601079543117
	pesos_i(6091) := b"0000000000000000_0000000000000000_0000110110000101_0001100101101111"; -- 0.052812184830276825
	pesos_i(6092) := b"0000000000000000_0000000000000000_0001001110011100_0000111000110011"; -- 0.07659996737687903
	pesos_i(6093) := b"1111111111111111_1111111111111111_1101100111001100_0110111101011111"; -- -0.14922431890610227
	pesos_i(6094) := b"0000000000000000_0000000000000000_0000010011001100_1000000110101110"; -- 0.018745522581779903
	pesos_i(6095) := b"1111111111111111_1111111111111111_1111111011111000_0110110011101111"; -- -0.00402182747491306
	pesos_i(6096) := b"1111111111111111_1111111111111111_1101110000101010_1110101000110000"; -- -0.1399701721309614
	pesos_i(6097) := b"0000000000000000_0000000000000000_0000000101001110_0001010011011110"; -- 0.005097679345452491
	pesos_i(6098) := b"1111111111111111_1111111111111111_1110101011001010_0000010101101111"; -- -0.08285490067186342
	pesos_i(6099) := b"1111111111111111_1111111111111111_1101100111001000_1101001101011000"; -- -0.1492793950347417
	pesos_i(6100) := b"1111111111111111_1111111111111111_1111101010010101_1100011101111000"; -- -0.021152051081496887
	pesos_i(6101) := b"0000000000000000_0000000000000000_0000000110110110_1111010010101100"; -- 0.006697933215503347
	pesos_i(6102) := b"0000000000000000_0000000000000000_0000111000101000_1010100111011110"; -- 0.0553079764918376
	pesos_i(6103) := b"0000000000000000_0000000000000000_0011010000100000_1011100101110100"; -- 0.20362433501934518
	pesos_i(6104) := b"1111111111111111_1111111111111111_1101100000000011_0000101011100000"; -- -0.1562035753828788
	pesos_i(6105) := b"1111111111111111_1111111111111111_1110010110000010_1000110001000010"; -- -0.10347674745743596
	pesos_i(6106) := b"1111111111111111_1111111111111111_1111101110110011_0010010010011010"; -- -0.01679774517101418
	pesos_i(6107) := b"0000000000000000_0000000000000000_0000111100100010_0000100100001100"; -- 0.05911308807362572
	pesos_i(6108) := b"0000000000000000_0000000000000000_0000111001110111_0101010111011111"; -- 0.05650841409907404
	pesos_i(6109) := b"0000000000000000_0000000000000000_0000111001011111_1110110101111000"; -- 0.056151239269213386
	pesos_i(6110) := b"0000000000000000_0000000000000000_0010010111011100_0111011101011001"; -- 0.1478952973775536
	pesos_i(6111) := b"0000000000000000_0000000000000000_0010101111111001_0001011000111111"; -- 0.17176951437508473
	pesos_i(6112) := b"0000000000000000_0000000000000000_0000011001110111_0000010010010001"; -- 0.025253568085902567
	pesos_i(6113) := b"0000000000000000_0000000000000000_0010000001000011_0000011111111100"; -- 0.12602281487824596
	pesos_i(6114) := b"1111111111111111_1111111111111111_1110110111010111_1011101111100111"; -- -0.07092691041181629
	pesos_i(6115) := b"1111111111111111_1111111111111111_1111010010001010_1000011111101111"; -- -0.044761184938204884
	pesos_i(6116) := b"0000000000000000_0000000000000000_0000001011100000_0100011011111000"; -- 0.011234698721336913
	pesos_i(6117) := b"1111111111111111_1111111111111111_1110111100001111_1011110110111010"; -- -0.06616605967233238
	pesos_i(6118) := b"1111111111111111_1111111111111111_1110100111010001_1001000101011110"; -- -0.08664599857345996
	pesos_i(6119) := b"0000000000000000_0000000000000000_0001101100011001_0111000010010110"; -- 0.10585693028467788
	pesos_i(6120) := b"0000000000000000_0000000000000000_0010100100101010_1101111001001011"; -- 0.16081036880783703
	pesos_i(6121) := b"1111111111111111_1111111111111111_1110011001001111_0110110000111001"; -- -0.1003506051068889
	pesos_i(6122) := b"1111111111111111_1111111111111111_1100111111001000_0101110111010110"; -- -0.1883488991700622
	pesos_i(6123) := b"0000000000000000_0000000000000000_0000011001101011_0111101011101110"; -- 0.025077517502650068
	pesos_i(6124) := b"1111111111111111_1111111111111111_1111111000100101_1111001000000111"; -- -0.007233498873206428
	pesos_i(6125) := b"0000000000000000_0000000000000000_0000100001100101_0000010100011111"; -- 0.0327914429265203
	pesos_i(6126) := b"1111111111111111_1111111111111111_1111011011101110_1111101101110110"; -- -0.03541591999503265
	pesos_i(6127) := b"0000000000000000_0000000000000000_0001101011100011_1000001010100010"; -- 0.10503403142981832
	pesos_i(6128) := b"1111111111111111_1111111111111111_1101010110100001_0001011001010101"; -- -0.16551075378804295
	pesos_i(6129) := b"1111111111111111_1111111111111111_1101010010010101_0010001110110001"; -- -0.16959931305857104
	pesos_i(6130) := b"1111111111111111_1111111111111111_1101111010010000_1101111111001100"; -- -0.13060189497294336
	pesos_i(6131) := b"0000000000000000_0000000000000000_0000101101010110_0010000001000011"; -- 0.04428292886622528
	pesos_i(6132) := b"1111111111111111_1111111111111111_1110101110100001_1110111010110000"; -- -0.07956035796871787
	pesos_i(6133) := b"1111111111111111_1111111111111111_1110001000010111_1011001011010110"; -- -0.11682588846785329
	pesos_i(6134) := b"0000000000000000_0000000000000000_0010100000000111_1011111111100001"; -- 0.15636824842776886
	pesos_i(6135) := b"0000000000000000_0000000000000000_0010111110100110_1110000101100111"; -- 0.18614014393299164
	pesos_i(6136) := b"1111111111111111_1111111111111111_1110000100110110_0010111000011111"; -- -0.12026702626232716
	pesos_i(6137) := b"1111111111111111_1111111111111111_1101110010011000_0010101010111001"; -- -0.13830311749154228
	pesos_i(6138) := b"1111111111111111_1111111111111111_1111110100011010_0011010100100000"; -- -0.011318854958343219
	pesos_i(6139) := b"0000000000000000_0000000000000000_0000000001101001_0101010110010010"; -- 0.001607273158269274
	pesos_i(6140) := b"0000000000000000_0000000000000000_0010110001111001_0010110110011011"; -- 0.17372403185211538
	pesos_i(6141) := b"0000000000000000_0000000000000000_0010100011101111_0010101111100111"; -- 0.15989946738011598
	pesos_i(6142) := b"1111111111111111_1111111111111111_1110000100011110_1000011011000110"; -- -0.1206279532878545
	pesos_i(6143) := b"1111111111111111_1111111111111111_1110111011111110_0011110101011111"; -- -0.0664331096484965
	pesos_i(6144) := b"0000000000000000_0000000000000000_0000001111001100_1110100010000100"; -- 0.014845402028003052
	pesos_i(6145) := b"0000000000000000_0000000000000000_0001101011110101_1110111000100001"; -- 0.1053150970114295
	pesos_i(6146) := b"1111111111111111_1111111111111111_1101110001010111_1100111000000100"; -- -0.13928520590388482
	pesos_i(6147) := b"1111111111111111_1111111111111111_1110010000011001_0010111000000000"; -- -0.10899078836245209
	pesos_i(6148) := b"0000000000000000_0000000000000000_0001011011110010_1110001100101010"; -- 0.0896436670255256
	pesos_i(6149) := b"0000000000000000_0000000000000000_0001110011011110_1100111110010010"; -- 0.112774823298275
	pesos_i(6150) := b"0000000000000000_0000000000000000_0000011011111000_0011110111011111"; -- 0.0272253674562347
	pesos_i(6151) := b"0000000000000000_0000000000000000_0010010000001100_0000011001100110"; -- 0.140808486805865
	pesos_i(6152) := b"0000000000000000_0000000000000000_0010111010101111_0110011101010110"; -- 0.18236394733190875
	pesos_i(6153) := b"0000000000000000_0000000000000000_0000111100001101_0100011011110001"; -- 0.058796342705817184
	pesos_i(6154) := b"0000000000000000_0000000000000000_0001010111110001_0011010000111010"; -- 0.08571173118135593
	pesos_i(6155) := b"0000000000000000_0000000000000000_0001101010110011_1010000100011011"; -- 0.10430342583720265
	pesos_i(6156) := b"1111111111111111_1111111111111111_1110001010100101_1001111111000010"; -- -0.11466027756768238
	pesos_i(6157) := b"1111111111111111_1111111111111111_1111100111001000_1001101010101011"; -- -0.024282773343182764
	pesos_i(6158) := b"0000000000000000_0000000000000000_0000000010011110_0010110011001111"; -- 0.0024135595181990076
	pesos_i(6159) := b"1111111111111111_1111111111111111_1111010100111100_0000110111010010"; -- -0.04205239887895036
	pesos_i(6160) := b"0000000000000000_0000000000000000_0010011011110001_0100010000011111"; -- 0.15211892852885248
	pesos_i(6161) := b"0000000000000000_0000000000000000_0001000101000111_1110011101111000"; -- 0.06750342056464281
	pesos_i(6162) := b"0000000000000000_0000000000000000_0010100100101101_0000111110100000"; -- 0.1608438268965561
	pesos_i(6163) := b"1111111111111111_1111111111111111_1101001111111110_0111101100001011"; -- -0.1718981837440287
	pesos_i(6164) := b"0000000000000000_0000000000000000_0000100000101001_1101011001100100"; -- 0.031888389123873644
	pesos_i(6165) := b"1111111111111111_1111111111111111_1110011010111110_1011001101001010"; -- -0.09865264358144757
	pesos_i(6166) := b"0000000000000000_0000000000000000_0000001111000110_0001011001110001"; -- 0.014741327915768333
	pesos_i(6167) := b"1111111111111111_1111111111111111_1110001010100110_0010000010001100"; -- -0.11465260096624204
	pesos_i(6168) := b"0000000000000000_0000000000000000_0000011010010000_1011101000111100"; -- 0.025645866023168314
	pesos_i(6169) := b"0000000000000000_0000000000000000_0010000100011000_1101011111000100"; -- 0.1292853215442168
	pesos_i(6170) := b"0000000000000000_0000000000000000_0000100000000111_0101001101101000"; -- 0.031361782996982716
	pesos_i(6171) := b"1111111111111111_1111111111111111_1110011000110011_1001100100010001"; -- -0.10077517824565772
	pesos_i(6172) := b"0000000000000000_0000000000000000_0001101110010010_0111001011100010"; -- 0.10770338078736666
	pesos_i(6173) := b"0000000000000000_0000000000000000_0001110101111110_0000101000111100"; -- 0.11520446737026079
	pesos_i(6174) := b"1111111111111111_1111111111111111_1110000101011110_1100001001100010"; -- -0.11964783760780061
	pesos_i(6175) := b"0000000000000000_0000000000000000_0000010111100111_0101001011001111"; -- 0.023060966141205647
	pesos_i(6176) := b"1111111111111111_1111111111111111_1101010101000000_1100010001010101"; -- -0.16698048517868494
	pesos_i(6177) := b"0000000000000000_0000000000000000_0000101111000011_1010100101110111"; -- 0.045954314765354796
	pesos_i(6178) := b"1111111111111111_1111111111111111_1110010000111000_1000001001000011"; -- -0.1085127437068985
	pesos_i(6179) := b"1111111111111111_1111111111111111_1111010100011100_1110110010111101"; -- -0.042527393315021034
	pesos_i(6180) := b"1111111111111111_1111111111111111_1110110001110011_0100011111010001"; -- -0.0763659586658278
	pesos_i(6181) := b"0000000000000000_0000000000000000_0000110111111111_1101010100100011"; -- 0.05468494513286405
	pesos_i(6182) := b"1111111111111111_1111111111111111_1111101101101111_0010110110111010"; -- -0.0178347989792054
	pesos_i(6183) := b"1111111111111111_1111111111111111_1111010110110001_0110101011111100"; -- -0.040261567468350856
	pesos_i(6184) := b"1111111111111111_1111111111111111_1110101001001001_1111011101000110"; -- -0.08480886977757257
	pesos_i(6185) := b"1111111111111111_1111111111111111_1101111101110101_0011110110000111"; -- -0.12711730445952057
	pesos_i(6186) := b"0000000000000000_0000000000000000_0000010101000101_1110110011000100"; -- 0.02059821866163068
	pesos_i(6187) := b"1111111111111111_1111111111111111_1110011011110101_0000111110010000"; -- -0.0978231689933031
	pesos_i(6188) := b"0000000000000000_0000000000000000_0000111001101110_0011110001110001"; -- 0.05636956932892481
	pesos_i(6189) := b"0000000000000000_0000000000000000_0000010110111111_0010101101100011"; -- 0.022448264660276003
	pesos_i(6190) := b"0000000000000000_0000000000000000_0010000011110110_0101100011111101"; -- 0.12875896630863345
	pesos_i(6191) := b"1111111111111111_1111111111111111_1101111010011100_0000100110110010"; -- -0.13043155098147505
	pesos_i(6192) := b"0000000000000000_0000000000000000_0001001000111100_0011011010110101"; -- 0.07123128814526469
	pesos_i(6193) := b"0000000000000000_0000000000000000_0001011110100000_0100000100101011"; -- 0.09228904058465272
	pesos_i(6194) := b"1111111111111111_1111111111111111_1110101100100101_0111000101000011"; -- -0.08145992392908263
	pesos_i(6195) := b"0000000000000000_0000000000000000_0010000100010100_0010000000000111"; -- 0.12921333473620805
	pesos_i(6196) := b"1111111111111111_1111111111111111_1111101001110101_1100010001000001"; -- -0.02164052410286511
	pesos_i(6197) := b"1111111111111111_1111111111111111_1101110100100011_1011000000100011"; -- -0.13617419373512735
	pesos_i(6198) := b"1111111111111111_1111111111111111_1110011110100111_1011110100011010"; -- -0.09509676093931191
	pesos_i(6199) := b"1111111111111111_1111111111111111_1101011000010101_1011001011100001"; -- -0.16373140332861105
	pesos_i(6200) := b"1111111111111111_1111111111111111_1110000101111101_0101100000101100"; -- -0.11918114581113248
	pesos_i(6201) := b"1111111111111111_1111111111111111_1111011000010101_1110001000110101"; -- -0.03872858244240478
	pesos_i(6202) := b"0000000000000000_0000000000000000_0001000111010011_0011110110100000"; -- 0.06962952770999649
	pesos_i(6203) := b"0000000000000000_0000000000000000_0001010010101000_0100101110110110"; -- 0.08069298925362522
	pesos_i(6204) := b"1111111111111111_1111111111111111_1110000111010011_0100110100111110"; -- -0.1178695414551017
	pesos_i(6205) := b"1111111111111111_1111111111111111_1101110001001001_1011001000011000"; -- -0.13950049314600949
	pesos_i(6206) := b"1111111111111111_1111111111111111_1111001111101100_1010010110010100"; -- -0.047170306450221564
	pesos_i(6207) := b"0000000000000000_0000000000000000_0000010101010100_1010111110100010"; -- 0.020823456881770928
	pesos_i(6208) := b"1111111111111111_1111111111111111_1101010100100100_1000011110111111"; -- -0.1674113423947027
	pesos_i(6209) := b"0000000000000000_0000000000000000_0010010110111111_1110011100101000"; -- 0.14745945680797837
	pesos_i(6210) := b"1111111111111111_1111111111111111_1111111000000010_1000100100010111"; -- -0.00777381118643296
	pesos_i(6211) := b"0000000000000000_0000000000000000_0000100100110101_1011000101111011"; -- 0.0359755444117985
	pesos_i(6212) := b"0000000000000000_0000000000000000_0010000011111111_0010000011100111"; -- 0.12889295242136833
	pesos_i(6213) := b"1111111111111111_1111111111111111_1101111110000011_0000000000101110"; -- -0.12690733782967364
	pesos_i(6214) := b"0000000000000000_0000000000000000_0000110010001101_1000001111100011"; -- 0.049034350273348744
	pesos_i(6215) := b"1111111111111111_1111111111111111_1111101001100010_0001010001100101"; -- -0.021940923038897296
	pesos_i(6216) := b"0000000000000000_0000000000000000_0011001101111101_1101011001000111"; -- 0.20113887064405006
	pesos_i(6217) := b"1111111111111111_1111111111111111_1111000100011000_0011101001001111"; -- -0.05822406357276655
	pesos_i(6218) := b"1111111111111111_1111111111111111_1110110011000011_0001011110101010"; -- -0.07514812569459614
	pesos_i(6219) := b"1111111111111111_1111111111111111_1111010001010101_0010101111101100"; -- -0.045575385003155645
	pesos_i(6220) := b"1111111111111111_1111111111111111_1110110010101100_0101101111001011"; -- -0.07549501703469921
	pesos_i(6221) := b"1111111111111111_1111111111111111_1111000011110111_1100100111101100"; -- -0.058719043721434896
	pesos_i(6222) := b"0000000000000000_0000000000000000_0001000011011001_0011110000000000"; -- 0.06581473357504079
	pesos_i(6223) := b"1111111111111111_1111111111111111_1101100001001011_0101110101110110"; -- -0.15510002020532787
	pesos_i(6224) := b"0000000000000000_0000000000000000_0010011111111001_0100010101101010"; -- 0.15614732588837768
	pesos_i(6225) := b"1111111111111111_1111111111111111_1101110000111101_1111100100011110"; -- -0.13967936536918935
	pesos_i(6226) := b"0000000000000000_0000000000000000_0000100010011101_1000000011100001"; -- 0.033653311755965795
	pesos_i(6227) := b"0000000000000000_0000000000000000_0001000001111011_0111001100011010"; -- 0.06438369166768657
	pesos_i(6228) := b"1111111111111111_1111111111111111_1110101001110001_0101001111111000"; -- -0.0842082519228667
	pesos_i(6229) := b"1111111111111111_1111111111111111_1111100011001101_1110010110001101"; -- -0.02810826593203745
	pesos_i(6230) := b"0000000000000000_0000000000000000_0000001011101011_0101000110010110"; -- 0.011403178409770249
	pesos_i(6231) := b"0000000000000000_0000000000000000_0010001011011110_1110000110011110"; -- 0.13621339893993942
	pesos_i(6232) := b"0000000000000000_0000000000000000_0001000111010000_0100001010100001"; -- 0.06958404941378563
	pesos_i(6233) := b"0000000000000000_0000000000000000_0001110100101001_1001000001000001"; -- 0.113915458490862
	pesos_i(6234) := b"1111111111111111_1111111111111111_1111110011101001_0111000101111000"; -- -0.012062938851889301
	pesos_i(6235) := b"1111111111111111_1111111111111111_1111000010110000_0011101101100101"; -- -0.05981091293489679
	pesos_i(6236) := b"1111111111111111_1111111111111111_1101110101010101_1100000111101101"; -- -0.135410194138669
	pesos_i(6237) := b"0000000000000000_0000000000000000_0000011001111000_1100100100110000"; -- 0.025280546397133043
	pesos_i(6238) := b"1111111111111111_1111111111111111_1110101110100001_1110100001011000"; -- -0.07956073609124192
	pesos_i(6239) := b"1111111111111111_1111111111111111_1101110100111011_0101010011000110"; -- -0.1358134285969413
	pesos_i(6240) := b"1111111111111111_1111111111111111_1111001110111011_0111111101111100"; -- -0.047920257813736405
	pesos_i(6241) := b"1111111111111111_1111111111111111_1111101000110110_1011101111100010"; -- -0.022602326666008955
	pesos_i(6242) := b"1111111111111111_1111111111111111_1111010000011111_1101000111001100"; -- -0.046389472662830014
	pesos_i(6243) := b"0000000000000000_0000000000000000_0010001110110100_0010011011111111"; -- 0.13946765647932388
	pesos_i(6244) := b"0000000000000000_0000000000000000_0000111100011101_1101101100110010"; -- 0.05904931989441815
	pesos_i(6245) := b"0000000000000000_0000000000000000_0001010100010000_1010000000011000"; -- 0.08228493289989272
	pesos_i(6246) := b"1111111111111111_1111111111111111_1111110111001000_0111000111101111"; -- -0.008660201216403937
	pesos_i(6247) := b"0000000000000000_0000000000000000_0010101101000110_1010001110100010"; -- 0.16904661851004785
	pesos_i(6248) := b"0000000000000000_0000000000000000_0010100010010000_0100011101110011"; -- 0.1584515242751077
	pesos_i(6249) := b"0000000000000000_0000000000000000_0010001110011100_0101011100110100"; -- 0.13910431889366526
	pesos_i(6250) := b"0000000000000000_0000000000000000_0010011101111001_1011011010101001"; -- 0.15420095081050317
	pesos_i(6251) := b"1111111111111111_1111111111111111_1110011011110010_0111001110010111"; -- -0.09786298345997436
	pesos_i(6252) := b"0000000000000000_0000000000000000_0010000001001001_1000101100001011"; -- 0.12612217912502588
	pesos_i(6253) := b"0000000000000000_0000000000000000_0001110110110111_0100100110010011"; -- 0.11607799379152413
	pesos_i(6254) := b"1111111111111111_1111111111111111_1101010111010101_1101010011100001"; -- -0.16470593946121395
	pesos_i(6255) := b"0000000000000000_0000000000000000_0000111000000011_0111110011000110"; -- 0.05474071346804993
	pesos_i(6256) := b"1111111111111111_1111111111111111_1111001010001001_0101101000100001"; -- -0.05259167382112444
	pesos_i(6257) := b"1111111111111111_1111111111111111_1110101101000010_0011000100010111"; -- -0.08102124396033401
	pesos_i(6258) := b"0000000000000000_0000000000000000_0000000100010010_1111100000100011"; -- 0.004195698352307222
	pesos_i(6259) := b"1111111111111111_1111111111111111_1110001110010110_0001101001100100"; -- -0.11099085854286703
	pesos_i(6260) := b"1111111111111111_1111111111111111_1111000111011001_0001110101101101"; -- -0.05528083885844586
	pesos_i(6261) := b"0000000000000000_0000000000000000_0010101100101110_0111101111011011"; -- 0.16867803670778322
	pesos_i(6262) := b"0000000000000000_0000000000000000_0001010101011010_1010001010111111"; -- 0.08341424153078215
	pesos_i(6263) := b"1111111111111111_1111111111111111_1101101001111100_1011000011000011"; -- -0.14653487429060869
	pesos_i(6264) := b"1111111111111111_1111111111111111_1111011111011111_1111101011010111"; -- -0.031738588756078545
	pesos_i(6265) := b"1111111111111111_1111111111111111_1110010011110010_1111110011101110"; -- -0.10566729729348537
	pesos_i(6266) := b"0000000000000000_0000000000000000_0001100011000100_0100001110000001"; -- 0.09674474611721848
	pesos_i(6267) := b"1111111111111111_1111111111111111_1110001100001110_0110111110110011"; -- -0.11306096908386921
	pesos_i(6268) := b"1111111111111111_1111111111111111_1111011011111000_1110100101110000"; -- -0.03526440626711821
	pesos_i(6269) := b"0000000000000000_0000000000000000_0010001100111110_0100001011110100"; -- 0.1376687855318232
	pesos_i(6270) := b"1111111111111111_1111111111111111_1101011011101011_0000011010100111"; -- -0.1604762880087976
	pesos_i(6271) := b"0000000000000000_0000000000000000_0000010010000001_0001111111001111"; -- 0.017595279810053686
	pesos_i(6272) := b"0000000000000000_0000000000000000_0000001111110000_1111101000010111"; -- 0.015395765838610798
	pesos_i(6273) := b"0000000000000000_0000000000000000_0010000000000111_0011001001000110"; -- 0.12510980799394344
	pesos_i(6274) := b"1111111111111111_1111111111111111_1110101111001001_1001010111100000"; -- -0.07895530023299145
	pesos_i(6275) := b"1111111111111111_1111111111111111_1110101001001110_0010000110111101"; -- -0.08474530345104088
	pesos_i(6276) := b"1111111111111111_1111111111111111_1101010101010001_0100000101011010"; -- -0.16672889280683628
	pesos_i(6277) := b"1111111111111111_1111111111111111_1110011010000010_0111001111100011"; -- -0.09957195009743612
	pesos_i(6278) := b"1111111111111111_1111111111111111_1110011100001100_0111111111100000"; -- -0.09746552266071334
	pesos_i(6279) := b"0000000000000000_0000000000000000_0001011001001110_0111000110110100"; -- 0.08713446271847888
	pesos_i(6280) := b"0000000000000000_0000000000000000_0000101011001000_0111111110111011"; -- 0.04212187106081642
	pesos_i(6281) := b"0000000000000000_0000000000000000_0010010000011101_0000111000011000"; -- 0.14106834484344694
	pesos_i(6282) := b"0000000000000000_0000000000000000_0000111111001110_1110001101011000"; -- 0.0617506112627785
	pesos_i(6283) := b"1111111111111111_1111111111111111_1110111101000010_1010001011101111"; -- -0.06538945825040518
	pesos_i(6284) := b"0000000000000000_0000000000000000_0000111010010000_1001110011110110"; -- 0.056894121187540246
	pesos_i(6285) := b"0000000000000000_0000000000000000_0001111100010000_1110011001110101"; -- 0.1213516269393833
	pesos_i(6286) := b"1111111111111111_1111111111111111_1111101011101001_0010010001100100"; -- -0.019880033047594295
	pesos_i(6287) := b"0000000000000000_0000000000000000_0011001111101111_1011000010010011"; -- 0.20287612524960422
	pesos_i(6288) := b"1111111111111111_1111111111111111_1110001101111010_0100010001101110"; -- -0.11141559890117489
	pesos_i(6289) := b"1111111111111111_1111111111111111_1111111001110011_0001001001111111"; -- -0.006056636827787033
	pesos_i(6290) := b"1111111111111111_1111111111111111_1111111000001100_1010011110001000"; -- -0.007619408793228819
	pesos_i(6291) := b"0000000000000000_0000000000000000_0010101010101111_1100010110011110"; -- 0.16674456687216477
	pesos_i(6292) := b"0000000000000000_0000000000000000_0001100111011001_1110111010100001"; -- 0.10098163069065134
	pesos_i(6293) := b"0000000000000000_0000000000000000_0010010011101111_0011010010011110"; -- 0.14427498670385833
	pesos_i(6294) := b"1111111111111111_1111111111111111_1110110100000011_0110110000010011"; -- -0.07416653199004963
	pesos_i(6295) := b"1111111111111111_1111111111111111_1110001000111010_0101011110111100"; -- -0.11629726094184176
	pesos_i(6296) := b"0000000000000000_0000000000000000_0010011110000101_0010011011001111"; -- 0.1543754820358234
	pesos_i(6297) := b"1111111111111111_1111111111111111_1111011000011010_0101010010001000"; -- -0.0386607329399448
	pesos_i(6298) := b"0000000000000000_0000000000000000_0001001100110011_0100100110110111"; -- 0.07500134190285333
	pesos_i(6299) := b"1111111111111111_1111111111111111_1111010000100111_0110100110000000"; -- -0.046273618942588066
	pesos_i(6300) := b"0000000000000000_0000000000000000_0000011100000101_0111001001100110"; -- 0.02742686267730627
	pesos_i(6301) := b"1111111111111111_1111111111111111_1110000000110011_0101111001101011"; -- -0.12421617399830456
	pesos_i(6302) := b"0000000000000000_0000000000000000_0000111010001101_1000101001001010"; -- 0.056847231910052705
	pesos_i(6303) := b"0000000000000000_0000000000000000_0001010001010101_0011010011101011"; -- 0.07942515118231533
	pesos_i(6304) := b"1111111111111111_1111111111111111_1110111101000100_1100000100001000"; -- -0.06535714669576385
	pesos_i(6305) := b"1111111111111111_1111111111111111_1111001001110001_0001001100110001"; -- -0.052962112977026674
	pesos_i(6306) := b"0000000000000000_0000000000000000_0010011101000011_0100011001010000"; -- 0.15337027973884534
	pesos_i(6307) := b"0000000000000000_0000000000000000_0001001001001111_1010000100100011"; -- 0.07152754883312086
	pesos_i(6308) := b"0000000000000000_0000000000000000_0000100110001001_0101100000001010"; -- 0.03725195164129146
	pesos_i(6309) := b"0000000000000000_0000000000000000_0001010001001001_0101011011110100"; -- 0.0792440743856195
	pesos_i(6310) := b"1111111111111111_1111111111111111_1110001111110100_1010000001000001"; -- -0.10954855357848595
	pesos_i(6311) := b"1111111111111111_1111111111111111_1101011111000011_1101111001100010"; -- -0.15716753107410472
	pesos_i(6312) := b"1111111111111111_1111111111111111_1101100100001101_1011001001111000"; -- -0.15213474820814868
	pesos_i(6313) := b"0000000000000000_0000000000000000_0000110100011010_1011101011101101"; -- 0.051189120049938794
	pesos_i(6314) := b"1111111111111111_1111111111111111_1111101000000101_0011110101101110"; -- -0.02335754465078727
	pesos_i(6315) := b"1111111111111111_1111111111111111_1111101001101101_0001001101010010"; -- -0.021773140359547114
	pesos_i(6316) := b"1111111111111111_1111111111111111_1101100000100101_1000101110010011"; -- -0.15567710542551996
	pesos_i(6317) := b"0000000000000000_0000000000000000_0001000101101111_1000011011011101"; -- 0.06810801409650014
	pesos_i(6318) := b"1111111111111111_1111111111111111_1111100110000000_0001011000001011"; -- -0.025389311170252997
	pesos_i(6319) := b"0000000000000000_0000000000000000_0001001010011001_0110111101010011"; -- 0.07265373008840602
	pesos_i(6320) := b"1111111111111111_1111111111111111_1110011011011110_0000100100010000"; -- -0.098174508695349
	pesos_i(6321) := b"0000000000000000_0000000000000000_0010001101101001_0010110110000100"; -- 0.13832363585590446
	pesos_i(6322) := b"0000000000000000_0000000000000000_0000110101011001_1011001111010100"; -- 0.05215000087179421
	pesos_i(6323) := b"1111111111111111_1111111111111111_1101100010111111_1000110010000000"; -- -0.15332719693523156
	pesos_i(6324) := b"0000000000000000_0000000000000000_0010010011010011_1100010100101010"; -- 0.14385635627283175
	pesos_i(6325) := b"0000000000000000_0000000000000000_0000000010110010_0111111010110111"; -- 0.0027236173019695776
	pesos_i(6326) := b"0000000000000000_0000000000000000_0000111101100100_0010000101111000"; -- 0.0601216237220516
	pesos_i(6327) := b"0000000000000000_0000000000000000_0001010011111111_1101100100110010"; -- 0.08202893704879367
	pesos_i(6328) := b"0000000000000000_0000000000000000_0000101101101110_1110000111011001"; -- 0.04466067833752774
	pesos_i(6329) := b"1111111111111111_1111111111111111_1110001010001111_0000111001010110"; -- -0.11500463876257488
	pesos_i(6330) := b"0000000000000000_0000000000000000_0010000011101101_1000101000110111"; -- 0.12862457132411925
	pesos_i(6331) := b"0000000000000000_0000000000000000_0000100001001100_1110001110010100"; -- 0.03242323273631001
	pesos_i(6332) := b"1111111111111111_1111111111111111_1110100011011011_1111110010000011"; -- -0.09039327443875565
	pesos_i(6333) := b"0000000000000000_0000000000000000_0001111010100001_0000011010001100"; -- 0.1196445551730935
	pesos_i(6334) := b"1111111111111111_1111111111111111_1111010100001010_0010000110001111"; -- -0.0428141619649319
	pesos_i(6335) := b"0000000000000000_0000000000000000_0000100010011111_0010101000100110"; -- 0.0336786596155574
	pesos_i(6336) := b"1111111111111111_1111111111111111_1110101101001110_0110111011010010"; -- -0.08083445907088002
	pesos_i(6337) := b"0000000000000000_0000000000000000_0001000000010110_1101101011101001"; -- 0.06284874152654114
	pesos_i(6338) := b"0000000000000000_0000000000000000_0000101010010000_0001001111000001"; -- 0.041260943152588256
	pesos_i(6339) := b"1111111111111111_1111111111111111_1101100111000111_0101110011110111"; -- -0.14930170992605402
	pesos_i(6340) := b"0000000000000000_0000000000000000_0000110000011000_0111111001010110"; -- 0.04724874116556135
	pesos_i(6341) := b"1111111111111111_1111111111111111_1111110110000011_1110000100011001"; -- -0.009706431851022743
	pesos_i(6342) := b"0000000000000000_0000000000000000_0010011010001011_1101111011010111"; -- 0.15057175396716568
	pesos_i(6343) := b"0000000000000000_0000000000000000_0000000100011011_1100101111010110"; -- 0.004330386935938057
	pesos_i(6344) := b"1111111111111111_1111111111111111_1111000000010101_1000100001110100"; -- -0.0621714322611894
	pesos_i(6345) := b"1111111111111111_1111111111111111_1111001101111011_0100110111000010"; -- -0.04889978424034993
	pesos_i(6346) := b"1111111111111111_1111111111111111_1110111001010101_1001000000010111"; -- -0.06900691439258817
	pesos_i(6347) := b"0000000000000000_0000000000000000_0000000111000100_1111011010101011"; -- 0.0069116752402535505
	pesos_i(6348) := b"1111111111111111_1111111111111111_1101101111011110_0011001101010110"; -- -0.14114073906910543
	pesos_i(6349) := b"1111111111111111_1111111111111111_1110000010011101_0001111001101101"; -- -0.12260255653281792
	pesos_i(6350) := b"0000000000000000_0000000000000000_0010010111100000_1001111000111000"; -- 0.14795864932944885
	pesos_i(6351) := b"1111111111111111_1111111111111111_1110001110000000_1001111101101001"; -- -0.11131862337452027
	pesos_i(6352) := b"0000000000000000_0000000000000000_0010010100100001_1011100010000100"; -- 0.14504578805231474
	pesos_i(6353) := b"1111111111111111_1111111111111111_1110001101110110_0111011000110100"; -- -0.11147366739959666
	pesos_i(6354) := b"1111111111111111_1111111111111111_1110000001110000_1011110001011010"; -- -0.12327978899145885
	pesos_i(6355) := b"0000000000000000_0000000000000000_0010100110111110_1111111111010111"; -- 0.163070669252306
	pesos_i(6356) := b"1111111111111111_1111111111111111_1111100111101010_0010011100100011"; -- -0.023770860556198
	pesos_i(6357) := b"0000000000000000_0000000000000000_0010101101001001_0100011101001001"; -- 0.16908689060357102
	pesos_i(6358) := b"1111111111111111_1111111111111111_1110011001010010_1111011001010110"; -- -0.10029659643727729
	pesos_i(6359) := b"0000000000000000_0000000000000000_0000111011000110_0110000010101100"; -- 0.057714502428191344
	pesos_i(6360) := b"1111111111111111_1111111111111111_1111110011101100_0100001011011010"; -- -0.012019941200298962
	pesos_i(6361) := b"0000000000000000_0000000000000000_0010001101010111_0101000001100000"; -- 0.13805105540451582
	pesos_i(6362) := b"1111111111111111_1111111111111111_1101011111101010_0110000000110101"; -- -0.15657995904461108
	pesos_i(6363) := b"1111111111111111_1111111111111111_1111110011110111_1001000010001101"; -- -0.011847463245133248
	pesos_i(6364) := b"1111111111111111_1111111111111111_1111110110000000_0001010001000101"; -- -0.009764416762197584
	pesos_i(6365) := b"1111111111111111_1111111111111111_1101110101100000_0011110010000001"; -- -0.13525029985185272
	pesos_i(6366) := b"1111111111111111_1111111111111111_1110101011100111_1111010111111100"; -- -0.08239805790673273
	pesos_i(6367) := b"0000000000000000_0000000000000000_0000110100101011_0110011100100011"; -- 0.051443525439092114
	pesos_i(6368) := b"0000000000000000_0000000000000000_0010001010100100_1000101110001000"; -- 0.13532325821411026
	pesos_i(6369) := b"1111111111111111_1111111111111111_1101100110011011_1010010111111011"; -- -0.14996874449936068
	pesos_i(6370) := b"0000000000000000_0000000000000000_0000111111100101_1101011000000101"; -- 0.06210076934905064
	pesos_i(6371) := b"1111111111111111_1111111111111111_1110110110011101_0000011111010000"; -- -0.07182265446794747
	pesos_i(6372) := b"1111111111111111_1111111111111111_1101011100001111_1000011001011010"; -- -0.15991936015624025
	pesos_i(6373) := b"1111111111111111_1111111111111111_1111111110000001_0100011001010000"; -- -0.0019336751856528006
	pesos_i(6374) := b"0000000000000000_0000000000000000_0000010011000011_0001101110011111"; -- 0.018602110100377395
	pesos_i(6375) := b"0000000000000000_0000000000000000_0010010011011111_0110011010101110"; -- 0.1440338302545651
	pesos_i(6376) := b"0000000000000000_0000000000000000_0010001101010101_1110100110110000"; -- 0.13802967590695878
	pesos_i(6377) := b"1111111111111111_1111111111111111_1110001000101100_0000011010110111"; -- -0.11651571314866561
	pesos_i(6378) := b"0000000000000000_0000000000000000_0000000100001101_1001010000010110"; -- 0.004113440913754388
	pesos_i(6379) := b"1111111111111111_1111111111111111_1111111110001000_1000111101110010"; -- -0.0018225047792389411
	pesos_i(6380) := b"1111111111111111_1111111111111111_1110010000111111_0100000001110010"; -- -0.10840985494740127
	pesos_i(6381) := b"0000000000000000_0000000000000000_0000111101100101_0110001000110001"; -- 0.06014074037610461
	pesos_i(6382) := b"0000000000000000_0000000000000000_0001000111110110_1101101111010110"; -- 0.07017301546747777
	pesos_i(6383) := b"0000000000000000_0000000000000000_0000100111001010_1000101100001110"; -- 0.038246813650569235
	pesos_i(6384) := b"0000000000000000_0000000000000000_0001000000101111_1001000111011011"; -- 0.06322585678128331
	pesos_i(6385) := b"1111111111111111_1111111111111111_1111001110110000_1001100010000101"; -- -0.04808661225926918
	pesos_i(6386) := b"1111111111111111_1111111111111111_1111100101110011_0001111111011100"; -- -0.0255870903285447
	pesos_i(6387) := b"0000000000000000_0000000000000000_0000101000100001_0100011100110101"; -- 0.03957028431147687
	pesos_i(6388) := b"0000000000000000_0000000000000000_0001100111111000_0100101001100100"; -- 0.10144486375961245
	pesos_i(6389) := b"0000000000000000_0000000000000000_0000111001110100_0000000100011011"; -- 0.05645758531668357
	pesos_i(6390) := b"1111111111111111_1111111111111111_1110001110011010_0101111010100010"; -- -0.11092575590256934
	pesos_i(6391) := b"1111111111111111_1111111111111111_1110000000011011_0111101000110010"; -- -0.12458072929159288
	pesos_i(6392) := b"0000000000000000_0000000000000000_0000111110110101_1001101000110101"; -- 0.061364782172193655
	pesos_i(6393) := b"1111111111111111_1111111111111111_1111011111010100_1001010111111110"; -- -0.03191244652511939
	pesos_i(6394) := b"1111111111111111_1111111111111111_1110110010100100_0100001110111110"; -- -0.07561852093642003
	pesos_i(6395) := b"0000000000000000_0000000000000000_0000000000010010_0100100100001000"; -- 0.00027901110590366953
	pesos_i(6396) := b"0000000000000000_0000000000000000_0010010111010001_1010010110110101"; -- 0.14773021384759114
	pesos_i(6397) := b"0000000000000000_0000000000000000_0010011101110011_0001101101100100"; -- 0.1541001433210215
	pesos_i(6398) := b"0000000000000000_0000000000000000_0001010010001010_0110111001111110"; -- 0.08023729863308499
	pesos_i(6399) := b"1111111111111111_1111111111111111_1110010011111000_1000111100111001"; -- -0.1055822835252606
	pesos_i(6400) := b"1111111111111111_1111111111111111_1110001100011111_0100000001011110"; -- -0.11280439090999132
	pesos_i(6401) := b"0000000000000000_0000000000000000_0001011011100011_1111000000010110"; -- 0.08941555527978358
	pesos_i(6402) := b"0000000000000000_0000000000000000_0010100101101100_1110011110000010"; -- 0.16181799816847403
	pesos_i(6403) := b"0000000000000000_0000000000000000_0000010011110000_0110100100001011"; -- 0.019293370375544284
	pesos_i(6404) := b"0000000000000000_0000000000000000_0000010001010110_0011100100000010"; -- 0.0169406538415959
	pesos_i(6405) := b"0000000000000000_0000000000000000_0001101111000000_1011100001011000"; -- 0.10840942525136915
	pesos_i(6406) := b"1111111111111111_1111111111111111_1111010000101001_0001111010110001"; -- -0.04624756032308063
	pesos_i(6407) := b"0000000000000000_0000000000000000_0000110111011000_0001110001000110"; -- 0.05407883375172727
	pesos_i(6408) := b"1111111111111111_1111111111111111_1111100000000101_1100100010110110"; -- -0.031161742665203856
	pesos_i(6409) := b"1111111111111111_1111111111111111_1110100101101110_1000001110100001"; -- -0.08815743759120126
	pesos_i(6410) := b"1111111111111111_1111111111111111_1101110111110110_1001100001110101"; -- -0.13295600063195112
	pesos_i(6411) := b"1111111111111111_1111111111111111_1110110100110001_0011111001000000"; -- -0.07346735905864923
	pesos_i(6412) := b"0000000000000000_0000000000000000_0000110011001000_1000000100011100"; -- 0.04993445331070982
	pesos_i(6413) := b"1111111111111111_1111111111111111_1111111111101110_0110111111000010"; -- -0.0002679969727515218
	pesos_i(6414) := b"1111111111111111_1111111111111111_1110001110111100_1101110001001011"; -- -0.11039946723944967
	pesos_i(6415) := b"0000000000000000_0000000000000000_0000101100010011_1010010101010111"; -- 0.043268522106155956
	pesos_i(6416) := b"1111111111111111_1111111111111111_1111111011010111_1110100111001110"; -- -0.004517924501894477
	pesos_i(6417) := b"0000000000000000_0000000000000000_0001111010000000_1001000100001001"; -- 0.11914926974890057
	pesos_i(6418) := b"1111111111111111_1111111111111111_1110111000011010_0101100100101000"; -- -0.06991045740113078
	pesos_i(6419) := b"0000000000000000_0000000000000000_0001001000010110_1101101011001011"; -- 0.07066123450208045
	pesos_i(6420) := b"0000000000000000_0000000000000000_0000101101110000_0000010011100000"; -- 0.04467802494607973
	pesos_i(6421) := b"0000000000000000_0000000000000000_0001011011000110_0001111011110000"; -- 0.08896058423646537
	pesos_i(6422) := b"0000000000000000_0000000000000000_0000010010010111_0101100100011111"; -- 0.01793438913419282
	pesos_i(6423) := b"0000000000000000_0000000000000000_0001000111111011_0101110001100100"; -- 0.07024171293355036
	pesos_i(6424) := b"0000000000000000_0000000000000000_0001011011101100_0001010010011100"; -- 0.08953980254386751
	pesos_i(6425) := b"0000000000000000_0000000000000000_0010001111011111_1000010100000100"; -- 0.1401293881964371
	pesos_i(6426) := b"1111111111111111_1111111111111111_1111000001111010_0101010111111010"; -- -0.06063330324631619
	pesos_i(6427) := b"1111111111111111_1111111111111111_1110000001111010_0100110101100010"; -- -0.12313381539829843
	pesos_i(6428) := b"0000000000000000_0000000000000000_0001101010000101_1010110101100011"; -- 0.10360225359637067
	pesos_i(6429) := b"1111111111111111_1111111111111111_1111000001011000_0001001100000111"; -- -0.061156092342129265
	pesos_i(6430) := b"1111111111111111_1111111111111111_1110100101010000_1111010011111011"; -- -0.08860844480380514
	pesos_i(6431) := b"1111111111111111_1111111111111111_1101100010110001_1000111100111100"; -- -0.15354065701224667
	pesos_i(6432) := b"1111111111111111_1111111111111111_1111110011000001_1011001111010011"; -- -0.012669335375701613
	pesos_i(6433) := b"1111111111111111_1111111111111111_1110001110100111_0110000001111001"; -- -0.11072728210569638
	pesos_i(6434) := b"1111111111111111_1111111111111111_1110001111000000_0001101010010011"; -- -0.11034997849192668
	pesos_i(6435) := b"0000000000000000_0000000000000000_0001101010011111_0111111101000000"; -- 0.10399623204102033
	pesos_i(6436) := b"0000000000000000_0000000000000000_0000011110011010_1111111111011100"; -- 0.02970885388101823
	pesos_i(6437) := b"0000000000000000_0000000000000000_0010100001101010_0110111010110110"; -- 0.15787403058786464
	pesos_i(6438) := b"0000000000000000_0000000000000000_0001111110011000_1110111110011001"; -- 0.12342736702744316
	pesos_i(6439) := b"0000000000000000_0000000000000000_0001001010100100_0001111100000110"; -- 0.07281679064346178
	pesos_i(6440) := b"0000000000000000_0000000000000000_0000100101100011_0001100110110001"; -- 0.03666840138612107
	pesos_i(6441) := b"1111111111111111_1111111111111111_1110100011111111_1101001001011000"; -- -0.08984647133377602
	pesos_i(6442) := b"0000000000000000_0000000000000000_0000100001100101_0001110011000100"; -- 0.032792852299110824
	pesos_i(6443) := b"1111111111111111_1111111111111111_1110001010000010_0011001000000110"; -- -0.11520087578475718
	pesos_i(6444) := b"1111111111111111_1111111111111111_1110100000000000_1101101110011111"; -- -0.09373690959393022
	pesos_i(6445) := b"1111111111111111_1111111111111111_1110100100001100_1000011100111110"; -- -0.08965258355795733
	pesos_i(6446) := b"1111111111111111_1111111111111111_1101000100110010_1111111011000000"; -- -0.18281562624939834
	pesos_i(6447) := b"1111111111111111_1111111111111111_1111110001000111_0111110001011101"; -- -0.014534213304574491
	pesos_i(6448) := b"0000000000000000_0000000000000000_0010010010110110_1010000000101101"; -- 0.1434116468819621
	pesos_i(6449) := b"1111111111111111_1111111111111111_1111111011100100_0101100001011010"; -- -0.0043282298859376005
	pesos_i(6450) := b"1111111111111111_1111111111111111_1110010111011001_1001010100000111"; -- -0.10214871003285839
	pesos_i(6451) := b"0000000000000000_0000000000000000_0010100110110110_1000111001010111"; -- 0.1629418337757048
	pesos_i(6452) := b"1111111111111111_1111111111111111_1111111110010101_0011010000000000"; -- -0.0016295908739696007
	pesos_i(6453) := b"1111111111111111_1111111111111111_1111011101110110_0010110100100110"; -- -0.033353021868798696
	pesos_i(6454) := b"0000000000000000_0000000000000000_0001011011001101_1100011110011110"; -- 0.08907744981892411
	pesos_i(6455) := b"1111111111111111_1111111111111111_1111000001000101_0011100111010000"; -- -0.06144369761064413
	pesos_i(6456) := b"0000000000000000_0000000000000000_0000010001001100_1100011011111110"; -- 0.016796528749059486
	pesos_i(6457) := b"0000000000000000_0000000000000000_0001000010001101_0000100111011011"; -- 0.06465207671740453
	pesos_i(6458) := b"1111111111111111_1111111111111111_1111010000011011_1010010000101101"; -- -0.04645322714076431
	pesos_i(6459) := b"1111111111111111_1111111111111111_1110000010111111_1100001010111000"; -- -0.12207396526134598
	pesos_i(6460) := b"1111111111111111_1111111111111111_1111110111000000_1000010101100101"; -- -0.008781111650877041
	pesos_i(6461) := b"0000000000000000_0000000000000000_0001011000110000_0111101000011101"; -- 0.0866772003130749
	pesos_i(6462) := b"1111111111111111_1111111111111111_1101111100111101_1010010011101000"; -- -0.127965634756774
	pesos_i(6463) := b"0000000000000000_0000000000000000_0000011011111000_0000011110010001"; -- 0.027222130630248618
	pesos_i(6464) := b"1111111111111111_1111111111111111_1110101111011111_1100101001000000"; -- -0.07861648489137307
	pesos_i(6465) := b"0000000000000000_0000000000000000_0000001011110111_0100110010111010"; -- 0.011585994269261272
	pesos_i(6466) := b"1111111111111111_1111111111111111_1110010110101000_0010110101000111"; -- -0.10290257466544349
	pesos_i(6467) := b"1111111111111111_1111111111111111_1101101100101011_0001001111100110"; -- -0.1438739360475336
	pesos_i(6468) := b"1111111111111111_1111111111111111_1110110100000100_0001100101111000"; -- -0.0741561968783765
	pesos_i(6469) := b"1111111111111111_1111111111111111_1110111000011101_1100001101110111"; -- -0.06985834450487938
	pesos_i(6470) := b"0000000000000000_0000000000000000_0001101110100100_0001000111000101"; -- 0.10797225046346232
	pesos_i(6471) := b"1111111111111111_1111111111111111_1111000001101111_0111011000010101"; -- -0.06079923611804461
	pesos_i(6472) := b"0000000000000000_0000000000000000_0001011111111001_0110110101100001"; -- 0.09364970785715611
	pesos_i(6473) := b"0000000000000000_0000000000000000_0001001011001101_1010110110101100"; -- 0.07345090331479566
	pesos_i(6474) := b"0000000000000000_0000000000000000_0001001110100111_1100000010111011"; -- 0.07677845530388437
	pesos_i(6475) := b"0000000000000000_0000000000000000_0001000100001011_0101110100101011"; -- 0.06657965000812387
	pesos_i(6476) := b"0000000000000000_0000000000000000_0010101100101001_0110100100110000"; -- 0.16860063008782836
	pesos_i(6477) := b"1111111111111111_1111111111111111_1110100101101011_0111101110111111"; -- -0.08820368366734439
	pesos_i(6478) := b"0000000000000000_0000000000000000_0010110001110110_0111010101111101"; -- 0.17368254006393946
	pesos_i(6479) := b"1111111111111111_1111111111111111_1110010000010111_0100010000100010"; -- -0.10901998672488554
	pesos_i(6480) := b"1111111111111111_1111111111111111_1111111011000000_0101010011110111"; -- -0.004877748284667943
	pesos_i(6481) := b"0000000000000000_0000000000000000_0000010101011011_0111011100010100"; -- 0.020926897373601365
	pesos_i(6482) := b"1111111111111111_1111111111111111_1110100101001001_1101011000111111"; -- -0.08871708831810704
	pesos_i(6483) := b"1111111111111111_1111111111111111_1110000111111111_1011000010111001"; -- -0.11719222538252701
	pesos_i(6484) := b"1111111111111111_1111111111111111_1110000111110000_1101011100101000"; -- -0.11741881635640679
	pesos_i(6485) := b"1111111111111111_1111111111111111_1110110100101100_0111000001101010"; -- -0.07354066295622372
	pesos_i(6486) := b"0000000000000000_0000000000000000_0001001010100001_0100010011000110"; -- 0.07277326417493661
	pesos_i(6487) := b"0000000000000000_0000000000000000_0001111001010011_0011001001010011"; -- 0.1184569790229299
	pesos_i(6488) := b"0000000000000000_0000000000000000_0000100100100001_0100010001101001"; -- 0.035663867601267774
	pesos_i(6489) := b"0000000000000000_0000000000000000_0010010110100011_0110110000101010"; -- 0.14702487975628842
	pesos_i(6490) := b"0000000000000000_0000000000000000_0010010011001011_0100101000011001"; -- 0.14372695068619873
	pesos_i(6491) := b"0000000000000000_0000000000000000_0001111010100101_1111001100010001"; -- 0.11971968811680327
	pesos_i(6492) := b"0000000000000000_0000000000000000_0001100110001111_1001010110101100"; -- 0.09984717791275487
	pesos_i(6493) := b"1111111111111111_1111111111111111_1110100011000110_1101111100000110"; -- -0.09071546658617168
	pesos_i(6494) := b"1111111111111111_1111111111111111_1110101001100101_1011001111000011"; -- -0.08438564776943636
	pesos_i(6495) := b"1111111111111111_1111111111111111_1111001010000001_0101101000110111"; -- -0.05271373893265492
	pesos_i(6496) := b"0000000000000000_0000000000000000_0000110010111000_0011111100000000"; -- 0.0496863722143539
	pesos_i(6497) := b"0000000000000000_0000000000000000_0000111101000110_0110000010111010"; -- 0.05966763058791902
	pesos_i(6498) := b"1111111111111111_1111111111111111_1101100110100111_1111010100000010"; -- -0.14978092871155252
	pesos_i(6499) := b"0000000000000000_0000000000000000_0001000110100001_0000101111101111"; -- 0.06886362644900378
	pesos_i(6500) := b"1111111111111111_1111111111111111_1111010011001010_0110000111111001"; -- -0.04378688489790138
	pesos_i(6501) := b"1111111111111111_1111111111111111_1111111001010101_1000010001101111"; -- -0.00650760923882849
	pesos_i(6502) := b"0000000000000000_0000000000000000_0001010010100011_1100100101010000"; -- 0.08062418180772371
	pesos_i(6503) := b"1111111111111111_1111111111111111_1111000010010100_0101101101110011"; -- -0.06023624852772484
	pesos_i(6504) := b"1111111111111111_1111111111111111_1110001101010000_0110101111000100"; -- -0.11205412363078737
	pesos_i(6505) := b"1111111111111111_1111111111111111_1111111001011011_0100011001110101"; -- -0.006419750731049043
	pesos_i(6506) := b"1111111111111111_1111111111111111_1111011100101100_1011001111100101"; -- -0.0344741407785533
	pesos_i(6507) := b"0000000000000000_0000000000000000_0010010011100111_1101101111101010"; -- 0.14416288812868555
	pesos_i(6508) := b"0000000000000000_0000000000000000_0000111101010110_0110100101011111"; -- 0.059912286429684665
	pesos_i(6509) := b"0000000000000000_0000000000000000_0000010001001010_1001110001100000"; -- 0.016763471114112596
	pesos_i(6510) := b"0000000000000000_0000000000000000_0000010011101011_0111011110001010"; -- 0.019217940499291646
	pesos_i(6511) := b"0000000000000000_0000000000000000_0001110101110100_0111010000111100"; -- 0.11505819762759087
	pesos_i(6512) := b"1111111111111111_1111111111111111_1101110011000000_1000000010011011"; -- -0.1376876469862273
	pesos_i(6513) := b"0000000000000000_0000000000000000_0010101000011011_1001110001101111"; -- 0.1644838114903665
	pesos_i(6514) := b"0000000000000000_0000000000000000_0001100100001100_0000011011101010"; -- 0.09783976765237837
	pesos_i(6515) := b"0000000000000000_0000000000000000_0010011100000111_0110001010011101"; -- 0.1524564392346399
	pesos_i(6516) := b"0000000000000000_0000000000000000_0001110001100110_1010111111100111"; -- 0.11094188114302746
	pesos_i(6517) := b"0000000000000000_0000000000000000_0010001110101101_0000011000100011"; -- 0.13935888625791584
	pesos_i(6518) := b"1111111111111111_1111111111111111_1110100110010001_0011111111110111"; -- -0.08762741309309945
	pesos_i(6519) := b"1111111111111111_1111111111111111_1111111001100011_0000001110000000"; -- -0.006301671197026771
	pesos_i(6520) := b"1111111111111111_1111111111111111_1101101111100011_1000010110110111"; -- -0.14105953480253874
	pesos_i(6521) := b"1111111111111111_1111111111111111_1110100111110001_0000100011101000"; -- -0.08616585106277672
	pesos_i(6522) := b"0000000000000000_0000000000000000_0001011111000101_0011100001011011"; -- 0.09285309059721268
	pesos_i(6523) := b"0000000000000000_0000000000000000_0010000111010001_1100011011000110"; -- 0.13210718479146022
	pesos_i(6524) := b"1111111111111111_1111111111111111_1110000000011110_1111101000011011"; -- -0.12452732897888662
	pesos_i(6525) := b"1111111111111111_1111111111111111_1111110101111110_1111101001010001"; -- -0.009781222631921613
	pesos_i(6526) := b"0000000000000000_0000000000000000_0001000001100000_1000000101000100"; -- 0.06397254855578231
	pesos_i(6527) := b"1111111111111111_1111111111111111_1111001001110000_1010000001001011"; -- -0.05296896136843386
	pesos_i(6528) := b"0000000000000000_0000000000000000_0010110100001001_0101010000000100"; -- 0.17592358693580792
	pesos_i(6529) := b"0000000000000000_0000000000000000_0010010100001010_1011101101000111"; -- 0.14469500048012118
	pesos_i(6530) := b"1111111111111111_1111111111111111_1111110000101011_1001001011000100"; -- -0.01496012405961953
	pesos_i(6531) := b"1111111111111111_1111111111111111_1111111101000111_1100100111001111"; -- -0.002810847281283882
	pesos_i(6532) := b"0000000000000000_0000000000000000_0001101110011001_1111010011100111"; -- 0.1078179420900932
	pesos_i(6533) := b"0000000000000000_0000000000000000_0010001110100010_1101100011111001"; -- 0.1392036064939929
	pesos_i(6534) := b"0000000000000000_0000000000000000_0000100000011101_0110100110111000"; -- 0.03169880625846948
	pesos_i(6535) := b"1111111111111111_1111111111111111_1111011000100111_0101000001111110"; -- -0.0384626095864651
	pesos_i(6536) := b"1111111111111111_1111111111111111_1111111011000001_0000110000101100"; -- -0.004866828182311259
	pesos_i(6537) := b"0000000000000000_0000000000000000_0000101101011011_0010001011110101"; -- 0.04435938336546679
	pesos_i(6538) := b"1111111111111111_1111111111111111_1101100101010110_1100101011101101"; -- -0.1510193988862949
	pesos_i(6539) := b"0000000000000000_0000000000000000_0000110000000011_1111111101101001"; -- 0.046936000015114034
	pesos_i(6540) := b"1111111111111111_1111111111111111_1101100010101010_1101110011001001"; -- -0.15364284612623938
	pesos_i(6541) := b"0000000000000000_0000000000000000_0001100010110010_1100010110001001"; -- 0.09647783854319165
	pesos_i(6542) := b"0000000000000000_0000000000000000_0001000110100101_0010000001111110"; -- 0.06892588680150913
	pesos_i(6543) := b"1111111111111111_1111111111111111_1111111001010110_1111111010101001"; -- -0.006485065196623991
	pesos_i(6544) := b"0000000000000000_0000000000000000_0010011110110000_0000101111010000"; -- 0.1550300009635173
	pesos_i(6545) := b"0000000000000000_0000000000000000_0010010001000001_1010010111011000"; -- 0.14162670642718816
	pesos_i(6546) := b"0000000000000000_0000000000000000_0010001000010010_0111111110100010"; -- 0.13309476563041392
	pesos_i(6547) := b"1111111111111111_1111111111111111_1110010010001100_0101111111101100"; -- -0.10723305206555989
	pesos_i(6548) := b"0000000000000000_0000000000000000_0010000100000000_0100100011010001"; -- 0.12891059023389953
	pesos_i(6549) := b"1111111111111111_1111111111111111_1110110001001011_0111100100100001"; -- -0.07697337097504175
	pesos_i(6550) := b"0000000000000000_0000000000000000_0001011011101101_1101101011111110"; -- 0.08956688587822309
	pesos_i(6551) := b"0000000000000000_0000000000000000_0001000001010110_1110101101011000"; -- 0.06382628346278589
	pesos_i(6552) := b"0000000000000000_0000000000000000_0001111101111011_1111101000010001"; -- 0.12298548611924517
	pesos_i(6553) := b"0000000000000000_0000000000000000_0010000010100001_1110100110001001"; -- 0.12747058486464963
	pesos_i(6554) := b"0000000000000000_0000000000000000_0000010110111001_0111001101101101"; -- 0.022361005949437518
	pesos_i(6555) := b"1111111111111111_1111111111111111_1111101010111000_1110010000110001"; -- -0.02061628161037941
	pesos_i(6556) := b"1111111111111111_1111111111111111_1101010100000001_0000100010101111"; -- -0.16795297371323673
	pesos_i(6557) := b"1111111111111111_1111111111111111_1101001010011111_1010001111000110"; -- -0.17725159090261977
	pesos_i(6558) := b"0000000000000000_0000000000000000_0001101011111101_0110010110100101"; -- 0.10542903221156612
	pesos_i(6559) := b"0000000000000000_0000000000000000_0010000011101001_1000101110111000"; -- 0.12856362583850564
	pesos_i(6560) := b"1111111111111111_1111111111111111_1101100001110101_0011101111001100"; -- -0.15446115754910453
	pesos_i(6561) := b"1111111111111111_1111111111111111_1101011111011110_1110011011100101"; -- -0.15675503632560853
	pesos_i(6562) := b"1111111111111111_1111111111111111_1110011110100010_1001100111000111"; -- -0.09517516035839764
	pesos_i(6563) := b"1111111111111111_1111111111111111_1101101000010110_1001010100110001"; -- -0.148092914165238
	pesos_i(6564) := b"0000000000000000_0000000000000000_0000011111011010_1100101100111111"; -- 0.030682280397988353
	pesos_i(6565) := b"0000000000000000_0000000000000000_0000000100111000_0100111011100111"; -- 0.0047654452330024655
	pesos_i(6566) := b"1111111111111111_1111111111111111_1110001011010001_0010100110101111"; -- -0.11399592853338777
	pesos_i(6567) := b"1111111111111111_1111111111111111_1110101011000111_1011101011101110"; -- -0.08288985906990606
	pesos_i(6568) := b"0000000000000000_0000000000000000_0010000000101110_1010111011110001"; -- 0.12571233165678883
	pesos_i(6569) := b"1111111111111111_1111111111111111_1110010010001101_1101111110111101"; -- -0.10721017494653934
	pesos_i(6570) := b"0000000000000000_0000000000000000_0010011000001111_1011100010001011"; -- 0.14867738140684514
	pesos_i(6571) := b"1111111111111111_1111111111111111_1111100110111100_0001000001110111"; -- -0.02447411625760058
	pesos_i(6572) := b"0000000000000000_0000000000000000_0010101110011001_0010000110010001"; -- 0.17030534533363512
	pesos_i(6573) := b"0000000000000000_0000000000000000_0001010001010010_0100100001001001"; -- 0.07938052921268243
	pesos_i(6574) := b"0000000000000000_0000000000000000_0010100000000011_1000000111010010"; -- 0.15630351420491181
	pesos_i(6575) := b"1111111111111111_1111111111111111_1110100010101101_0111100110110111"; -- -0.09110297482817006
	pesos_i(6576) := b"0000000000000000_0000000000000000_0000001010010000_0110010001000101"; -- 0.010015742190377153
	pesos_i(6577) := b"0000000000000000_0000000000000000_0000111000001011_0110101000111100"; -- 0.05486167867349629
	pesos_i(6578) := b"1111111111111111_1111111111111111_1110000000010000_1000000010010011"; -- -0.12474819581504752
	pesos_i(6579) := b"0000000000000000_0000000000000000_0000101110111101_1000011000101110"; -- 0.045860658926524064
	pesos_i(6580) := b"0000000000000000_0000000000000000_0001010101101001_1001001000001000"; -- 0.08364212705745842
	pesos_i(6581) := b"0000000000000000_0000000000000000_0000111010101101_0001111101001001"; -- 0.057329135298912426
	pesos_i(6582) := b"1111111111111111_1111111111111111_1111010011011010_1111110110001001"; -- -0.04353347206315362
	pesos_i(6583) := b"1111111111111111_1111111111111111_1101111000110100_1101001100010101"; -- -0.13200646139026412
	pesos_i(6584) := b"1111111111111111_1111111111111111_1111010000000111_1101000000001001"; -- -0.04675578861268945
	pesos_i(6585) := b"1111111111111111_1111111111111111_1101111011010101_0100011101010010"; -- -0.12955812699139052
	pesos_i(6586) := b"1111111111111111_1111111111111111_1101100110111010_1101100110011111"; -- -0.1494926440219271
	pesos_i(6587) := b"0000000000000000_0000000000000000_0001000100000110_0110000101111100"; -- 0.0665036132422269
	pesos_i(6588) := b"1111111111111111_1111111111111111_1110111100101001_0010101011111100"; -- -0.06577807747106316
	pesos_i(6589) := b"0000000000000000_0000000000000000_0001101111011111_1110101101000110"; -- 0.10888548326200331
	pesos_i(6590) := b"0000000000000000_0000000000000000_0001000000110111_0100111101100111"; -- 0.06334396619633795
	pesos_i(6591) := b"0000000000000000_0000000000000000_0010100000100100_0001010110101101"; -- 0.156800608393338
	pesos_i(6592) := b"0000000000000000_0000000000000000_0001011101001011_1011100100111101"; -- 0.09099920027811378
	pesos_i(6593) := b"0000000000000000_0000000000000000_0000111111000010_0101110001100110"; -- 0.06155946248546343
	pesos_i(6594) := b"0000000000000000_0000000000000000_0010010110011101_0110011010011011"; -- 0.14693299569041973
	pesos_i(6595) := b"0000000000000000_0000000000000000_0001011010011010_0001100000001111"; -- 0.0882887875913605
	pesos_i(6596) := b"1111111111111111_1111111111111111_1110010111001000_1001010110100000"; -- -0.10240807383270535
	pesos_i(6597) := b"1111111111111111_1111111111111111_1101101101101010_0110111101001000"; -- -0.14290718541398542
	pesos_i(6598) := b"1111111111111111_1111111111111111_1110111010110111_0000001111000000"; -- -0.06751991804621714
	pesos_i(6599) := b"0000000000000000_0000000000000000_0001101100010010_0101110000001011"; -- 0.10574889447276939
	pesos_i(6600) := b"0000000000000000_0000000000000000_0001100100010101_0001011001100001"; -- 0.0979780183467041
	pesos_i(6601) := b"0000000000000000_0000000000000000_0010010000111010_0110001101100010"; -- 0.14151593339334348
	pesos_i(6602) := b"0000000000000000_0000000000000000_0001100110000101_1001111010111000"; -- 0.09969512933729488
	pesos_i(6603) := b"1111111111111111_1111111111111111_1111001011011000_0001100111010101"; -- -0.05139006184890629
	pesos_i(6604) := b"0000000000000000_0000000000000000_0000101100001111_1110001000010100"; -- 0.04321110714297511
	pesos_i(6605) := b"0000000000000000_0000000000000000_0010000001110000_0101101010011101"; -- 0.12671438535986396
	pesos_i(6606) := b"1111111111111111_1111111111111111_1111010000011110_1011001011010101"; -- -0.046406577147672504
	pesos_i(6607) := b"1111111111111111_1111111111111111_1101100000001000_1010110000001011"; -- -0.15611767510095106
	pesos_i(6608) := b"1111111111111111_1111111111111111_1111101011010110_0100000010011000"; -- -0.020168269076203782
	pesos_i(6609) := b"1111111111111111_1111111111111111_1111000011101011_1110101111111001"; -- -0.05890011960700857
	pesos_i(6610) := b"1111111111111111_1111111111111111_1110011100001111_0001010010000001"; -- -0.0974261459671187
	pesos_i(6611) := b"1111111111111111_1111111111111111_1101111100110010_0000001110100100"; -- -0.12814309353443262
	pesos_i(6612) := b"0000000000000000_0000000000000000_0001110010111000_0110111110100000"; -- 0.11218927056935414
	pesos_i(6613) := b"1111111111111111_1111111111111111_1110001101001001_0111100111011011"; -- -0.11216009523570095
	pesos_i(6614) := b"0000000000000000_0000000000000000_0000100011011001_1100001010010100"; -- 0.03457275498178438
	pesos_i(6615) := b"0000000000000000_0000000000000000_0001100000101100_0111011011010100"; -- 0.09442846953346366
	pesos_i(6616) := b"0000000000000000_0000000000000000_0001101000011110_0110101011011011"; -- 0.10202663271793107
	pesos_i(6617) := b"0000000000000000_0000000000000000_0001101100100101_1101000011100100"; -- 0.10604577600495821
	pesos_i(6618) := b"0000000000000000_0000000000000000_0001111000000110_1000010001011110"; -- 0.11728694238661486
	pesos_i(6619) := b"0000000000000000_0000000000000000_0001010000101101_1010101101010111"; -- 0.07882185805394606
	pesos_i(6620) := b"1111111111111111_1111111111111111_1101001001101010_1101111010100101"; -- -0.17805679782273837
	pesos_i(6621) := b"1111111111111111_1111111111111111_1111110111100110_0100010010111100"; -- -0.008205131608746674
	pesos_i(6622) := b"1111111111111111_1111111111111111_1110110000001011_0001101010111110"; -- -0.0779555593075759
	pesos_i(6623) := b"0000000000000000_0000000000000000_0010101110111001_1011001101011010"; -- 0.17080231613009408
	pesos_i(6624) := b"0000000000000000_0000000000000000_0001001011000010_1000000010101100"; -- 0.07328037445005411
	pesos_i(6625) := b"1111111111111111_1111111111111111_1110100110110111_0111011011001111"; -- -0.08704431011087352
	pesos_i(6626) := b"1111111111111111_1111111111111111_1110110101001011_1001000110011001"; -- -0.07306566249527381
	pesos_i(6627) := b"0000000000000000_0000000000000000_0010011101101111_1101000101101111"; -- 0.1540499588464466
	pesos_i(6628) := b"0000000000000000_0000000000000000_0001001110011010_1011001111100110"; -- 0.07657932619300026
	pesos_i(6629) := b"0000000000000000_0000000000000000_0001000011110001_0101011100100001"; -- 0.06618256146320861
	pesos_i(6630) := b"0000000000000000_0000000000000000_0001010111110000_1111000100110010"; -- 0.08570773577924655
	pesos_i(6631) := b"0000000000000000_0000000000000000_0001001101111001_0001101011101111"; -- 0.07606666884404203
	pesos_i(6632) := b"0000000000000000_0000000000000000_0000010001011011_0011001011010001"; -- 0.017016578594275633
	pesos_i(6633) := b"1111111111111111_1111111111111111_1101100101100111_1100110001000110"; -- -0.15075991912728928
	pesos_i(6634) := b"1111111111111111_1111111111111111_1101010111010100_0110010101111101"; -- -0.16472783761087342
	pesos_i(6635) := b"0000000000000000_0000000000000000_0001011110010011_1000101000001001"; -- 0.09209501953410912
	pesos_i(6636) := b"1111111111111111_1111111111111111_1111010100011011_0001000000001011"; -- -0.0425558065246999
	pesos_i(6637) := b"1111111111111111_1111111111111111_1111111000000101_0110110001010001"; -- -0.007729749985671474
	pesos_i(6638) := b"1111111111111111_1111111111111111_1101111010010110_0110010101001110"; -- -0.13051764336313962
	pesos_i(6639) := b"0000000000000000_0000000000000000_0000001010100010_0000000000110111"; -- 0.01028443667366096
	pesos_i(6640) := b"0000000000000000_0000000000000000_0000101101101111_0100111011110110"; -- 0.044667182030835834
	pesos_i(6641) := b"0000000000000000_0000000000000000_0001110011000001_0011110011001110"; -- 0.11232357059692595
	pesos_i(6642) := b"0000000000000000_0000000000000000_0000101110000111_1110011101010101"; -- 0.04504247496330552
	pesos_i(6643) := b"0000000000000000_0000000000000000_0000011000011011_0001000000110110"; -- 0.023850453495066197
	pesos_i(6644) := b"0000000000000000_0000000000000000_0001000000100101_1010110101100010"; -- 0.06307490966832359
	pesos_i(6645) := b"0000000000000000_0000000000000000_0010100010000111_1001001000011000"; -- 0.15831864449726496
	pesos_i(6646) := b"0000000000000000_0000000000000000_0000000011100010_0010001001101110"; -- 0.0034505383953931613
	pesos_i(6647) := b"0000000000000000_0000000000000000_0000111101100111_1000010000011111"; -- 0.06017328020800116
	pesos_i(6648) := b"1111111111111111_1111111111111111_1110001000011101_0010110100011010"; -- -0.11674230682721778
	pesos_i(6649) := b"0000000000000000_0000000000000000_0000100101000000_1010111101011000"; -- 0.03614326377363154
	pesos_i(6650) := b"1111111111111111_1111111111111111_1110100011100000_1001100101011101"; -- -0.09032289000981963
	pesos_i(6651) := b"0000000000000000_0000000000000000_0000001001100110_0111010010110111"; -- 0.009375853286636773
	pesos_i(6652) := b"1111111111111111_1111111111111111_1101010010100010_0010100010000101"; -- -0.1694006610182174
	pesos_i(6653) := b"1111111111111111_1111111111111111_1110111101111110_0101010100110110"; -- -0.06447856362026191
	pesos_i(6654) := b"1111111111111111_1111111111111111_1101110001101101_0000111000000100"; -- -0.1389609566877938
	pesos_i(6655) := b"1111111111111111_1111111111111111_1101000110111100_1011101110101110"; -- -0.1807139111267598
	pesos_i(6656) := b"0000000000000000_0000000000000000_0000110100110111_0101000101111100"; -- 0.051625340172021944
	pesos_i(6657) := b"0000000000000000_0000000000000000_0001100001110000_1110111010101001"; -- 0.095473209582928
	pesos_i(6658) := b"0000000000000000_0000000000000000_0001111011010110_0001101101110111"; -- 0.12045451792592084
	pesos_i(6659) := b"0000000000000000_0000000000000000_0001000011111101_1000100100101100"; -- 0.06636864961403312
	pesos_i(6660) := b"1111111111111111_1111111111111111_1101101001000000_0010110110000101"; -- -0.1474582243662921
	pesos_i(6661) := b"1111111111111111_1111111111111111_1110001100111001_1101001100100101"; -- -0.11239891388130421
	pesos_i(6662) := b"0000000000000000_0000000000000000_0000101000111011_0001111101101011"; -- 0.0399646412204543
	pesos_i(6663) := b"1111111111111111_1111111111111111_1110010110000111_0111010010001110"; -- -0.10340186622413283
	pesos_i(6664) := b"1111111111111111_1111111111111111_1101110100000100_1100110001111101"; -- -0.1366455263043837
	pesos_i(6665) := b"1111111111111111_1111111111111111_1101001111111111_1110011000111000"; -- -0.171876536708862
	pesos_i(6666) := b"0000000000000000_0000000000000000_0010000010000110_0000011000101010"; -- 0.12704504508288947
	pesos_i(6667) := b"1111111111111111_1111111111111111_1111100110000100_0100001111011110"; -- -0.025325544546988123
	pesos_i(6668) := b"0000000000000000_0000000000000000_0010011010110011_0101110100110110"; -- 0.15117437906020914
	pesos_i(6669) := b"0000000000000000_0000000000000000_0010001110011011_0010011101100101"; -- 0.13908621032702598
	pesos_i(6670) := b"1111111111111111_1111111111111111_1110101111101110_1111011110000110"; -- -0.07838490460030333
	pesos_i(6671) := b"1111111111111111_1111111111111111_1101111000011001_1101000111001100"; -- -0.13241852541536042
	pesos_i(6672) := b"1111111111111111_1111111111111111_1111101010100001_0111100101011010"; -- -0.020973601869579472
	pesos_i(6673) := b"0000000000000000_0000000000000000_0000001101011000_0110101110010011"; -- 0.013067935390597562
	pesos_i(6674) := b"0000000000000000_0000000000000000_0000000010001011_0001100001101111"; -- 0.0021224279954302574
	pesos_i(6675) := b"1111111111111111_1111111111111111_1111100011010100_0101010001011110"; -- -0.028010107926741867
	pesos_i(6676) := b"0000000000000000_0000000000000000_0010101000000000_1100010111110110"; -- 0.16407429932782971
	pesos_i(6677) := b"1111111111111111_1111111111111111_1110011101111000_0101110101111000"; -- -0.09581962415511268
	pesos_i(6678) := b"1111111111111111_1111111111111111_1110000100011100_1000111110011010"; -- -0.12065794450292765
	pesos_i(6679) := b"0000000000000000_0000000000000000_0010100111010011_0000010111000111"; -- 0.1633761987565794
	pesos_i(6680) := b"1111111111111111_1111111111111111_1111010111111001_1110110000011111"; -- -0.039155237685413166
	pesos_i(6681) := b"1111111111111111_1111111111111111_1111110111000101_1001110101001100"; -- -0.00870339294045451
	pesos_i(6682) := b"1111111111111111_1111111111111111_1101000011001010_1000010100100111"; -- -0.1844097880884582
	pesos_i(6683) := b"1111111111111111_1111111111111111_1110111011010101_1100011001000110"; -- -0.06705056000303564
	pesos_i(6684) := b"0000000000000000_0000000000000000_0001101011111001_1010111011101100"; -- 0.10537236471160012
	pesos_i(6685) := b"0000000000000000_0000000000000000_0010011001011110_0011000000100101"; -- 0.14987469589087102
	pesos_i(6686) := b"0000000000000000_0000000000000000_0001111010011001_0111110110111110"; -- 0.11952958946390194
	pesos_i(6687) := b"1111111111111111_1111111111111111_1110110101110110_0101001001010100"; -- -0.07241330563696431
	pesos_i(6688) := b"0000000000000000_0000000000000000_0010110000011001_1001101110001010"; -- 0.17226574057918267
	pesos_i(6689) := b"0000000000000000_0000000000000000_0001110111111001_1001101111101011"; -- 0.11708998201710584
	pesos_i(6690) := b"1111111111111111_1111111111111111_1110110110011110_1101111101010110"; -- -0.07179454946508766
	pesos_i(6691) := b"1111111111111111_1111111111111111_1110100000011000_0001100100000111"; -- -0.09338229733355029
	pesos_i(6692) := b"0000000000000000_0000000000000000_0000110010010011_0000010000100111"; -- 0.049118289466156186
	pesos_i(6693) := b"1111111111111111_1111111111111111_1101100100101101_1100111010011001"; -- -0.15164479031719047
	pesos_i(6694) := b"0000000000000000_0000000000000000_0000001010101110_1011101100110111"; -- 0.010478688161747086
	pesos_i(6695) := b"1111111111111111_1111111111111111_1110001010010000_1000101111000000"; -- -0.11498190468039336
	pesos_i(6696) := b"1111111111111111_1111111111111111_1101110100001111_1001000000101110"; -- -0.13648127449963549
	pesos_i(6697) := b"1111111111111111_1111111111111111_1111010000101001_0111010000010110"; -- -0.046242470401375024
	pesos_i(6698) := b"0000000000000000_0000000000000000_0010000000100011_0001100110111100"; -- 0.12553559139298825
	pesos_i(6699) := b"1111111111111111_1111111111111111_1101111101111011_1010110101000100"; -- -0.12701909140264725
	pesos_i(6700) := b"0000000000000000_0000000000000000_0000110111101100_0101011101111011"; -- 0.054387538395074056
	pesos_i(6701) := b"1111111111111111_1111111111111111_1111011111101000_1111111011001000"; -- -0.03160102475615289
	pesos_i(6702) := b"1111111111111111_1111111111111111_1110110010111001_1100110001001001"; -- -0.07528994775638942
	pesos_i(6703) := b"1111111111111111_1111111111111111_1111101000000101_1001010101001011"; -- -0.023352307419490417
	pesos_i(6704) := b"1111111111111111_1111111111111111_1111100010010101_1101100111110000"; -- -0.028963450419732722
	pesos_i(6705) := b"0000000000000000_0000000000000000_0000010001010100_1011100000100101"; -- 0.016917714052962055
	pesos_i(6706) := b"0000000000000000_0000000000000000_0000001101101100_0001110111101000"; -- 0.013368481883509184
	pesos_i(6707) := b"1111111111111111_1111111111111111_1111111100000001_0101110011111001"; -- -0.0038854496545426896
	pesos_i(6708) := b"1111111111111111_1111111111111111_1101100000010010_1011111001110110"; -- -0.15596398949524298
	pesos_i(6709) := b"1111111111111111_1111111111111111_1111100011110011_0110111101100100"; -- -0.027535474793558785
	pesos_i(6710) := b"0000000000000000_0000000000000000_0001010000010011_1100111101101110"; -- 0.07842728082704796
	pesos_i(6711) := b"0000000000000000_0000000000000000_0001000110111100_1011110100000110"; -- 0.06928616908544873
	pesos_i(6712) := b"0000000000000000_0000000000000000_0001011100100100_0100111101111101"; -- 0.09039780420724566
	pesos_i(6713) := b"0000000000000000_0000000000000000_0000111010010000_1001111011100101"; -- 0.056894236592001345
	pesos_i(6714) := b"0000000000000000_0000000000000000_0010110111111011_1100011101110100"; -- 0.17962309441170168
	pesos_i(6715) := b"0000000000000000_0000000000000000_0001110100100010_1011111110001001"; -- 0.11381146519582203
	pesos_i(6716) := b"1111111111111111_1111111111111111_1110111010110010_1001100010101011"; -- -0.06758733583733983
	pesos_i(6717) := b"0000000000000000_0000000000000000_0000001100001111_0100100101111100"; -- 0.011952011883220065
	pesos_i(6718) := b"1111111111111111_1111111111111111_1111111101001100_0111010000111000"; -- -0.002739654896100127
	pesos_i(6719) := b"1111111111111111_1111111111111111_1101111000000101_0011101110010110"; -- -0.13273265434445392
	pesos_i(6720) := b"1111111111111111_1111111111111111_1110111100010010_1101111001010100"; -- -0.06611833995259161
	pesos_i(6721) := b"1111111111111111_1111111111111111_1111010100110111_1100100001110001"; -- -0.042117569370473125
	pesos_i(6722) := b"0000000000000000_0000000000000000_0001111000001011_1101100001000110"; -- 0.11736823752394922
	pesos_i(6723) := b"0000000000000000_0000000000000000_0000001111011011_0110000100110011"; -- 0.01506621840853426
	pesos_i(6724) := b"1111111111111111_1111111111111111_1110011110111011_1010000101101100"; -- -0.09479323506028448
	pesos_i(6725) := b"0000000000000000_0000000000000000_0010100001001001_0100101001001101"; -- 0.15736832016161015
	pesos_i(6726) := b"1111111111111111_1111111111111111_1110011111101100_0110001100100101"; -- -0.0940492662234199
	pesos_i(6727) := b"0000000000000000_0000000000000000_0001001010010110_1001111010010101"; -- 0.0726107706732847
	pesos_i(6728) := b"0000000000000000_0000000000000000_0000100110011010_0010111010111011"; -- 0.03750888893345486
	pesos_i(6729) := b"1111111111111111_1111111111111111_1110110111010110_0010110111111111"; -- -0.07095062766736895
	pesos_i(6730) := b"1111111111111111_1111111111111111_1111001000011101_1011000100011100"; -- -0.05423443862027859
	pesos_i(6731) := b"0000000000000000_0000000000000000_0010010001100111_1111110100111001"; -- 0.14221174843402415
	pesos_i(6732) := b"1111111111111111_1111111111111111_1111010010011001_1100101100011111"; -- -0.044528298258659955
	pesos_i(6733) := b"0000000000000000_0000000000000000_0001100011101001_0001001001010010"; -- 0.09730638974351088
	pesos_i(6734) := b"1111111111111111_1111111111111111_1110010110100111_0001111010110101"; -- -0.10291870194188335
	pesos_i(6735) := b"0000000000000000_0000000000000000_0010100001101110_0000101011111111"; -- 0.15792912219976246
	pesos_i(6736) := b"0000000000000000_0000000000000000_0010011010001110_0001101111100101"; -- 0.15060591071162502
	pesos_i(6737) := b"1111111111111111_1111111111111111_1101101110111101_1010101101111100"; -- -0.14163711763665923
	pesos_i(6738) := b"0000000000000000_0000000000000000_0001011000000101_1101010110111101"; -- 0.08602653382732056
	pesos_i(6739) := b"1111111111111111_1111111111111111_1101011001000101_1000111001010001"; -- -0.16300116080357366
	pesos_i(6740) := b"1111111111111111_1111111111111111_1110100111100101_0000010010101000"; -- -0.08634920982487813
	pesos_i(6741) := b"0000000000000000_0000000000000000_0000110100000110_0010000110010101"; -- 0.05087480439093933
	pesos_i(6742) := b"0000000000000000_0000000000000000_0001000010011101_0010000000110110"; -- 0.06489754981680783
	pesos_i(6743) := b"0000000000000000_0000000000000000_0001010010000010_1100111001111001"; -- 0.08012094937663848
	pesos_i(6744) := b"1111111111111111_1111111111111111_1101010010001111_0101000100111010"; -- -0.16968815168802856
	pesos_i(6745) := b"1111111111111111_1111111111111111_1111110111010111_1101100101100110"; -- -0.008425152354033252
	pesos_i(6746) := b"0000000000000000_0000000000000000_0000010110000100_0010010111110000"; -- 0.02154767151893193
	pesos_i(6747) := b"0000000000000000_0000000000000000_0001011101110000_1011111101011010"; -- 0.09156413991271829
	pesos_i(6748) := b"0000000000000000_0000000000000000_0001110010001101_1011111001011101"; -- 0.11153783578652753
	pesos_i(6749) := b"0000000000000000_0000000000000000_0010101110101100_1111111100100010"; -- 0.1706084688663908
	pesos_i(6750) := b"1111111111111111_1111111111111111_1110101010110000_1100111010100001"; -- -0.08323963710503642
	pesos_i(6751) := b"1111111111111111_1111111111111111_1110100100111010_1100000001100100"; -- -0.08894727293801613
	pesos_i(6752) := b"0000000000000000_0000000000000000_0010110010110111_0110001010100101"; -- 0.17467323803401022
	pesos_i(6753) := b"0000000000000000_0000000000000000_0010101110110110_1011001011010110"; -- 0.17075650897385933
	pesos_i(6754) := b"1111111111111111_1111111111111111_1101110101010011_1001011001010100"; -- -0.1354433102730822
	pesos_i(6755) := b"1111111111111111_1111111111111111_1110001011100001_1011101000110111"; -- -0.11374317326945556
	pesos_i(6756) := b"1111111111111111_1111111111111111_1101100110110101_1000110110100010"; -- -0.14957346710175423
	pesos_i(6757) := b"1111111111111111_1111111111111111_1110000110001001_0111101100100000"; -- -0.11899595711294697
	pesos_i(6758) := b"1111111111111111_1111111111111111_1110100011011101_1000010100100001"; -- -0.09036987260359158
	pesos_i(6759) := b"1111111111111111_1111111111111111_1110000000101110_1000011111001101"; -- -0.12429000142820965
	pesos_i(6760) := b"0000000000000000_0000000000000000_0000110001110100_1001010010000101"; -- 0.048653871883511834
	pesos_i(6761) := b"0000000000000000_0000000000000000_0010001001110111_1011110101000011"; -- 0.1346395768437139
	pesos_i(6762) := b"0000000000000000_0000000000000000_0000111010000000_0110111001001000"; -- 0.05664719836543238
	pesos_i(6763) := b"1111111111111111_1111111111111111_1101100001000001_1010111111110111"; -- -0.1552476904265245
	pesos_i(6764) := b"0000000000000000_0000000000000000_0000001100100110_0110110110110000"; -- 0.012305121941587263
	pesos_i(6765) := b"0000000000000000_0000000000000000_0000011010001100_1001111101111011"; -- 0.025583236224900878
	pesos_i(6766) := b"0000000000000000_0000000000000000_0000111001111011_1001111101100100"; -- 0.05657383147050086
	pesos_i(6767) := b"1111111111111111_1111111111111111_1110000100000000_0011111110110001"; -- -0.1210899535959196
	pesos_i(6768) := b"0000000000000000_0000000000000000_0000100010000001_1100000100101100"; -- 0.03322989766958562
	pesos_i(6769) := b"0000000000000000_0000000000000000_0010000111111110_1011101110001000"; -- 0.13279316025909957
	pesos_i(6770) := b"0000000000000000_0000000000000000_0001111100001101_0011100101011010"; -- 0.12129553275269948
	pesos_i(6771) := b"0000000000000000_0000000000000000_0001110101111010_0110011101110011"; -- 0.11514898836614874
	pesos_i(6772) := b"0000000000000000_0000000000000000_0000001010011010_0000101101000001"; -- 0.01016302419128106
	pesos_i(6773) := b"0000000000000000_0000000000000000_0000001000100010_1101001111100001"; -- 0.008343927881981066
	pesos_i(6774) := b"0000000000000000_0000000000000000_0010001001001011_0110111001000100"; -- 0.1339634815077089
	pesos_i(6775) := b"0000000000000000_0000000000000000_0000110101110111_1000100001101000"; -- 0.05260517641728948
	pesos_i(6776) := b"1111111111111111_1111111111111111_1110000101011100_0000111000011100"; -- -0.11968910033128496
	pesos_i(6777) := b"1111111111111111_1111111111111111_1110101111101111_1010110110011111"; -- -0.07837405081796045
	pesos_i(6778) := b"0000000000000000_0000000000000000_0000011001101011_0110001010011110"; -- 0.02507606849062842
	pesos_i(6779) := b"0000000000000000_0000000000000000_0001010101001110_1001000110111011"; -- 0.0832301217096801
	pesos_i(6780) := b"0000000000000000_0000000000000000_0001001101010100_0111000110100011"; -- 0.07550726152688694
	pesos_i(6781) := b"0000000000000000_0000000000000000_0001101111100001_0010111101111101"; -- 0.10890480795104944
	pesos_i(6782) := b"0000000000000000_0000000000000000_0010100110010111_1101011011111010"; -- 0.16247314068558885
	pesos_i(6783) := b"0000000000000000_0000000000000000_0010011010000111_1011001001000000"; -- 0.1505080609793538
	pesos_i(6784) := b"0000000000000000_0000000000000000_0010101100101111_1111011101011100"; -- 0.1687006567498968
	pesos_i(6785) := b"0000000000000000_0000000000000000_0000010110100111_1011110011111100"; -- 0.022090732094862692
	pesos_i(6786) := b"1111111111111111_1111111111111111_1111100011011001_1011101011010000"; -- -0.027927707784996425
	pesos_i(6787) := b"0000000000000000_0000000000000000_0010011111010001_1100100110010010"; -- 0.155544851512785
	pesos_i(6788) := b"1111111111111111_1111111111111111_1111001000100101_0010000011101010"; -- -0.05412096286902077
	pesos_i(6789) := b"0000000000000000_0000000000000000_0000101111110011_1100010100001001"; -- 0.04668838003853501
	pesos_i(6790) := b"1111111111111111_1111111111111111_1110111110000101_0101111111010010"; -- -0.06437111970111652
	pesos_i(6791) := b"0000000000000000_0000000000000000_0001001110110101_0000111010100010"; -- 0.07698146306214139
	pesos_i(6792) := b"1111111111111111_1111111111111111_1110001010001010_1100011010100000"; -- -0.11506994806414213
	pesos_i(6793) := b"0000000000000000_0000000000000000_0001010101010101_1100011010101101"; -- 0.08334008908482662
	pesos_i(6794) := b"0000000000000000_0000000000000000_0010001110100011_0011110101101110"; -- 0.13920959408904646
	pesos_i(6795) := b"0000000000000000_0000000000000000_0000100100000000_1110100000010111"; -- 0.03517008369987058
	pesos_i(6796) := b"0000000000000000_0000000000000000_0000011000011101_1101001011000101"; -- 0.023892567743980637
	pesos_i(6797) := b"0000000000000000_0000000000000000_0000101110010110_1010101101110000"; -- 0.045267786898066854
	pesos_i(6798) := b"1111111111111111_1111111111111111_1110000110111010_1111000101000001"; -- -0.11824123548171107
	pesos_i(6799) := b"1111111111111111_1111111111111111_1100111011111000_0011111100000001"; -- -0.19152456497732911
	pesos_i(6800) := b"0000000000000000_0000000000000000_0001101110101111_0001110001000111"; -- 0.10814072348956502
	pesos_i(6801) := b"0000000000000000_0000000000000000_0001100111101101_1110000111110011"; -- 0.1012860505283289
	pesos_i(6802) := b"1111111111111111_1111111111111111_1110111011110101_1111111111100100"; -- -0.0665588443466826
	pesos_i(6803) := b"0000000000000000_0000000000000000_0010111110111001_1100001111001001"; -- 0.18642829576382816
	pesos_i(6804) := b"0000000000000000_0000000000000000_0001000101100000_0010010111110100"; -- 0.06787335590726985
	pesos_i(6805) := b"0000000000000000_0000000000000000_0001101110011010_1000011001010111"; -- 0.10782661082713903
	pesos_i(6806) := b"0000000000000000_0000000000000000_0001111011011110_1100000001010011"; -- 0.12058641467977346
	pesos_i(6807) := b"1111111111111111_1111111111111111_1101001111001001_1111011000001111"; -- -0.17269956727151464
	pesos_i(6808) := b"0000000000000000_0000000000000000_0000001000000000_1011010100000111"; -- 0.007823289978620557
	pesos_i(6809) := b"1111111111111111_1111111111111111_1110001100111010_1100001011000001"; -- -0.11238463192049364
	pesos_i(6810) := b"1111111111111111_1111111111111111_1110110100110011_1110001011110101"; -- -0.07342702412878857
	pesos_i(6811) := b"1111111111111111_1111111111111111_1110011011101000_0100110001101000"; -- -0.09801790673080792
	pesos_i(6812) := b"1111111111111111_1111111111111111_1110110011110110_1010100001110110"; -- -0.0743612968338519
	pesos_i(6813) := b"1111111111111111_1111111111111111_1110000111110100_0100010101101011"; -- -0.11736646784470073
	pesos_i(6814) := b"1111111111111111_1111111111111111_1110011011010011_0110001110010111"; -- -0.09833695939375982
	pesos_i(6815) := b"1111111111111111_1111111111111111_1111010001100110_0010100001010011"; -- -0.045316200026340986
	pesos_i(6816) := b"1111111111111111_1111111111111111_1101100111101110_0001000010100100"; -- -0.14871116628941594
	pesos_i(6817) := b"0000000000000000_0000000000000000_0000011001111111_0111111110000110"; -- 0.0253829672684645
	pesos_i(6818) := b"1111111111111111_1111111111111111_1110001000000001_1001111000101101"; -- -0.11716281327081543
	pesos_i(6819) := b"0000000000000000_0000000000000000_0000011010100110_0000010100101011"; -- 0.02597076707591367
	pesos_i(6820) := b"0000000000000000_0000000000000000_0010010001011011_1111101110011101"; -- 0.14202854702787254
	pesos_i(6821) := b"0000000000000000_0000000000000000_0000111010000010_0001101001101110"; -- 0.05667271792375177
	pesos_i(6822) := b"1111111111111111_1111111111111111_1101101011111110_0110111101000101"; -- -0.14455513534067624
	pesos_i(6823) := b"1111111111111111_1111111111111111_1111011000101111_0110110110011001"; -- -0.038338804399614346
	pesos_i(6824) := b"0000000000000000_0000000000000000_0001011010111110_0010010111000011"; -- 0.08883892062254081
	pesos_i(6825) := b"1111111111111111_1111111111111111_1110010010011011_1111100100100000"; -- -0.1069950386611695
	pesos_i(6826) := b"1111111111111111_1111111111111111_1110100010111010_0110110110011011"; -- -0.09090533215837303
	pesos_i(6827) := b"0000000000000000_0000000000000000_0001111101011111_0110111101011010"; -- 0.12254997204986912
	pesos_i(6828) := b"0000000000000000_0000000000000000_0000001101111001_0001110111010101"; -- 0.013566841690747672
	pesos_i(6829) := b"1111111111111111_1111111111111111_1101111010001000_1010010001010000"; -- -0.13072751082101833
	pesos_i(6830) := b"1111111111111111_1111111111111111_1101100101111111_0001111011000011"; -- -0.1504040501513162
	pesos_i(6831) := b"0000000000000000_0000000000000000_0010001010001010_0011000000101110"; -- 0.13492108467039174
	pesos_i(6832) := b"0000000000000000_0000000000000000_0001100000110100_0111101111001101"; -- 0.09455083612902601
	pesos_i(6833) := b"0000000000000000_0000000000000000_0001111100000010_0110100110100111"; -- 0.12113056506162953
	pesos_i(6834) := b"0000000000000000_0000000000000000_0001110101101100_1110110011101001"; -- 0.11494332009706698
	pesos_i(6835) := b"1111111111111111_1111111111111111_1111110011100011_1011101001000101"; -- -0.012150152423468303
	pesos_i(6836) := b"1111111111111111_1111111111111111_1111100111010101_1101111011001111"; -- -0.02408034745259791
	pesos_i(6837) := b"0000000000000000_0000000000000000_0000100101000101_1111001000101110"; -- 0.03622354143118122
	pesos_i(6838) := b"0000000000000000_0000000000000000_0000111101111110_0010101100010110"; -- 0.060518925569061806
	pesos_i(6839) := b"0000000000000000_0000000000000000_0001001101100101_1110101110110000"; -- 0.07577393584463833
	pesos_i(6840) := b"1111111111111111_1111111111111111_1111101000011100_1110111111000000"; -- -0.022995963591865176
	pesos_i(6841) := b"0000000000000000_0000000000000000_0010000011110110_1010011100100110"; -- 0.12876362495788585
	pesos_i(6842) := b"1111111111111111_1111111111111111_1110101110111011_0110100001111010"; -- -0.07917162920109205
	pesos_i(6843) := b"0000000000000000_0000000000000000_0001111100100110_1111100010000101"; -- 0.12168839685413256
	pesos_i(6844) := b"1111111111111111_1111111111111111_1111010101010111_1110111111110011"; -- -0.04162693329266119
	pesos_i(6845) := b"1111111111111111_1111111111111111_1110001001101000_0000100011110000"; -- -0.1156000531335551
	pesos_i(6846) := b"1111111111111111_1111111111111111_1110011101111110_1110100101010000"; -- -0.09571973617919255
	pesos_i(6847) := b"1111111111111111_1111111111111111_1110000111011111_0000100000010001"; -- -0.11769055916518592
	pesos_i(6848) := b"1111111111111111_1111111111111111_1110001010111011_0111011100111111"; -- -0.11432699888514
	pesos_i(6849) := b"1111111111111111_1111111111111111_1110010101101111_0111000001010011"; -- -0.10376832925898923
	pesos_i(6850) := b"1111111111111111_1111111111111111_1101100111110110_1101101000111111"; -- -0.14857707945236925
	pesos_i(6851) := b"1111111111111111_1111111111111111_1111000111011111_1101010101011010"; -- -0.05517832335133314
	pesos_i(6852) := b"1111111111111111_1111111111111111_1101011001100010_0001111111011001"; -- -0.16256524041582643
	pesos_i(6853) := b"0000000000000000_0000000000000000_0000011001010001_1000110101010001"; -- 0.02468188497619175
	pesos_i(6854) := b"1111111111111111_1111111111111111_1110100100011011_1101010111100101"; -- -0.08941901369120019
	pesos_i(6855) := b"0000000000000000_0000000000000000_0001110001010101_0101011101010011"; -- 0.11067720209321623
	pesos_i(6856) := b"0000000000000000_0000000000000000_0001000000110111_1111010011100101"; -- 0.06335383022386318
	pesos_i(6857) := b"0000000000000000_0000000000000000_0010010001101110_1111111111001010"; -- 0.14231871312799463
	pesos_i(6858) := b"1111111111111111_1111111111111111_1101100111011011_0001111111001110"; -- -0.1490001795654643
	pesos_i(6859) := b"1111111111111111_1111111111111111_1110100100100110_0011111100100100"; -- -0.0892601525349127
	pesos_i(6860) := b"1111111111111111_1111111111111111_1110001000010100_0101011110011011"; -- -0.11687710257127414
	pesos_i(6861) := b"0000000000000000_0000000000000000_0000000110011011_0001110110011110"; -- 0.006273127546373962
	pesos_i(6862) := b"0000000000000000_0000000000000000_0001110011111011_0110011111101011"; -- 0.11321114995677072
	pesos_i(6863) := b"0000000000000000_0000000000000000_0010011111001000_1000000010000000"; -- 0.15540316695167514
	pesos_i(6864) := b"0000000000000000_0000000000000000_0001000010100100_1111010001000111"; -- 0.065017001458196
	pesos_i(6865) := b"0000000000000000_0000000000000000_0010100100000110_1001111000110011"; -- 0.16025723220151797
	pesos_i(6866) := b"0000000000000000_0000000000000000_0000010001011010_0111111011110111"; -- 0.017005858599453267
	pesos_i(6867) := b"1111111111111111_1111111111111111_1111011100000010_1010101010111100"; -- -0.03511555594468049
	pesos_i(6868) := b"1111111111111111_1111111111111111_1110001010110011_0101111101001111"; -- -0.1144504959760419
	pesos_i(6869) := b"1111111111111111_1111111111111111_1111001011000110_1000011100001111"; -- -0.051658209597364085
	pesos_i(6870) := b"0000000000000000_0000000000000000_0000100000011110_1011001101101101"; -- 0.03171845825446309
	pesos_i(6871) := b"0000000000000000_0000000000000000_0000010010011100_1010001000010011"; -- 0.018015031381288196
	pesos_i(6872) := b"0000000000000000_0000000000000000_0011011100010110_1111011111010010"; -- 0.21519421463979652
	pesos_i(6873) := b"0000000000000000_0000000000000000_0000000100000100_0100111000000011"; -- 0.003971935001357867
	pesos_i(6874) := b"0000000000000000_0000000000000000_0001000000001101_1100001011111110"; -- 0.06270998661248464
	pesos_i(6875) := b"0000000000000000_0000000000000000_0001011011101111_1011100110000010"; -- 0.08959540766664231
	pesos_i(6876) := b"1111111111111111_1111111111111111_1101111110010001_0101010001111000"; -- -0.12668869079178813
	pesos_i(6877) := b"0000000000000000_0000000000000000_0000011010010000_1101010000010100"; -- 0.025647406366972835
	pesos_i(6878) := b"1111111111111111_1111111111111111_1110101000101000_1010110010111001"; -- -0.08531685336257204
	pesos_i(6879) := b"1111111111111111_1111111111111111_1101001100000101_0101100001010011"; -- -0.1756996915138437
	pesos_i(6880) := b"1111111111111111_1111111111111111_1111110001110001_0001101000010111"; -- -0.013899201746225998
	pesos_i(6881) := b"1111111111111111_1111111111111111_1100110111001010_1100101000010000"; -- -0.19612443072188793
	pesos_i(6882) := b"0000000000000000_0000000000000000_0010000101011000_1000011110110100"; -- 0.1302571120175403
	pesos_i(6883) := b"0000000000000000_0000000000000000_0000000110100011_1010101100011001"; -- 0.006403630906549251
	pesos_i(6884) := b"1111111111111111_1111111111111111_1111001101011011_1010100111000101"; -- -0.049382581116563344
	pesos_i(6885) := b"0000000000000000_0000000000000000_0001111011110001_0010110111011011"; -- 0.12086760142522596
	pesos_i(6886) := b"0000000000000000_0000000000000000_0010010111110000_1100111010100110"; -- 0.14820567646813126
	pesos_i(6887) := b"1111111111111111_1111111111111111_1110110100000011_1110110001000100"; -- -0.07415889115877922
	pesos_i(6888) := b"0000000000000000_0000000000000000_0001001010100100_0100010100110000"; -- 0.07281906536908142
	pesos_i(6889) := b"1111111111111111_1111111111111111_1111001011001101_1111111110000000"; -- -0.051544219284860755
	pesos_i(6890) := b"1111111111111111_1111111111111111_1101010011111101_1110101000010110"; -- -0.16800057375407584
	pesos_i(6891) := b"0000000000000000_0000000000000000_0001010001111001_0011111110010001"; -- 0.07997510235669147
	pesos_i(6892) := b"1111111111111111_1111111111111111_1110010011100011_0010001100011011"; -- -0.10590916232981742
	pesos_i(6893) := b"0000000000000000_0000000000000000_0000011000110000_1001101000100100"; -- 0.02417910930586012
	pesos_i(6894) := b"1111111111111111_1111111111111111_1101111001111010_1000010101100100"; -- -0.13094297713634453
	pesos_i(6895) := b"1111111111111111_1111111111111111_1111001101001110_0111100100000110"; -- -0.049583850919522526
	pesos_i(6896) := b"0000000000000000_0000000000000000_0010100011000010_0001111110100011"; -- 0.15921209074266954
	pesos_i(6897) := b"0000000000000000_0000000000000000_0001111000100001_0111010010111011"; -- 0.11769799774846888
	pesos_i(6898) := b"1111111111111111_1111111111111111_1111000100110010_0001011011010000"; -- -0.057829450931365774
	pesos_i(6899) := b"0000000000000000_0000000000000000_0001110001111010_0001010011100100"; -- 0.11123781733833478
	pesos_i(6900) := b"1111111111111111_1111111111111111_1110101010100000_0110101100101000"; -- -0.08348970671205647
	pesos_i(6901) := b"0000000000000000_0000000000000000_0010000001111001_0111110001111000"; -- 0.12685373239799427
	pesos_i(6902) := b"0000000000000000_0000000000000000_0001100101100111_1111101001011101"; -- 0.09924282814058273
	pesos_i(6903) := b"1111111111111111_1111111111111111_1101011100010110_0100000111111001"; -- -0.15981662432225816
	pesos_i(6904) := b"1111111111111111_1111111111111111_1110010000001101_1000110011011110"; -- -0.10916823945107261
	pesos_i(6905) := b"0000000000000000_0000000000000000_0010010111001110_0101010110110011"; -- 0.14767966855494688
	pesos_i(6906) := b"1111111111111111_1111111111111111_1110001110010101_1011111011010100"; -- -0.11099631629360036
	pesos_i(6907) := b"0000000000000000_0000000000000000_0000110011111000_1001111111010101"; -- 0.050668706366475996
	pesos_i(6908) := b"1111111111111111_1111111111111111_1110100101100111_0100101001111100"; -- -0.08826765517165962
	pesos_i(6909) := b"1111111111111111_1111111111111111_1111101010100010_0111010111011011"; -- -0.020958551551474303
	pesos_i(6910) := b"1111111111111111_1111111111111111_1101100110011001_0101010111111101"; -- -0.15000402986838005
	pesos_i(6911) := b"1111111111111111_1111111111111111_1110110010110110_1000010001011010"; -- -0.07534001163028613
	pesos_i(6912) := b"1111111111111111_1111111111111111_1101011101101011_1000100011011010"; -- -0.1585154026314254
	pesos_i(6913) := b"1111111111111111_1111111111111111_1111011000011100_0110110111001101"; -- -0.038628709360886394
	pesos_i(6914) := b"0000000000000000_0000000000000000_0001101110000010_0100010001101001"; -- 0.10745647012756115
	pesos_i(6915) := b"0000000000000000_0000000000000000_0000110001101111_0000000111001001"; -- 0.04856883205866276
	pesos_i(6916) := b"1111111111111111_1111111111111111_1110111111110111_1010010101001011"; -- -0.06262747687873757
	pesos_i(6917) := b"1111111111111111_1111111111111111_1111101101001100_0111110010001001"; -- -0.018364159052025413
	pesos_i(6918) := b"1111111111111111_1111111111111111_1110110110000100_0100110010101010"; -- -0.0722000203891083
	pesos_i(6919) := b"1111111111111111_1111111111111111_1111010100011101_0110010001010001"; -- -0.042520265756236374
	pesos_i(6920) := b"1111111111111111_1111111111111111_1110111011010110_0001001111110001"; -- -0.06704593044326007
	pesos_i(6921) := b"0000000000000000_0000000000000000_0010001001010001_0110011010010011"; -- 0.13405457592895567
	pesos_i(6922) := b"0000000000000000_0000000000000000_0010011110110111_1110110100001110"; -- 0.15515023790454732
	pesos_i(6923) := b"1111111111111111_1111111111111111_1111110010100110_0110110101011110"; -- -0.013085522259159347
	pesos_i(6924) := b"0000000000000000_0000000000000000_0001011010000011_0101001101110101"; -- 0.08794137581547465
	pesos_i(6925) := b"0000000000000000_0000000000000000_0000011010000101_0001000011001001"; -- 0.025467919414928278
	pesos_i(6926) := b"0000000000000000_0000000000000000_0000000011000011_0110110100010001"; -- 0.002981964784450442
	pesos_i(6927) := b"1111111111111111_1111111111111111_1101111100100000_1111111101000111"; -- -0.1284027531206186
	pesos_i(6928) := b"1111111111111111_1111111111111111_1101111110101101_1101000000001001"; -- -0.1262540797465577
	pesos_i(6929) := b"0000000000000000_0000000000000000_0001101101001101_1010010101111111"; -- 0.1066535411454273
	pesos_i(6930) := b"1111111111111111_1111111111111111_1101010110011111_1101110100000101"; -- -0.16552942877891197
	pesos_i(6931) := b"0000000000000000_0000000000000000_0001110000110111_1000101101011100"; -- 0.11022253980451056
	pesos_i(6932) := b"1111111111111111_1111111111111111_1110010000110100_0011000110010110"; -- -0.10857858745785318
	pesos_i(6933) := b"1111111111111111_1111111111111111_1111011100110101_0101101110001001"; -- -0.034342078183299526
	pesos_i(6934) := b"1111111111111111_1111111111111111_1101011000110010_1000010011011000"; -- -0.1632916425195402
	pesos_i(6935) := b"0000000000000000_0000000000000000_0010100111101011_1011001111110011"; -- 0.16375279121614214
	pesos_i(6936) := b"1111111111111111_1111111111111111_1111100001101110_1001000011110110"; -- -0.02956289284535522
	pesos_i(6937) := b"0000000000000000_0000000000000000_0010100000101110_1101111111111011"; -- 0.15696525450541882
	pesos_i(6938) := b"1111111111111111_1111111111111111_1110010010110111_1001110100010001"; -- -0.10657327982455449
	pesos_i(6939) := b"0000000000000000_0000000000000000_0010101000111100_1110101110001011"; -- 0.16499206679359596
	pesos_i(6940) := b"0000000000000000_0000000000000000_0000001101100110_1001110000101011"; -- 0.013284454788492455
	pesos_i(6941) := b"1111111111111111_1111111111111111_1111011111010000_1001110101001100"; -- -0.031973046156012354
	pesos_i(6942) := b"0000000000000000_0000000000000000_0010001001110000_0111100101111101"; -- 0.13452872568124066
	pesos_i(6943) := b"0000000000000000_0000000000000000_0010100101101001_1000100010011000"; -- 0.16176656451031432
	pesos_i(6944) := b"0000000000000000_0000000000000000_0001001010110011_0001110101110100"; -- 0.07304557886732271
	pesos_i(6945) := b"1111111111111111_1111111111111111_1101100100110011_0101001011111111"; -- -0.151560604769648
	pesos_i(6946) := b"0000000000000000_0000000000000000_0000010111000101_0111000100111110"; -- 0.022543981209567993
	pesos_i(6947) := b"0000000000000000_0000000000000000_0010101011100011_0010111011111010"; -- 0.1675290450799719
	pesos_i(6948) := b"0000000000000000_0000000000000000_0000010011111011_1001001010110010"; -- 0.019463699859810862
	pesos_i(6949) := b"1111111111111111_1111111111111111_1111010110000111_1000011111110000"; -- -0.040900710875012236
	pesos_i(6950) := b"1111111111111111_1111111111111111_1110100001001011_1011111110111010"; -- -0.09259416291434505
	pesos_i(6951) := b"1111111111111111_1111111111111111_1111011111000011_0000010101000101"; -- -0.032180472107844776
	pesos_i(6952) := b"0000000000000000_0000000000000000_0010011001100111_0000010110101011"; -- 0.15000949305095398
	pesos_i(6953) := b"0000000000000000_0000000000000000_0010010001110110_0010000000110101"; -- 0.14242745675666552
	pesos_i(6954) := b"1111111111111111_1111111111111111_1111001001011111_0010001000000000"; -- -0.05323588853834443
	pesos_i(6955) := b"1111111111111111_1111111111111111_1111100111010011_1001101110010011"; -- -0.024114872629878156
	pesos_i(6956) := b"1111111111111111_1111111111111111_1110101001111011_1111000000111111"; -- -0.0840463492114164
	pesos_i(6957) := b"0000000000000000_0000000000000000_0000010001101000_0101100100000011"; -- 0.01721721951974664
	pesos_i(6958) := b"1111111111111111_1111111111111111_1101011110011100_1111111110010101"; -- -0.1577606449433575
	pesos_i(6959) := b"1111111111111111_1111111111111111_1111001110000001_0001111001011011"; -- -0.048811056809356795
	pesos_i(6960) := b"1111111111111111_1111111111111111_1111110101010100_0011010110001000"; -- -0.010433820905573432
	pesos_i(6961) := b"0000000000000000_0000000000000000_0001110111111000_0110101010010001"; -- 0.1170717814761939
	pesos_i(6962) := b"1111111111111111_1111111111111111_1111101001101111_0101101110000000"; -- -0.021738320554100684
	pesos_i(6963) := b"0000000000000000_0000000000000000_0000000111100100_0000110100000100"; -- 0.0073860296211441
	pesos_i(6964) := b"0000000000000000_0000000000000000_0010010011010001_1111101100001101"; -- 0.14382905076696462
	pesos_i(6965) := b"1111111111111111_1111111111111111_1111110100110011_0100111111100010"; -- -0.01093579035662982
	pesos_i(6966) := b"1111111111111111_1111111111111111_1111111101001110_1100101100100010"; -- -0.0027039568311055732
	pesos_i(6967) := b"0000000000000000_0000000000000000_0000001010001000_1011001101101110"; -- 0.009898390105240521
	pesos_i(6968) := b"0000000000000000_0000000000000000_0001000111011010_0011111101100110"; -- 0.06973644493290485
	pesos_i(6969) := b"0000000000000000_0000000000000000_0000111010011111_1010100111000111"; -- 0.05712376693705276
	pesos_i(6970) := b"0000000000000000_0000000000000000_0001101001100110_0110100110011001"; -- 0.10312519066783676
	pesos_i(6971) := b"1111111111111111_1111111111111111_1101101101000001_1100111111100110"; -- -0.14352703708630293
	pesos_i(6972) := b"1111111111111111_1111111111111111_1111011010000101_1101100111110101"; -- -0.03702008975059259
	pesos_i(6973) := b"0000000000000000_0000000000000000_0010000110111110_1101001000011100"; -- 0.1318179433799334
	pesos_i(6974) := b"1111111111111111_1111111111111111_1111111011001001_0001010011010101"; -- -0.004744241652587921
	pesos_i(6975) := b"1111111111111111_1111111111111111_1110001011110111_1101100101001110"; -- -0.11340562668861301
	pesos_i(6976) := b"0000000000000000_0000000000000000_0001011110011100_1011111001110101"; -- 0.09223547311824018
	pesos_i(6977) := b"1111111111111111_1111111111111111_1111111111010010_0001101101101100"; -- -0.0007002699284905194
	pesos_i(6978) := b"0000000000000000_0000000000000000_0001111101010111_1000001111100010"; -- 0.12242912540698993
	pesos_i(6979) := b"0000000000000000_0000000000000000_0001010111101010_0111010000110110"; -- 0.08560873324404056
	pesos_i(6980) := b"0000000000000000_0000000000000000_0000011011111001_0101010110110100"; -- 0.0272420466965569
	pesos_i(6981) := b"1111111111111111_1111111111111111_1110101111111110_0000011000110101"; -- -0.07815514753246561
	pesos_i(6982) := b"1111111111111111_1111111111111111_1111101101110101_0001111110101110"; -- -0.017744083450754133
	pesos_i(6983) := b"0000000000000000_0000000000000000_0000001100000110_1000010001000101"; -- 0.01181818669951538
	pesos_i(6984) := b"1111111111111111_1111111111111111_1110110001110110_0000000100100001"; -- -0.07632439567060935
	pesos_i(6985) := b"0000000000000000_0000000000000000_0000110000001010_1001010111011011"; -- 0.04703651989992251
	pesos_i(6986) := b"0000000000000000_0000000000000000_0001111011010110_0000101100001010"; -- 0.12045353874570776
	pesos_i(6987) := b"0000000000000000_0000000000000000_0001000000010011_1000110111111010"; -- 0.06279837942171589
	pesos_i(6988) := b"1111111111111111_1111111111111111_1110010001011100_1101011010010100"; -- -0.10795840161271182
	pesos_i(6989) := b"1111111111111111_1111111111111111_1101110000000101_1001101101101010"; -- -0.14053944257440454
	pesos_i(6990) := b"1111111111111111_1111111111111111_1110110011101010_1100111011101000"; -- -0.07454211079577203
	pesos_i(6991) := b"0000000000000000_0000000000000000_0000001001011010_1010100100010000"; -- 0.009195867945183832
	pesos_i(6992) := b"0000000000000000_0000000000000000_0001011010111000_1100101100001001"; -- 0.08875721890969837
	pesos_i(6993) := b"1111111111111111_1111111111111111_1110100001010110_1111000001011010"; -- -0.09242341811898455
	pesos_i(6994) := b"0000000000000000_0000000000000000_0010000111100010_1011100010110111"; -- 0.13236574614192628
	pesos_i(6995) := b"0000000000000000_0000000000000000_0000110000011111_1000010110011010"; -- 0.04735598582105621
	pesos_i(6996) := b"1111111111111111_1111111111111111_1111111011000000_1101100000000000"; -- -0.004869937995367968
	pesos_i(6997) := b"1111111111111111_1111111111111111_1100111011010100_0000100101011111"; -- -0.1920770781539347
	pesos_i(6998) := b"0000000000000000_0000000000000000_0001001010110001_0001110111001011"; -- 0.07301508136875026
	pesos_i(6999) := b"1111111111111111_1111111111111111_1110111010011111_1010000011101001"; -- -0.06787676154386267
	pesos_i(7000) := b"1111111111111111_1111111111111111_1111110010000010_0011001011110111"; -- -0.01363831969795046
	pesos_i(7001) := b"1111111111111111_1111111111111111_1101010110111101_1010100001010011"; -- -0.1650748059480347
	pesos_i(7002) := b"0000000000000000_0000000000000000_0001110110011000_0001001100110010"; -- 0.11560173014001135
	pesos_i(7003) := b"0000000000000000_0000000000000000_0000100010101010_1000001000010111"; -- 0.033851748022955465
	pesos_i(7004) := b"1111111111111111_1111111111111111_1110100100001100_1110010111001101"; -- -0.08964694730019968
	pesos_i(7005) := b"0000000000000000_0000000000000000_0000011001111111_1100001010000001"; -- 0.02538695959561565
	pesos_i(7006) := b"1111111111111111_1111111111111111_1111000001110100_1001101100111100"; -- -0.06072072789010069
	pesos_i(7007) := b"1111111111111111_1111111111111111_1110101001000001_0011001001110001"; -- -0.08494267208396575
	pesos_i(7008) := b"0000000000000000_0000000000000000_0000100111001001_1010001010101011"; -- 0.03823296244973817
	pesos_i(7009) := b"1111111111111111_1111111111111111_1110110101010011_1110011110001000"; -- -0.07293847006781932
	pesos_i(7010) := b"0000000000000000_0000000000000000_0000010010011001_1111001110111100"; -- 0.017974122346343917
	pesos_i(7011) := b"1111111111111111_1111111111111111_1101101111000100_0101101000011100"; -- -0.14153515643161127
	pesos_i(7012) := b"0000000000000000_0000000000000000_0010010000111111_0000010010111101"; -- 0.14158658623232154
	pesos_i(7013) := b"0000000000000000_0000000000000000_0010011010011010_0011010101001101"; -- 0.15079053039038184
	pesos_i(7014) := b"1111111111111111_1111111111111111_1110101011101011_0110100011111001"; -- -0.08234542776477108
	pesos_i(7015) := b"1111111111111111_1111111111111111_1111001001001010_1111101101100110"; -- -0.05354336520595297
	pesos_i(7016) := b"1111111111111111_1111111111111111_1101110001011011_1111000010011111"; -- -0.1392221080932192
	pesos_i(7017) := b"0000000000000000_0000000000000000_0001101110110101_1111111111010001"; -- 0.10824583868650677
	pesos_i(7018) := b"0000000000000000_0000000000000000_0001010101110100_0111100111000001"; -- 0.08380852661372382
	pesos_i(7019) := b"0000000000000000_0000000000000000_0000100010001011_1100101010100101"; -- 0.03338305017513029
	pesos_i(7020) := b"0000000000000000_0000000000000000_0001100101011010_1101001101001011"; -- 0.09904213502389252
	pesos_i(7021) := b"0000000000000000_0000000000000000_0010000001001101_0011101010101001"; -- 0.12617842308243649
	pesos_i(7022) := b"1111111111111111_1111111111111111_1101111110001010_1000101001100100"; -- -0.1267922884718196
	pesos_i(7023) := b"1111111111111111_1111111111111111_1110011010001011_0001101110011110"; -- -0.09943988219063087
	pesos_i(7024) := b"1111111111111111_1111111111111111_1110101001110001_1110100101110010"; -- -0.08419934247321362
	pesos_i(7025) := b"0000000000000000_0000000000000000_0000100001110010_0100011000011101"; -- 0.03299368092651278
	pesos_i(7026) := b"1111111111111111_1111111111111111_1101010100011101_1001101010000100"; -- -0.16751703527114323
	pesos_i(7027) := b"1111111111111111_1111111111111111_1110010101110110_0000000101101000"; -- -0.10366812900508515
	pesos_i(7028) := b"0000000000000000_0000000000000000_0001001010110000_1111101110100011"; -- 0.07301304569328963
	pesos_i(7029) := b"1111111111111111_1111111111111111_1111101010101000_1001000111100001"; -- -0.020865328340482603
	pesos_i(7030) := b"1111111111111111_1111111111111111_1110100100111010_0010001110101110"; -- -0.08895661364987727
	pesos_i(7031) := b"0000000000000000_0000000000000000_0010011110100000_1110001110110000"; -- 0.15479872743984804
	pesos_i(7032) := b"1111111111111111_1111111111111111_1101011100010101_0000110110010110"; -- -0.15983500559816563
	pesos_i(7033) := b"1111111111111111_1111111111111111_1110110010100001_1111111010000000"; -- -0.07565316556074772
	pesos_i(7034) := b"1111111111111111_1111111111111111_1101110110010000_1110100000001111"; -- -0.13450765267495549
	pesos_i(7035) := b"0000000000000000_0000000000000000_0001101001000101_1111100111000100"; -- 0.1026302436748199
	pesos_i(7036) := b"0000000000000000_0000000000000000_0010010011000001_0010001000011100"; -- 0.14357197940066574
	pesos_i(7037) := b"1111111111111111_1111111111111111_1111100001011011_0101011100001000"; -- -0.029856262738049446
	pesos_i(7038) := b"0000000000000000_0000000000000000_0000010101110110_0101110101101011"; -- 0.02133735535496913
	pesos_i(7039) := b"1111111111111111_1111111111111111_1111011100010101_0110101100100100"; -- -0.0348294293803781
	pesos_i(7040) := b"0000000000000000_0000000000000000_0001001001110110_0100100011000010"; -- 0.07211737384579878
	pesos_i(7041) := b"1111111111111111_1111111111111111_1111110101110000_1100101111111001"; -- -0.009997607844253
	pesos_i(7042) := b"1111111111111111_1111111111111111_1101011100111110_0011011110101011"; -- -0.15920688701114655
	pesos_i(7043) := b"0000000000000000_0000000000000000_0010000010010000_0111110001001000"; -- 0.12720467333007027
	pesos_i(7044) := b"0000000000000000_0000000000000000_0001110001000100_0010101010100101"; -- 0.11041513939123222
	pesos_i(7045) := b"0000000000000000_0000000000000000_0000101100100101_0111010000110001"; -- 0.043540250683993455
	pesos_i(7046) := b"0000000000000000_0000000000000000_0010011101000010_1010110010000000"; -- 0.1533611118636299
	pesos_i(7047) := b"0000000000000000_0000000000000000_0010010110001100_1010101101110010"; -- 0.14667769940360698
	pesos_i(7048) := b"0000000000000000_0000000000000000_0001000010100100_0010110110011110"; -- 0.06500516043249938
	pesos_i(7049) := b"0000000000000000_0000000000000000_0000010100011100_0001100001010010"; -- 0.019959945715416965
	pesos_i(7050) := b"0000000000000000_0000000000000000_0000010110101111_0010110110110010"; -- 0.02220426177246946
	pesos_i(7051) := b"0000000000000000_0000000000000000_0000110100101101_1001000111000011"; -- 0.05147658363658186
	pesos_i(7052) := b"1111111111111111_1111111111111111_1111110100110100_1111000111010001"; -- -0.010910879471792822
	pesos_i(7053) := b"1111111111111111_1111111111111111_1101110100101000_1001001101110001"; -- -0.13609961020842148
	pesos_i(7054) := b"0000000000000000_0000000000000000_0001011011010011_1001110111100111"; -- 0.08916651624282808
	pesos_i(7055) := b"1111111111111111_1111111111111111_1111010001011110_1110010011010001"; -- -0.045427035420651345
	pesos_i(7056) := b"1111111111111111_1111111111111111_1111110000111011_1010001100001101"; -- -0.014715012925543391
	pesos_i(7057) := b"0000000000000000_0000000000000000_0001011001110000_1010011101111110"; -- 0.08765646778746353
	pesos_i(7058) := b"0000000000000000_0000000000000000_0001101110000101_1000111010011101"; -- 0.10750666930657791
	pesos_i(7059) := b"1111111111111111_1111111111111111_1101101000111101_0101001100111110"; -- -0.14750175225718587
	pesos_i(7060) := b"0000000000000000_0000000000000000_0001001101011100_1001110110100110"; -- 0.0756319551358126
	pesos_i(7061) := b"1111111111111111_1111111111111111_1110001000111011_0111110011101101"; -- -0.11627978537504012
	pesos_i(7062) := b"0000000000000000_0000000000000000_0010111000110001_1100001001011110"; -- 0.18044676590791386
	pesos_i(7063) := b"0000000000000000_0000000000000000_0001011001000100_1011101010101111"; -- 0.0869862248404137
	pesos_i(7064) := b"0000000000000000_0000000000000000_0000100011000000_1001100001001000"; -- 0.03418876417243175
	pesos_i(7065) := b"0000000000000000_0000000000000000_0000000010001011_0101110110001001"; -- 0.0021265466980680027
	pesos_i(7066) := b"0000000000000000_0000000000000000_0001110011011101_1011100100001000"; -- 0.11275822099471042
	pesos_i(7067) := b"0000000000000000_0000000000000000_0010010010001000_1001000100111101"; -- 0.14270885214154555
	pesos_i(7068) := b"1111111111111111_1111111111111111_1110101101110000_0000101101000101"; -- -0.08032159398032335
	pesos_i(7069) := b"0000000000000000_0000000000000000_0001110000110000_1101101011011011"; -- 0.11012046676547045
	pesos_i(7070) := b"0000000000000000_0000000000000000_0001101000101000_1110110110010110"; -- 0.10218701288005927
	pesos_i(7071) := b"0000000000000000_0000000000000000_0000001011011000_1010110100011101"; -- 0.011118716747520074
	pesos_i(7072) := b"0000000000000000_0000000000000000_0010100101000101_0001000010110100"; -- 0.16121010206166633
	pesos_i(7073) := b"1111111111111111_1111111111111111_1110100110100101_0101111111001000"; -- -0.08732034086455776
	pesos_i(7074) := b"0000000000000000_0000000000000000_0001111011101100_0101010110110100"; -- 0.12079368246878054
	pesos_i(7075) := b"1111111111111111_1111111111111111_1111010001010001_1100111110000110"; -- -0.04562666861455838
	pesos_i(7076) := b"1111111111111111_1111111111111111_1101010111000011_1100110101001000"; -- -0.16498105031147114
	pesos_i(7077) := b"1111111111111111_1111111111111111_1111101001011111_1001110001110101"; -- -0.021978589419631468
	pesos_i(7078) := b"1111111111111111_1111111111111111_1101011010100101_0010000010110100"; -- -0.16154285046965292
	pesos_i(7079) := b"0000000000000000_0000000000000000_0001001011010111_1001011101011110"; -- 0.07360216185204135
	pesos_i(7080) := b"0000000000000000_0000000000000000_0000011001101011_0101111110010100"; -- 0.0250758874135886
	pesos_i(7081) := b"0000000000000000_0000000000000000_0000111110000010_1101101000000000"; -- 0.06059038645767855
	pesos_i(7082) := b"1111111111111111_1111111111111111_1101011011101101_1010010101000001"; -- -0.16043631718512236
	pesos_i(7083) := b"0000000000000000_0000000000000000_0000110100111011_0110111010000000"; -- 0.05168810484549025
	pesos_i(7084) := b"1111111111111111_1111111111111111_1110110100001000_1100011111110110"; -- -0.07408476101430081
	pesos_i(7085) := b"0000000000000000_0000000000000000_0001110111100001_1111010011100010"; -- 0.11672907377037414
	pesos_i(7086) := b"1111111111111111_1111111111111111_1110110010110100_1100001010101110"; -- -0.07536681426916532
	pesos_i(7087) := b"1111111111111111_1111111111111111_1110100100010101_0001000111111101"; -- -0.08952224322307364
	pesos_i(7088) := b"0000000000000000_0000000000000000_0001001011010001_0010010011010100"; -- 0.0735037819609913
	pesos_i(7089) := b"1111111111111111_1111111111111111_1101011000010000_0010011111111000"; -- -0.1638159769752674
	pesos_i(7090) := b"0000000000000000_0000000000000000_0001011100101101_0000111100010100"; -- 0.0905312942663345
	pesos_i(7091) := b"0000000000000000_0000000000000000_0000110111000010_1110110010001000"; -- 0.053755553381328605
	pesos_i(7092) := b"0000000000000000_0000000000000000_0001010010111111_1010011100011110"; -- 0.08104938960027767
	pesos_i(7093) := b"1111111111111111_1111111111111111_1111001010010001_1000010011100100"; -- -0.052467054637601145
	pesos_i(7094) := b"1111111111111111_1111111111111111_1111111010011010_0010101100011111"; -- -0.00546007620210628
	pesos_i(7095) := b"0000000000000000_0000000000000000_0011101001000111_1111111000010100"; -- 0.22766101817954126
	pesos_i(7096) := b"0000000000000000_0000000000000000_0010110001111101_0110111001101001"; -- 0.17378892960185685
	pesos_i(7097) := b"0000000000000000_0000000000000000_0011010100100101_1101000111011011"; -- 0.20760833365422862
	pesos_i(7098) := b"0000000000000000_0000000000000000_0001110011011100_1101110111101001"; -- 0.11274516045668677
	pesos_i(7099) := b"0000000000000000_0000000000000000_0001001010111100_1111010100101000"; -- 0.07319576476868174
	pesos_i(7100) := b"1111111111111111_1111111111111111_1110011101000100_0101111001001100"; -- -0.09661303173627099
	pesos_i(7101) := b"1111111111111111_1111111111111111_1101111010011001_0000101001011110"; -- -0.13047728722880064
	pesos_i(7102) := b"1111111111111111_1111111111111111_1111101000001100_0000101000011000"; -- -0.023253792946408804
	pesos_i(7103) := b"0000000000000000_0000000000000000_0010011100110111_1110000010111000"; -- 0.15319637763234678
	pesos_i(7104) := b"0000000000000000_0000000000000000_0001011100111001_0010101101101110"; -- 0.09071608954349755
	pesos_i(7105) := b"1111111111111111_1111111111111111_1111000110001110_1010000100111110"; -- -0.05641739113822814
	pesos_i(7106) := b"1111111111111111_1111111111111111_1101111101010110_0111101011000111"; -- -0.12758667610303498
	pesos_i(7107) := b"0000000000000000_0000000000000000_0010101100001010_0100100011111110"; -- 0.168125688625898
	pesos_i(7108) := b"1111111111111111_1111111111111111_1110101111111011_1010011100100101"; -- -0.07819133138518926
	pesos_i(7109) := b"1111111111111111_1111111111111111_1101110101011101_1011011001010110"; -- -0.1352888144759174
	pesos_i(7110) := b"0000000000000000_0000000000000000_0000011011010010_1000000111010000"; -- 0.026649583174590534
	pesos_i(7111) := b"1111111111111111_1111111111111111_1111000101110101_0001101111100101"; -- -0.056806809107684424
	pesos_i(7112) := b"1111111111111111_1111111111111111_1111001110011001_1000101001111000"; -- -0.04843840186307158
	pesos_i(7113) := b"1111111111111111_1111111111111111_1101101100100010_0100110101010000"; -- -0.14400784295744049
	pesos_i(7114) := b"0000000000000000_0000000000000000_0001001010010001_0100110101001011"; -- 0.07252963145509664
	pesos_i(7115) := b"0000000000000000_0000000000000000_0000010110110111_0100010110011111"; -- 0.022327758085067137
	pesos_i(7116) := b"0000000000000000_0000000000000000_0000100010110011_0110101110010010"; -- 0.03398773496844772
	pesos_i(7117) := b"0000000000000000_0000000000000000_0001100000000100_1010000110010111"; -- 0.0938206666246475
	pesos_i(7118) := b"1111111111111111_1111111111111111_1101101110101100_0111001010100011"; -- -0.14189990532859484
	pesos_i(7119) := b"1111111111111111_1111111111111111_1111000110001001_1001000001001101"; -- -0.056494694831710775
	pesos_i(7120) := b"0000000000000000_0000000000000000_0000000001011010_1111011001101101"; -- 0.0013879791491054616
	pesos_i(7121) := b"0000000000000000_0000000000000000_0000111010100011_1110001010110110"; -- 0.05718819554564284
	pesos_i(7122) := b"0000000000000000_0000000000000000_0000010110001011_0100110111000110"; -- 0.021656857297899193
	pesos_i(7123) := b"0000000000000000_0000000000000000_0000101011000100_0110100111100001"; -- 0.04205953353387664
	pesos_i(7124) := b"0000000000000000_0000000000000000_0000000010100110_1100011010001011"; -- 0.0025447929627547116
	pesos_i(7125) := b"0000000000000000_0000000000000000_0000111111001000_1100101010101010"; -- 0.06165758762847931
	pesos_i(7126) := b"0000000000000000_0000000000000000_0000110101101100_1001001100001100"; -- 0.05243796393909011
	pesos_i(7127) := b"1111111111111111_1111111111111111_1101011101110011_1111001000000111"; -- -0.15838706336745983
	pesos_i(7128) := b"1111111111111111_1111111111111111_1110101110111001_1000011000100111"; -- -0.07920037790820007
	pesos_i(7129) := b"0000000000000000_0000000000000000_0001110110010100_0110110001001010"; -- 0.11554600540206779
	pesos_i(7130) := b"0000000000000000_0000000000000000_0010110111010000_1111110110011110"; -- 0.17897019497314004
	pesos_i(7131) := b"1111111111111111_1111111111111111_1111010000111101_1100000001001111"; -- -0.045932751285528615
	pesos_i(7132) := b"0000000000000000_0000000000000000_0000011010010000_0100011010110111"; -- 0.025638980539052645
	pesos_i(7133) := b"1111111111111111_1111111111111111_1110101110010011_0010010001011101"; -- -0.07978604067270585
	pesos_i(7134) := b"1111111111111111_1111111111111111_1110000110010111_0010001111100100"; -- -0.11878753351448793
	pesos_i(7135) := b"0000000000000000_0000000000000000_0000111001101100_1111000100100111"; -- 0.05634982312729317
	pesos_i(7136) := b"0000000000000000_0000000000000000_0000100010111000_1110011000101000"; -- 0.034071335500539535
	pesos_i(7137) := b"0000000000000000_0000000000000000_0001001110001001_0010101111100010"; -- 0.07631181983076286
	pesos_i(7138) := b"1111111111111111_1111111111111111_1111001101001100_1110001100110101"; -- -0.04960803954759131
	pesos_i(7139) := b"1111111111111111_1111111111111111_1110101001111011_0011000111001011"; -- -0.08405770104832194
	pesos_i(7140) := b"1111111111111111_1111111111111111_1101010111100001_1100111001011000"; -- -0.16452322348969844
	pesos_i(7141) := b"1111111111111111_1111111111111111_1101110110011100_1111111001110100"; -- -0.13432321220989046
	pesos_i(7142) := b"0000000000000000_0000000000000000_0000101000000111_0110011001111011"; -- 0.039175419798289285
	pesos_i(7143) := b"0000000000000000_0000000000000000_0000100100000011_1110100000110011"; -- 0.03521586645041083
	pesos_i(7144) := b"1111111111111111_1111111111111111_1111100010001010_1000011111011000"; -- -0.02913619025274744
	pesos_i(7145) := b"1111111111111111_1111111111111111_1110111011110001_0110111110111010"; -- -0.06662847239993873
	pesos_i(7146) := b"0000000000000000_0000000000000000_0000111001001000_1001100111100011"; -- 0.05579530510269128
	pesos_i(7147) := b"0000000000000000_0000000000000000_0010110010100010_1111000110101100"; -- 0.1743613286549406
	pesos_i(7148) := b"1111111111111111_1111111111111111_1110010001111101_0101111111101110"; -- -0.10746193345090746
	pesos_i(7149) := b"0000000000000000_0000000000000000_0001100000110111_1000001000110011"; -- 0.09459699393572045
	pesos_i(7150) := b"0000000000000000_0000000000000000_0001111100100011_1101100001010110"; -- 0.12164070235279607
	pesos_i(7151) := b"0000000000000000_0000000000000000_0000011011101010_0011011100010101"; -- 0.02701133980212487
	pesos_i(7152) := b"0000000000000000_0000000000000000_0000011001111010_1000000111110101"; -- 0.02530681840887633
	pesos_i(7153) := b"0000000000000000_0000000000000000_0000111101011000_0110101010001101"; -- 0.059942874321117695
	pesos_i(7154) := b"0000000000000000_0000000000000000_0010000010111111_0001000101011111"; -- 0.12791546406011753
	pesos_i(7155) := b"1111111111111111_1111111111111111_1101010011010111_1111000111101000"; -- -0.16857994170694102
	pesos_i(7156) := b"1111111111111111_1111111111111111_1101101010011000_1011001100011101"; -- -0.14610748807893834
	pesos_i(7157) := b"0000000000000000_0000000000000000_0000100010001110_1100101010010111"; -- 0.033428823431275664
	pesos_i(7158) := b"0000000000000000_0000000000000000_0000111011100101_0010011111111111"; -- 0.05818414665514693
	pesos_i(7159) := b"0000000000000000_0000000000000000_0000001111110101_0111110000001111"; -- 0.015464547842157329
	pesos_i(7160) := b"1111111111111111_1111111111111111_1111110000110110_0000111101000000"; -- -0.014800116373649919
	pesos_i(7161) := b"0000000000000000_0000000000000000_0001111001100101_1101101100110011"; -- 0.11874170295583224
	pesos_i(7162) := b"1111111111111111_1111111111111111_1110111111010000_1001011110000010"; -- -0.06322339139139256
	pesos_i(7163) := b"0000000000000000_0000000000000000_0001101110111101_0110111100011010"; -- 0.1083592832814737
	pesos_i(7164) := b"1111111111111111_1111111111111111_1101101011000101_1001100001110101"; -- -0.14542243139213207
	pesos_i(7165) := b"1111111111111111_1111111111111111_1110100001110101_1010001101110111"; -- -0.09195497844177601
	pesos_i(7166) := b"1111111111111111_1111111111111111_1111111001011000_0011001000111101"; -- -0.006466732179870117
	pesos_i(7167) := b"1111111111111111_1111111111111111_1111111110010000_1101000101010101"; -- -0.0016965073012276263
	pesos_i(7168) := b"0000000000000000_0000000000000000_0000010100001001_1101001010100010"; -- 0.019681133704712944
	pesos_i(7169) := b"0000000000000000_0000000000000000_0001110011111111_1000100011100110"; -- 0.11327415095979382
	pesos_i(7170) := b"1111111111111111_1111111111111111_1101101010000001_1100100010101000"; -- -0.1464571561251826
	pesos_i(7171) := b"1111111111111111_1111111111111111_1111010010111001_1110011001001101"; -- -0.044038396968885465
	pesos_i(7172) := b"1111111111111111_1111111111111111_1110100001010110_1100000101101100"; -- -0.09242621526363128
	pesos_i(7173) := b"1111111111111111_1111111111111111_1110110100001111_1011101000111111"; -- -0.07397876709640074
	pesos_i(7174) := b"0000000000000000_0000000000000000_0000111001101001_0000000010011010"; -- 0.0562897086985327
	pesos_i(7175) := b"1111111111111111_1111111111111111_1111001000000101_0010000111111011"; -- -0.05460918076178311
	pesos_i(7176) := b"0000000000000000_0000000000000000_0001001010110100_0101110100010100"; -- 0.07306462992581032
	pesos_i(7177) := b"1111111111111111_1111111111111111_1111101000111111_1011010110010001"; -- -0.022465374200776104
	pesos_i(7178) := b"1111111111111111_1111111111111111_1111100110010101_1100111100000111"; -- -0.025057850713381895
	pesos_i(7179) := b"1111111111111111_1111111111111111_1101111001000100_1101010101101001"; -- -0.13176218219626432
	pesos_i(7180) := b"0000000000000000_0000000000000000_0001110100110111_1100110111000110"; -- 0.11413274850837031
	pesos_i(7181) := b"0000000000000000_0000000000000000_0001101000000010_1010101010100010"; -- 0.10160318798785485
	pesos_i(7182) := b"0000000000000000_0000000000000000_0000110100101010_0010000011011001"; -- 0.05142407700631968
	pesos_i(7183) := b"0000000000000000_0000000000000000_0010100000011100_1100110000110100"; -- 0.15668941746109122
	pesos_i(7184) := b"0000000000000000_0000000000000000_0000011010011101_0010000111000000"; -- 0.025835141445944343
	pesos_i(7185) := b"0000000000000000_0000000000000000_0000001000111011_1110111100010111"; -- 0.00872701936100987
	pesos_i(7186) := b"1111111111111111_1111111111111111_1111000011110100_0100100110111011"; -- -0.058772460871613176
	pesos_i(7187) := b"0000000000000000_0000000000000000_0000100101010110_0100001010101100"; -- 0.03647247988612902
	pesos_i(7188) := b"1111111111111111_1111111111111111_1111000111000001_0001110111001110"; -- -0.055647027292006296
	pesos_i(7189) := b"0000000000000000_0000000000000000_0000001011100011_1111000001111100"; -- 0.011290579129716889
	pesos_i(7190) := b"1111111111111111_1111111111111111_1110100001101000_1101101001000100"; -- -0.09215007621827652
	pesos_i(7191) := b"0000000000000000_0000000000000000_0000110100100110_0101011100100101"; -- 0.05136627822561951
	pesos_i(7192) := b"1111111111111111_1111111111111111_1111110100000101_1111011111001110"; -- -0.01162768577982852
	pesos_i(7193) := b"0000000000000000_0000000000000000_0000111110100100_1001011111101110"; -- 0.061105247059293426
	pesos_i(7194) := b"1111111111111111_1111111111111111_1111110010000101_0101110010101000"; -- -0.01359005834806441
	pesos_i(7195) := b"1111111111111111_1111111111111111_1110111101011010_1010100001001010"; -- -0.06502292817005563
	pesos_i(7196) := b"0000000000000000_0000000000000000_0001010011011101_1001110010100111"; -- 0.08150652962182953
	pesos_i(7197) := b"0000000000000000_0000000000000000_0010010000000111_0010101010001100"; -- 0.14073434756865658
	pesos_i(7198) := b"1111111111111111_1111111111111111_1111101000100001_0010110100010100"; -- -0.022931273158316275
	pesos_i(7199) := b"0000000000000000_0000000000000000_0000010101111001_1001010010111010"; -- 0.021386428271390256
	pesos_i(7200) := b"0000000000000000_0000000000000000_0001000000101111_1110100111101110"; -- 0.06323110636205526
	pesos_i(7201) := b"0000000000000000_0000000000000000_0010010000111111_1110000100111110"; -- 0.1415997293029706
	pesos_i(7202) := b"0000000000000000_0000000000000000_0010010110111000_0110100101101000"; -- 0.1473451498704406
	pesos_i(7203) := b"0000000000000000_0000000000000000_0001010110001110_1101110010100000"; -- 0.08421114833354504
	pesos_i(7204) := b"1111111111111111_1111111111111111_1110001000101001_0010011111100001"; -- -0.1165595126027611
	pesos_i(7205) := b"0000000000000000_0000000000000000_0000100110100010_1100110010100111"; -- 0.03764037202207985
	pesos_i(7206) := b"0000000000000000_0000000000000000_0010011000101101_0101000000111001"; -- 0.1491289271134549
	pesos_i(7207) := b"1111111111111111_1111111111111111_1111011110100111_0101100000010001"; -- -0.03260278315153045
	pesos_i(7208) := b"0000000000000000_0000000000000000_0001100101010110_0011110001010000"; -- 0.09897210083600458
	pesos_i(7209) := b"0000000000000000_0000000000000000_0001100110010010_1101100000100101"; -- 0.09989691636234777
	pesos_i(7210) := b"0000000000000000_0000000000000000_0001010110011110_0001001110111101"; -- 0.08444331521786595
	pesos_i(7211) := b"1111111111111111_1111111111111111_1101001101111000_1001110101010010"; -- -0.17394081834974176
	pesos_i(7212) := b"0000000000000000_0000000000000000_0000001111111111_0011101000000010"; -- 0.015613198763775281
	pesos_i(7213) := b"0000000000000000_0000000000000000_0001011101011100_0000100101111101"; -- 0.09124812407972312
	pesos_i(7214) := b"0000000000000000_0000000000000000_0001001100001100_1110100000101101"; -- 0.07441569429468034
	pesos_i(7215) := b"0000000000000000_0000000000000000_0000010010111001_1100100011011000"; -- 0.01845984712974398
	pesos_i(7216) := b"1111111111111111_1111111111111111_1110010100111000_0010101100000100"; -- -0.10461169399119377
	pesos_i(7217) := b"1111111111111111_1111111111111111_1110000000100011_0010000100101011"; -- -0.12446396543946452
	pesos_i(7218) := b"0000000000000000_0000000000000000_0001000111100100_0100101100101111"; -- 0.06988973513924489
	pesos_i(7219) := b"0000000000000000_0000000000000000_0000111011001000_1111001110111110"; -- 0.057753786053169456
	pesos_i(7220) := b"0000000000000000_0000000000000000_0000101011111010_1000111111100001"; -- 0.04288577310047403
	pesos_i(7221) := b"1111111111111111_1111111111111111_1110000010100011_1110101000100101"; -- -0.12249886121582193
	pesos_i(7222) := b"0000000000000000_0000000000000000_0000010111110100_0000010100110000"; -- 0.023254703635939084
	pesos_i(7223) := b"1111111111111111_1111111111111111_1111011111111110_1000011010101000"; -- -0.031272491327652335
	pesos_i(7224) := b"1111111111111111_1111111111111111_1101101000111111_1000100110101110"; -- -0.14746798983495624
	pesos_i(7225) := b"0000000000000000_0000000000000000_0001110100001111_1001010101000111"; -- 0.11351902954436142
	pesos_i(7226) := b"0000000000000000_0000000000000000_0001100010110011_1011001010111110"; -- 0.0964919771276896
	pesos_i(7227) := b"1111111111111111_1111111111111111_1111101011010101_1100101001011100"; -- -0.020175316428162567
	pesos_i(7228) := b"0000000000000000_0000000000000000_0010000101000101_0010111001011010"; -- 0.12996186927117462
	pesos_i(7229) := b"1111111111111111_1111111111111111_1110110110011001_1011011011110111"; -- -0.07187324966758125
	pesos_i(7230) := b"1111111111111111_1111111111111111_1111001100001101_0010011010110110"; -- -0.05058057840528269
	pesos_i(7231) := b"1111111111111111_1111111111111111_1111110001110100_0111101101000101"; -- -0.013847632915836024
	pesos_i(7232) := b"0000000000000000_0000000000000000_0010100101111111_0111011001110011"; -- 0.16210117627288015
	pesos_i(7233) := b"1111111111111111_1111111111111111_1111001011011100_1111101011000001"; -- -0.051315620284929385
	pesos_i(7234) := b"0000000000000000_0000000000000000_0010011001111110_1111111001001101"; -- 0.15037526499459297
	pesos_i(7235) := b"0000000000000000_0000000000000000_0010011011001010_0001111010100000"; -- 0.15152160069686135
	pesos_i(7236) := b"0000000000000000_0000000000000000_0000100011100010_0101101111111100"; -- 0.03470396899509881
	pesos_i(7237) := b"1111111111111111_1111111111111111_1111101111010000_1010011101011010"; -- -0.016347447009081303
	pesos_i(7238) := b"1111111111111111_1111111111111111_1101100111110010_0010011111000010"; -- -0.1486487532074595
	pesos_i(7239) := b"0000000000000000_0000000000000000_0000110100111000_0101101110100101"; -- 0.05164120466232088
	pesos_i(7240) := b"1111111111111111_1111111111111111_1101111011011001_1011001011101101"; -- -0.12949067806172285
	pesos_i(7241) := b"0000000000000000_0000000000000000_0000100101100001_1100011001101100"; -- 0.03664817939780125
	pesos_i(7242) := b"0000000000000000_0000000000000000_0001110000010110_0001011001010110"; -- 0.10971202472152175
	pesos_i(7243) := b"1111111111111111_1111111111111111_1101011101100001_1110000101000001"; -- -0.15866272123232947
	pesos_i(7244) := b"1111111111111111_1111111111111111_1101100000010100_0101010001110010"; -- -0.15593979095316848
	pesos_i(7245) := b"0000000000000000_0000000000000000_0001010100000100_1110010000111010"; -- 0.08210588840630473
	pesos_i(7246) := b"1111111111111111_1111111111111111_1101011001111011_1011011100000011"; -- -0.162174760532663
	pesos_i(7247) := b"0000000000000000_0000000000000000_0001011010101111_0100011000000100"; -- 0.0886119613031503
	pesos_i(7248) := b"0000000000000000_0000000000000000_0001000111000101_1101101011001011"; -- 0.06942527251254735
	pesos_i(7249) := b"1111111111111111_1111111111111111_1101011101100010_1101000010111011"; -- -0.1586484473674965
	pesos_i(7250) := b"0000000000000000_0000000000000000_0000101100001001_1111011110111111"; -- 0.04312084598739895
	pesos_i(7251) := b"1111111111111111_1111111111111111_1111000001110011_0101100011001011"; -- -0.060739946811745
	pesos_i(7252) := b"0000000000000000_0000000000000000_0000111011110000_0101110011001111"; -- 0.058355141131881914
	pesos_i(7253) := b"0000000000000000_0000000000000000_0001011000010101_1000011111100110"; -- 0.08626603469551719
	pesos_i(7254) := b"0000000000000000_0000000000000000_0000111010110100_0001000110011110"; -- 0.05743513208414553
	pesos_i(7255) := b"1111111111111111_1111111111111111_1110110010110101_1011010000110111"; -- -0.07535241765111049
	pesos_i(7256) := b"0000000000000000_0000000000000000_0001001010011010_0011011110011000"; -- 0.07266566714967591
	pesos_i(7257) := b"1111111111111111_1111111111111111_1110011100001001_0001010001101011"; -- -0.0975177039179404
	pesos_i(7258) := b"0000000000000000_0000000000000000_0000101110011011_0111010100111001"; -- 0.045340849361096905
	pesos_i(7259) := b"1111111111111111_1111111111111111_1111010101000100_0011011010001110"; -- -0.04192790070824299
	pesos_i(7260) := b"1111111111111111_1111111111111111_1101100101011101_1010101100010000"; -- -0.1509144865940118
	pesos_i(7261) := b"0000000000000000_0000000000000000_0001011100000010_0001110101000110"; -- 0.08987601234435037
	pesos_i(7262) := b"1111111111111111_1111111111111111_1111001100110011_1101000110000101"; -- -0.04999056348327774
	pesos_i(7263) := b"0000000000000000_0000000000000000_0000001100111001_0001011101101101"; -- 0.012589897243994258
	pesos_i(7264) := b"1111111111111111_1111111111111111_1101100010100101_1111100001001111"; -- -0.15371749948229285
	pesos_i(7265) := b"0000000000000000_0000000000000000_0001100011110011_0110010000011111"; -- 0.09746385339685007
	pesos_i(7266) := b"0000000000000000_0000000000000000_0000111011100011_1011011000011000"; -- 0.05816209867424788
	pesos_i(7267) := b"1111111111111111_1111111111111111_1101100100111001_1110110100111101"; -- -0.1514598585722758
	pesos_i(7268) := b"1111111111111111_1111111111111111_1101100001011010_1110010000011000"; -- -0.15486311356514318
	pesos_i(7269) := b"1111111111111111_1111111111111111_1111000010100010_1110101000101000"; -- -0.060014119436119964
	pesos_i(7270) := b"1111111111111111_1111111111111111_1110001001101001_1100110101110100"; -- -0.11557308117743961
	pesos_i(7271) := b"1111111111111111_1111111111111111_1111011000111001_0101101100111101"; -- -0.03818731079898652
	pesos_i(7272) := b"1111111111111111_1111111111111111_1110110111101100_1100011010000000"; -- -0.07060584415539295
	pesos_i(7273) := b"0000000000000000_0000000000000000_0001101000011101_1011101001111011"; -- 0.10201612010090938
	pesos_i(7274) := b"1111111111111111_1111111111111111_1111010011110110_1110010011011100"; -- -0.04310769670724933
	pesos_i(7275) := b"1111111111111111_1111111111111111_1101000000111000_1101011100111011"; -- -0.18663267904063546
	pesos_i(7276) := b"0000000000000000_0000000000000000_0000111101011110_0100101000001000"; -- 0.060032488770772004
	pesos_i(7277) := b"0000000000000000_0000000000000000_0000011110011011_1110101100111010"; -- 0.029722882865484433
	pesos_i(7278) := b"0000000000000000_0000000000000000_0010101011010110_1001101011111101"; -- 0.16733711882586136
	pesos_i(7279) := b"0000000000000000_0000000000000000_0001100100010111_0100101011000110"; -- 0.09801165889832673
	pesos_i(7280) := b"0000000000000000_0000000000000000_0001010000101100_0110110010011110"; -- 0.07880286087661934
	pesos_i(7281) := b"0000000000000000_0000000000000000_0000111011110000_0011011010010101"; -- 0.058352862643442485
	pesos_i(7282) := b"1111111111111111_1111111111111111_1111111011000000_0001100001000100"; -- -0.004881366170711039
	pesos_i(7283) := b"0000000000000000_0000000000000000_0001000101101010_1111110001111010"; -- 0.06803873032608977
	pesos_i(7284) := b"0000000000000000_0000000000000000_0010001100100101_0100101101011000"; -- 0.137287815948474
	pesos_i(7285) := b"0000000000000000_0000000000000000_0010001111011111_0100011000111111"; -- 0.14012564693321547
	pesos_i(7286) := b"0000000000000000_0000000000000000_0001101000110000_1010011011101011"; -- 0.1023048710279634
	pesos_i(7287) := b"0000000000000000_0000000000000000_0000000010101111_0100101010110000"; -- 0.002674739799714783
	pesos_i(7288) := b"1111111111111111_1111111111111111_1111110110101110_1111111000101100"; -- -0.009048570885301144
	pesos_i(7289) := b"1111111111111111_1111111111111111_1110000110101010_0001001001110000"; -- -0.11849865680339386
	pesos_i(7290) := b"1111111111111111_1111111111111111_1111001001010110_1011101101001111"; -- -0.053364079699053546
	pesos_i(7291) := b"1111111111111111_1111111111111111_1111001110001000_1111010001000011"; -- -0.04869149554242176
	pesos_i(7292) := b"1111111111111111_1111111111111111_1110111001110001_0011000010111000"; -- -0.06858535298863008
	pesos_i(7293) := b"0000000000000000_0000000000000000_0001110111110111_1000001000010101"; -- 0.11705792447981808
	pesos_i(7294) := b"0000000000000000_0000000000000000_0010101010000011_0100110110000000"; -- 0.1660660207987696
	pesos_i(7295) := b"0000000000000000_0000000000000000_0011011010000110_0111001010010001"; -- 0.21298900647814506
	pesos_i(7296) := b"1111111111111111_1111111111111111_1110010111010011_1110110111000111"; -- -0.10223497290504927
	pesos_i(7297) := b"1111111111111111_1111111111111111_1111001100111110_0010110101001001"; -- -0.049832505795249706
	pesos_i(7298) := b"0000000000000000_0000000000000000_0001110101010010_1001000000111101"; -- 0.11454106795898013
	pesos_i(7299) := b"0000000000000000_0000000000000000_0001101000110000_1001110110010001"; -- 0.10230431353271725
	pesos_i(7300) := b"1111111111111111_1111111111111111_1111010110110010_0000110101000011"; -- -0.040251895150617875
	pesos_i(7301) := b"1111111111111111_1111111111111111_1101110101101100_1001100001001110"; -- -0.13506172276164252
	pesos_i(7302) := b"1111111111111111_1111111111111111_1111011100001010_1001111111100100"; -- -0.03499413185859607
	pesos_i(7303) := b"0000000000000000_0000000000000000_0010011100001110_0001111010010011"; -- 0.15255919532320278
	pesos_i(7304) := b"0000000000000000_0000000000000000_0000101101000101_0011101100001011"; -- 0.04402512571184226
	pesos_i(7305) := b"0000000000000000_0000000000000000_0000111000110101_0011011110000110"; -- 0.05549952525750424
	pesos_i(7306) := b"1111111111111111_1111111111111111_1101111001001111_0101100001110101"; -- -0.13160178316607485
	pesos_i(7307) := b"0000000000000000_0000000000000000_0010010011000101_1000101011101000"; -- 0.14363926091047588
	pesos_i(7308) := b"0000000000000000_0000000000000000_0000011110100100_1110001111100000"; -- 0.02985977372053422
	pesos_i(7309) := b"0000000000000000_0000000000000000_0001001100110100_0010111010001000"; -- 0.07501498044515768
	pesos_i(7310) := b"1111111111111111_1111111111111111_1110101111101100_1010101101000010"; -- -0.07841996796007883
	pesos_i(7311) := b"1111111111111111_1111111111111111_1101100011111111_0101111101001111"; -- -0.15235332800192458
	pesos_i(7312) := b"1111111111111111_1111111111111111_1111011010001011_0010010111010101"; -- -0.03693927333681296
	pesos_i(7313) := b"1111111111111111_1111111111111111_1101111001110110_0000001000001100"; -- -0.13101184087148923
	pesos_i(7314) := b"0000000000000000_0000000000000000_0001011000100111_0011111011111011"; -- 0.0865363467125698
	pesos_i(7315) := b"1111111111111111_1111111111111111_1101101010100110_0110011010001100"; -- -0.14589842879434373
	pesos_i(7316) := b"0000000000000000_0000000000000000_0000100110110110_1110001000101100"; -- 0.037946830586652026
	pesos_i(7317) := b"0000000000000000_0000000000000000_0010001101001111_1001111100010010"; -- 0.13793367555203337
	pesos_i(7318) := b"1111111111111111_1111111111111111_1110100011000001_0110110101001000"; -- -0.09079854012812233
	pesos_i(7319) := b"1111111111111111_1111111111111111_1111101011101010_0000110010100101"; -- -0.01986618960646893
	pesos_i(7320) := b"0000000000000000_0000000000000000_0000000010111010_1101010100111100"; -- 0.002850844549442003
	pesos_i(7321) := b"1111111111111111_1111111111111111_1100111011001001_0100100110011001"; -- -0.19224109664161002
	pesos_i(7322) := b"0000000000000000_0000000000000000_0010011100101000_1100111000011001"; -- 0.15296638593727072
	pesos_i(7323) := b"0000000000000000_0000000000000000_0001001111110110_0100001011110001"; -- 0.07797640213803678
	pesos_i(7324) := b"1111111111111111_1111111111111111_1110010010110110_1100100111011001"; -- -0.10658586944717928
	pesos_i(7325) := b"0000000000000000_0000000000000000_0000100000011010_1111111001000100"; -- 0.03166188381194069
	pesos_i(7326) := b"0000000000000000_0000000000000000_0001111001011101_0001110011000011"; -- 0.11860828172409203
	pesos_i(7327) := b"1111111111111111_1111111111111111_1101100000011010_1101010101000101"; -- -0.1558405595564116
	pesos_i(7328) := b"0000000000000000_0000000000000000_0000110000101000_1001010111101110"; -- 0.04749428795339036
	pesos_i(7329) := b"1111111111111111_1111111111111111_1111010100000001_0101111111001001"; -- -0.04294778208151374
	pesos_i(7330) := b"0000000000000000_0000000000000000_0001001110001010_0000001001100100"; -- 0.07632460533054504
	pesos_i(7331) := b"1111111111111111_1111111111111111_1101011000011110_1101001001110011"; -- -0.16359219266784017
	pesos_i(7332) := b"0000000000000000_0000000000000000_0010100000000011_0101111000101011"; -- 0.15630138912158528
	pesos_i(7333) := b"1111111111111111_1111111111111111_1100111111010010_1011100001011010"; -- -0.18819091599853802
	pesos_i(7334) := b"0000000000000000_0000000000000000_0001000100100000_1111010100111001"; -- 0.06690914758600337
	pesos_i(7335) := b"1111111111111111_1111111111111111_1101010001111010_0110011111001110"; -- -0.17000724052918328
	pesos_i(7336) := b"0000000000000000_0000000000000000_0000011101110100_0101110111011101"; -- 0.029119364186277974
	pesos_i(7337) := b"0000000000000000_0000000000000000_0000110100000011_0001010100101000"; -- 0.050828287332008136
	pesos_i(7338) := b"0000000000000000_0000000000000000_0000110101110001_0110010101100110"; -- 0.052511537061728314
	pesos_i(7339) := b"0000000000000000_0000000000000000_0000010001011000_1000011011101111"; -- 0.016975816081653536
	pesos_i(7340) := b"0000000000000000_0000000000000000_0001010111010000_1110110101111011"; -- 0.08521923304987213
	pesos_i(7341) := b"0000000000000000_0000000000000000_0010001101110100_0101100010000011"; -- 0.13849404517486327
	pesos_i(7342) := b"1111111111111111_1111111111111111_1111011011011001_0000110000011010"; -- -0.03575062141271958
	pesos_i(7343) := b"1111111111111111_1111111111111111_1101011101110101_0101011111110101"; -- -0.1583657290871084
	pesos_i(7344) := b"0000000000000000_0000000000000000_0001100010010111_0101000100100101"; -- 0.09605891378892192
	pesos_i(7345) := b"0000000000000000_0000000000000000_0000111101010000_1111100101001100"; -- 0.059829312391218775
	pesos_i(7346) := b"1111111111111111_1111111111111111_1110111000111010_1111010010011111"; -- -0.06941290956484404
	pesos_i(7347) := b"0000000000000000_0000000000000000_0010100110010100_1011110010100011"; -- 0.16242579434013024
	pesos_i(7348) := b"1111111111111111_1111111111111111_1101011011011000_1001101111111111"; -- -0.16075730345104228
	pesos_i(7349) := b"1111111111111111_1111111111111111_1110111000101110_1100100011110010"; -- -0.06959861836329718
	pesos_i(7350) := b"0000000000000000_0000000000000000_0001011010101001_1110100001000011"; -- 0.08853007922083277
	pesos_i(7351) := b"1111111111111111_1111111111111111_1111001011000111_0000010101010101"; -- -0.05165068315424009
	pesos_i(7352) := b"1111111111111111_1111111111111111_1111101010010100_1100110100111110"; -- -0.021166965838508356
	pesos_i(7353) := b"0000000000000000_0000000000000000_0000101000101000_0011010101011111"; -- 0.03967603264209638
	pesos_i(7354) := b"1111111111111111_1111111111111111_1101111000001100_1001100110111101"; -- -0.1326202309861381
	pesos_i(7355) := b"1111111111111111_1111111111111111_1111111111100011_1100001000110111"; -- -0.0004309288687389046
	pesos_i(7356) := b"1111111111111111_1111111111111111_1111001101110001_1010100100111001"; -- -0.04904692048913072
	pesos_i(7357) := b"1111111111111111_1111111111111111_1110101111110001_1011010011110001"; -- -0.07834309685014913
	pesos_i(7358) := b"0000000000000000_0000000000000000_0000110001110011_0000001111011010"; -- 0.04862999020186956
	pesos_i(7359) := b"1111111111111111_1111111111111111_1110100001010101_0011101101010110"; -- -0.09244946627879448
	pesos_i(7360) := b"0000000000000000_0000000000000000_0001001000011011_0001011110000100"; -- 0.07072588893665299
	pesos_i(7361) := b"1111111111111111_1111111111111111_1110000111000001_1110011011011000"; -- -0.11813504439345057
	pesos_i(7362) := b"1111111111111111_1111111111111111_1101011010101011_0111010110111110"; -- -0.1614462291246934
	pesos_i(7363) := b"0000000000000000_0000000000000000_0000101100011011_1101110101010111"; -- 0.04339393010916429
	pesos_i(7364) := b"1111111111111111_1111111111111111_1101100010011000_0010011011011010"; -- -0.15392834829231475
	pesos_i(7365) := b"0000000000000000_0000000000000000_0010111010110000_1101001011100001"; -- 0.18238561631296926
	pesos_i(7366) := b"1111111111111111_1111111111111111_1110100011101110_1101101000101000"; -- -0.09010540507859231
	pesos_i(7367) := b"1111111111111111_1111111111111111_1111010001110001_1100010000001101"; -- -0.045139071211760695
	pesos_i(7368) := b"1111111111111111_1111111111111111_1110011100110100_0011010110111001"; -- -0.09685959082783936
	pesos_i(7369) := b"1111111111111111_1111111111111111_1110000010001111_1001001100011100"; -- -0.12280922468292133
	pesos_i(7370) := b"1111111111111111_1111111111111111_1110010001111101_1100100001001100"; -- -0.10745571270070359
	pesos_i(7371) := b"0000000000000000_0000000000000000_0001101000011010_0001010100111010"; -- 0.1019604936229959
	pesos_i(7372) := b"1111111111111111_1111111111111111_1101110011001111_1100001100000000"; -- -0.13745480776435087
	pesos_i(7373) := b"1111111111111111_1111111111111111_1110110010010001_0011010100011001"; -- -0.07590931068182384
	pesos_i(7374) := b"1111111111111111_1111111111111111_1101100010100101_1000101110100001"; -- -0.15372397729022363
	pesos_i(7375) := b"1111111111111111_1111111111111111_1110000010100010_1101110011110000"; -- -0.12251490719992818
	pesos_i(7376) := b"1111111111111111_1111111111111111_1111000100111101_1001100000001101"; -- -0.057653900820160586
	pesos_i(7377) := b"1111111111111111_1111111111111111_1111110010011010_0101101110101001"; -- -0.013269683137994138
	pesos_i(7378) := b"1111111111111111_1111111111111111_1110011100001101_0000011101000101"; -- -0.09745745247339731
	pesos_i(7379) := b"1111111111111111_1111111111111111_1111100001111111_0101011010110100"; -- -0.029306965769984244
	pesos_i(7380) := b"1111111111111111_1111111111111111_1111010110010100_0010011110000001"; -- -0.04070809468731077
	pesos_i(7381) := b"1111111111111111_1111111111111111_1111111000001111_0011110001110101"; -- -0.007580014588874251
	pesos_i(7382) := b"1111111111111111_1111111111111111_1110100111001000_1011001101011110"; -- -0.0867813009952308
	pesos_i(7383) := b"1111111111111111_1111111111111111_1110011011111011_0111000011000100"; -- -0.09772582250744526
	pesos_i(7384) := b"0000000000000000_0000000000000000_0000000101000100_1111010100010010"; -- 0.004958455017994455
	pesos_i(7385) := b"1111111111111111_1111111111111111_1110111000111110_1110001100101111"; -- -0.0693529138140938
	pesos_i(7386) := b"1111111111111111_1111111111111111_1101100101100000_0000100100100110"; -- -0.15087836107074326
	pesos_i(7387) := b"0000000000000000_0000000000000000_0010011100101000_0100011100001100"; -- 0.15295833618173216
	pesos_i(7388) := b"1111111111111111_1111111111111111_1101111100101011_1100001000010011"; -- -0.1282385542643068
	pesos_i(7389) := b"0000000000000000_0000000000000000_0010010000100111_0011000010110100"; -- 0.14122299562976992
	pesos_i(7390) := b"0000000000000000_0000000000000000_0001000101101010_1101001101000110"; -- 0.068036274560042
	pesos_i(7391) := b"1111111111111111_1111111111111111_1110011010101100_0000000110100110"; -- -0.09893788997205928
	pesos_i(7392) := b"1111111111111111_1111111111111111_1111110111110110_1110011011000101"; -- -0.007951332985123155
	pesos_i(7393) := b"1111111111111111_1111111111111111_1111111110100101_0100010011001011"; -- -0.0013844494414845092
	pesos_i(7394) := b"1111111111111111_1111111111111111_1111010000101100_1100000001100101"; -- -0.04619214560643727
	pesos_i(7395) := b"1111111111111111_1111111111111111_1101011100101010_0001010110100010"; -- -0.1595140913366086
	pesos_i(7396) := b"1111111111111111_1111111111111111_1101110101110100_0010000101001100"; -- -0.13494674587391656
	pesos_i(7397) := b"1111111111111111_1111111111111111_1110100010010010_1001001001110000"; -- -0.09151348853689252
	pesos_i(7398) := b"1111111111111111_1111111111111111_1110001000101111_0000011010000101"; -- -0.11646994821305033
	pesos_i(7399) := b"1111111111111111_1111111111111111_1110001001011001_1000001100111000"; -- -0.11582164646432483
	pesos_i(7400) := b"0000000000000000_0000000000000000_0010000101100101_1001101011010110"; -- 0.13045661673130174
	pesos_i(7401) := b"1111111111111111_1111111111111111_1110100011010100_0000101111011011"; -- -0.09051443016520426
	pesos_i(7402) := b"0000000000000000_0000000000000000_0000010101101110_0000011111010101"; -- 0.021210183653288302
	pesos_i(7403) := b"1111111111111111_1111111111111111_1111110101111010_1000110100111011"; -- -0.009848759840553086
	pesos_i(7404) := b"0000000000000000_0000000000000000_0010110100000010_0110010111000100"; -- 0.17581783335755238
	pesos_i(7405) := b"1111111111111111_1111111111111111_1111001011101010_1111000011110110"; -- -0.05110258100180506
	pesos_i(7406) := b"0000000000000000_0000000000000000_0001011110011010_0111001101110011"; -- 0.09220048479917647
	pesos_i(7407) := b"0000000000000000_0000000000000000_0000110010101111_0010101000111101"; -- 0.049547805663412325
	pesos_i(7408) := b"1111111111111111_1111111111111111_1111101010011010_0100101011110001"; -- -0.021083179529864132
	pesos_i(7409) := b"0000000000000000_0000000000000000_0000101001110101_0011100000101011"; -- 0.04085112611006615
	pesos_i(7410) := b"1111111111111111_1111111111111111_1111100110101000_0100001001101101"; -- -0.02477631406534268
	pesos_i(7411) := b"0000000000000000_0000000000000000_0000001100110010_1100101101011011"; -- 0.012493810343454736
	pesos_i(7412) := b"0000000000000000_0000000000000000_0000111011110011_0100101101010011"; -- 0.058399875431856776
	pesos_i(7413) := b"0000000000000000_0000000000000000_0000010101111001_1111100010111001"; -- 0.021392388423337325
	pesos_i(7414) := b"1111111111111111_1111111111111111_1110000100001000_1111101110001001"; -- -0.12095668705176593
	pesos_i(7415) := b"0000000000000000_0000000000000000_0000101000100110_0011010001101111"; -- 0.03964545916214459
	pesos_i(7416) := b"1111111111111111_1111111111111111_1101011011110001_0010110000000111"; -- -0.1603825076670986
	pesos_i(7417) := b"1111111111111111_1111111111111111_1110101011100001_0001010100111101"; -- -0.08250300655469132
	pesos_i(7418) := b"1111111111111111_1111111111111111_1111100100100000_1001111010110111"; -- -0.026846008550445565
	pesos_i(7419) := b"0000000000000000_0000000000000000_0010001011100011_0101010010100010"; -- 0.13628128966249206
	pesos_i(7420) := b"1111111111111111_1111111111111111_1110000110001010_1011000000001101"; -- -0.11897754355387873
	pesos_i(7421) := b"0000000000000000_0000000000000000_0010101000011101_0100000010010100"; -- 0.16450885405567606
	pesos_i(7422) := b"1111111111111111_1111111111111111_1110110110011110_0011101100100010"; -- -0.07180433681122342
	pesos_i(7423) := b"1111111111111111_1111111111111111_1111111111101111_0110110000011101"; -- -0.00025295539690426176
	pesos_i(7424) := b"0000000000000000_0000000000000000_0001111001110001_0100111001101111"; -- 0.11891641808362599
	pesos_i(7425) := b"0000000000000000_0000000000000000_0000110110011110_1010010100001001"; -- 0.053201975447658686
	pesos_i(7426) := b"1111111111111111_1111111111111111_1111000011101111_0110101111101001"; -- -0.05884671752182278
	pesos_i(7427) := b"0000000000000000_0000000000000000_0010100111011010_1100000110001101"; -- 0.16349420248282415
	pesos_i(7428) := b"1111111111111111_1111111111111111_1111011011111101_0010100010100101"; -- -0.03519960387671071
	pesos_i(7429) := b"1111111111111111_1111111111111111_1101100101111001_0111101101000010"; -- -0.1504900897059627
	pesos_i(7430) := b"0000000000000000_0000000000000000_0000111110100110_1011100110001000"; -- 0.06113776749324015
	pesos_i(7431) := b"1111111111111111_1111111111111111_1101110011111101_1101110100111010"; -- -0.13675134019812993
	pesos_i(7432) := b"0000000000000000_0000000000000000_0000011110110001_0010100111101111"; -- 0.030047055009793395
	pesos_i(7433) := b"0000000000000000_0000000000000000_0001100101001111_1110001111001010"; -- 0.09887527167721331
	pesos_i(7434) := b"0000000000000000_0000000000000000_0000100111110010_0011010001110110"; -- 0.038852003762688166
	pesos_i(7435) := b"1111111111111111_1111111111111111_1111011000011011_1011011110100011"; -- -0.03863956711062472
	pesos_i(7436) := b"0000000000000000_0000000000000000_0001000011111011_0111001100101011"; -- 0.0663368204898439
	pesos_i(7437) := b"0000000000000000_0000000000000000_0010101001010010_0111111100010110"; -- 0.1653212956318691
	pesos_i(7438) := b"1111111111111111_1111111111111111_1111001001011111_1001110000001100"; -- -0.05322861400323831
	pesos_i(7439) := b"1111111111111111_1111111111111111_1110110001010111_1101101100000111"; -- -0.07678443026674989
	pesos_i(7440) := b"1111111111111111_1111111111111111_1111100110101111_0111101111111101"; -- -0.024666071679013024
	pesos_i(7441) := b"1111111111111111_1111111111111111_1111100011101000_1010101110100101"; -- -0.0276997300718575
	pesos_i(7442) := b"0000000000000000_0000000000000000_0001011011101011_1001001000010110"; -- 0.08953202275408491
	pesos_i(7443) := b"1111111111111111_1111111111111111_1101001111101001_0100110111101110"; -- -0.17222130722741133
	pesos_i(7444) := b"1111111111111111_1111111111111111_1110011101101000_0010010011010010"; -- -0.09606714136444203
	pesos_i(7445) := b"0000000000000000_0000000000000000_0001111111011110_0110111100100001"; -- 0.1244878248947544
	pesos_i(7446) := b"1111111111111111_1111111111111111_1111001110001100_0111001000000000"; -- -0.04863822457814978
	pesos_i(7447) := b"0000000000000000_0000000000000000_0000110010101011_0110011110101010"; -- 0.0494904318690462
	pesos_i(7448) := b"1111111111111111_1111111111111111_1101111010011101_0001000100000100"; -- -0.1304158559328034
	pesos_i(7449) := b"0000000000000000_0000000000000000_0010000000000001_0010000001001000"; -- 0.12501718297302322
	pesos_i(7450) := b"0000000000000000_0000000000000000_0000101010110110_1000110111000011"; -- 0.04184804924239784
	pesos_i(7451) := b"1111111111111111_1111111111111111_1110001100010010_0101010100100010"; -- -0.11300151746555899
	pesos_i(7452) := b"0000000000000000_0000000000000000_0001110100011000_1000011000111011"; -- 0.11365546167048991
	pesos_i(7453) := b"0000000000000000_0000000000000000_0000100010100100_0111010100111001"; -- 0.033759428497485734
	pesos_i(7454) := b"0000000000000000_0000000000000000_0001110111010011_0011111000101000"; -- 0.11650455930407395
	pesos_i(7455) := b"0000000000000000_0000000000000000_0001001110010111_1100111001000000"; -- 0.07653512065816978
	pesos_i(7456) := b"1111111111111111_1111111111111111_1111010100011010_0001101101000101"; -- -0.04257039618156919
	pesos_i(7457) := b"0000000000000000_0000000000000000_0001101110000111_1110001000110010"; -- 0.10754216876569798
	pesos_i(7458) := b"0000000000000000_0000000000000000_0001001100100110_1110001100101011"; -- 0.07481212429228071
	pesos_i(7459) := b"0000000000000000_0000000000000000_0010101100011011_0100010101110000"; -- 0.16838487607837782
	pesos_i(7460) := b"0000000000000000_0000000000000000_0000110100001000_0011111110100011"; -- 0.05090711339815413
	pesos_i(7461) := b"1111111111111111_1111111111111111_1110111011101101_0001011010011011"; -- -0.06669481948783335
	pesos_i(7462) := b"1111111111111111_1111111111111111_1101101001111101_1001110001010010"; -- -0.14652083402877009
	pesos_i(7463) := b"0000000000000000_0000000000000000_0010110100111100_0000111110100011"; -- 0.1766977093491948
	pesos_i(7464) := b"0000000000000000_0000000000000000_0000110110010100_1110010101010110"; -- 0.0530532202583853
	pesos_i(7465) := b"0000000000000000_0000000000000000_0000111101100101_0010110100001001"; -- 0.06013757210078842
	pesos_i(7466) := b"1111111111111111_1111111111111111_1110101110101010_1101110000101111"; -- -0.07942413186786146
	pesos_i(7467) := b"0000000000000000_0000000000000000_0010000110111001_1111100111000100"; -- 0.13174401319390658
	pesos_i(7468) := b"1111111111111111_1111111111111111_1110011000011000_1000001000011101"; -- -0.10118853360662225
	pesos_i(7469) := b"1111111111111111_1111111111111111_1110111001011110_1011111100011101"; -- -0.06886678268735152
	pesos_i(7470) := b"1111111111111111_1111111111111111_1111000111010001_0110000110010010"; -- -0.05539884739383747
	pesos_i(7471) := b"1111111111111111_1111111111111111_1111100101110101_0111010101001100"; -- -0.02555148035644086
	pesos_i(7472) := b"0000000000000000_0000000000000000_0010001101001000_1011000011001110"; -- 0.1378279212332252
	pesos_i(7473) := b"1111111111111111_1111111111111111_1111010101000110_1010100100100001"; -- -0.04189055378941243
	pesos_i(7474) := b"0000000000000000_0000000000000000_0001100100111110_0000011100100100"; -- 0.09860272061566852
	pesos_i(7475) := b"1111111111111111_1111111111111111_1111001100100001_1000010100000110"; -- -0.05026978110182509
	pesos_i(7476) := b"1111111111111111_1111111111111111_1111110001101011_1111000110101110"; -- -0.013977904335489861
	pesos_i(7477) := b"1111111111111111_1111111111111111_1111111000110111_0000001011101000"; -- -0.006973093411858123
	pesos_i(7478) := b"1111111111111111_1111111111111111_1101010101101111_0000100111111001"; -- -0.16627443005141465
	pesos_i(7479) := b"0000000000000000_0000000000000000_0010111111111010_1000000100110001"; -- 0.1874161475768395
	pesos_i(7480) := b"0000000000000000_0000000000000000_0001010101011000_0100101100100111"; -- 0.08337850282188583
	pesos_i(7481) := b"1111111111111111_1111111111111111_1111101010000100_0001011101111101"; -- -0.02142193974413791
	pesos_i(7482) := b"1111111111111111_1111111111111111_1110101011011110_1100010001101010"; -- -0.08253834163254008
	pesos_i(7483) := b"1111111111111111_1111111111111111_1111111001100001_1100111111111000"; -- -0.006320001500212425
	pesos_i(7484) := b"0000000000000000_0000000000000000_0001011100001011_0110100111100101"; -- 0.09001790839493494
	pesos_i(7485) := b"0000000000000000_0000000000000000_0010101100101111_0111001001000001"; -- 0.1686927231527023
	pesos_i(7486) := b"0000000000000000_0000000000000000_0010110001100111_1111111011111111"; -- 0.1734618541701562
	pesos_i(7487) := b"1111111111111111_1111111111111111_1110001010110111_1111101000011001"; -- -0.11438023465485364
	pesos_i(7488) := b"0000000000000000_0000000000000000_0000111001111100_1101101100101101"; -- 0.05659265362716526
	pesos_i(7489) := b"0000000000000000_0000000000000000_0000000101010011_1101110001011110"; -- 0.005185864446175993
	pesos_i(7490) := b"1111111111111111_1111111111111111_1110101010111101_1010010101100001"; -- -0.0830437315368631
	pesos_i(7491) := b"0000000000000000_0000000000000000_0010010000100011_1001001100011010"; -- 0.1411678256125947
	pesos_i(7492) := b"1111111111111111_1111111111111111_1111001111000110_0101011011101101"; -- -0.047754828681716044
	pesos_i(7493) := b"0000000000000000_0000000000000000_0001010010110001_1100010000011001"; -- 0.08083749391100578
	pesos_i(7494) := b"1111111111111111_1111111111111111_1101111110101100_0111010110101110"; -- -0.12627472409425003
	pesos_i(7495) := b"1111111111111111_1111111111111111_1111100110110010_1111101011010110"; -- -0.024612734639926442
	pesos_i(7496) := b"0000000000000000_0000000000000000_0010110000100001_1101111001100101"; -- 0.17239179580802033
	pesos_i(7497) := b"0000000000000000_0000000000000000_0001111111000110_1000101100001101"; -- 0.12412327839988553
	pesos_i(7498) := b"1111111111111111_1111111111111111_1101101011011011_0101011001000001"; -- -0.14509068416000462
	pesos_i(7499) := b"1111111111111111_1111111111111111_1111100010100011_0111110101100101"; -- -0.028755343393336602
	pesos_i(7500) := b"1111111111111111_1111111111111111_1111101000110000_0100100001011000"; -- -0.02270076612919854
	pesos_i(7501) := b"1111111111111111_1111111111111111_1111101100010011_0110011111011111"; -- -0.019235141720589762
	pesos_i(7502) := b"0000000000000000_0000000000000000_0000100011011111_0101011110001111"; -- 0.034657928749140865
	pesos_i(7503) := b"0000000000000000_0000000000000000_0001100100000010_1100000000000111"; -- 0.09769821338663026
	pesos_i(7504) := b"1111111111111111_1111111111111111_1111100001000110_0010000001110100"; -- -0.030179950510106995
	pesos_i(7505) := b"0000000000000000_0000000000000000_0010011011100101_1010110100111111"; -- 0.15194208891922023
	pesos_i(7506) := b"0000000000000000_0000000000000000_0001100011100011_1101110001110010"; -- 0.09722688457425156
	pesos_i(7507) := b"1111111111111111_1111111111111111_1110010000111011_1011011010011111"; -- -0.10846384647753013
	pesos_i(7508) := b"1111111111111111_1111111111111111_1101010010101000_0100100000010111"; -- -0.16930722644104776
	pesos_i(7509) := b"0000000000000000_0000000000000000_0010101001100010_0010101100000011"; -- 0.16556042514144204
	pesos_i(7510) := b"0000000000000000_0000000000000000_0001111110110010_0000010101110001"; -- 0.12381013873409585
	pesos_i(7511) := b"1111111111111111_1111111111111111_1101100011100000_1001101011111001"; -- -0.15282279426339854
	pesos_i(7512) := b"1111111111111111_1111111111111111_1101000001100110_0110110100001000"; -- -0.18593710471633176
	pesos_i(7513) := b"0000000000000000_0000000000000000_0000010010111100_0110000000111111"; -- 0.018499389164232112
	pesos_i(7514) := b"1111111111111111_1111111111111111_1111001110110001_1011000011100000"; -- -0.04806990184441784
	pesos_i(7515) := b"1111111111111111_1111111111111111_1111111001000001_1110110101010001"; -- -0.006806533486906862
	pesos_i(7516) := b"0000000000000000_0000000000000000_0001010011101110_1111110000001110"; -- 0.08177161546354571
	pesos_i(7517) := b"1111111111111111_1111111111111111_1111001111111011_0110101011011101"; -- -0.046944924333752865
	pesos_i(7518) := b"0000000000000000_0000000000000000_0010011000011011_1101110011000011"; -- 0.14886264568329663
	pesos_i(7519) := b"1111111111111111_1111111111111111_1110011111110111_0000111010010000"; -- -0.09388646111806437
	pesos_i(7520) := b"1111111111111111_1111111111111111_1101011100100100_0000010100010010"; -- -0.15960663129520086
	pesos_i(7521) := b"0000000000000000_0000000000000000_0001000000000100_1000010010001000"; -- 0.06256893452148467
	pesos_i(7522) := b"0000000000000000_0000000000000000_0000111011111100_0000000111001001"; -- 0.05853282117028192
	pesos_i(7523) := b"0000000000000000_0000000000000000_0010101010001010_0111101111000101"; -- 0.16617559021126665
	pesos_i(7524) := b"1111111111111111_1111111111111111_1110001000011011_0111001011110101"; -- -0.11676866064867308
	pesos_i(7525) := b"1111111111111111_1111111111111111_1110011010101011_1110000001101101"; -- -0.0989398702011251
	pesos_i(7526) := b"0000000000000000_0000000000000000_0010011011001000_1001001001110000"; -- 0.15149798609872325
	pesos_i(7527) := b"0000000000000000_0000000000000000_0000001000100011_0111100000011011"; -- 0.008353716472679545
	pesos_i(7528) := b"1111111111111111_1111111111111111_1110101000111101_0011110111111011"; -- -0.08500301945687619
	pesos_i(7529) := b"1111111111111111_1111111111111111_1110001011111100_1111001010011001"; -- -0.11332782518209801
	pesos_i(7530) := b"1111111111111111_1111111111111111_1101010101001011_1100100000101111"; -- -0.16681240897135363
	pesos_i(7531) := b"0000000000000000_0000000000000000_0001101100100000_0010010000010001"; -- 0.10595918104118329
	pesos_i(7532) := b"1111111111111111_1111111111111111_1110011010100101_0011111111000110"; -- -0.09904099859697461
	pesos_i(7533) := b"1111111111111111_1111111111111111_1111101100100010_1001100010101001"; -- -0.019003351989075063
	pesos_i(7534) := b"0000000000000000_0000000000000000_0010101001111110_1111011010000011"; -- 0.16599980060025119
	pesos_i(7535) := b"0000000000000000_0000000000000000_0001111010011010_1001001111001001"; -- 0.11954616220135268
	pesos_i(7536) := b"0000000000000000_0000000000000000_0001000010110010_0010110100100011"; -- 0.06521875475483022
	pesos_i(7537) := b"0000000000000000_0000000000000000_0001011000110010_1110000000000111"; -- 0.08671379260284436
	pesos_i(7538) := b"0000000000000000_0000000000000000_0000110011000011_0101100101011001"; -- 0.04985578942343631
	pesos_i(7539) := b"1111111111111111_1111111111111111_1110101011100011_1001110010011111"; -- -0.08246441957843159
	pesos_i(7540) := b"0000000000000000_0000000000000000_0000111001000011_0000010000001100"; -- 0.055710080035712595
	pesos_i(7541) := b"0000000000000000_0000000000000000_0010000111100111_0000011100011010"; -- 0.13243145349607643
	pesos_i(7542) := b"1111111111111111_1111111111111111_1110110111001110_0101010010110110"; -- -0.07107039031683969
	pesos_i(7543) := b"0000000000000000_0000000000000000_0011000011111111_0010110000010000"; -- 0.19139361754998577
	pesos_i(7544) := b"1111111111111111_1111111111111111_1111010011100100_1101110010110100"; -- -0.043382841183189524
	pesos_i(7545) := b"0000000000000000_0000000000000000_0001010100111011_0110100110011101"; -- 0.08293781354948154
	pesos_i(7546) := b"0000000000000000_0000000000000000_0000111111100110_0101111110010111"; -- 0.062108968994407585
	pesos_i(7547) := b"1111111111111111_1111111111111111_1110010011111000_0000001010010011"; -- -0.10559066684347537
	pesos_i(7548) := b"1111111111111111_1111111111111111_1110111100101011_1100011011110000"; -- -0.06573826451050037
	pesos_i(7549) := b"0000000000000000_0000000000000000_0010101000010011_0101100010100011"; -- 0.16435770023229762
	pesos_i(7550) := b"0000000000000000_0000000000000000_0000001001000101_1010110010000101"; -- 0.008875639445757736
	pesos_i(7551) := b"0000000000000000_0000000000000000_0010001010100110_1111110110111111"; -- 0.13536058347304253
	pesos_i(7552) := b"0000000000000000_0000000000000000_0010000010101010_0001101100111100"; -- 0.12759561751523582
	pesos_i(7553) := b"0000000000000000_0000000000000000_0010100000100111_0100011010110011"; -- 0.15684930666995867
	pesos_i(7554) := b"0000000000000000_0000000000000000_0010110011000010_1011111011110010"; -- 0.17484658624098098
	pesos_i(7555) := b"1111111111111111_1111111111111111_1110000101101011_1010000110011010"; -- -0.11945142733218439
	pesos_i(7556) := b"0000000000000000_0000000000000000_0000110101011101_1001010100111110"; -- 0.052209212848865164
	pesos_i(7557) := b"1111111111111111_1111111111111111_1111100011111010_0100111011000001"; -- -0.027430608696307746
	pesos_i(7558) := b"0000000000000000_0000000000000000_0000111111111101_0000100000110001"; -- 0.06245471182080577
	pesos_i(7559) := b"0000000000000000_0000000000000000_0010011101000101_1011000110010001"; -- 0.15340719016251708
	pesos_i(7560) := b"1111111111111111_1111111111111111_1110011000110100_1010101011101000"; -- -0.10075885606446108
	pesos_i(7561) := b"1111111111111111_1111111111111111_1101111010011100_1110011001010111"; -- -0.13041839955810833
	pesos_i(7562) := b"1111111111111111_1111111111111111_1101011011010011_0001011011010001"; -- -0.16084153557410605
	pesos_i(7563) := b"1111111111111111_1111111111111111_1111101101011000_0001011100000100"; -- -0.018187104830476072
	pesos_i(7564) := b"0000000000000000_0000000000000000_0010001111110101_0111010101100110"; -- 0.1404641507390022
	pesos_i(7565) := b"0000000000000000_0000000000000000_0010001010110001_0001111011001001"; -- 0.13551514066709106
	pesos_i(7566) := b"1111111111111111_1111111111111111_1110111001111100_0111001011010110"; -- -0.068413565324138
	pesos_i(7567) := b"1111111111111111_1111111111111111_1101101100011000_0110111000101001"; -- -0.14415847294314693
	pesos_i(7568) := b"1111111111111111_1111111111111111_1101011100101011_0101110010111101"; -- -0.15949459439937622
	pesos_i(7569) := b"1111111111111111_1111111111111111_1110100000101000_0011001001110011"; -- -0.09313664138535728
	pesos_i(7570) := b"1111111111111111_1111111111111111_1110000011100101_0010011100111100"; -- -0.12150339866418745
	pesos_i(7571) := b"1111111111111111_1111111111111111_1110110110000100_0001101100100110"; -- -0.07220297163221472
	pesos_i(7572) := b"0000000000000000_0000000000000000_0001011010011011_0010001011110100"; -- 0.08830469575857135
	pesos_i(7573) := b"1111111111111111_1111111111111111_1110001100100100_0001110000111011"; -- -0.11273025082482252
	pesos_i(7574) := b"0000000000000000_0000000000000000_0010000000011010_0101100110111001"; -- 0.1254020763255574
	pesos_i(7575) := b"1111111111111111_1111111111111111_1110110100101001_0001110100111011"; -- -0.0735913972731716
	pesos_i(7576) := b"0000000000000000_0000000000000000_0000101000110100_0101100011111101"; -- 0.039861261082421565
	pesos_i(7577) := b"1111111111111111_1111111111111111_1111111010011001_0101001111101110"; -- -0.005472902633711093
	pesos_i(7578) := b"1111111111111111_1111111111111111_1111011011111111_1110000001110101"; -- -0.03515813005369885
	pesos_i(7579) := b"1111111111111111_1111111111111111_1110100100010101_1000101000100010"; -- -0.08951508217688775
	pesos_i(7580) := b"0000000000000000_0000000000000000_0010001010011011_1111101000011011"; -- 0.1351925197954273
	pesos_i(7581) := b"1111111111111111_1111111111111111_1111101010000010_1111100000010000"; -- -0.021439071857062363
	pesos_i(7582) := b"0000000000000000_0000000000000000_0000010100101000_0011111111000110"; -- 0.020145402670643447
	pesos_i(7583) := b"1111111111111111_1111111111111111_1110111011101001_1011001011001000"; -- -0.06674654584451302
	pesos_i(7584) := b"1111111111111111_1111111111111111_1101101111111001_0100010110100011"; -- -0.14072766085596022
	pesos_i(7585) := b"1111111111111111_1111111111111111_1111100000111001_0111100010110001"; -- -0.03037305532517368
	pesos_i(7586) := b"0000000000000000_0000000000000000_0000110010111101_1110000001100110"; -- 0.04977228624633995
	pesos_i(7587) := b"1111111111111111_1111111111111111_1110101011001100_0001101100111110"; -- -0.08282308320341972
	pesos_i(7588) := b"0000000000000000_0000000000000000_0010010011101111_1010110111000101"; -- 0.1442822080445867
	pesos_i(7589) := b"1111111111111111_1111111111111111_1111001110000110_0101101111111100"; -- -0.04873108954634873
	pesos_i(7590) := b"0000000000000000_0000000000000000_0010101010110010_1100100001110000"; -- 0.16679051147918528
	pesos_i(7591) := b"1111111111111111_1111111111111111_1110111000100001_1100101001011101"; -- -0.0697968981455448
	pesos_i(7592) := b"1111111111111111_1111111111111111_1110011001111110_0011001111101100"; -- -0.09963679782919906
	pesos_i(7593) := b"1111111111111111_1111111111111111_1110011101011101_0010010101010101"; -- -0.09623495738487307
	pesos_i(7594) := b"0000000000000000_0000000000000000_0000000111010101_1000011101101011"; -- 0.007164443600808127
	pesos_i(7595) := b"0000000000000000_0000000000000000_0000000101011000_1110100100100001"; -- 0.005262918896109282
	pesos_i(7596) := b"1111111111111111_1111111111111111_1101010010111111_0001000100111001"; -- -0.1689595447013195
	pesos_i(7597) := b"1111111111111111_1111111111111111_1110101101101110_0110101101111001"; -- -0.08034637729093566
	pesos_i(7598) := b"0000000000000000_0000000000000000_0010011101100010_1000100001011100"; -- 0.15384723892188237
	pesos_i(7599) := b"0000000000000000_0000000000000000_0000000101001011_1110000011100001"; -- 0.00506406291600366
	pesos_i(7600) := b"1111111111111111_1111111111111111_1110001111101001_1101101011100110"; -- -0.10971290489259816
	pesos_i(7601) := b"0000000000000000_0000000000000000_0001111000111010_0000000010001010"; -- 0.11807254201069156
	pesos_i(7602) := b"1111111111111111_1111111111111111_1111110000110010_1001101100010100"; -- -0.014852817140996146
	pesos_i(7603) := b"0000000000000000_0000000000000000_0001111011110001_0100101100111100"; -- 0.12086935250904005
	pesos_i(7604) := b"0000000000000000_0000000000000000_0000110011000110_1101010100101100"; -- 0.04990894621860037
	pesos_i(7605) := b"0000000000000000_0000000000000000_0000010100000010_1111100001000001"; -- 0.0195765646871558
	pesos_i(7606) := b"0000000000000000_0000000000000000_0001111001000111_1101111101011010"; -- 0.11828418679265397
	pesos_i(7607) := b"0000000000000000_0000000000000000_0010100111010000_1010000000000010"; -- 0.16333961522761836
	pesos_i(7608) := b"1111111111111111_1111111111111111_1111101100101001_0101011110111000"; -- -0.01890041115278393
	pesos_i(7609) := b"0000000000000000_0000000000000000_0001010111100100_0101001011101010"; -- 0.08551519587026778
	pesos_i(7610) := b"0000000000000000_0000000000000000_0000110010010010_0111010100011011"; -- 0.049109763179895155
	pesos_i(7611) := b"1111111111111111_1111111111111111_1111001111111111_1101001000100001"; -- -0.04687773423171974
	pesos_i(7612) := b"0000000000000000_0000000000000000_0010100001100001_0011100011010100"; -- 0.15773348974404444
	pesos_i(7613) := b"1111111111111111_1111111111111111_1110010101001000_0101001011110001"; -- -0.10436517359754614
	pesos_i(7614) := b"0000000000000000_0000000000000000_0010100110011011_0000001101010000"; -- 0.16252155971017518
	pesos_i(7615) := b"0000000000000000_0000000000000000_0001001010100000_0001101011011100"; -- 0.07275550723772015
	pesos_i(7616) := b"0000000000000000_0000000000000000_0001000110111000_0011101100100010"; -- 0.06921739187854731
	pesos_i(7617) := b"1111111111111111_1111111111111111_1110111011010101_0011100111001010"; -- -0.0670589334732456
	pesos_i(7618) := b"0000000000000000_0000000000000000_0001010010101111_0110110000011100"; -- 0.08080173186720102
	pesos_i(7619) := b"1111111111111111_1111111111111111_1110101111101000_1111001100110100"; -- -0.07847671484983362
	pesos_i(7620) := b"1111111111111111_1111111111111111_1110010011000000_0101001000000100"; -- -0.10644042394884624
	pesos_i(7621) := b"1111111111111111_1111111111111111_1101011100011100_0101000001000011"; -- -0.15972421998231348
	pesos_i(7622) := b"0000000000000000_0000000000000000_0010011100100110_1000000000111011"; -- 0.152931227029705
	pesos_i(7623) := b"1111111111111111_1111111111111111_1111101001100010_0110000011110001"; -- -0.0219363605571344
	pesos_i(7624) := b"0000000000000000_0000000000000000_0011110101111000_0011011010110010"; -- 0.24011556489758584
	pesos_i(7625) := b"0000000000000000_0000000000000000_0010110101011101_0111001001100101"; -- 0.1772071358537169
	pesos_i(7626) := b"1111111111111111_1111111111111111_1101101111000101_1100010000110011"; -- -0.14151357417081814
	pesos_i(7627) := b"1111111111111111_1111111111111111_1110010100110100_1100011100000111"; -- -0.1046634299403001
	pesos_i(7628) := b"1111111111111111_1111111111111111_1111010101000010_1111000101010010"; -- -0.041947286170079416
	pesos_i(7629) := b"0000000000000000_0000000000000000_0001110000000110_0000001001001000"; -- 0.10946668860000512
	pesos_i(7630) := b"1111111111111111_1111111111111111_1110011110010010_1011110101011000"; -- -0.09541718097925925
	pesos_i(7631) := b"1111111111111111_1111111111111111_1111100001011010_0101010111000011"; -- -0.029871597166460227
	pesos_i(7632) := b"1111111111111111_1111111111111111_1110100000001111_0111001111111101"; -- -0.09351420466837694
	pesos_i(7633) := b"0000000000000000_0000000000000000_0001001110001111_0101011001100001"; -- 0.07640590541265053
	pesos_i(7634) := b"1111111111111111_1111111111111111_1111101100011111_1110001000111010"; -- -0.019044743348198813
	pesos_i(7635) := b"0000000000000000_0000000000000000_0000100000110011_0001101111000000"; -- 0.032029852306726614
	pesos_i(7636) := b"1111111111111111_1111111111111111_1101100000111101_0111110000111001"; -- -0.15531180970605393
	pesos_i(7637) := b"1111111111111111_1111111111111111_1101010100100110_0011001110001001"; -- -0.1673858443363147
	pesos_i(7638) := b"0000000000000000_0000000000000000_0001011000000000_1010101010000001"; -- 0.08594766275897502
	pesos_i(7639) := b"1111111111111111_1111111111111111_1110100101110110_1110110011100011"; -- -0.08802909333844848
	pesos_i(7640) := b"0000000000000000_0000000000000000_0010001000110100_0110101111101000"; -- 0.13361238866391756
	pesos_i(7641) := b"0000000000000000_0000000000000000_0000001001011111_1110100011100001"; -- 0.00927596568367177
	pesos_i(7642) := b"1111111111111111_1111111111111111_1110101110110100_0000011100000100"; -- -0.07928424987511835
	pesos_i(7643) := b"1111111111111111_1111111111111111_1101100010110110_0111111100010001"; -- -0.15346532674142221
	pesos_i(7644) := b"0000000000000000_0000000000000000_0001011100100000_1011100101001001"; -- 0.09034307510974826
	pesos_i(7645) := b"1111111111111111_1111111111111111_1111110000101000_0001100000101010"; -- -0.015013208092102038
	pesos_i(7646) := b"0000000000000000_0000000000000000_0000000011000011_1111110100000110"; -- 0.002990545312752688
	pesos_i(7647) := b"0000000000000000_0000000000000000_0001011001111011_1110000101101101"; -- 0.08782776757192115
	pesos_i(7648) := b"1111111111111111_1111111111111111_1101001110110101_1100001110101111"; -- -0.17300774556539805
	pesos_i(7649) := b"1111111111111111_1111111111111111_1111001110010110_1011011110011001"; -- -0.048481488384501364
	pesos_i(7650) := b"0000000000000000_0000000000000000_0010110011000111_0110111011110000"; -- 0.17491811151724163
	pesos_i(7651) := b"0000000000000000_0000000000000000_0001100110010110_0100001000111111"; -- 0.09994901701724375
	pesos_i(7652) := b"0000000000000000_0000000000000000_0010101110101101_1011111101101010"; -- 0.1706199296922027
	pesos_i(7653) := b"1111111111111111_1111111111111111_1110101010111010_1101101010000110"; -- -0.08308634012684323
	pesos_i(7654) := b"1111111111111111_1111111111111111_1101101011101001_1100100100110110"; -- -0.14487020903800735
	pesos_i(7655) := b"0000000000000000_0000000000000000_0001100001100011_0110111000001001"; -- 0.09526717878227445
	pesos_i(7656) := b"0000000000000000_0000000000000000_0001000011001100_1000001001100110"; -- 0.06562056535577601
	pesos_i(7657) := b"0000000000000000_0000000000000000_0000111111100110_1010111110001100"; -- 0.06211373482505481
	pesos_i(7658) := b"0000000000000000_0000000000000000_0010101000011100_1010011110000001"; -- 0.164499730196445
	pesos_i(7659) := b"1111111111111111_1111111111111111_1110110110101000_0101110011010010"; -- -0.07164974089765201
	pesos_i(7660) := b"1111111111111111_1111111111111111_1111100111011010_0000011010100011"; -- -0.02401693837935113
	pesos_i(7661) := b"0000000000000000_0000000000000000_0001010100101110_0100110111100010"; -- 0.08273779639512022
	pesos_i(7662) := b"0000000000000000_0000000000000000_0001101100000101_1110110001100011"; -- 0.10555913359265873
	pesos_i(7663) := b"1111111111111111_1111111111111111_1110011011010100_1100000010011011"; -- -0.09831615648528022
	pesos_i(7664) := b"0000000000000000_0000000000000000_0000001000000101_0110000110011100"; -- 0.007894612020082459
	pesos_i(7665) := b"1111111111111111_1111111111111111_1110001111010110_1111110000000000"; -- -0.11000084882624146
	pesos_i(7666) := b"1111111111111111_1111111111111111_1111010101001100_0111100101000010"; -- -0.04180185441102271
	pesos_i(7667) := b"0000000000000000_0000000000000000_0010001011100010_0000001101010011"; -- 0.13626118453188796
	pesos_i(7668) := b"0000000000000000_0000000000000000_0001001011011001_1110000010101110"; -- 0.07363704912005362
	pesos_i(7669) := b"1111111111111111_1111111111111111_1110100010001010_1101110101111101"; -- -0.09163108532119689
	pesos_i(7670) := b"0000000000000000_0000000000000000_0001100100001100_0110111100111101"; -- 0.09784598568217302
	pesos_i(7671) := b"0000000000000000_0000000000000000_0010100101000001_0101111001001111"; -- 0.16115369250655104
	pesos_i(7672) := b"0000000000000000_0000000000000000_0000010011000100_1111001111001110"; -- 0.018630254574748567
	pesos_i(7673) := b"1111111111111111_1111111111111111_1101000011001101_1111111100011000"; -- -0.18435674339882344
	pesos_i(7674) := b"0000000000000000_0000000000000000_0001000000110100_0100010011010010"; -- 0.06329755915747193
	pesos_i(7675) := b"1111111111111111_1111111111111111_1101110110100010_0111101110100111"; -- -0.13423945600777998
	pesos_i(7676) := b"0000000000000000_0000000000000000_0000110111111110_0101010110001110"; -- 0.054662081833892553
	pesos_i(7677) := b"1111111111111111_1111111111111111_1111010011101111_0010000010000010"; -- -0.04322621179989279
	pesos_i(7678) := b"1111111111111111_1111111111111111_1101100101100011_0101010101101011"; -- -0.1508280385213313
	pesos_i(7679) := b"0000000000000000_0000000000000000_0010100100001011_0101101111011101"; -- 0.1603295722077184
	pesos_i(7680) := b"1111111111111111_1111111111111111_1110001010000010_1110000100010010"; -- -0.11519044217202343
	pesos_i(7681) := b"1111111111111111_1111111111111111_1101010101110010_0110111111000010"; -- -0.16622258676012935
	pesos_i(7682) := b"0000000000000000_0000000000000000_0001001010110100_1001100000101001"; -- 0.07306815146428537
	pesos_i(7683) := b"1111111111111111_1111111111111111_1111111101101101_0000110011001101"; -- -0.0022422789124416803
	pesos_i(7684) := b"1111111111111111_1111111111111111_1110011100011100_0000110110110000"; -- -0.09722818802824555
	pesos_i(7685) := b"1111111111111111_1111111111111111_1101111100110001_1111000000110001"; -- -0.12814425290731912
	pesos_i(7686) := b"0000000000000000_0000000000000000_0000010111100100_0011100001000111"; -- 0.023013608285041412
	pesos_i(7687) := b"0000000000000000_0000000000000000_0010011011011101_0111100001101011"; -- 0.15181686988734397
	pesos_i(7688) := b"1111111111111111_1111111111111111_1110110101000001_1100111011011011"; -- -0.07321459926149747
	pesos_i(7689) := b"1111111111111111_1111111111111111_1111000001001001_0010110011000010"; -- -0.06138344064759118
	pesos_i(7690) := b"1111111111111111_1111111111111111_1111000110000101_1011101000011011"; -- -0.056553238292559274
	pesos_i(7691) := b"0000000000000000_0000000000000000_0010101110000110_1110111011000001"; -- 0.17002765862792485
	pesos_i(7692) := b"1111111111111111_1111111111111111_1110000111011110_1001110001000001"; -- -0.11769698532952146
	pesos_i(7693) := b"0000000000000000_0000000000000000_0010000111101010_0100011001000000"; -- 0.1324809938859068
	pesos_i(7694) := b"0000000000000000_0000000000000000_0000111000010010_0000111100101011"; -- 0.054963062297619956
	pesos_i(7695) := b"1111111111111111_1111111111111111_1111010000011010_0011111101111101"; -- -0.04647448719254171
	pesos_i(7696) := b"0000000000000000_0000000000000000_0001110000001010_1111111011000100"; -- 0.10954277309888319
	pesos_i(7697) := b"0000000000000000_0000000000000000_0000001100010110_0111010000011000"; -- 0.012061362998101325
	pesos_i(7698) := b"1111111111111111_1111111111111111_1111001000101000_0101111010111011"; -- -0.05407150198757286
	pesos_i(7699) := b"0000000000000000_0000000000000000_0010010001011010_0000001010010011"; -- 0.14199844448843907
	pesos_i(7700) := b"1111111111111111_1111111111111111_1110011100111110_1011111100010001"; -- -0.09669881655980901
	pesos_i(7701) := b"1111111111111111_1111111111111111_1101110000110100_0111010101100101"; -- -0.13982454574464062
	pesos_i(7702) := b"0000000000000000_0000000000000000_0001101100000101_1101011110010111"; -- 0.10555789412447425
	pesos_i(7703) := b"0000000000000000_0000000000000000_0000100011001000_0100100110000011"; -- 0.03430613936677425
	pesos_i(7704) := b"1111111111111111_1111111111111111_1111000011011100_0010101000110110"; -- -0.05914055048861465
	pesos_i(7705) := b"0000000000000000_0000000000000000_0001100010010001_1100000000111101"; -- 0.095973982729065
	pesos_i(7706) := b"1111111111111111_1111111111111111_1110000001011001_1111111001100111"; -- -0.12362680413391772
	pesos_i(7707) := b"0000000000000000_0000000000000000_0010101110100100_1011100110101110"; -- 0.17048225871027323
	pesos_i(7708) := b"0000000000000000_0000000000000000_0000101000000011_1011011101110001"; -- 0.039119210416428254
	pesos_i(7709) := b"0000000000000000_0000000000000000_0001011110011100_1111100000111001"; -- 0.09223891641027744
	pesos_i(7710) := b"1111111111111111_1111111111111111_1111000101000000_1110000001101101"; -- -0.05760381063515929
	pesos_i(7711) := b"1111111111111111_1111111111111111_1111000101111010_0011110101001111"; -- -0.05672852357278052
	pesos_i(7712) := b"1111111111111111_1111111111111111_1101110010111001_0000110010000010"; -- -0.1378013784732799
	pesos_i(7713) := b"0000000000000000_0000000000000000_0001001001110001_0100000100100011"; -- 0.07204062551866008
	pesos_i(7714) := b"1111111111111111_1111111111111111_1101110101101101_0100001111101111"; -- -0.1350514928025385
	pesos_i(7715) := b"0000000000000000_0000000000000000_0001010111101001_1010011101011101"; -- 0.08559652350892655
	pesos_i(7716) := b"1111111111111111_1111111111111111_1110011110101000_0011110010001100"; -- -0.09508916464403427
	pesos_i(7717) := b"0000000000000000_0000000000000000_0001111011011000_1100111001001000"; -- 0.1204956936903845
	pesos_i(7718) := b"1111111111111111_1111111111111111_1101110001111000_1010110010110010"; -- -0.13878365186654035
	pesos_i(7719) := b"1111111111111111_1111111111111111_1110100100000110_0011000010001100"; -- -0.08974930367115289
	pesos_i(7720) := b"0000000000000000_0000000000000000_0000000111110111_0101000001011000"; -- 0.00767995981531544
	pesos_i(7721) := b"1111111111111111_1111111111111111_1111110111100101_0000111111101010"; -- -0.008223538666960859
	pesos_i(7722) := b"1111111111111111_1111111111111111_1110001110110011_0110011000110101"; -- -0.11054383479466151
	pesos_i(7723) := b"1111111111111111_1111111111111111_1101110100001101_1000111110100100"; -- -0.1365118240113571
	pesos_i(7724) := b"1111111111111111_1111111111111111_1111010101000110_0010011000001101"; -- -0.04189836678664757
	pesos_i(7725) := b"0000000000000000_0000000000000000_0001010100011101_0011010100100010"; -- 0.0824769218852449
	pesos_i(7726) := b"0000000000000000_0000000000000000_0010000010000011_0011000010111100"; -- 0.12700180606931966
	pesos_i(7727) := b"0000000000000000_0000000000000000_0010011111101011_1010000010001101"; -- 0.15593913502800952
	pesos_i(7728) := b"0000000000000000_0000000000000000_0010100101101110_1111001011011111"; -- 0.16184919311724663
	pesos_i(7729) := b"0000000000000000_0000000000000000_0000111011001000_0010000100001101"; -- 0.05774122774231759
	pesos_i(7730) := b"1111111111111111_1111111111111111_1101101100000110_1100010110100101"; -- -0.1444279168466258
	pesos_i(7731) := b"0000000000000000_0000000000000000_0010010110110111_0010110100010110"; -- 0.1473262957873473
	pesos_i(7732) := b"0000000000000000_0000000000000000_0001010110100100_1001111000110010"; -- 0.08454312069463273
	pesos_i(7733) := b"1111111111111111_1111111111111111_1110000100111011_1110000001100011"; -- -0.1201801069516181
	pesos_i(7734) := b"1111111111111111_1111111111111111_1110111111110001_1110110011101000"; -- -0.06271476111804658
	pesos_i(7735) := b"0000000000000000_0000000000000000_0001000010111101_0000011000001001"; -- 0.06538427089112069
	pesos_i(7736) := b"1111111111111111_1111111111111111_1101111111100111_0010010010110011"; -- -0.12537928221727843
	pesos_i(7737) := b"0000000000000000_0000000000000000_0000001000000010_0100110010000111"; -- 0.00784757898979296
	pesos_i(7738) := b"0000000000000000_0000000000000000_0000101001011010_0001011010010001"; -- 0.04043713609275159
	pesos_i(7739) := b"1111111111111111_1111111111111111_1101111111101001_0000001001101011"; -- -0.12535080811073623
	pesos_i(7740) := b"1111111111111111_1111111111111111_1110010111101000_0110001011101111"; -- -0.10192281408358275
	pesos_i(7741) := b"1111111111111111_1111111111111111_1111010111011111_0010100010011101"; -- -0.03956361933159998
	pesos_i(7742) := b"1111111111111111_1111111111111111_1111100110100010_0101111110001010"; -- -0.024866131521133306
	pesos_i(7743) := b"1111111111111111_1111111111111111_1101010010100111_1100110010010111"; -- -0.16931458783786152
	pesos_i(7744) := b"0000000000000000_0000000000000000_0000101001111000_0100101001101010"; -- 0.04089799020028115
	pesos_i(7745) := b"1111111111111111_1111111111111111_1110100000010011_0001111100010110"; -- -0.09345823003252451
	pesos_i(7746) := b"1111111111111111_1111111111111111_1110101010110010_0110001010110111"; -- -0.0832155517502442
	pesos_i(7747) := b"0000000000000000_0000000000000000_0010101010110100_1110000000111101"; -- 0.16682244774216098
	pesos_i(7748) := b"1111111111111111_1111111111111111_1110100111110001_0101100111101100"; -- -0.0861610221308566
	pesos_i(7749) := b"1111111111111111_1111111111111111_1101101111101111_1110000100001110"; -- -0.14087098505480614
	pesos_i(7750) := b"0000000000000000_0000000000000000_0000101010010101_1000111010101011"; -- 0.04134456316517433
	pesos_i(7751) := b"0000000000000000_0000000000000000_0001110110001110_0001110110010010"; -- 0.11544976059055229
	pesos_i(7752) := b"1111111111111111_1111111111111111_1100111011001011_0101011011001011"; -- -0.1922097926623249
	pesos_i(7753) := b"1111111111111111_1111111111111111_1101110010111101_0011011001001010"; -- -0.1377378529942467
	pesos_i(7754) := b"1111111111111111_1111111111111111_1110011101101000_1101011110011000"; -- -0.09605648546340566
	pesos_i(7755) := b"0000000000000000_0000000000000000_0001101000100101_0010111110001110"; -- 0.10212990976582104
	pesos_i(7756) := b"1111111111111111_1111111111111111_1110111010001111_1001011000011101"; -- -0.0681215456449221
	pesos_i(7757) := b"0000000000000000_0000000000000000_0000101100000111_0000001010111001"; -- 0.04307572390983683
	pesos_i(7758) := b"1111111111111111_1111111111111111_1100111111000010_0010100010011010"; -- -0.18844362498867312
	pesos_i(7759) := b"0000000000000000_0000000000000000_0001110101000110_0001101101001010"; -- 0.11435099178212926
	pesos_i(7760) := b"0000000000000000_0000000000000000_0000001011011110_0101111011100000"; -- 0.011205606159357201
	pesos_i(7761) := b"1111111111111111_1111111111111111_1110011110110101_0101001000111100"; -- -0.09488950774077666
	pesos_i(7762) := b"1111111111111111_1111111111111111_1110010101111010_1001010110100101"; -- -0.10359825824086841
	pesos_i(7763) := b"0000000000000000_0000000000000000_0000101110010000_1001011101000001"; -- 0.04517503113964636
	pesos_i(7764) := b"1111111111111111_1111111111111111_1111001111100001_0011000101011100"; -- -0.04734508045895164
	pesos_i(7765) := b"0000000000000000_0000000000000000_0001101010100001_1011111110101001"; -- 0.10403058893878568
	pesos_i(7766) := b"0000000000000000_0000000000000000_0001111001000001_1001111011111101"; -- 0.11818879773632508
	pesos_i(7767) := b"0000000000000000_0000000000000000_0010000101100111_1011100110100000"; -- 0.130488969285397
	pesos_i(7768) := b"1111111111111111_1111111111111111_1101111001000010_1100101011110100"; -- -0.1317933230815996
	pesos_i(7769) := b"0000000000000000_0000000000000000_0001101011001010_0110101000111110"; -- 0.10465110799623846
	pesos_i(7770) := b"1111111111111111_1111111111111111_1111001001101000_0100101011100000"; -- -0.05309612310764444
	pesos_i(7771) := b"1111111111111111_1111111111111111_1101011010001000_1011100100000000"; -- -0.16197627785314855
	pesos_i(7772) := b"1111111111111111_1111111111111111_1110000000101111_1000001111101111"; -- -0.12427497299698391
	pesos_i(7773) := b"1111111111111111_1111111111111111_1101011110010010_0010111101010000"; -- -0.15792564670703926
	pesos_i(7774) := b"1111111111111111_1111111111111111_1111000011110010_0100001000110110"; -- -0.05880342661626311
	pesos_i(7775) := b"0000000000000000_0000000000000000_0000010000110011_0001111100001000"; -- 0.016405047853000676
	pesos_i(7776) := b"0000000000000000_0000000000000000_0010100110000001_1000000100010000"; -- 0.16213232651752504
	pesos_i(7777) := b"0000000000000000_0000000000000000_0010010001100000_1010110011011001"; -- 0.1421001462537383
	pesos_i(7778) := b"1111111111111111_1111111111111111_1110101001001100_1101001010001001"; -- -0.08476528323226466
	pesos_i(7779) := b"1111111111111111_1111111111111111_1111010100110010_0111100010100110"; -- -0.04219861934024311
	pesos_i(7780) := b"0000000000000000_0000000000000000_0010010001010101_1111011010010010"; -- 0.14193669376465282
	pesos_i(7781) := b"1111111111111111_1111111111111111_1110101010110001_0010111111110111"; -- -0.08323383545781889
	pesos_i(7782) := b"0000000000000000_0000000000000000_0010000001101111_0101111000101111"; -- 0.12669933933398667
	pesos_i(7783) := b"0000000000000000_0000000000000000_0010100011111110_0011001000111000"; -- 0.16012872559127775
	pesos_i(7784) := b"1111111111111111_1111111111111111_1111010010000101_1011101011010110"; -- -0.04483444485174057
	pesos_i(7785) := b"0000000000000000_0000000000000000_0000000111011110_0111101100111001"; -- 0.0073010457864318735
	pesos_i(7786) := b"0000000000000000_0000000000000000_0000001100111001_1000001110010100"; -- 0.012596343605143473
	pesos_i(7787) := b"0000000000000000_0000000000000000_0000011110100000_0100110111010101"; -- 0.029789795355548647
	pesos_i(7788) := b"0000000000000000_0000000000000000_0010010100101101_1001101110110011"; -- 0.1452271758800204
	pesos_i(7789) := b"0000000000000000_0000000000000000_0000110110010100_0100011000011111"; -- 0.05304373043744213
	pesos_i(7790) := b"1111111111111111_1111111111111111_1110011000110011_0110100001101111"; -- -0.10077807698366258
	pesos_i(7791) := b"0000000000000000_0000000000000000_0011110110000011_1101001111110001"; -- 0.24029278404243748
	pesos_i(7792) := b"0000000000000000_0000000000000000_0000110001001101_0011101010011001"; -- 0.048053419458793156
	pesos_i(7793) := b"0000000000000000_0000000000000000_0000010111001000_0010100011011110"; -- 0.022585443615858368
	pesos_i(7794) := b"0000000000000000_0000000000000000_0000111111111110_1001010101011100"; -- 0.06247838501879516
	pesos_i(7795) := b"1111111111111111_1111111111111111_1101011111111010_0011111100011001"; -- -0.1563377918607002
	pesos_i(7796) := b"1111111111111111_1111111111111111_1111110001111001_1101010011101011"; -- -0.013765995628900202
	pesos_i(7797) := b"1111111111111111_1111111111111111_1110001000011011_0110010100000100"; -- -0.11676949178856093
	pesos_i(7798) := b"0000000000000000_0000000000000000_0000010001111001_0110011110001100"; -- 0.01747748539796494
	pesos_i(7799) := b"1111111111111111_1111111111111111_1110100010001001_0010101011010001"; -- -0.09165699390313603
	pesos_i(7800) := b"1111111111111111_1111111111111111_1111101011101111_0010010101110011"; -- -0.019788417344010656
	pesos_i(7801) := b"1111111111111111_1111111111111111_1110011000100101_0101000001101010"; -- -0.1009931317290048
	pesos_i(7802) := b"1111111111111111_1111111111111111_1101101110100000_1100100010101110"; -- -0.1420778823108977
	pesos_i(7803) := b"1111111111111111_1111111111111111_1110100100000001_0111000011101110"; -- -0.0898217600193294
	pesos_i(7804) := b"1111111111111111_1111111111111111_1111000011101001_1100101000110110"; -- -0.058932649363189454
	pesos_i(7805) := b"1111111111111111_1111111111111111_1111110110110100_1110011011111011"; -- -0.008958400358086547
	pesos_i(7806) := b"0000000000000000_0000000000000000_0000110000001001_1000101010001110"; -- 0.04702058768333598
	pesos_i(7807) := b"0000000000000000_0000000000000000_0010010001110011_0010010011010000"; -- 0.14238195502493384
	pesos_i(7808) := b"1111111111111111_1111111111111111_1110110111110111_0000011010000100"; -- -0.07044944076300456
	pesos_i(7809) := b"0000000000000000_0000000000000000_0001110000000011_0110010101011011"; -- 0.10942681758745654
	pesos_i(7810) := b"1111111111111111_1111111111111111_1110011100110010_0101011111110100"; -- -0.09688806821542137
	pesos_i(7811) := b"1111111111111111_1111111111111111_1111000101010001_0011100010000100"; -- -0.05735441941783352
	pesos_i(7812) := b"1111111111111111_1111111111111111_1101110100100001_1110011100101100"; -- -0.13620143109170393
	pesos_i(7813) := b"1111111111111111_1111111111111111_1110101010001111_1000010011111101"; -- -0.0837475664908933
	pesos_i(7814) := b"1111111111111111_1111111111111111_1110111100101101_0110010000001010"; -- -0.06571364174658602
	pesos_i(7815) := b"1111111111111111_1111111111111111_1111000100001111_0010100001011000"; -- -0.05836246339728884
	pesos_i(7816) := b"0000000000000000_0000000000000000_0000010000000111_1110000010000111"; -- 0.015745194394994787
	pesos_i(7817) := b"1111111111111111_1111111111111111_1110101111111010_0101110000111010"; -- -0.07821105559298866
	pesos_i(7818) := b"0000000000000000_0000000000000000_0000011000111000_1011001000011111"; -- 0.024302608984120927
	pesos_i(7819) := b"0000000000000000_0000000000000000_0000011101001100_1100100011011101"; -- 0.028515390323846885
	pesos_i(7820) := b"1111111111111111_1111111111111111_1111111110110111_0100100100101111"; -- -0.0011095294734640593
	pesos_i(7821) := b"0000000000000000_0000000000000000_0010001010001110_0001010111101100"; -- 0.13498055475466583
	pesos_i(7822) := b"0000000000000000_0000000000000000_0010011111010010_0111111101011010"; -- 0.15555568655444088
	pesos_i(7823) := b"1111111111111111_1111111111111111_1111101101101101_1000001100000011"; -- -0.017860233177440028
	pesos_i(7824) := b"1111111111111111_1111111111111111_1101101000111010_1011100110110111"; -- -0.14754142085249636
	pesos_i(7825) := b"1111111111111111_1111111111111111_1110100100010001_1100101011011101"; -- -0.08957225900552639
	pesos_i(7826) := b"0000000000000000_0000000000000000_0010100111011101_0011010100001001"; -- 0.16353160348094015
	pesos_i(7827) := b"0000000000000000_0000000000000000_0001010100001101_1010101001110100"; -- 0.0822397740155652
	pesos_i(7828) := b"0000000000000000_0000000000000000_0010001110001011_0110001010101100"; -- 0.13884560302759386
	pesos_i(7829) := b"0000000000000000_0000000000000000_0000111001011010_1000110100000000"; -- 0.05606919523605191
	pesos_i(7830) := b"1111111111111111_1111111111111111_1111111001110100_1001010101110100"; -- -0.006033572289001044
	pesos_i(7831) := b"0000000000000000_0000000000000000_0010010111101111_0111111110101111"; -- 0.1481857111494118
	pesos_i(7832) := b"0000000000000000_0000000000000000_0001011010100100_0110011000011011"; -- 0.08844602745603751
	pesos_i(7833) := b"0000000000000000_0000000000000000_0010001110100000_0100001011110000"; -- 0.13916414597169632
	pesos_i(7834) := b"0000000000000000_0000000000000000_0010110000111111_1010100001010100"; -- 0.1728463367898294
	pesos_i(7835) := b"1111111111111111_1111111111111111_1111001011000101_1011111011101011"; -- -0.051670138863629145
	pesos_i(7836) := b"0000000000000000_0000000000000000_0000010011110110_1111111011100101"; -- 0.01939385498557314
	pesos_i(7837) := b"1111111111111111_1111111111111111_1111110110111111_0110110010010111"; -- -0.00879784876777811
	pesos_i(7838) := b"1111111111111111_1111111111111111_1111011101001101_0110100101111100"; -- -0.03397503584925437
	pesos_i(7839) := b"0000000000000000_0000000000000000_0010000100101011_1010101001110101"; -- 0.12957253792432452
	pesos_i(7840) := b"1111111111111111_1111111111111111_1111111110001010_1010101010000011"; -- -0.0017903737502543149
	pesos_i(7841) := b"1111111111111111_1111111111111111_1101011111001001_0111110100011011"; -- -0.15708177646168192
	pesos_i(7842) := b"1111111111111111_1111111111111111_1111111111010010_0111101000000101"; -- -0.0006946314413419616
	pesos_i(7843) := b"1111111111111111_1111111111111111_1101101111000110_0000010000110001"; -- -0.1415097599029124
	pesos_i(7844) := b"0000000000000000_0000000000000000_0010001001000101_0100101100011000"; -- 0.13386983229933389
	pesos_i(7845) := b"0000000000000000_0000000000000000_0000111101101111_0011011000010111"; -- 0.06029069958492422
	pesos_i(7846) := b"0000000000000000_0000000000000000_0010010101101110_1111100010001111"; -- 0.1462245319642704
	pesos_i(7847) := b"0000000000000000_0000000000000000_0001010001101000_0000001000111111"; -- 0.0797120478881467
	pesos_i(7848) := b"1111111111111111_1111111111111111_1101001101111001_1011110001100111"; -- -0.1739237069339202
	pesos_i(7849) := b"1111111111111111_1111111111111111_1111001100001000_1010101110100000"; -- -0.050648950038022486
	pesos_i(7850) := b"0000000000000000_0000000000000000_0000010010010001_1011110001000110"; -- 0.017848746407426147
	pesos_i(7851) := b"0000000000000000_0000000000000000_0010011111011010_1101111010010001"; -- 0.15568343207172958
	pesos_i(7852) := b"0000000000000000_0000000000000000_0000110111111010_1101110100000000"; -- 0.05460911994029051
	pesos_i(7853) := b"1111111111111111_1111111111111111_1110001101110000_0001100001010010"; -- -0.11157081613033754
	pesos_i(7854) := b"0000000000000000_0000000000000000_0001100011101111_1101001101110001"; -- 0.09740945350617769
	pesos_i(7855) := b"0000000000000000_0000000000000000_0001010110101001_1110101100011010"; -- 0.08462399852999765
	pesos_i(7856) := b"1111111111111111_1111111111111111_1110000101101000_1010000011100110"; -- -0.1194972456901418
	pesos_i(7857) := b"1111111111111111_1111111111111111_1101001100100001_1110101111011001"; -- -0.17526365233489574
	pesos_i(7858) := b"0000000000000000_0000000000000000_0001101010011011_0110010100001000"; -- 0.10393363435159099
	pesos_i(7859) := b"1111111111111111_1111111111111111_1110111010101100_0110111110111001"; -- -0.06768132912884367
	pesos_i(7860) := b"1111111111111111_1111111111111111_1110011111100010_0000010010111110"; -- -0.09420748112699662
	pesos_i(7861) := b"0000000000000000_0000000000000000_0010010000100100_1011011001001000"; -- 0.14118518124764992
	pesos_i(7862) := b"1111111111111111_1111111111111111_1111010010111000_1000011001011111"; -- -0.04405937377568328
	pesos_i(7863) := b"0000000000000000_0000000000000000_0001011111000001_1100101010000111"; -- 0.09280076781903915
	pesos_i(7864) := b"1111111111111111_1111111111111111_1110110110000100_1101011110000000"; -- -0.07219174495808182
	pesos_i(7865) := b"1111111111111111_1111111111111111_1111100110100010_1100010011100010"; -- -0.024860091134946177
	pesos_i(7866) := b"0000000000000000_0000000000000000_0000111110101001_0100001001000001"; -- 0.06117643432137169
	pesos_i(7867) := b"1111111111111111_1111111111111111_1101100110000100_0100001110000010"; -- -0.15032556595113977
	pesos_i(7868) := b"1111111111111111_1111111111111111_1110101110101011_1111111110110001"; -- -0.07940675662845739
	pesos_i(7869) := b"1111111111111111_1111111111111111_1101010101101011_0010110011110001"; -- -0.16633338089036842
	pesos_i(7870) := b"0000000000000000_0000000000000000_0001111111110011_1101011110101110"; -- 0.12481449124092854
	pesos_i(7871) := b"0000000000000000_0000000000000000_0010100110000110_0100101111011000"; -- 0.16220544848349042
	pesos_i(7872) := b"0000000000000000_0000000000000000_0000111100101111_1010111001111000"; -- 0.059321312234013907
	pesos_i(7873) := b"0000000000000000_0000000000000000_0000100011101011_1111100100011100"; -- 0.03485066347149701
	pesos_i(7874) := b"1111111111111111_1111111111111111_1101110101000011_1100110011010011"; -- -0.13568420269694342
	pesos_i(7875) := b"1111111111111111_1111111111111111_1110010001100010_1011010011011010"; -- -0.1078688590351952
	pesos_i(7876) := b"1111111111111111_1111111111111111_1111010101100101_1000001011110110"; -- -0.041419806538127414
	pesos_i(7877) := b"1111111111111111_1111111111111111_1111000000000101_1100111000101000"; -- -0.06241141816618571
	pesos_i(7878) := b"0000000000000000_0000000000000000_0001001011001000_1011101101010110"; -- 0.073375423949282
	pesos_i(7879) := b"1111111111111111_1111111111111111_1111110010000010_1011110001111001"; -- -0.013630123602821407
	pesos_i(7880) := b"0000000000000000_0000000000000000_0000001001000111_1101000111011100"; -- 0.008908382620720459
	pesos_i(7881) := b"0000000000000000_0000000000000000_0001110101010011_0011001001111011"; -- 0.11455073834716045
	pesos_i(7882) := b"1111111111111111_1111111111111111_1110101000010001_1100000101101001"; -- -0.08566657247678094
	pesos_i(7883) := b"0000000000000000_0000000000000000_0001011110100111_1100111000010100"; -- 0.09240425095777148
	pesos_i(7884) := b"0000000000000000_0000000000000000_0001001000100010_1111100000100100"; -- 0.07084608908748827
	pesos_i(7885) := b"0000000000000000_0000000000000000_0010010001010110_1100010110111110"; -- 0.14194904217505058
	pesos_i(7886) := b"1111111111111111_1111111111111111_1110000110000000_0001101101000011"; -- -0.11913900009724068
	pesos_i(7887) := b"1111111111111111_1111111111111111_1111000100101000_0011011001010000"; -- -0.05798016113046213
	pesos_i(7888) := b"0000000000000000_0000000000000000_0000000101010011_0100111110001001"; -- 0.005177470063894157
	pesos_i(7889) := b"0000000000000000_0000000000000000_0000100010110110_1111000011000100"; -- 0.03404145032732647
	pesos_i(7890) := b"1111111111111111_1111111111111111_1111110010100000_1101001111010011"; -- -0.013170968061671876
	pesos_i(7891) := b"0000000000000000_0000000000000000_0001110110001011_1111010101001010"; -- 0.11541684203956305
	pesos_i(7892) := b"0000000000000000_0000000000000000_0001110100011000_1000010001100011"; -- 0.11365535186989811
	pesos_i(7893) := b"1111111111111111_1111111111111111_1101100000111111_0011101111100101"; -- -0.15528512636283906
	pesos_i(7894) := b"1111111111111111_1111111111111111_1110001101111011_1101000100011101"; -- -0.11139195484645406
	pesos_i(7895) := b"0000000000000000_0000000000000000_0010101101100101_0000100010001100"; -- 0.16951039718300098
	pesos_i(7896) := b"0000000000000000_0000000000000000_0001100101111010_0110001101111011"; -- 0.09952375164817685
	pesos_i(7897) := b"0000000000000000_0000000000000000_0000010010011000_1001110000110111"; -- 0.017953647085297834
	pesos_i(7898) := b"1111111111111111_1111111111111111_1111100001111100_0010100000000001"; -- -0.02935552563200456
	pesos_i(7899) := b"1111111111111111_1111111111111111_1111100000000101_0011011110010011"; -- -0.031170393594269645
	pesos_i(7900) := b"1111111111111111_1111111111111111_1110110100010110_1001010001111011"; -- -0.07387420656214257
	pesos_i(7901) := b"1111111111111111_1111111111111111_1110111101101001_0100110010110100"; -- -0.06479950526513752
	pesos_i(7902) := b"1111111111111111_1111111111111111_1101111111010000_1000000110011111"; -- -0.12572469584621726
	pesos_i(7903) := b"0000000000000000_0000000000000000_0010101000100001_0010001101011011"; -- 0.1645681473701853
	pesos_i(7904) := b"0000000000000000_0000000000000000_0010000100000010_1001010011010001"; -- 0.12894563775065046
	pesos_i(7905) := b"1111111111111111_1111111111111111_1110101001101101_1010011110100010"; -- -0.08426430035998309
	pesos_i(7906) := b"0000000000000000_0000000000000000_0001011110101111_0011000100011000"; -- 0.09251696436117535
	pesos_i(7907) := b"1111111111111111_1111111111111111_1101010011111010_1100100001100100"; -- -0.1680483584604963
	pesos_i(7908) := b"0000000000000000_0000000000000000_0010001000100101_0001011101011000"; -- 0.13337846649637977
	pesos_i(7909) := b"0000000000000000_0000000000000000_0000011110100101_1010100001000101"; -- 0.0298714798453363
	pesos_i(7910) := b"0000000000000000_0000000000000000_0001111101011000_1110100100010111"; -- 0.12245041678313305
	pesos_i(7911) := b"1111111111111111_1111111111111111_1110010101111001_1001100000100000"; -- -0.10361336911680875
	pesos_i(7912) := b"0000000000000000_0000000000000000_0001010101100000_1101100010001010"; -- 0.083509000597529
	pesos_i(7913) := b"0000000000000000_0000000000000000_0000000101001110_1110111000110001"; -- 0.005110632975711975
	pesos_i(7914) := b"0000000000000000_0000000000000000_0010000100011110_1110110101010110"; -- 0.1293781600274912
	pesos_i(7915) := b"1111111111111111_1111111111111111_1101110001101111_1111111001000011"; -- -0.1389161192349729
	pesos_i(7916) := b"1111111111111111_1111111111111111_1110101001010010_1110000100101000"; -- -0.08467285895273177
	pesos_i(7917) := b"0000000000000000_0000000000000000_0010000100000101_1110011111011110"; -- 0.12899636440564896
	pesos_i(7918) := b"1111111111111111_1111111111111111_1110000010001110_1101001101111010"; -- -0.12282064703311961
	pesos_i(7919) := b"0000000000000000_0000000000000000_0001110111110010_1000000010101010"; -- 0.11698154597179443
	pesos_i(7920) := b"1111111111111111_1111111111111111_1101110110000111_0000111100110001"; -- -0.13465790793582227
	pesos_i(7921) := b"1111111111111111_1111111111111111_1100111100001000_0011110111111001"; -- -0.19128048575674642
	pesos_i(7922) := b"0000000000000000_0000000000000000_0000101000110011_1000111010001000"; -- 0.039849193751748696
	pesos_i(7923) := b"1111111111111111_1111111111111111_1101100001011101_0010101101000001"; -- -0.1548283544292602
	pesos_i(7924) := b"0000000000000000_0000000000000000_0000010111101100_1101010011011000"; -- 0.02314501066743293
	pesos_i(7925) := b"0000000000000000_0000000000000000_0001101100010011_1111111011010111"; -- 0.10577385673427155
	pesos_i(7926) := b"1111111111111111_1111111111111111_1111010001001100_0001101010110001"; -- -0.045713741053513744
	pesos_i(7927) := b"1111111111111111_1111111111111111_1111100110101011_1111010001101000"; -- -0.024719929287596542
	pesos_i(7928) := b"0000000000000000_0000000000000000_0001101110000001_1001111100010011"; -- 0.10744661527035296
	pesos_i(7929) := b"0000000000000000_0000000000000000_0010000111010101_0000101001000010"; -- 0.13215698359832848
	pesos_i(7930) := b"1111111111111111_1111111111111111_1101011100000100_0000001111101111"; -- -0.1600949803151799
	pesos_i(7931) := b"0000000000000000_0000000000000000_0000001110100111_1101101101111111"; -- 0.01428005081944695
	pesos_i(7932) := b"0000000000000000_0000000000000000_0001000100100110_0010100010111100"; -- 0.06698851185919263
	pesos_i(7933) := b"1111111111111111_1111111111111111_1111110100011111_0011011010001111"; -- -0.011242475673636612
	pesos_i(7934) := b"1111111111111111_1111111111111111_1111010000010001_1100001010011010"; -- -0.046604001318851514
	pesos_i(7935) := b"0000000000000000_0000000000000000_0010011101100001_1010110001010101"; -- 0.15383412427760715
	pesos_i(7936) := b"0000000000000000_0000000000000000_0001110100111011_1001011100100001"; -- 0.11419052655282194
	pesos_i(7937) := b"0000000000000000_0000000000000000_0010110101011110_1011011110111010"; -- 0.1772265272012333
	pesos_i(7938) := b"0000000000000000_0000000000000000_0001001111100101_0101011010101101"; -- 0.0777181788643791
	pesos_i(7939) := b"1111111111111111_1111111111111111_1110110010111010_1111011011011101"; -- -0.07527215110722528
	pesos_i(7940) := b"0000000000000000_0000000000000000_0000001100001010_0110111110011111"; -- 0.011877990920995547
	pesos_i(7941) := b"0000000000000000_0000000000000000_0000000010010000_1000111000010000"; -- 0.002205733230810124
	pesos_i(7942) := b"0000000000000000_0000000000000000_0000000111010110_1100011110001000"; -- 0.007183523762432509
	pesos_i(7943) := b"1111111111111111_1111111111111111_1111010001101000_1000000111000110"; -- -0.04528035080664027
	pesos_i(7944) := b"0000000000000000_0000000000000000_0000010110110101_1001111110011110"; -- 0.022302604828599353
	pesos_i(7945) := b"1111111111111111_1111111111111111_1110100010000010_1011100101011110"; -- -0.09175530856695013
	pesos_i(7946) := b"1111111111111111_1111111111111111_1111000111001011_1010000101111101"; -- -0.05548659033428485
	pesos_i(7947) := b"0000000000000000_0000000000000000_0000011000100100_1101110100110100"; -- 0.024000001132236284
	pesos_i(7948) := b"0000000000000000_0000000000000000_0000100000011101_1010011111000001"; -- 0.03170250371210643
	pesos_i(7949) := b"0000000000000000_0000000000000000_0000101110111011_1011110010000010"; -- 0.045833379540513086
	pesos_i(7950) := b"1111111111111111_1111111111111111_1110000100010110_1110001001111010"; -- -0.12074455750724257
	pesos_i(7951) := b"1111111111111111_1111111111111111_1101010111100000_1100100010110101"; -- -0.16453881809358736
	pesos_i(7952) := b"0000000000000000_0000000000000000_0010011000010010_1001101000000011"; -- 0.14872133809158336
	pesos_i(7953) := b"1111111111111111_1111111111111111_1110101100110001_0100011000001010"; -- -0.08127939461819184
	pesos_i(7954) := b"1111111111111111_1111111111111111_1110011000010001_1101001110111101"; -- -0.10129047990412211
	pesos_i(7955) := b"0000000000000000_0000000000000000_0000010000111010_0111010110011001"; -- 0.016517019070350004
	pesos_i(7956) := b"0000000000000000_0000000000000000_0000101011111101_0111110000110001"; -- 0.042930375972374465
	pesos_i(7957) := b"1111111111111111_1111111111111111_1110101011101001_0000000011101101"; -- -0.08238214701350165
	pesos_i(7958) := b"1111111111111111_1111111111111111_1110010001110011_0110001011011100"; -- -0.1076143468086197
	pesos_i(7959) := b"0000000000000000_0000000000000000_0000101101010011_0001101110101100"; -- 0.04423687887003238
	pesos_i(7960) := b"1111111111111111_1111111111111111_1100101100111001_0010111000010101"; -- -0.20615875240482234
	pesos_i(7961) := b"0000000000000000_0000000000000000_0001101000000110_0100000011011100"; -- 0.10165791876082024
	pesos_i(7962) := b"1111111111111111_1111111111111111_1111001111111001_0000011111110001"; -- -0.04698133819102124
	pesos_i(7963) := b"0000000000000000_0000000000000000_0000100100100111_1101111000101100"; -- 0.03576458524687472
	pesos_i(7964) := b"1111111111111111_1111111111111111_1110011001000101_1000010110110111"; -- -0.10050167354527033
	pesos_i(7965) := b"1111111111111111_1111111111111111_1110000011000110_0101110011100100"; -- -0.12197322299975062
	pesos_i(7966) := b"1111111111111111_1111111111111111_1111100011000100_1010111100001000"; -- -0.0282488447212588
	pesos_i(7967) := b"0000000000000000_0000000000000000_0010010001111011_0101100101101100"; -- 0.14250716103272734
	pesos_i(7968) := b"0000000000000000_0000000000000000_0001010010100110_0001010001010011"; -- 0.08065917032561234
	pesos_i(7969) := b"0000000000000000_0000000000000000_0001111010001011_0110010101100010"; -- 0.11931451461600417
	pesos_i(7970) := b"1111111111111111_1111111111111111_1110100111101001_1110010010101111"; -- -0.08627482155500861
	pesos_i(7971) := b"0000000000000000_0000000000000000_0001000011010011_0111111011110101"; -- 0.06572717174992283
	pesos_i(7972) := b"0000000000000000_0000000000000000_0000101000110000_1110110001111101"; -- 0.039809017605382586
	pesos_i(7973) := b"0000000000000000_0000000000000000_0001100111110000_1110011110101100"; -- 0.1013321681006906
	pesos_i(7974) := b"0000000000000000_0000000000000000_0001010101010010_1010101001101111"; -- 0.08329262933907415
	pesos_i(7975) := b"0000000000000000_0000000000000000_0000111100111110_0100111010111010"; -- 0.0595444874275316
	pesos_i(7976) := b"1111111111111111_1111111111111111_1111100100011011_0001000010010010"; -- -0.026930774997283496
	pesos_i(7977) := b"1111111111111111_1111111111111111_1111001010110111_1011000100001010"; -- -0.051884589347286826
	pesos_i(7978) := b"1111111111111111_1111111111111111_1111100011010110_1110100011110000"; -- -0.02797073487230218
	pesos_i(7979) := b"0000000000000000_0000000000000000_0001001000010001_1011001000010010"; -- 0.07058251316921593
	pesos_i(7980) := b"1111111111111111_1111111111111111_1111001110011101_1100101001000110"; -- -0.04837356374711472
	pesos_i(7981) := b"1111111111111111_1111111111111111_1101010000101111_0010110101110000"; -- -0.17115512870177557
	pesos_i(7982) := b"1111111111111111_1111111111111111_1111100000110110_0011001101010010"; -- -0.030422966512464008
	pesos_i(7983) := b"1111111111111111_1111111111111111_1110011101011111_1000101110101100"; -- -0.09619833992469151
	pesos_i(7984) := b"1111111111111111_1111111111111111_1110101010001111_1101010101101111"; -- -0.08374277153666537
	pesos_i(7985) := b"0000000000000000_0000000000000000_0000000111000101_0000100001100110"; -- 0.006912732139338426
	pesos_i(7986) := b"0000000000000000_0000000000000000_0000101010010100_0001110011111111"; -- 0.04132252897997294
	pesos_i(7987) := b"0000000000000000_0000000000000000_0010011111111100_0110000010111011"; -- 0.15619473039892318
	pesos_i(7988) := b"1111111111111111_1111111111111111_1111111011010000_0001111010010111"; -- -0.004636848534796457
	pesos_i(7989) := b"1111111111111111_1111111111111111_1110000100000010_1011010000011101"; -- -0.121052496827461
	pesos_i(7990) := b"0000000000000000_0000000000000000_0000110101110010_0000101100001010"; -- 0.05252140993784338
	pesos_i(7991) := b"1111111111111111_1111111111111111_1111111000100010_0001100110110111"; -- -0.007292168396667407
	pesos_i(7992) := b"1111111111111111_1111111111111111_1110100100110101_1100011011001110"; -- -0.08902318451799371
	pesos_i(7993) := b"1111111111111111_1111111111111111_1110011111101101_1100001011100001"; -- -0.09402830139917828
	pesos_i(7994) := b"0000000000000000_0000000000000000_0010100011001010_0101101110010110"; -- 0.15933773443427995
	pesos_i(7995) := b"1111111111111111_1111111111111111_1101110100011001_1011100000110000"; -- -0.1363263019108461
	pesos_i(7996) := b"0000000000000000_0000000000000000_0001000101101011_0000001100010101"; -- 0.06803912421750491
	pesos_i(7997) := b"0000000000000000_0000000000000000_0001110101100000_1000101001001110"; -- 0.11475433733586463
	pesos_i(7998) := b"0000000000000000_0000000000000000_0001011010110001_0010101111110100"; -- 0.08864092548232594
	pesos_i(7999) := b"0000000000000000_0000000000000000_0010000011000111_0000010110100011"; -- 0.12803683491859294
	pesos_i(8000) := b"0000000000000000_0000000000000000_0010101110110111_0100001000111011"; -- 0.17076505615596396
	pesos_i(8001) := b"1111111111111111_1111111111111111_1101100010011101_0111110000111110"; -- -0.15384696464916967
	pesos_i(8002) := b"0000000000000000_0000000000000000_0010011000111010_0011010110010100"; -- 0.14932570325870492
	pesos_i(8003) := b"0000000000000000_0000000000000000_0010010000011011_0100010001000010"; -- 0.14104105576908602
	pesos_i(8004) := b"1111111111111111_1111111111111111_1110110101100111_1010011010000101"; -- -0.07263716927398116
	pesos_i(8005) := b"0000000000000000_0000000000000000_0001110100100000_0001010111110100"; -- 0.11377083979697816
	pesos_i(8006) := b"0000000000000000_0000000000000000_0010001001000101_1011011100110011"; -- 0.1338762759976061
	pesos_i(8007) := b"0000000000000000_0000000000000000_0000101010111011_0011111101110111"; -- 0.041919676428381174
	pesos_i(8008) := b"0000000000000000_0000000000000000_0010011011010111_0111110111001100"; -- 0.1517256376130593
	pesos_i(8009) := b"0000000000000000_0000000000000000_0010001011101010_1000001101110010"; -- 0.13639089138866764
	pesos_i(8010) := b"1111111111111111_1111111111111111_1111010111000000_0000110111110111"; -- -0.040038230222881686
	pesos_i(8011) := b"1111111111111111_1111111111111111_1110011100111110_0001001101000011"; -- -0.09670905690629031
	pesos_i(8012) := b"0000000000000000_0000000000000000_0001100111000101_1001001111100011"; -- 0.10067104608954637
	pesos_i(8013) := b"0000000000000000_0000000000000000_0000101111101101_1110010110100010"; -- 0.046598770118882984
	pesos_i(8014) := b"1111111111111111_1111111111111111_1101101100111101_1011100111000000"; -- -0.14358939222481362
	pesos_i(8015) := b"0000000000000000_0000000000000000_0000010111111010_1001000100010000"; -- 0.0233545936197396
	pesos_i(8016) := b"1111111111111111_1111111111111111_1111011010111100_0100100100011100"; -- -0.036189489910250894
	pesos_i(8017) := b"0000000000000000_0000000000000000_0010010110010101_0100101101011010"; -- 0.14680930090624178
	pesos_i(8018) := b"1111111111111111_1111111111111111_1111001111110101_0011111011100101"; -- -0.04703909788618161
	pesos_i(8019) := b"0000000000000000_0000000000000000_0001110110001000_1110111110110011"; -- 0.11537073252272874
	pesos_i(8020) := b"0000000000000000_0000000000000000_0000011110001010_0111001111100111"; -- 0.029456371118550213
	pesos_i(8021) := b"1111111111111111_1111111111111111_1111111001100110_0010101010000101"; -- -0.006253569146536477
	pesos_i(8022) := b"1111111111111111_1111111111111111_1110000000111001_0000111110100001"; -- -0.12412931755659803
	pesos_i(8023) := b"1111111111111111_1111111111111111_1111101000100010_0101110110001111"; -- -0.02291312462743983
	pesos_i(8024) := b"1111111111111111_1111111111111111_1110100011000100_0100111010000010"; -- -0.09075459783842664
	pesos_i(8025) := b"0000000000000000_0000000000000000_0000010001000100_1001001101101001"; -- 0.01667138389831054
	pesos_i(8026) := b"0000000000000000_0000000000000000_0000111001111110_0001011100110110"; -- 0.056611490931829885
	pesos_i(8027) := b"1111111111111111_1111111111111111_1111010011100000_0011110111011011"; -- -0.0434533444135963
	pesos_i(8028) := b"0000000000000000_0000000000000000_0010000110111101_0110110000001010"; -- 0.13179660086113232
	pesos_i(8029) := b"1111111111111111_1111111111111111_1101110001001010_1011111000110100"; -- -0.13948451255287125
	pesos_i(8030) := b"1111111111111111_1111111111111111_1101011100011010_1010110001111001"; -- -0.15974924133063464
	pesos_i(8031) := b"1111111111111111_1111111111111111_1101100011111000_0111000100110001"; -- -0.1524590736566228
	pesos_i(8032) := b"0000000000000000_0000000000000000_0001100101010000_0000000010100000"; -- 0.09887699033079148
	pesos_i(8033) := b"0000000000000000_0000000000000000_0001001111110110_1000100010111101"; -- 0.07798056245149551
	pesos_i(8034) := b"1111111111111111_1111111111111111_1111111000100001_1001001111101100"; -- -0.007300143142268926
	pesos_i(8035) := b"0000000000000000_0000000000000000_0010001111001111_1101100111110100"; -- 0.13989031046112707
	pesos_i(8036) := b"0000000000000000_0000000000000000_0010001110011000_1110110100001001"; -- 0.13905221433911275
	pesos_i(8037) := b"0000000000000000_0000000000000000_0010001010110011_1010101100111110"; -- 0.1355540300282395
	pesos_i(8038) := b"0000000000000000_0000000000000000_0000101110001110_1100110100101011"; -- 0.0451477270358834
	pesos_i(8039) := b"0000000000000000_0000000000000000_0001110001110001_0110010001010010"; -- 0.11110522260694025
	pesos_i(8040) := b"0000000000000000_0000000000000000_0000000101010101_1101001111001100"; -- 0.005215871066186206
	pesos_i(8041) := b"1111111111111111_1111111111111111_1110001101110011_0000110110110000"; -- -0.11152567341247445
	pesos_i(8042) := b"1111111111111111_1111111111111111_1101101001010011_1011100110100011"; -- -0.14715995561862036
	pesos_i(8043) := b"0000000000000000_0000000000000000_0010101110110110_0111000110101010"; -- 0.17075262446506018
	pesos_i(8044) := b"1111111111111111_1111111111111111_1110011010010000_0101100110111010"; -- -0.09935988635629678
	pesos_i(8045) := b"1111111111111111_1111111111111111_1111010001100001_0110110111010010"; -- -0.045388351568092615
	pesos_i(8046) := b"1111111111111111_1111111111111111_1110100010100010_0100010110011011"; -- -0.09127392736780564
	pesos_i(8047) := b"1111111111111111_1111111111111111_1110011111100010_1001111000100001"; -- -0.09419833841641308
	pesos_i(8048) := b"0000000000000000_0000000000000000_0000101111001000_0010001010001101"; -- 0.046022567173584106
	pesos_i(8049) := b"1111111111111111_1111111111111111_1110000010110110_0111000101110011"; -- -0.12221613830594356
	pesos_i(8050) := b"0000000000000000_0000000000000000_0010010100001110_1110000100001110"; -- 0.1447582874111407
	pesos_i(8051) := b"0000000000000000_0000000000000000_0001010110001001_0101010100101010"; -- 0.08412678032025804
	pesos_i(8052) := b"0000000000000000_0000000000000000_0000111100010111_1011111101011010"; -- 0.058956107579877015
	pesos_i(8053) := b"1111111111111111_1111111111111111_1111001000100011_0000111100111110"; -- -0.054152533952973154
	pesos_i(8054) := b"0000000000000000_0000000000000000_0010101100010111_0111000001011001"; -- 0.16832639868916802
	pesos_i(8055) := b"1111111111111111_1111111111111111_1101000000101100_0101111011011100"; -- -0.18682295916137207
	pesos_i(8056) := b"0000000000000000_0000000000000000_0000001101001100_1110011011001000"; -- 0.012892173714110722
	pesos_i(8057) := b"1111111111111111_1111111111111111_1101101011011111_0110101110010010"; -- -0.14502837824584966
	pesos_i(8058) := b"1111111111111111_1111111111111111_1111101101000111_1010000101100001"; -- -0.018438256949304458
	pesos_i(8059) := b"1111111111111111_1111111111111111_1110100100011111_1011010111101000"; -- -0.08935988501878459
	pesos_i(8060) := b"0000000000000000_0000000000000000_0000110111010010_0110011111011100"; -- 0.05399178629290297
	pesos_i(8061) := b"1111111111111111_1111111111111111_1110000101010000_0110101001011001"; -- -0.11986670796790273
	pesos_i(8062) := b"0000000000000000_0000000000000000_0000010010011011_1100110000011001"; -- 0.018002277457829716
	pesos_i(8063) := b"1111111111111111_1111111111111111_1111111001101100_1000110001100001"; -- -0.006156183494669205
	pesos_i(8064) := b"1111111111111111_1111111111111111_1111001001001100_0001000010100000"; -- -0.05352684113159384
	pesos_i(8065) := b"0000000000000000_0000000000000000_0010101101001101_1000101101100110"; -- 0.16915198563509837
	pesos_i(8066) := b"0000000000000000_0000000000000000_0010101000100110_1111001000111011"; -- 0.16465677194021044
	pesos_i(8067) := b"1111111111111111_1111111111111111_1111101101100110_1000101110011011"; -- -0.017966532354175595
	pesos_i(8068) := b"1111111111111111_1111111111111111_1101111010000100_1010001111111000"; -- -0.13078856660496807
	pesos_i(8069) := b"1111111111111111_1111111111111111_1110100000001110_0101111001001100"; -- -0.09353075630791831
	pesos_i(8070) := b"0000000000000000_0000000000000000_0010101000000110_1110011010001101"; -- 0.16416779473332282
	pesos_i(8071) := b"0000000000000000_0000000000000000_0000000100100000_1011010011011111"; -- 0.004405311895889657
	pesos_i(8072) := b"0000000000000000_0000000000000000_0001011010000011_1100011110001111"; -- 0.0879482960405156
	pesos_i(8073) := b"0000000000000000_0000000000000000_0000010110111101_0110100100010001"; -- 0.022421423685309957
	pesos_i(8074) := b"1111111111111111_1111111111111111_1111101100110001_0111110011010101"; -- -0.018776128701304733
	pesos_i(8075) := b"1111111111111111_1111111111111111_1111001110011011_1001101111111100"; -- -0.04840684032480915
	pesos_i(8076) := b"1111111111111111_1111111111111111_1110010011010110_1010111110001101"; -- -0.10609915549825907
	pesos_i(8077) := b"1111111111111111_1111111111111111_1101011111010001_0010001000110011"; -- -0.15696512474216884
	pesos_i(8078) := b"1111111111111111_1111111111111111_1101101000101100_1010010000100001"; -- -0.14775633037952424
	pesos_i(8079) := b"0000000000000000_0000000000000000_0000000101001100_0000110001001110"; -- 0.005066651269526562
	pesos_i(8080) := b"1111111111111111_1111111111111111_1111111111111110_0000000000110101"; -- -3.0505160765165185e-05
	pesos_i(8081) := b"1111111111111111_1111111111111111_1110000100001111_1111011111100010"; -- -0.12085009315750558
	pesos_i(8082) := b"1111111111111111_1111111111111111_1111010111110001_0110011001001010"; -- -0.039285284921294614
	pesos_i(8083) := b"1111111111111111_1111111111111111_1110110111110011_1001101111011110"; -- -0.0705015739130868
	pesos_i(8084) := b"1111111111111111_1111111111111111_1111100111001010_0010011101001101"; -- -0.024259132181617262
	pesos_i(8085) := b"1111111111111111_1111111111111111_1110001011110010_1101101111110000"; -- -0.11348176372393261
	pesos_i(8086) := b"0000000000000000_0000000000000000_0001100011100010_0001110110010101"; -- 0.09720024965711938
	pesos_i(8087) := b"1111111111111111_1111111111111111_1101000001100000_1101010010000110"; -- -0.18602248876525895
	pesos_i(8088) := b"0000000000000000_0000000000000000_0010110000011001_1111100111011011"; -- 0.17227136217354005
	pesos_i(8089) := b"1111111111111111_1111111111111111_1110100001000000_1101011111111011"; -- -0.09276056397479163
	pesos_i(8090) := b"0000000000000000_0000000000000000_0001011110101001_0010010101001101"; -- 0.09242470858654743
	pesos_i(8091) := b"1111111111111111_1111111111111111_1101111100100011_1100011110100011"; -- -0.12836029311361555
	pesos_i(8092) := b"1111111111111111_1111111111111111_1110110100110110_1001111001010111"; -- -0.07338533749065265
	pesos_i(8093) := b"1111111111111111_1111111111111111_1111111000110110_0011001111110111"; -- -0.006985427984924516
	pesos_i(8094) := b"1111111111111111_1111111111111111_1111011101000101_0001100000100011"; -- -0.03410195483842693
	pesos_i(8095) := b"1111111111111111_1111111111111111_1101111100001000_0010101110101001"; -- -0.12878157724430245
	pesos_i(8096) := b"0000000000000000_0000000000000000_0000111001000010_1001101001100010"; -- 0.05570378204946988
	pesos_i(8097) := b"0000000000000000_0000000000000000_0010011111111001_1001001000111000"; -- 0.1561519037184478
	pesos_i(8098) := b"0000000000000000_0000000000000000_0000011111111101_0100110011110100"; -- 0.03120881033870887
	pesos_i(8099) := b"0000000000000000_0000000000000000_0001111110111000_0110000110000010"; -- 0.12390717906423206
	pesos_i(8100) := b"0000000000000000_0000000000000000_0010100100101111_1010000000001000"; -- 0.16088295159552948
	pesos_i(8101) := b"0000000000000000_0000000000000000_0010011010011001_1001111010011110"; -- 0.15078154908216782
	pesos_i(8102) := b"0000000000000000_0000000000000000_0001110011010101_1000100010100101"; -- 0.11263326667718665
	pesos_i(8103) := b"0000000000000000_0000000000000000_0010001001101111_1111101001100000"; -- 0.13452114906374693
	pesos_i(8104) := b"1111111111111111_1111111111111111_1110111101111110_1101010100110100"; -- -0.06447093472109645
	pesos_i(8105) := b"0000000000000000_0000000000000000_0010000101001000_0011011101111011"; -- 0.13000818967956151
	pesos_i(8106) := b"0000000000000000_0000000000000000_0001011111010001_0101101101001000"; -- 0.09303827767073916
	pesos_i(8107) := b"0000000000000000_0000000000000000_0001000100110000_1100010100010001"; -- 0.06715041787411669
	pesos_i(8108) := b"0000000000000000_0000000000000000_0000100011011110_1001101011001100"; -- 0.03464667775054024
	pesos_i(8109) := b"0000000000000000_0000000000000000_0010011110010101_1000000111010000"; -- 0.15462504703645039
	pesos_i(8110) := b"0000000000000000_0000000000000000_0010100000100000_0111110100111101"; -- 0.1567457460839058
	pesos_i(8111) := b"1111111111111111_1111111111111111_1111110010101001_0111110000110110"; -- -0.013038861031526548
	pesos_i(8112) := b"1111111111111111_1111111111111111_1111011010110100_1111111101111110"; -- -0.03630068945922443
	pesos_i(8113) := b"1111111111111111_1111111111111111_1110100101010010_1001110100111010"; -- -0.08858315790985871
	pesos_i(8114) := b"1111111111111111_1111111111111111_1110001110001110_1110101010010100"; -- -0.11110052005844336
	pesos_i(8115) := b"0000000000000000_0000000000000000_0010010010000101_1011111100000101"; -- 0.14266580453300015
	pesos_i(8116) := b"1111111111111111_1111111111111111_1111000101110100_0001111100111100"; -- -0.05682186865359424
	pesos_i(8117) := b"1111111111111111_1111111111111111_1111101010111110_1100100000111000"; -- -0.020526396076004826
	pesos_i(8118) := b"1111111111111111_1111111111111111_1110100000010010_1110010110010100"; -- -0.09346165787548721
	pesos_i(8119) := b"1111111111111111_1111111111111111_1101010101000011_0011000100011001"; -- -0.16694348464366823
	pesos_i(8120) := b"0000000000000000_0000000000000000_0001000100011010_0111000110110001"; -- 0.06680975494955446
	pesos_i(8121) := b"0000000000000000_0000000000000000_0010010100101110_0001010101000010"; -- 0.14523442138435944
	pesos_i(8122) := b"1111111111111111_1111111111111111_1111010011100101_1001101100001001"; -- -0.0433714964258345
	pesos_i(8123) := b"1111111111111111_1111111111111111_1101001110000000_0100111111011000"; -- -0.1738233658612755
	pesos_i(8124) := b"1111111111111111_1111111111111111_1111101101001100_1001000111110100"; -- -0.01836288260085989
	pesos_i(8125) := b"0000000000000000_0000000000000000_0010111010110111_1010001001001101"; -- 0.1824895322458092
	pesos_i(8126) := b"0000000000000000_0000000000000000_0001010100111111_1110110011110011"; -- 0.08300667700620334
	pesos_i(8127) := b"0000000000000000_0000000000000000_0001001100010111_0100011000001111"; -- 0.07457387791860061
	pesos_i(8128) := b"0000000000000000_0000000000000000_0000111010001010_0000111010010011"; -- 0.056794081619896186
	pesos_i(8129) := b"0000000000000000_0000000000000000_0000000011000010_1010000111010010"; -- 0.002969850211969275
	pesos_i(8130) := b"1111111111111111_1111111111111111_1111010111010100_1001100001110011"; -- -0.03972479996471994
	pesos_i(8131) := b"0000000000000000_0000000000000000_0000111101110101_1011111000101010"; -- 0.060390362908459144
	pesos_i(8132) := b"1111111111111111_1111111111111111_1101101110110000_0000101110000110"; -- -0.14184501632125346
	pesos_i(8133) := b"1111111111111111_1111111111111111_1110000111101110_1000011000010101"; -- -0.11745416634780316
	pesos_i(8134) := b"1111111111111111_1111111111111111_1110001111010100_0110010001010010"; -- -0.11004040713797329
	pesos_i(8135) := b"1111111111111111_1111111111111111_1111011110001011_1100011011010011"; -- -0.033023427551208795
	pesos_i(8136) := b"1111111111111111_1111111111111111_1110011111111101_0111101101010010"; -- -0.09378842583254561
	pesos_i(8137) := b"0000000000000000_0000000000000000_0010001000001011_1111001111110100"; -- 0.13299488737563742
	pesos_i(8138) := b"1111111111111111_1111111111111111_1111001010100010_1101001001010010"; -- -0.05220304016364432
	pesos_i(8139) := b"1111111111111111_1111111111111111_1110110111110001_0000101010010001"; -- -0.07054075212339277
	pesos_i(8140) := b"0000000000000000_0000000000000000_0001100000011110_0001111001010111"; -- 0.09420957214801597
	pesos_i(8141) := b"0000000000000000_0000000000000000_0001100100011111_1011000100100001"; -- 0.09813983016436618
	pesos_i(8142) := b"0000000000000000_0000000000000000_0001011111000001_0000011000000011"; -- 0.09278905450586189
	pesos_i(8143) := b"0000000000000000_0000000000000000_0011011010101000_0011011100011101"; -- 0.21350426148253326
	pesos_i(8144) := b"0000000000000000_0000000000000000_0010101011111001_0100010011001100"; -- 0.16786603897353328
	pesos_i(8145) := b"1111111111111111_1111111111111111_1111111111000110_0000100100000010"; -- -0.0008844728679662324
	pesos_i(8146) := b"1111111111111111_1111111111111111_1111011111010010_0110010111111001"; -- -0.03194582626855434
	pesos_i(8147) := b"0000000000000000_0000000000000000_0001100011011000_1100010011111110"; -- 0.09705763998915487
	pesos_i(8148) := b"0000000000000000_0000000000000000_0001101101001000_1000001101100101"; -- 0.10657521448431694
	pesos_i(8149) := b"1111111111111111_1111111111111111_1111111110100001_1000110111001010"; -- -0.0014411336322620873
	pesos_i(8150) := b"1111111111111111_1111111111111111_1111001010101010_1101101001100001"; -- -0.052080489447969086
	pesos_i(8151) := b"1111111111111111_1111111111111111_1101110101110101_1111101010101111"; -- -0.1349185298640992
	pesos_i(8152) := b"1111111111111111_1111111111111111_1111010000111000_0110100011111110"; -- -0.04601424971447842
	pesos_i(8153) := b"1111111111111111_1111111111111111_1111110100001111_0000001101010111"; -- -0.011489668984641257
	pesos_i(8154) := b"0000000000000000_0000000000000000_0001100110000000_0110111011010000"; -- 0.09961597988582402
	pesos_i(8155) := b"1111111111111111_1111111111111111_1110010000000011_1110100010111000"; -- -0.10931535251525946
	pesos_i(8156) := b"0000000000000000_0000000000000000_0010101100111000_1011000100011111"; -- 0.1688337994124348
	pesos_i(8157) := b"0000000000000000_0000000000000000_0000001000011111_1011001110011101"; -- 0.00829622836264174
	pesos_i(8158) := b"1111111111111111_1111111111111111_1111001001010110_0010101010001100"; -- -0.053372708204472735
	pesos_i(8159) := b"1111111111111111_1111111111111111_1101101010111010_1100100010000110"; -- -0.145587413056598
	pesos_i(8160) := b"1111111111111111_1111111111111111_1110110110011110_1101101101100000"; -- -0.07179478560720128
	pesos_i(8161) := b"0000000000000000_0000000000000000_0001010111000100_1110101100011101"; -- 0.08503598642718717
	pesos_i(8162) := b"0000000000000000_0000000000000000_0000001001001111_0101001011000101"; -- 0.009022877810732294
	pesos_i(8163) := b"1111111111111111_1111111111111111_1110110110100110_0000010111110111"; -- -0.07168543550783235
	pesos_i(8164) := b"0000000000000000_0000000000000000_0010000000111100_0110011000110111"; -- 0.1259216197553756
	pesos_i(8165) := b"1111111111111111_1111111111111111_1101011011101010_1110010010011110"; -- -0.16047831660157114
	pesos_i(8166) := b"1111111111111111_1111111111111111_1101010011011111_1101100011000001"; -- -0.16845937057231974
	pesos_i(8167) := b"1111111111111111_1111111111111111_1111000110011011_1000101001100100"; -- -0.05622038892375851
	pesos_i(8168) := b"1111111111111111_1111111111111111_1101001101110110_1110111001000100"; -- -0.17396651111391492
	pesos_i(8169) := b"1111111111111111_1111111111111111_1101011110100101_0000000100010110"; -- -0.15763848514880757
	pesos_i(8170) := b"1111111111111111_1111111111111111_1111011110000001_1011111010010001"; -- -0.033176507587023986
	pesos_i(8171) := b"0000000000000000_0000000000000000_0000011001011001_1100000011001001"; -- 0.024807023042962333
	pesos_i(8172) := b"0000000000000000_0000000000000000_0010011000110001_0011000010000000"; -- 0.14918807146180435
	pesos_i(8173) := b"0000000000000000_0000000000000000_0010011111000100_1011010001100010"; -- 0.15534522432473427
	pesos_i(8174) := b"1111111111111111_1111111111111111_1101110110010011_0100111100101010"; -- -0.13447098956523218
	pesos_i(8175) := b"0000000000000000_0000000000000000_0010010101011101_0110011110100110"; -- 0.14595649524908488
	pesos_i(8176) := b"0000000000000000_0000000000000000_0010001100110001_1001101001100001"; -- 0.13747563243742253
	pesos_i(8177) := b"1111111111111111_1111111111111111_1110111001100010_0011111001110000"; -- -0.0688134170355151
	pesos_i(8178) := b"1111111111111111_1111111111111111_1111011111011011_1000010111100010"; -- -0.03180659523690498
	pesos_i(8179) := b"0000000000000000_0000000000000000_0010101101010110_0010001101101001"; -- 0.16928311644829494
	pesos_i(8180) := b"1111111111111111_1111111111111111_1110110110000100_1111100001111001"; -- -0.07218977981736147
	pesos_i(8181) := b"0000000000000000_0000000000000000_0000111000001100_1011011110001011"; -- 0.05488154555032549
	pesos_i(8182) := b"0000000000000000_0000000000000000_0000001011000001_0001011100100010"; -- 0.010758825042192057
	pesos_i(8183) := b"0000000000000000_0000000000000000_0001111001011110_0101101001100101"; -- 0.11862721417999973
	pesos_i(8184) := b"1111111111111111_1111111111111111_1101100100000001_0011101111111010"; -- -0.1523249162252211
	pesos_i(8185) := b"0000000000000000_0000000000000000_0001111111111101_1101011010010011"; -- 0.12496701333795253
	pesos_i(8186) := b"0000000000000000_0000000000000000_0000000001000011_1110011111011001"; -- 0.0010361579627236543
	pesos_i(8187) := b"0000000000000000_0000000000000000_0010010001011001_0010011101010110"; -- 0.141985376812935
	pesos_i(8188) := b"1111111111111111_1111111111111111_1110011000011100_1010000100110000"; -- -0.10112564626884576
	pesos_i(8189) := b"0000000000000000_0000000000000000_0000010001010110_1101100011110111"; -- 0.016950187981346492
	pesos_i(8190) := b"0000000000000000_0000000000000000_0000001001000011_1101000001100001"; -- 0.008847259258953879
	pesos_i(8191) := b"1111111111111111_1111111111111111_1111011100101101_0000001110001111"; -- -0.03446939235325384
	pesos_i(8192) := b"0000000000000000_0000000000000000_0010101001100111_1011101100111000"; -- 0.16564531432245638
	pesos_i(8193) := b"1111111111111111_1111111111111111_1111110111100101_0000011100010010"; -- -0.00822406596582874
	pesos_i(8194) := b"1111111111111111_1111111111111111_1110110101000000_0001101110110001"; -- -0.07324053692437141
	pesos_i(8195) := b"1111111111111111_1111111111111111_1101101010101000_1000101000100000"; -- -0.14586579047324852
	pesos_i(8196) := b"1111111111111111_1111111111111111_1101110100101001_1110000101110011"; -- -0.13607970192685107
	pesos_i(8197) := b"1111111111111111_1111111111111111_1110000101010001_1111001000111000"; -- -0.11984335067507895
	pesos_i(8198) := b"1111111111111111_1111111111111111_1111101100111111_0011010000111011"; -- -0.018566833126337137
	pesos_i(8199) := b"1111111111111111_1111111111111111_1101111100001000_0001001011010000"; -- -0.12878305835293058
	pesos_i(8200) := b"1111111111111111_1111111111111111_1111111000000101_1101001110101111"; -- -0.007723588806590715
	pesos_i(8201) := b"0000000000000000_0000000000000000_0000110011111000_0000100111011000"; -- 0.05065976642383683
	pesos_i(8202) := b"0000000000000000_0000000000000000_0000110100101110_1100111101010110"; -- 0.051495512505101614
	pesos_i(8203) := b"0000000000000000_0000000000000000_0010100001001011_0001100101111010"; -- 0.15739592774777794
	pesos_i(8204) := b"1111111111111111_1111111111111111_1101101100010111_1011111100100100"; -- -0.14416890499160095
	pesos_i(8205) := b"1111111111111111_1111111111111111_1111110111001110_0110011000101110"; -- -0.0085693491199213
	pesos_i(8206) := b"0000000000000000_0000000000000000_0001010111010100_1000010111110000"; -- 0.08527409651060926
	pesos_i(8207) := b"1111111111111111_1111111111111111_1110100000111011_1100110010101000"; -- -0.09283753289968805
	pesos_i(8208) := b"1111111111111111_1111111111111111_1101111010010011_1001011111110111"; -- -0.13056040024129814
	pesos_i(8209) := b"0000000000000000_0000000000000000_0001111000001001_1111011001111100"; -- 0.11733952061234976
	pesos_i(8210) := b"0000000000000000_0000000000000000_0001000010100000_0111001001010010"; -- 0.06494822028626615
	pesos_i(8211) := b"0000000000000000_0000000000000000_0010000101101100_0101100110010001"; -- 0.13055953777532175
	pesos_i(8212) := b"0000000000000000_0000000000000000_0001101001011011_0101010001101010"; -- 0.10295608118185046
	pesos_i(8213) := b"0000000000000000_0000000000000000_0001111111111001_0101011110100001"; -- 0.12489841159356371
	pesos_i(8214) := b"1111111111111111_1111111111111111_1110111100110011_0001110010100010"; -- -0.06562634515162605
	pesos_i(8215) := b"0000000000000000_0000000000000000_0000001100011010_0001000100111001"; -- 0.012116505041937876
	pesos_i(8216) := b"1111111111111111_1111111111111111_1101010101111001_0110110100111101"; -- -0.16611592533593864
	pesos_i(8217) := b"0000000000000000_0000000000000000_0001100101011100_0011110111110100"; -- 0.09906375133494225
	pesos_i(8218) := b"0000000000000000_0000000000000000_0000100001101000_0110110110111100"; -- 0.03284345468264708
	pesos_i(8219) := b"0000000000000000_0000000000000000_0001100100001111_1001101000000000"; -- 0.09789431096944415
	pesos_i(8220) := b"0000000000000000_0000000000000000_0001111101101101_0101010011111110"; -- 0.12276202395746984
	pesos_i(8221) := b"1111111111111111_1111111111111111_1111100100011110_1010111001101010"; -- -0.026875590357765485
	pesos_i(8222) := b"0000000000000000_0000000000000000_0000000110000111_0101101000111010"; -- 0.005971564369969871
	pesos_i(8223) := b"0000000000000000_0000000000000000_0001001100101101_1100101111100111"; -- 0.07491754900986293
	pesos_i(8224) := b"1111111111111111_1111111111111111_1101100110000101_1010011110110011"; -- -0.15030433542126884
	pesos_i(8225) := b"0000000000000000_0000000000000000_0000001010100101_1110111110110000"; -- 0.010344486793838523
	pesos_i(8226) := b"0000000000000000_0000000000000000_0000011000100100_0010011111100011"; -- 0.023989193885384993
	pesos_i(8227) := b"1111111111111111_1111111111111111_1101111100111011_0111001100000010"; -- -0.12799912638636543
	pesos_i(8228) := b"1111111111111111_1111111111111111_1101101001001010_0011010100110010"; -- -0.14730517897498155
	pesos_i(8229) := b"1111111111111111_1111111111111111_1111111101010001_0111101100110000"; -- -0.0026629455672788466
	pesos_i(8230) := b"0000000000000000_0000000000000000_0001010010101000_1101100101110010"; -- 0.08070143742216994
	pesos_i(8231) := b"0000000000000000_0000000000000000_0001110011000110_0001010110111110"; -- 0.11239753617066567
	pesos_i(8232) := b"1111111111111111_1111111111111111_1111001100010001_1111101010011101"; -- -0.05050691296814061
	pesos_i(8233) := b"1111111111111111_1111111111111111_1111000000101101_0011000101111101"; -- -0.061810404838970934
	pesos_i(8234) := b"0000000000000000_0000000000000000_0000100101001111_0000000111010000"; -- 0.036361802458645155
	pesos_i(8235) := b"1111111111111111_1111111111111111_1111010101010000_1100110111011110"; -- -0.04173577632986293
	pesos_i(8236) := b"1111111111111111_1111111111111111_1110001000010101_0011110101001110"; -- -0.1168634112903996
	pesos_i(8237) := b"0000000000000000_0000000000000000_0001100011100010_0011101111110101"; -- 0.09720206008816071
	pesos_i(8238) := b"0000000000000000_0000000000000000_0010010001100010_1101100000011101"; -- 0.14213324277858208
	pesos_i(8239) := b"1111111111111111_1111111111111111_1111100001110100_0111000000110001"; -- -0.02947329341267432
	pesos_i(8240) := b"0000000000000000_0000000000000000_0001011101111110_0100101101000100"; -- 0.0917708436332593
	pesos_i(8241) := b"1111111111111111_1111111111111111_1101101001111011_1000000010011101"; -- -0.14655300291888285
	pesos_i(8242) := b"1111111111111111_1111111111111111_1110010101100011_1000010111100101"; -- -0.10395014908709048
	pesos_i(8243) := b"0000000000000000_0000000000000000_0001111010111100_0001110100110111"; -- 0.12005789359355021
	pesos_i(8244) := b"0000000000000000_0000000000000000_0001100001010001_1011000010110110"; -- 0.09499649470727232
	pesos_i(8245) := b"0000000000000000_0000000000000000_0010011111101010_0101100100010000"; -- 0.1559196152606022
	pesos_i(8246) := b"1111111111111111_1111111111111111_1110010011111111_1000001010011100"; -- -0.10547622378688225
	pesos_i(8247) := b"0000000000000000_0000000000000000_0000001110001000_1010001000011100"; -- 0.013803607848157725
	pesos_i(8248) := b"1111111111111111_1111111111111111_1110010111001110_1101111001100110"; -- -0.10231218339796304
	pesos_i(8249) := b"0000000000000000_0000000000000000_0010001000000011_1111101001101100"; -- 0.13287320259296528
	pesos_i(8250) := b"0000000000000000_0000000000000000_0000100101100000_1111101000100111"; -- 0.0366360041058222
	pesos_i(8251) := b"0000000000000000_0000000000000000_0000100110000110_0010010100110111"; -- 0.03720314590054272
	pesos_i(8252) := b"0000000000000000_0000000000000000_0001100001011100_1001110100111111"; -- 0.09516318111121913
	pesos_i(8253) := b"1111111111111111_1111111111111111_1110011110011000_1010011010111100"; -- -0.09532697581195686
	pesos_i(8254) := b"1111111111111111_1111111111111111_1111111010111100_1101000110100110"; -- -0.004931351591038474
	pesos_i(8255) := b"1111111111111111_1111111111111111_1111000111110111_0011011101110001"; -- -0.0548215245187525
	pesos_i(8256) := b"1111111111111111_1111111111111111_1111010111001011_1000000001011111"; -- -0.03986356425350784
	pesos_i(8257) := b"1111111111111111_1111111111111111_1110100110101100_1110100111110100"; -- -0.08720529347252254
	pesos_i(8258) := b"0000000000000000_0000000000000000_0001001011010010_1010010010101100"; -- 0.0735266608303439
	pesos_i(8259) := b"1111111111111111_1111111111111111_1111101100100000_1111100001110110"; -- -0.019028159231725364
	pesos_i(8260) := b"0000000000000000_0000000000000000_0000110011001101_0011101001010101"; -- 0.05000652859527654
	pesos_i(8261) := b"1111111111111111_1111111111111111_1111100010000011_1101110100100101"; -- -0.029237917417292817
	pesos_i(8262) := b"0000000000000000_0000000000000000_0000000111100011_1111000011000100"; -- 0.007384345770645302
	pesos_i(8263) := b"0000000000000000_0000000000000000_0000000110110001_0011111100101000"; -- 0.0066108201423229285
	pesos_i(8264) := b"0000000000000000_0000000000000000_0000000110111011_1100111011110101"; -- 0.006771979169541984
	pesos_i(8265) := b"0000000000000000_0000000000000000_0001000010110110_1111101011110111"; -- 0.0652920583661525
	pesos_i(8266) := b"1111111111111111_1111111111111111_1110010011101011_0110101111000101"; -- -0.1057827610320368
	pesos_i(8267) := b"1111111111111111_1111111111111111_1110010111111001_0011001001000010"; -- -0.10166631603296986
	pesos_i(8268) := b"0000000000000000_0000000000000000_0000101100111110_0111001100000110"; -- 0.0439216507753781
	pesos_i(8269) := b"0000000000000000_0000000000000000_0001111010000011_0000101101000110"; -- 0.11918707340759067
	pesos_i(8270) := b"1111111111111111_1111111111111111_1110101111100000_1000001111000000"; -- -0.07860542827519752
	pesos_i(8271) := b"0000000000000000_0000000000000000_0001010011100010_1011010010111111"; -- 0.08158425958747496
	pesos_i(8272) := b"1111111111111111_1111111111111111_1110011100101100_1111111000011110"; -- -0.0969697166412017
	pesos_i(8273) := b"1111111111111111_1111111111111111_1110000000010111_0111100011001001"; -- -0.12464184859954988
	pesos_i(8274) := b"0000000000000000_0000000000000000_0001000111000111_1111001100000000"; -- 0.06945723300971103
	pesos_i(8275) := b"1111111111111111_1111111111111111_1111111100100000_1101110100010000"; -- -0.0034047924089506245
	pesos_i(8276) := b"0000000000000000_0000000000000000_0000101011001101_1110111111110111"; -- 0.04220485469284001
	pesos_i(8277) := b"0000000000000000_0000000000000000_0001000011110011_0101100100011111"; -- 0.06621319777517659
	pesos_i(8278) := b"1111111111111111_1111111111111111_1111111101111000_1111100000101100"; -- -0.0020604031785076845
	pesos_i(8279) := b"1111111111111111_1111111111111111_1110011010111100_1111000100011011"; -- -0.09867947667777703
	pesos_i(8280) := b"1111111111111111_1111111111111111_1110101101111000_0101100111111100"; -- -0.08019483178415987
	pesos_i(8281) := b"0000000000000000_0000000000000000_0001011000101011_0100011111011101"; -- 0.08659791136453307
	pesos_i(8282) := b"1111111111111111_1111111111111111_1101100011100010_1010001011100111"; -- -0.1527918039328353
	pesos_i(8283) := b"1111111111111111_1111111111111111_1111011101001101_1100111001101100"; -- -0.033969019558543256
	pesos_i(8284) := b"0000000000000000_0000000000000000_0001101101000011_1111000101111001"; -- 0.10650548184109355
	pesos_i(8285) := b"0000000000000000_0000000000000000_0010001111010001_1101111001100011"; -- 0.13992109222895657
	pesos_i(8286) := b"0000000000000000_0000000000000000_0010001011000101_0100111010110100"; -- 0.13582317258274723
	pesos_i(8287) := b"1111111111111111_1111111111111111_1111000011111101_1110100000011001"; -- -0.05862569235012451
	pesos_i(8288) := b"0000000000000000_0000000000000000_0010001110010100_1100110101000101"; -- 0.1389892856927408
	pesos_i(8289) := b"1111111111111111_1111111111111111_1111100110100011_1101001001001001"; -- -0.024844033351648094
	pesos_i(8290) := b"0000000000000000_0000000000000000_0000010001001011_1111111100000000"; -- 0.01678460847080797
	pesos_i(8291) := b"1111111111111111_1111111111111111_1111110011110011_1101000100100111"; -- -0.011904647790654935
	pesos_i(8292) := b"0000000000000000_0000000000000000_0010010101001111_1000000110101000"; -- 0.14574442243555355
	pesos_i(8293) := b"1111111111111111_1111111111111111_1110000010101101_1001101011000100"; -- -0.12235100468833623
	pesos_i(8294) := b"0000000000000000_0000000000000000_0001111010000101_1010110001001000"; -- 0.11922718767055726
	pesos_i(8295) := b"0000000000000000_0000000000000000_0001101010101101_0110011101010001"; -- 0.10420842868497875
	pesos_i(8296) := b"1111111111111111_1111111111111111_1111011111110111_0001101100010011"; -- -0.03138571534610242
	pesos_i(8297) := b"0000000000000000_0000000000000000_0001000111111000_0100101100100010"; -- 0.07019490795435958
	pesos_i(8298) := b"1111111111111111_1111111111111111_1111010101010000_1011111011001001"; -- -0.04173667524796692
	pesos_i(8299) := b"1111111111111111_1111111111111111_1110100101100110_0010010000001011"; -- -0.08828520521637245
	pesos_i(8300) := b"0000000000000000_0000000000000000_0000110011000100_1111110110001001"; -- 0.049880834551833
	pesos_i(8301) := b"1111111111111111_1111111111111111_1111100010101100_1110011111110110"; -- -0.02861166244691519
	pesos_i(8302) := b"1111111111111111_1111111111111111_1111101011101110_0101111110111101"; -- -0.019800201822578353
	pesos_i(8303) := b"0000000000000000_0000000000000000_0000110011000101_0011110010101111"; -- 0.049884598582100745
	pesos_i(8304) := b"1111111111111111_1111111111111111_1110101000011011_1000110011001100"; -- -0.08551712046996318
	pesos_i(8305) := b"1111111111111111_1111111111111111_1110111000101010_0000100111100100"; -- -0.06967104136309754
	pesos_i(8306) := b"0000000000000000_0000000000000000_0010000100101100_1100101111100110"; -- 0.1295897901210293
	pesos_i(8307) := b"1111111111111111_1111111111111111_1110110100000101_1010010101110010"; -- -0.07413259469843185
	pesos_i(8308) := b"1111111111111111_1111111111111111_1111100101111111_1010111000110001"; -- -0.025395501084005026
	pesos_i(8309) := b"0000000000000000_0000000000000000_0001101110011010_1000011001100000"; -- 0.10782661284349834
	pesos_i(8310) := b"1111111111111111_1111111111111111_1111111001111000_0110000101100110"; -- -0.005975639887905712
	pesos_i(8311) := b"0000000000000000_0000000000000000_0010001100000001_0101011100001000"; -- 0.13673919619651762
	pesos_i(8312) := b"1111111111111111_1111111111111111_1110011110101001_1111101100101001"; -- -0.09506254426158052
	pesos_i(8313) := b"0000000000000000_0000000000000000_0001111011100111_1111000001100101"; -- 0.12072660899163508
	pesos_i(8314) := b"1111111111111111_1111111111111111_1110101110110101_1110011010100101"; -- -0.07925566175107697
	pesos_i(8315) := b"1111111111111111_1111111111111111_1111001001111000_0111011011001111"; -- -0.052849363657691696
	pesos_i(8316) := b"1111111111111111_1111111111111111_1111110010011110_1100000100010100"; -- -0.013202603075893257
	pesos_i(8317) := b"1111111111111111_1111111111111111_1110011101010001_0110000001110110"; -- -0.0964145384598498
	pesos_i(8318) := b"1111111111111111_1111111111111111_1111110110101001_1010000101101100"; -- -0.009130393264055302
	pesos_i(8319) := b"0000000000000000_0000000000000000_0000100101101100_0110000001011011"; -- 0.03680994251794174
	pesos_i(8320) := b"0000000000000000_0000000000000000_0001111101101110_0010100111011000"; -- 0.12277471088204274
	pesos_i(8321) := b"1111111111111111_1111111111111111_1110110000100100_1001100011111010"; -- -0.0775665654690196
	pesos_i(8322) := b"0000000000000000_0000000000000000_0000111000110010_0110011100000010"; -- 0.05545657923543012
	pesos_i(8323) := b"0000000000000000_0000000000000000_0000000010111001_1000100001110010"; -- 0.0028310088612955686
	pesos_i(8324) := b"0000000000000000_0000000000000000_0000010001111101_1001100001011001"; -- 0.017541429211651603
	pesos_i(8325) := b"1111111111111111_1111111111111111_1110011011001100_0011110001010011"; -- -0.09844611151412146
	pesos_i(8326) := b"0000000000000000_0000000000000000_0000011011100011_1101100111100011"; -- 0.026914232261197494
	pesos_i(8327) := b"0000000000000000_0000000000000000_0000101010101001_0001011000000000"; -- 0.04164254675584536
	pesos_i(8328) := b"1111111111111111_1111111111111111_1110000110001110_1110100110111100"; -- -0.11891307022029227
	pesos_i(8329) := b"1111111111111111_1111111111111111_1111010101000111_1000000110010110"; -- -0.041877651997416186
	pesos_i(8330) := b"1111111111111111_1111111111111111_1110010101011111_1011111000111001"; -- -0.10400782684752818
	pesos_i(8331) := b"0000000000000000_0000000000000000_0001010100110110_1100001110110111"; -- 0.08286689004620125
	pesos_i(8332) := b"1111111111111111_1111111111111111_1111001001101101_0100000001100000"; -- -0.053020454924095316
	pesos_i(8333) := b"0000000000000000_0000000000000000_0001001000111100_0001101011100110"; -- 0.07122963064115574
	pesos_i(8334) := b"0000000000000000_0000000000000000_0000101010100101_0100101001100000"; -- 0.041584633188886944
	pesos_i(8335) := b"1111111111111111_1111111111111111_1110100011100111_1011100011100111"; -- -0.09021419877766972
	pesos_i(8336) := b"1111111111111111_1111111111111111_1110101111110000_1110110111010101"; -- -0.07835496477823788
	pesos_i(8337) := b"0000000000000000_0000000000000000_0010100001100111_0101110011111001"; -- 0.15782719677559903
	pesos_i(8338) := b"1111111111111111_1111111111111111_1111000011011000_1100001011011111"; -- -0.05919248622538347
	pesos_i(8339) := b"0000000000000000_0000000000000000_0001110010011100_0010110010010100"; -- 0.11175802809147967
	pesos_i(8340) := b"1111111111111111_1111111111111111_1111001110110100_0001010011111111"; -- -0.04803341648556754
	pesos_i(8341) := b"0000000000000000_0000000000000000_0010010000110101_1100000100100111"; -- 0.14144522849399688
	pesos_i(8342) := b"1111111111111111_1111111111111111_1110101101011111_1111100111100001"; -- -0.08056677110346838
	pesos_i(8343) := b"0000000000000000_0000000000000000_0010011000011101_1110011110110111"; -- 0.1488938160600423
	pesos_i(8344) := b"0000000000000000_0000000000000000_0001101111011100_1100101100010110"; -- 0.10883778853230427
	pesos_i(8345) := b"1111111111111111_1111111111111111_1110100110100011_0000010000101000"; -- -0.08735631970915224
	pesos_i(8346) := b"1111111111111111_1111111111111111_1110101100111110_1100001100011001"; -- -0.0810735763404493
	pesos_i(8347) := b"1111111111111111_1111111111111111_1111011011100100_1010001101011100"; -- -0.035573759180516744
	pesos_i(8348) := b"1111111111111111_1111111111111111_1110010100100101_0100010001111010"; -- -0.10490009319854994
	pesos_i(8349) := b"1111111111111111_1111111111111111_1111111011011001_1100001111110111"; -- -0.004489662330896275
	pesos_i(8350) := b"0000000000000000_0000000000000000_0000010101001111_0100011011110010"; -- 0.020740923121879033
	pesos_i(8351) := b"1111111111111111_1111111111111111_1110010101101010_1011011011111101"; -- -0.10384041144941236
	pesos_i(8352) := b"0000000000000000_0000000000000000_0010000010100011_0101011110101111"; -- 0.1274924088998817
	pesos_i(8353) := b"1111111111111111_1111111111111111_1111001111111110_1100011000011111"; -- -0.046893708694510414
	pesos_i(8354) := b"1111111111111111_1111111111111111_1111110111100110_1010000011001101"; -- -0.00819964415125378
	pesos_i(8355) := b"0000000000000000_0000000000000000_0000000000111100_1011010011010001"; -- 0.0009263048930607501
	pesos_i(8356) := b"1111111111111111_1111111111111111_1111000000111011_1010000000110010"; -- -0.06159018312779002
	pesos_i(8357) := b"1111111111111111_1111111111111111_1111010100111100_0010111110111010"; -- -0.04205037799484161
	pesos_i(8358) := b"0000000000000000_0000000000000000_0001111010100111_0110100010011100"; -- 0.11974195286271809
	pesos_i(8359) := b"0000000000000000_0000000000000000_0010000100101001_1000111100000011"; -- 0.12954038455948022
	pesos_i(8360) := b"1111111111111111_1111111111111111_1101110100001010_1110011010001010"; -- -0.13655242084865318
	pesos_i(8361) := b"1111111111111111_1111111111111111_1110000111010011_1011110001000110"; -- -0.11786292347938211
	pesos_i(8362) := b"1111111111111111_1111111111111111_1101101010110011_0110101000001101"; -- -0.14569985567139362
	pesos_i(8363) := b"0000000000000000_0000000000000000_0001110111100111_1110011100100100"; -- 0.11681980733868853
	pesos_i(8364) := b"1111111111111111_1111111111111111_1111001101111001_0001011111100001"; -- -0.04893351313195528
	pesos_i(8365) := b"1111111111111111_1111111111111111_1110100100011101_1101000111111110"; -- -0.08938872855064588
	pesos_i(8366) := b"0000000000000000_0000000000000000_0010001101001101_1111110001100000"; -- 0.13790871955110318
	pesos_i(8367) := b"0000000000000000_0000000000000000_0000110011110111_1101000101110000"; -- 0.0506564043368216
	pesos_i(8368) := b"1111111111111111_1111111111111111_1101110000010001_1111000100111110"; -- -0.14035122137517717
	pesos_i(8369) := b"1111111111111111_1111111111111111_1101101101000010_0010101011110000"; -- -0.1435216105326099
	pesos_i(8370) := b"0000000000000000_0000000000000000_0000111001000110_0111001110011000"; -- 0.05576250506454992
	pesos_i(8371) := b"0000000000000000_0000000000000000_0000100100101010_0100001100111011"; -- 0.03580112643574835
	pesos_i(8372) := b"0000000000000000_0000000000000000_0001101111010111_0110001001110001"; -- 0.10875525726621756
	pesos_i(8373) := b"0000000000000000_0000000000000000_0000111101010101_1001111001111011"; -- 0.05990019325924791
	pesos_i(8374) := b"0000000000000000_0000000000000000_0000001011101110_1111101010000001"; -- 0.011459022887726284
	pesos_i(8375) := b"1111111111111111_1111111111111111_1101101000110111_0110011001110000"; -- -0.14759216082768814
	pesos_i(8376) := b"0000000000000000_0000000000000000_0001001001010011_0011000011100100"; -- 0.07158189367074137
	pesos_i(8377) := b"0000000000000000_0000000000000000_0001001101100111_0010101010010111"; -- 0.07579294373462203
	pesos_i(8378) := b"0000000000000000_0000000000000000_0001000010100010_1001011010000110"; -- 0.06498089562280197
	pesos_i(8379) := b"0000000000000000_0000000000000000_0000000011001010_1001101100110101"; -- 0.003091526385531366
	pesos_i(8380) := b"0000000000000000_0000000000000000_0001010101111110_0010011001011100"; -- 0.08395614386516281
	pesos_i(8381) := b"0000000000000000_0000000000000000_0000001101001111_0000011000010100"; -- 0.01292455662072418
	pesos_i(8382) := b"0000000000000000_0000000000000000_0000101101101001_0001010110010101"; -- 0.04457220916407375
	pesos_i(8383) := b"0000000000000000_0000000000000000_0000100111001110_0110100111001101"; -- 0.03830586669880379
	pesos_i(8384) := b"0000000000000000_0000000000000000_0010000100000110_0111011000001000"; -- 0.12900483803158083
	pesos_i(8385) := b"1111111111111111_1111111111111111_1101111011011011_0110100011110011"; -- -0.12946456974063647
	pesos_i(8386) := b"0000000000000000_0000000000000000_0000001110100010_0011111000010001"; -- 0.014194373364240669
	pesos_i(8387) := b"0000000000000000_0000000000000000_0001110100111011_0100001010100111"; -- 0.11418549127539825
	pesos_i(8388) := b"0000000000000000_0000000000000000_0000000010110111_1001110010100010"; -- 0.0028016944284445715
	pesos_i(8389) := b"0000000000000000_0000000000000000_0010000011111100_0101010111010000"; -- 0.12885032969496146
	pesos_i(8390) := b"0000000000000000_0000000000000000_0000111010010111_0011100000101101"; -- 0.05699492555557444
	pesos_i(8391) := b"0000000000000000_0000000000000000_0001110011000100_0000110111000001"; -- 0.11236654249588043
	pesos_i(8392) := b"0000000000000000_0000000000000000_0000000110101000_1000110101001011"; -- 0.006478148312772376
	pesos_i(8393) := b"0000000000000000_0000000000000000_0010000101110000_0101101101000000"; -- 0.13062067332004876
	pesos_i(8394) := b"0000000000000000_0000000000000000_0001000111110111_1111100011001010"; -- 0.07018999985385783
	pesos_i(8395) := b"1111111111111111_1111111111111111_1110011111001000_1000110111101101"; -- -0.09459603275663743
	pesos_i(8396) := b"1111111111111111_1111111111111111_1111010001111011_1101000101111110"; -- -0.04498568226985629
	pesos_i(8397) := b"0000000000000000_0000000000000000_0001110010000010_0010010110111101"; -- 0.11136089202965994
	pesos_i(8398) := b"0000000000000000_0000000000000000_0000100011110010_1111110111001110"; -- 0.03495775482576185
	pesos_i(8399) := b"0000000000000000_0000000000000000_0001010111001111_1001011100011100"; -- 0.08519882616157207
	pesos_i(8400) := b"0000000000000000_0000000000000000_0001101011001001_1011100110010011"; -- 0.10464057779928371
	pesos_i(8401) := b"0000000000000000_0000000000000000_0001100010100100_1101100101110010"; -- 0.09626540220575207
	pesos_i(8402) := b"1111111111111111_1111111111111111_1110111001000101_0011001010001010"; -- -0.06925663111694395
	pesos_i(8403) := b"1111111111111111_1111111111111111_1110110100111010_0101000100101001"; -- -0.07332890271918338
	pesos_i(8404) := b"0000000000000000_0000000000000000_0001101110110111_1100011001101101"; -- 0.10827293558530388
	pesos_i(8405) := b"1111111111111111_1111111111111111_1111011011011111_1111010001101111"; -- -0.0356452206488828
	pesos_i(8406) := b"1111111111111111_1111111111111111_1101101010110011_0000001000011110"; -- -0.1457060506354567
	pesos_i(8407) := b"1111111111111111_1111111111111111_1110110111111001_1011011000011011"; -- -0.07040845724593355
	pesos_i(8408) := b"0000000000000000_0000000000000000_0001101011110100_0111001100111001"; -- 0.10529251225489736
	pesos_i(8409) := b"0000000000000000_0000000000000000_0010000010011011_1111111100011111"; -- 0.12738031881418962
	pesos_i(8410) := b"0000000000000000_0000000000000000_0000001011001011_0010001010110011"; -- 0.010912102362115416
	pesos_i(8411) := b"1111111111111111_1111111111111111_1111010100110001_1100001110111000"; -- -0.04220940370229374
	pesos_i(8412) := b"0000000000000000_0000000000000000_0000100010100101_1111100101010011"; -- 0.033782561163793204
	pesos_i(8413) := b"0000000000000000_0000000000000000_0010001011010111_1100001010001101"; -- 0.13610473570225365
	pesos_i(8414) := b"0000000000000000_0000000000000000_0000110011101101_1111001110100101"; -- 0.050505855404346295
	pesos_i(8415) := b"0000000000000000_0000000000000000_0001000101100110_1000001110100111"; -- 0.06797049360065892
	pesos_i(8416) := b"0000000000000000_0000000000000000_0000110011000011_1110010011100101"; -- 0.04986410693007883
	pesos_i(8417) := b"1111111111111111_1111111111111111_1111010101110100_0001101010110010"; -- -0.04119713929888877
	pesos_i(8418) := b"1111111111111111_1111111111111111_1110011101100100_1111110110010000"; -- -0.09611525760296183
	pesos_i(8419) := b"1111111111111111_1111111111111111_1111010111110010_1111111101001101"; -- -0.03926090596144971
	pesos_i(8420) := b"1111111111111111_1111111111111111_1101110110101100_1100011010000110"; -- -0.1340824053202323
	pesos_i(8421) := b"1111111111111111_1111111111111111_1110010010000011_0001001010110101"; -- -0.10737498355540011
	pesos_i(8422) := b"1111111111111111_1111111111111111_1111011111000001_1110110010101111"; -- -0.032197196163108066
	pesos_i(8423) := b"1111111111111111_1111111111111111_1111001000000101_1010111000011000"; -- -0.05460082915405293
	pesos_i(8424) := b"0000000000000000_0000000000000000_0000000001011101_0111000000111110"; -- 0.0014257574339791323
	pesos_i(8425) := b"1111111111111111_1111111111111111_1101100110011100_0001101010001100"; -- -0.1499617965657332
	pesos_i(8426) := b"0000000000000000_0000000000000000_0000110010000011_1010000110011110"; -- 0.0488835345549226
	pesos_i(8427) := b"0000000000000000_0000000000000000_0001111000110101_1010011011011010"; -- 0.11800616097456056
	pesos_i(8428) := b"1111111111111111_1111111111111111_1110110000111100_0010100001000111"; -- -0.07720707197863838
	pesos_i(8429) := b"0000000000000000_0000000000000000_0000100000000011_0111011001000001"; -- 0.03130282480705994
	pesos_i(8430) := b"1111111111111111_1111111111111111_1111110000111110_0110010110001110"; -- -0.01467290187305266
	pesos_i(8431) := b"1111111111111111_1111111111111111_1111110101000010_1101100011111010"; -- -0.010698737166002989
	pesos_i(8432) := b"1111111111111111_1111111111111111_1110101110110001_0100110100000111"; -- -0.07932585303947368
	pesos_i(8433) := b"1111111111111111_1111111111111111_1110110111000111_1010110011100011"; -- -0.07117194603507755
	pesos_i(8434) := b"0000000000000000_0000000000000000_0000001001111101_1010110100110101"; -- 0.009730172555782225
	pesos_i(8435) := b"0000000000000000_0000000000000000_0001111100011110_1110100101011010"; -- 0.12156542241885208
	pesos_i(8436) := b"1111111111111111_1111111111111111_1101111010101001_1010000110000100"; -- -0.13022413762211976
	pesos_i(8437) := b"1111111111111111_1111111111111111_1110000111011001_1011000100100001"; -- -0.11777203513905768
	pesos_i(8438) := b"1111111111111111_1111111111111111_1111100001001110_1010101101000110"; -- -0.030049605704877146
	pesos_i(8439) := b"1111111111111111_1111111111111111_1101101111000001_0111001101001110"; -- -0.1415794309785693
	pesos_i(8440) := b"0000000000000000_0000000000000000_0001110001010100_1010110010111101"; -- 0.11066703421049935
	pesos_i(8441) := b"1111111111111111_1111111111111111_1101111011111111_1011010100001011"; -- -0.12891071789109607
	pesos_i(8442) := b"1111111111111111_1111111111111111_1111011101000011_0001111010011101"; -- -0.0341320864349175
	pesos_i(8443) := b"0000000000000000_0000000000000000_0001011111001111_1011010001000000"; -- 0.09301306300754206
	pesos_i(8444) := b"0000000000000000_0000000000000000_0000111000011111_1010110100011010"; -- 0.05517084014732183
	pesos_i(8445) := b"0000000000000000_0000000000000000_0000110101001011_1100100011001110"; -- 0.05193762799818761
	pesos_i(8446) := b"1111111111111111_1111111111111111_1110100011101000_1011110100000111"; -- -0.09019869399655998
	pesos_i(8447) := b"0000000000000000_0000000000000000_0001110011110001_0111010011100011"; -- 0.11305933510847344
	pesos_i(8448) := b"1111111111111111_1111111111111111_1110000000110000_1011111010111101"; -- -0.12425620924832209
	pesos_i(8449) := b"0000000000000000_0000000000000000_0001101111101111_0010001110011011"; -- 0.10911772276211137
	pesos_i(8450) := b"0000000000000000_0000000000000000_0000110010001110_0100010101000011"; -- 0.0490458764460098
	pesos_i(8451) := b"1111111111111111_1111111111111111_1111011010110111_1110001010011001"; -- -0.03625663525129
	pesos_i(8452) := b"1111111111111111_1111111111111111_1111110001010011_1000001111011011"; -- -0.014350661359520296
	pesos_i(8453) := b"1111111111111111_1111111111111111_1101010001000101_1110101001001101"; -- -0.17080817818620642
	pesos_i(8454) := b"0000000000000000_0000000000000000_0000101001111000_1100100111111000"; -- 0.040905593047922684
	pesos_i(8455) := b"0000000000000000_0000000000000000_0000110011000001_1111110100010100"; -- 0.049835030911631495
	pesos_i(8456) := b"0000000000000000_0000000000000000_0001100001110100_0111111110011101"; -- 0.09552762594229766
	pesos_i(8457) := b"1111111111111111_1111111111111111_1110010010110001_1101010011000011"; -- -0.10666151275385992
	pesos_i(8458) := b"1111111111111111_1111111111111111_1111000110001110_1111011001100001"; -- -0.056412316709656476
	pesos_i(8459) := b"1111111111111111_1111111111111111_1110011100001111_0101011110111000"; -- -0.09742213970372048
	pesos_i(8460) := b"0000000000000000_0000000000000000_0001011101101101_0010011111001100"; -- 0.09150933011551374
	pesos_i(8461) := b"1111111111111111_1111111111111111_1101101001001010_0100110111000100"; -- -0.14730371447889334
	pesos_i(8462) := b"0000000000000000_0000000000000000_0010000111011001_1101101100010010"; -- 0.13223046477183428
	pesos_i(8463) := b"0000000000000000_0000000000000000_0000100011011110_0100100101001101"; -- 0.03464182012992944
	pesos_i(8464) := b"1111111111111111_1111111111111111_1111010011001011_0111101011000101"; -- -0.043770148078695836
	pesos_i(8465) := b"1111111111111111_1111111111111111_1110001011101011_0100000001110000"; -- -0.11359784381527481
	pesos_i(8466) := b"1111111111111111_1111111111111111_1110100110010000_0111111111000001"; -- -0.08763886962493493
	pesos_i(8467) := b"0000000000000000_0000000000000000_0010000010000100_0001001111000111"; -- 0.12701533899987033
	pesos_i(8468) := b"1111111111111111_1111111111111111_1111001110111111_1000100000101001"; -- -0.047858705514189456
	pesos_i(8469) := b"0000000000000000_0000000000000000_0001000110001111_0001111000001010"; -- 0.0685900472229935
	pesos_i(8470) := b"1111111111111111_1111111111111111_1111000001101001_0111101110011001"; -- -0.060890460068634966
	pesos_i(8471) := b"1111111111111111_1111111111111111_1111111010110000_1010100001011101"; -- -0.005116917903070071
	pesos_i(8472) := b"0000000000000000_0000000000000000_0001101011111001_0001101001010111"; -- 0.1053635084914108
	pesos_i(8473) := b"0000000000000000_0000000000000000_0010010110101011_1010110011000001"; -- 0.14715079985004534
	pesos_i(8474) := b"1111111111111111_1111111111111111_1110111100010100_1011011000001110"; -- -0.06609022296624485
	pesos_i(8475) := b"1111111111111111_1111111111111111_1110010111010110_0011001100111001"; -- -0.10220031603931372
	pesos_i(8476) := b"1111111111111111_1111111111111111_1111111101000100_0001011111110110"; -- -0.002867224262738009
	pesos_i(8477) := b"0000000000000000_0000000000000000_0010000111110000_1010000001000101"; -- 0.1325779121275649
	pesos_i(8478) := b"0000000000000000_0000000000000000_0001001111001100_1111011000011111"; -- 0.0773462129830875
	pesos_i(8479) := b"1111111111111111_1111111111111111_1111110110111111_0001101011001110"; -- -0.008802723579332332
	pesos_i(8480) := b"1111111111111111_1111111111111111_1111110111001000_0010101011011011"; -- -0.008664437790524237
	pesos_i(8481) := b"1111111111111111_1111111111111111_1110010011001001_1101001100000110"; -- -0.10629540533554378
	pesos_i(8482) := b"1111111111111111_1111111111111111_1111110000100000_0001110000011100"; -- -0.015135043251162718
	pesos_i(8483) := b"0000000000000000_0000000000000000_0000011111011101_1110010110001011"; -- 0.03072962412334534
	pesos_i(8484) := b"1111111111111111_1111111111111111_1101111111101000_0011100011110001"; -- -0.12536281697611215
	pesos_i(8485) := b"0000000000000000_0000000000000000_0010011000011000_1101000011010111"; -- 0.14881615879162566
	pesos_i(8486) := b"0000000000000000_0000000000000000_0001001010010011_1110110000000011"; -- 0.07256960927570152
	pesos_i(8487) := b"1111111111111111_1111111111111111_1110010110100011_0011010110110001"; -- -0.1029783670978952
	pesos_i(8488) := b"0000000000000000_0000000000000000_0010000110010001_0110101111110011"; -- 0.13112520873477507
	pesos_i(8489) := b"1111111111111111_1111111111111111_1111100111000010_1001101001100001"; -- -0.024374343159661832
	pesos_i(8490) := b"1111111111111111_1111111111111111_1111110100001010_0000011010101101"; -- -0.011565764245188946
	pesos_i(8491) := b"0000000000000000_0000000000000000_0001010011100010_0111111111010010"; -- 0.08158110505488503
	pesos_i(8492) := b"0000000000000000_0000000000000000_0001100011110011_1101001000001100"; -- 0.09747040540046117
	pesos_i(8493) := b"1111111111111111_1111111111111111_1110000100010010_1001100011110101"; -- -0.12080997487397818
	pesos_i(8494) := b"1111111111111111_1111111111111111_1110101010001000_0111111010000000"; -- -0.08385476462050538
	pesos_i(8495) := b"1111111111111111_1111111111111111_1111001101001101_1110110010100100"; -- -0.049592218296400245
	pesos_i(8496) := b"0000000000000000_0000000000000000_0001111110101100_0101101001011011"; -- 0.12372364739537868
	pesos_i(8497) := b"1111111111111111_1111111111111111_1111110011001101_0101001100100100"; -- -0.012491992743526923
	pesos_i(8498) := b"1111111111111111_1111111111111111_1111111100000100_1100111111010100"; -- -0.003832827391385922
	pesos_i(8499) := b"0000000000000000_0000000000000000_0000100100000111_1100100111100111"; -- 0.03527509575022446
	pesos_i(8500) := b"0000000000000000_0000000000000000_0010101001010001_0010111110110010"; -- 0.16530130477269714
	pesos_i(8501) := b"1111111111111111_1111111111111111_1110110101110011_1100010111111110"; -- -0.07245218797450194
	pesos_i(8502) := b"0000000000000000_0000000000000000_0000000010001100_1000100001010110"; -- 0.002144356746835467
	pesos_i(8503) := b"0000000000000000_0000000000000000_0000001100111110_1010001111111101"; -- 0.012674569378262763
	pesos_i(8504) := b"1111111111111111_1111111111111111_1101111011101100_1011100110110101"; -- -0.12920035686407572
	pesos_i(8505) := b"1111111111111111_1111111111111111_1101111110101110_1001101100101111"; -- -0.12624197110129118
	pesos_i(8506) := b"1111111111111111_1111111111111111_1110100101011101_1101000010110011"; -- -0.08841224313921224
	pesos_i(8507) := b"0000000000000000_0000000000000000_0000001101000011_1101100001110100"; -- 0.012753990374701048
	pesos_i(8508) := b"1111111111111111_1111111111111111_1101111010111100_0011011101110011"; -- -0.1299405425816284
	pesos_i(8509) := b"1111111111111111_1111111111111111_1111110101101100_1101000111011001"; -- -0.010058292858840226
	pesos_i(8510) := b"1111111111111111_1111111111111111_1111000110110010_1111011110010101"; -- -0.055862928539244135
	pesos_i(8511) := b"0000000000000000_0000000000000000_0000010001000110_1110000000110111"; -- 0.01670647940784631
	pesos_i(8512) := b"0000000000000000_0000000000000000_0001111110101101_0000001001001100"; -- 0.1237336573311115
	pesos_i(8513) := b"1111111111111111_1111111111111111_1110001110111101_1100110111101001"; -- -0.1103850656783234
	pesos_i(8514) := b"1111111111111111_1111111111111111_1111000001000101_1110011011001001"; -- -0.06143338763596575
	pesos_i(8515) := b"0000000000000000_0000000000000000_0001101101110111_1011110101000110"; -- 0.10729582751240983
	pesos_i(8516) := b"1111111111111111_1111111111111111_1111101010110100_0010010101001100"; -- -0.02068869492606318
	pesos_i(8517) := b"0000000000000000_0000000000000000_0000111111101111_1101100001101111"; -- 0.06225350108296182
	pesos_i(8518) := b"1111111111111111_1111111111111111_1111010110100010_1111000111011100"; -- -0.040482410308295906
	pesos_i(8519) := b"1111111111111111_1111111111111111_1110011110110111_1010100111010101"; -- -0.09485376871782919
	pesos_i(8520) := b"0000000000000000_0000000000000000_0000111000001001_1011111101011010"; -- 0.05483623461060075
	pesos_i(8521) := b"0000000000000000_0000000000000000_0010011000101000_0111011100000001"; -- 0.14905494477545833
	pesos_i(8522) := b"1111111111111111_1111111111111111_1111100001000011_1101001000010101"; -- -0.030215139357718683
	pesos_i(8523) := b"1111111111111111_1111111111111111_1111000101011000_0011101001101010"; -- -0.05724749481501308
	pesos_i(8524) := b"0000000000000000_0000000000000000_0000111110110010_1000100111001001"; -- 0.061318027160312975
	pesos_i(8525) := b"0000000000000000_0000000000000000_0010000010101010_1101101100010001"; -- 0.12760705160835997
	pesos_i(8526) := b"0000000000000000_0000000000000000_0000101011001110_1011000011111010"; -- 0.04221635909720834
	pesos_i(8527) := b"0000000000000000_0000000000000000_0010001001010110_0010000110110111"; -- 0.13412676550286565
	pesos_i(8528) := b"1111111111111111_1111111111111111_1110101110101011_1010110011011111"; -- -0.07941169316784423
	pesos_i(8529) := b"1111111111111111_1111111111111111_1110101001101101_1110101001100001"; -- -0.08426032191731445
	pesos_i(8530) := b"0000000000000000_0000000000000000_0000110110101110_0001000100101111"; -- 0.053437303511170056
	pesos_i(8531) := b"0000000000000000_0000000000000000_0010011101001101_0011100011101110"; -- 0.15352207000689783
	pesos_i(8532) := b"1111111111111111_1111111111111111_1110011100101110_1110101011001101"; -- -0.0969403504777242
	pesos_i(8533) := b"1111111111111111_1111111111111111_1110001001011100_1101100100110101"; -- -0.11577074478880288
	pesos_i(8534) := b"1111111111111111_1111111111111111_1101111000101011_0100010110010111"; -- -0.13215222429914042
	pesos_i(8535) := b"0000000000000000_0000000000000000_0000100111110110_1010001101110110"; -- 0.03891965519232001
	pesos_i(8536) := b"0000000000000000_0000000000000000_0001000110001001_0000000000111010"; -- 0.06849671756454467
	pesos_i(8537) := b"1111111111111111_1111111111111111_1111010100001011_1010010111011010"; -- -0.04279101786067191
	pesos_i(8538) := b"1111111111111111_1111111111111111_1111011110011011_0001100010011010"; -- -0.032789671286481206
	pesos_i(8539) := b"0000000000000000_0000000000000000_0010001001111110_0101110011110010"; -- 0.1347406474805127
	pesos_i(8540) := b"0000000000000000_0000000000000000_0000110101100010_1010000111000010"; -- 0.052286252857980414
	pesos_i(8541) := b"1111111111111111_1111111111111111_1101110000010110_1100011101011100"; -- -0.1402774239822258
	pesos_i(8542) := b"0000000000000000_0000000000000000_0000000001101100_1000100001101100"; -- 0.0016560806764865917
	pesos_i(8543) := b"1111111111111111_1111111111111111_1110101101110101_1011101011110100"; -- -0.08023482832362973
	pesos_i(8544) := b"0000000000000000_0000000000000000_0000110111100011_0000101000100111"; -- 0.05424560018590465
	pesos_i(8545) := b"0000000000000000_0000000000000000_0010001000100001_1001100000010111"; -- 0.13332510537922634
	pesos_i(8546) := b"1111111111111111_1111111111111111_1110001101100010_0001110100000000"; -- -0.11178416021537406
	pesos_i(8547) := b"0000000000000000_0000000000000000_0000100110001010_1011101101101010"; -- 0.037273133734824174
	pesos_i(8548) := b"1111111111111111_1111111111111111_1110000010011110_1101100011101111"; -- -0.12257618103301494
	pesos_i(8549) := b"1111111111111111_1111111111111111_1110000000111100_1010100111011100"; -- -0.12407434819547689
	pesos_i(8550) := b"1111111111111111_1111111111111111_1111010110000000_0110111010011000"; -- -0.04100903301075884
	pesos_i(8551) := b"0000000000000000_0000000000000000_0010001011110001_1001100101111100"; -- 0.13649901656091934
	pesos_i(8552) := b"1111111111111111_1111111111111111_1101110101110111_1110111001000011"; -- -0.1348887526867395
	pesos_i(8553) := b"1111111111111111_1111111111111111_1111110100101001_0110110010000101"; -- -0.011086671271755244
	pesos_i(8554) := b"1111111111111111_1111111111111111_1101100111001100_1011000111001100"; -- -0.1492203596242446
	pesos_i(8555) := b"1111111111111111_1111111111111111_1110001110001111_1111110111010111"; -- -0.11108411317763506
	pesos_i(8556) := b"0000000000000000_0000000000000000_0001110110101000_0011011100000100"; -- 0.11584800571312634
	pesos_i(8557) := b"1111111111111111_1111111111111111_1111011001101111_1101111001100000"; -- -0.037355519873205886
	pesos_i(8558) := b"1111111111111111_1111111111111111_1111001101101001_0111100101001010"; -- -0.04917184785573
	pesos_i(8559) := b"0000000000000000_0000000000000000_0010001011001000_0101101110001101"; -- 0.13586971465455394
	pesos_i(8560) := b"0000000000000000_0000000000000000_0000100111101110_0111101101111011"; -- 0.03879520180592854
	pesos_i(8561) := b"0000000000000000_0000000000000000_0010001111100101_1010011111010111"; -- 0.1402230168390255
	pesos_i(8562) := b"1111111111111111_1111111111111111_1110111001010010_0011110010101101"; -- -0.06905766271067415
	pesos_i(8563) := b"1111111111111111_1111111111111111_1110100110110100_0001110011000101"; -- -0.08709545305866495
	pesos_i(8564) := b"0000000000000000_0000000000000000_0001111100000000_1000111101101100"; -- 0.12110229851066386
	pesos_i(8565) := b"0000000000000000_0000000000000000_0001001010100101_1000000101101001"; -- 0.07283791372857652
	pesos_i(8566) := b"1111111111111111_1111111111111111_1111111110101111_0101100110000010"; -- -0.0012306269451816307
	pesos_i(8567) := b"0000000000000000_0000000000000000_0001011111101111_1010111010010111"; -- 0.09350100697348541
	pesos_i(8568) := b"1111111111111111_1111111111111111_1101101100111101_0001010101110100"; -- -0.143599185044922
	pesos_i(8569) := b"1111111111111111_1111111111111111_1101101100110110_1110111010111011"; -- -0.14369304595278506
	pesos_i(8570) := b"0000000000000000_0000000000000000_0000110111000100_1001100011000001"; -- 0.053781077382336805
	pesos_i(8571) := b"0000000000000000_0000000000000000_0001100110010001_1100011001111001"; -- 0.09988060431153312
	pesos_i(8572) := b"0000000000000000_0000000000000000_0001110110001100_1111001101111111"; -- 0.11543199385664824
	pesos_i(8573) := b"0000000000000000_0000000000000000_0010000101101000_1001110000110101"; -- 0.13050247462400477
	pesos_i(8574) := b"1111111111111111_1111111111111111_1111100001001100_0100111101001000"; -- -0.03008560647540961
	pesos_i(8575) := b"0000000000000000_0000000000000000_0000010101010010_0100110010010001"; -- 0.020787034374790746
	pesos_i(8576) := b"1111111111111111_1111111111111111_1111000001011011_0101000100101010"; -- -0.061106612390541895
	pesos_i(8577) := b"0000000000000000_0000000000000000_0001011011101110_1001101110100010"; -- 0.08957836831013201
	pesos_i(8578) := b"1111111111111111_1111111111111111_1111110101010100_0110000011010000"; -- -0.01043124119006301
	pesos_i(8579) := b"1111111111111111_1111111111111111_1110000011011100_0010001011111011"; -- -0.12164098136371154
	pesos_i(8580) := b"0000000000000000_0000000000000000_0001010110000011_1100101010101010"; -- 0.08404223119951036
	pesos_i(8581) := b"0000000000000000_0000000000000000_0010100111100111_0011010110100000"; -- 0.16368422657739554
	pesos_i(8582) := b"1111111111111111_1111111111111111_1110101011100110_0000000010101000"; -- -0.08242793941312829
	pesos_i(8583) := b"1111111111111111_1111111111111111_1111101010110010_0010011101101010"; -- -0.02071908632190406
	pesos_i(8584) := b"1111111111111111_1111111111111111_1111010111110101_1111100001111011"; -- -0.039215535994470516
	pesos_i(8585) := b"0000000000000000_0000000000000000_0010010000001001_0110000111010000"; -- 0.1407681592791672
	pesos_i(8586) := b"1111111111111111_1111111111111111_1101110110010111_0101110000101110"; -- -0.13440917858404913
	pesos_i(8587) := b"1111111111111111_1111111111111111_1110100011010010_1101110110110010"; -- -0.09053244019652279
	pesos_i(8588) := b"0000000000000000_0000000000000000_0000110111100011_1110010010011011"; -- 0.0542586210859839
	pesos_i(8589) := b"1111111111111111_1111111111111111_1110110101011010_0101010110011000"; -- -0.07284035726873062
	pesos_i(8590) := b"1111111111111111_1111111111111111_1110011101001001_1000000010000101"; -- -0.09653469809565636
	pesos_i(8591) := b"1111111111111111_1111111111111111_1101110110100110_1100100001100100"; -- -0.13417384675822108
	pesos_i(8592) := b"0000000000000000_0000000000000000_0000101010111010_1001110101100101"; -- 0.041910016146516196
	pesos_i(8593) := b"0000000000000000_0000000000000000_0010010011011000_1011000000010101"; -- 0.14393139376445913
	pesos_i(8594) := b"1111111111111111_1111111111111111_1111001101010100_0101100011000000"; -- -0.049494221716886874
	pesos_i(8595) := b"1111111111111111_1111111111111111_1110001000101100_1111101001011101"; -- -0.11650119045566666
	pesos_i(8596) := b"0000000000000000_0000000000000000_0001000000001110_1100110111011011"; -- 0.06272589293293311
	pesos_i(8597) := b"1111111111111111_1111111111111111_1110111110110100_1100010000111001"; -- -0.0636479722360679
	pesos_i(8598) := b"0000000000000000_0000000000000000_0001100010100101_0000000101110100"; -- 0.09626778675941085
	pesos_i(8599) := b"0000000000000000_0000000000000000_0000001001010010_0100010010110100"; -- 0.00906781561759587
	pesos_i(8600) := b"0000000000000000_0000000000000000_0001000001001101_0101000110110100"; -- 0.06367979670114203
	pesos_i(8601) := b"1111111111111111_1111111111111111_1111111000001111_1101011000111111"; -- -0.007570848059900142
	pesos_i(8602) := b"0000000000000000_0000000000000000_0001100101110001_1101111111011000"; -- 0.09939383529771285
	pesos_i(8603) := b"1111111111111111_1111111111111111_1110110111000010_0011010100011001"; -- -0.07125538013606662
	pesos_i(8604) := b"0000000000000000_0000000000000000_0000110110101011_0110010111010001"; -- 0.05339657163852768
	pesos_i(8605) := b"1111111111111111_1111111111111111_1110001011101001_1010001100011111"; -- -0.11362247941336213
	pesos_i(8606) := b"1111111111111111_1111111111111111_1101101101100011_1001011100101011"; -- -0.14301161948377006
	pesos_i(8607) := b"0000000000000000_0000000000000000_0000110110001100_0000101101111100"; -- 0.05291816500744302
	pesos_i(8608) := b"1111111111111111_1111111111111111_1110011001100110_0000001001011100"; -- -0.10000596293452707
	pesos_i(8609) := b"1111111111111111_1111111111111111_1101110010000000_0001001011010001"; -- -0.13867075333957754
	pesos_i(8610) := b"0000000000000000_0000000000000000_0010001000010011_1010100100100011"; -- 0.13311249827003033
	pesos_i(8611) := b"0000000000000000_0000000000000000_0001001011000011_0000011001001110"; -- 0.0732883396578623
	pesos_i(8612) := b"0000000000000000_0000000000000000_0010001001111110_0111110110111101"; -- 0.13474260203051053
	pesos_i(8613) := b"0000000000000000_0000000000000000_0001101010010011_0010000000010110"; -- 0.1038074544956567
	pesos_i(8614) := b"0000000000000000_0000000000000000_0010001100001100_1111101111001111"; -- 0.13691686442683892
	pesos_i(8615) := b"1111111111111111_1111111111111111_1101110101101111_1001101111000111"; -- -0.13501573933434036
	pesos_i(8616) := b"0000000000000000_0000000000000000_0001110111110011_1011010101110101"; -- 0.11699995149623722
	pesos_i(8617) := b"1111111111111111_1111111111111111_1110100010001100_0010110010010101"; -- -0.09161111226559487
	pesos_i(8618) := b"1111111111111111_1111111111111111_1111111110101111_1000111111110011"; -- -0.001227381848449655
	pesos_i(8619) := b"0000000000000000_0000000000000000_0001111100001000_0110101000101001"; -- 0.12122214785880722
	pesos_i(8620) := b"0000000000000000_0000000000000000_0010011011100000_0101000110101100"; -- 0.15186033675568375
	pesos_i(8621) := b"0000000000000000_0000000000000000_0010010011011010_0001101000000110"; -- 0.14395296716262557
	pesos_i(8622) := b"1111111111111111_1111111111111111_1110011001000110_0001001011010000"; -- -0.10049326336468563
	pesos_i(8623) := b"1111111111111111_1111111111111111_1110011111010001_0010111001001010"; -- -0.09446440410163838
	pesos_i(8624) := b"0000000000000000_0000000000000000_0010001101000011_1000011011101000"; -- 0.13774912998094493
	pesos_i(8625) := b"0000000000000000_0000000000000000_0010000100001010_1110011100001010"; -- 0.1290726087981393
	pesos_i(8626) := b"1111111111111111_1111111111111111_1110011011101011_1000101100000111"; -- -0.09796839782726137
	pesos_i(8627) := b"0000000000000000_0000000000000000_0000011011011000_1001011101111111"; -- 0.02674242821513941
	pesos_i(8628) := b"0000000000000000_0000000000000000_0000010101011011_1100011001110101"; -- 0.02093162884078623
	pesos_i(8629) := b"0000000000000000_0000000000000000_0001011011011000_1100111001111010"; -- 0.08924570529401575
	pesos_i(8630) := b"0000000000000000_0000000000000000_0001000100001111_0110001101100100"; -- 0.06664105597597009
	pesos_i(8631) := b"0000000000000000_0000000000000000_0000111110110101_0100010010011010"; -- 0.061359679716713425
	pesos_i(8632) := b"1111111111111111_1111111111111111_1110001010000111_1011011110100101"; -- -0.1151166174534143
	pesos_i(8633) := b"0000000000000000_0000000000000000_0001010010110011_0100101001010010"; -- 0.08086075300129855
	pesos_i(8634) := b"1111111111111111_1111111111111111_1110011110100001_1100101010100101"; -- -0.09518750631025287
	pesos_i(8635) := b"1111111111111111_1111111111111111_1111110010010110_1001010100010010"; -- -0.01332729637372804
	pesos_i(8636) := b"1111111111111111_1111111111111111_1101101011110010_0111001100001010"; -- -0.14473801621219437
	pesos_i(8637) := b"0000000000000000_0000000000000000_0000100001110101_0100000010111011"; -- 0.03303913659546165
	pesos_i(8638) := b"1111111111111111_1111111111111111_1101101011110011_0010000000001011"; -- -0.14472770424297227
	pesos_i(8639) := b"0000000000000000_0000000000000000_0010010001011011_1110000000101111"; -- 0.14202691211495225
	pesos_i(8640) := b"1111111111111111_1111111111111111_1111010100010100_1000000001111100"; -- -0.04265591597884014
	pesos_i(8641) := b"1111111111111111_1111111111111111_1111010010001101_1000101011111101"; -- -0.04471522637453727
	pesos_i(8642) := b"0000000000000000_0000000000000000_0001101001001010_1000000100000101"; -- 0.10269934057518268
	pesos_i(8643) := b"0000000000000000_0000000000000000_0001010101001011_0110011000111110"; -- 0.08318175338868972
	pesos_i(8644) := b"1111111111111111_1111111111111111_1111111000111010_1011101000100000"; -- -0.006916396301240446
	pesos_i(8645) := b"1111111111111111_1111111111111111_1110000111001010_1000100100001010"; -- -0.11800330638863855
	pesos_i(8646) := b"1111111111111111_1111111111111111_1110100010100010_1100001010101001"; -- -0.09126647356113965
	pesos_i(8647) := b"1111111111111111_1111111111111111_1111100011100111_1000101011011111"; -- -0.02771694239055694
	pesos_i(8648) := b"0000000000000000_0000000000000000_0010010001010000_0110011100101011"; -- 0.14185185236719133
	pesos_i(8649) := b"1111111111111111_1111111111111111_1110111111000011_0001000100000111"; -- -0.06342977115634625
	pesos_i(8650) := b"1111111111111111_1111111111111111_1111001000110111_1110101110110001"; -- -0.053834218242295825
	pesos_i(8651) := b"0000000000000000_0000000000000000_0000111111101111_1100101000011100"; -- 0.06225264720929114
	pesos_i(8652) := b"0000000000000000_0000000000000000_0001001000011010_0100001011001011"; -- 0.07071320976112266
	pesos_i(8653) := b"0000000000000000_0000000000000000_0000111010011011_0111000110010110"; -- 0.05705938260184316
	pesos_i(8654) := b"1111111111111111_1111111111111111_1111011110111100_1110111010010101"; -- -0.03227337711726756
	pesos_i(8655) := b"0000000000000000_0000000000000000_0000110100101110_0101000000000001"; -- 0.05148792292854542
	pesos_i(8656) := b"0000000000000000_0000000000000000_0000001110101000_1000111110111100"; -- 0.01429079386952332
	pesos_i(8657) := b"1111111111111111_1111111111111111_1111010001000001_0010100110100110"; -- -0.045880696163782334
	pesos_i(8658) := b"1111111111111111_1111111111111111_1111010100011111_0000101111000111"; -- -0.0424950255824738
	pesos_i(8659) := b"1111111111111111_1111111111111111_1110110000010000_0110000001010011"; -- -0.07787511805600818
	pesos_i(8660) := b"1111111111111111_1111111111111111_1110010100100111_0111011101111101"; -- -0.10486653524342103
	pesos_i(8661) := b"1111111111111111_1111111111111111_1101110101111001_0100100101100000"; -- -0.13486806306421567
	pesos_i(8662) := b"1111111111111111_1111111111111111_1110011111110001_1100110000001111"; -- -0.09396671896202062
	pesos_i(8663) := b"1111111111111111_1111111111111111_1111001011111010_1000110110010011"; -- -0.0508643641386832
	pesos_i(8664) := b"0000000000000000_0000000000000000_0000100101010010_0000010010101000"; -- 0.036407748313482445
	pesos_i(8665) := b"1111111111111111_1111111111111111_1110111001010000_1111010100001101"; -- -0.06907719071862568
	pesos_i(8666) := b"1111111111111111_1111111111111111_1110010000001111_1101000110101001"; -- -0.1091336213700332
	pesos_i(8667) := b"0000000000000000_0000000000000000_0001101111101011_1000010000011000"; -- 0.10906243871935004
	pesos_i(8668) := b"0000000000000000_0000000000000000_0001110100100101_1010011101100001"; -- 0.11385580177406901
	pesos_i(8669) := b"0000000000000000_0000000000000000_0000100111111011_1111111100010010"; -- 0.03900140931959068
	pesos_i(8670) := b"1111111111111111_1111111111111111_1111110010001101_0100000110001100"; -- -0.013469603850514279
	pesos_i(8671) := b"1111111111111111_1111111111111111_1111101001110111_1010000100111101"; -- -0.021612093647316845
	pesos_i(8672) := b"0000000000000000_0000000000000000_0000001010110010_0111000111101111"; -- 0.010535355461165873
	pesos_i(8673) := b"0000000000000000_0000000000000000_0010001011001100_0000011011010111"; -- 0.13592570069904952
	pesos_i(8674) := b"0000000000000000_0000000000000000_0000001101111011_1001101110011111"; -- 0.013604856876608602
	pesos_i(8675) := b"0000000000000000_0000000000000000_0000110000101100_0111011000000100"; -- 0.04755342098534913
	pesos_i(8676) := b"1111111111111111_1111111111111111_1111001110111100_1110111011010001"; -- -0.04789836311202828
	pesos_i(8677) := b"1111111111111111_1111111111111111_1110010001100101_1100111010010001"; -- -0.1078215500881344
	pesos_i(8678) := b"0000000000000000_0000000000000000_0000001101010110_0010101001010000"; -- 0.013033527912459904
	pesos_i(8679) := b"1111111111111111_1111111111111111_1111010110000110_1011000101111100"; -- -0.04091349337982289
	pesos_i(8680) := b"0000000000000000_0000000000000000_0000000000011111_1100000101100111"; -- 0.0004845502317881193
	pesos_i(8681) := b"1111111111111111_1111111111111111_1110100010001111_0110001111101101"; -- -0.09156203716394959
	pesos_i(8682) := b"1111111111111111_1111111111111111_1111001101001000_0110000000110000"; -- -0.04967688387700191
	pesos_i(8683) := b"1111111111111111_1111111111111111_1110000100111000_0010110010100000"; -- -0.1202365979898906
	pesos_i(8684) := b"1111111111111111_1111111111111111_1111101001001001_0110101100110100"; -- -0.022317218484125968
	pesos_i(8685) := b"1111111111111111_1111111111111111_1101100111100110_0010111111010010"; -- -0.14883137827743115
	pesos_i(8686) := b"0000000000000000_0000000000000000_0001111010011100_0101100111111011"; -- 0.11957323443769077
	pesos_i(8687) := b"1111111111111111_1111111111111111_1111111010010100_0011011010101001"; -- -0.005550941225481328
	pesos_i(8688) := b"1111111111111111_1111111111111111_1111111100000110_0000010001110101"; -- -0.0038144315250685772
	pesos_i(8689) := b"1111111111111111_1111111111111111_1101111001000000_1100100010011010"; -- -0.13182398069655896
	pesos_i(8690) := b"0000000000000000_0000000000000000_0001000001000110_0100110101000110"; -- 0.06357272113016459
	pesos_i(8691) := b"0000000000000000_0000000000000000_0000000010110000_1000011011110010"; -- 0.0026935902107454984
	pesos_i(8692) := b"0000000000000000_0000000000000000_0000010010000111_0100101010001101"; -- 0.017689380124496078
	pesos_i(8693) := b"0000000000000000_0000000000000000_0000010001000010_1010110110100010"; -- 0.016642429350042995
	pesos_i(8694) := b"0000000000000000_0000000000000000_0001000010100000_0000111111011110"; -- 0.06494235207257315
	pesos_i(8695) := b"0000000000000000_0000000000000000_0001011011001010_0100101110111011"; -- 0.08902428932471573
	pesos_i(8696) := b"1111111111111111_1111111111111111_1111101001101110_0111110110000100"; -- -0.02175155180101908
	pesos_i(8697) := b"0000000000000000_0000000000000000_0001111011110010_0010100111111011"; -- 0.12088262910984125
	pesos_i(8698) := b"0000000000000000_0000000000000000_0001000000010011_0010101111010111"; -- 0.06279253015622475
	pesos_i(8699) := b"1111111111111111_1111111111111111_1101111010100101_0001011100100101"; -- -0.13029342016909867
	pesos_i(8700) := b"0000000000000000_0000000000000000_0001100001011011_1011011010001010"; -- 0.0951494298849997
	pesos_i(8701) := b"0000000000000000_0000000000000000_0000011101011100_0110001100100111"; -- 0.028753468558145888
	pesos_i(8702) := b"0000000000000000_0000000000000000_0000111110101100_0011000100100000"; -- 0.06122118982216386
	pesos_i(8703) := b"0000000000000000_0000000000000000_0001101111101000_0100110011110100"; -- 0.10901337587250026
	pesos_i(8704) := b"1111111111111111_1111111111111111_1110110110010110_1110000000011111"; -- -0.07191657291235229
	pesos_i(8705) := b"1111111111111111_1111111111111111_1111010010100101_0000010010000101"; -- -0.04435703046620962
	pesos_i(8706) := b"0000000000000000_0000000000000000_0001111101111010_1000100011010011"; -- 0.12296347752460957
	pesos_i(8707) := b"0000000000000000_0000000000000000_0000001000101101_1110000001111101"; -- 0.008512525998435815
	pesos_i(8708) := b"0000000000000000_0000000000000000_0001111010001101_0000011000101100"; -- 0.11933935716347982
	pesos_i(8709) := b"1111111111111111_1111111111111111_1101010000011111_1011011111001111"; -- -0.17139102169678422
	pesos_i(8710) := b"1111111111111111_1111111111111111_1110011111101000_1110101011101000"; -- -0.09410220936966153
	pesos_i(8711) := b"0000000000000000_0000000000000000_0010000001010100_1101100000001000"; -- 0.12629461476847345
	pesos_i(8712) := b"0000000000000000_0000000000000000_0000111100100011_1111000101000110"; -- 0.059142188596634206
	pesos_i(8713) := b"1111111111111111_1111111111111111_1110010110110111_0011010111011111"; -- -0.10267318061452936
	pesos_i(8714) := b"1111111111111111_1111111111111111_1111101100110110_1111011010011011"; -- -0.01869257647863514
	pesos_i(8715) := b"1111111111111111_1111111111111111_1111110100111010_0010010001000000"; -- -0.010831579519441059
	pesos_i(8716) := b"0000000000000000_0000000000000000_0000001001000001_1110100001101011"; -- 0.008818174371683274
	pesos_i(8717) := b"1111111111111111_1111111111111111_1111110110101110_0001000000100111"; -- -0.009062757983107779
	pesos_i(8718) := b"1111111111111111_1111111111111111_1111110101011010_0110101001000001"; -- -0.010339125828049932
	pesos_i(8719) := b"1111111111111111_1111111111111111_1101110101111001_1001100010111100"; -- -0.1348633327320418
	pesos_i(8720) := b"0000000000000000_0000000000000000_0000001110100011_0010110010001010"; -- 0.014208587403930363
	pesos_i(8721) := b"0000000000000000_0000000000000000_0000110101011100_0010110101010100"; -- 0.05218776026896114
	pesos_i(8722) := b"0000000000000000_0000000000000000_0001111000001111_1000111101100001"; -- 0.11742492788407491
	pesos_i(8723) := b"1111111111111111_1111111111111111_1101101010100100_1010011100001110"; -- -0.14592510145011808
	pesos_i(8724) := b"1111111111111111_1111111111111111_1111100000110100_1000111011010111"; -- -0.030448028977114534
	pesos_i(8725) := b"0000000000000000_0000000000000000_0010010111000111_1000001110001111"; -- 0.14757559063960993
	pesos_i(8726) := b"1111111111111111_1111111111111111_1110001100001101_0101010000000010"; -- -0.11307787848523525
	pesos_i(8727) := b"1111111111111111_1111111111111111_1111100000010110_1111101111111001"; -- -0.030899287976028696
	pesos_i(8728) := b"1111111111111111_1111111111111111_1111000011011011_0000100100100101"; -- -0.059157780240774366
	pesos_i(8729) := b"0000000000000000_0000000000000000_0001111001010111_0101001111001001"; -- 0.11852000867973492
	pesos_i(8730) := b"1111111111111111_1111111111111111_1101100100101100_0011101101010111"; -- -0.15166882646159321
	pesos_i(8731) := b"1111111111111111_1111111111111111_1110001110101001_0000101011001010"; -- -0.11070187163521868
	pesos_i(8732) := b"0000000000000000_0000000000000000_0001010100010111_1001011001000000"; -- 0.08239115780688132
	pesos_i(8733) := b"0000000000000000_0000000000000000_0010011000011011_1100100000001010"; -- 0.148861410599684
	pesos_i(8734) := b"1111111111111111_1111111111111111_1110001111110010_1111110011010111"; -- -0.10957355264648183
	pesos_i(8735) := b"0000000000000000_0000000000000000_0001100000011001_1100110100111100"; -- 0.09414370254431428
	pesos_i(8736) := b"1111111111111111_1111111111111111_1111010000010111_0100110000010111"; -- -0.04651951264606363
	pesos_i(8737) := b"1111111111111111_1111111111111111_1110111000110000_1010001001001110"; -- -0.0695704040287178
	pesos_i(8738) := b"0000000000000000_0000000000000000_0001101011001000_1001111000110010"; -- 0.1046236868778044
	pesos_i(8739) := b"0000000000000000_0000000000000000_0001011101001011_0100011101010001"; -- 0.09099240986147354
	pesos_i(8740) := b"0000000000000000_0000000000000000_0001000001101101_0100010000111101"; -- 0.064167275397137
	pesos_i(8741) := b"1111111111111111_1111111111111111_1101111110010011_1001100001111101"; -- -0.1266541188845979
	pesos_i(8742) := b"1111111111111111_1111111111111111_1110110001001101_1000001011110001"; -- -0.07694226859559217
	pesos_i(8743) := b"0000000000000000_0000000000000000_0001010000011101_0000011001010011"; -- 0.07856788187182454
	pesos_i(8744) := b"0000000000000000_0000000000000000_0001101000111000_0100010001110111"; -- 0.10242107311336723
	pesos_i(8745) := b"1111111111111111_1111111111111111_1101110101010011_1011011110001101"; -- -0.13544133012228132
	pesos_i(8746) := b"0000000000000000_0000000000000000_0000011110000001_0000011110101111"; -- 0.029312591747119095
	pesos_i(8747) := b"1111111111111111_1111111111111111_1110010011010111_1100011010000000"; -- -0.10608252879515612
	pesos_i(8748) := b"1111111111111111_1111111111111111_1110000000111001_0011001110011011"; -- -0.12412717299023784
	pesos_i(8749) := b"1111111111111111_1111111111111111_1110101101101011_1110100001100110"; -- -0.08038470749212319
	pesos_i(8750) := b"0000000000000000_0000000000000000_0000011100000000_0100011101110000"; -- 0.02734800809608863
	pesos_i(8751) := b"0000000000000000_0000000000000000_0001011111001101_1011011010111000"; -- 0.09298269256052945
	pesos_i(8752) := b"1111111111111111_1111111111111111_1110100111011000_1011010010001111"; -- -0.08653708943690369
	pesos_i(8753) := b"0000000000000000_0000000000000000_0000001010000100_0111111000010101"; -- 0.009834175149941716
	pesos_i(8754) := b"0000000000000000_0000000000000000_0000111001001000_0011100000101101"; -- 0.055789481047589365
	pesos_i(8755) := b"0000000000000000_0000000000000000_0001111110010010_1100111100000010"; -- 0.12333387176040599
	pesos_i(8756) := b"1111111111111111_1111111111111111_1110010111001001_1101001011100111"; -- -0.1023891626536638
	pesos_i(8757) := b"0000000000000000_0000000000000000_0001010001011110_1010100101101011"; -- 0.07956942416001787
	pesos_i(8758) := b"0000000000000000_0000000000000000_0001110111110001_1001000000101110"; -- 0.11696721197278787
	pesos_i(8759) := b"1111111111111111_1111111111111111_1110000010011011_0000001100000100"; -- -0.12263470794388025
	pesos_i(8760) := b"1111111111111111_1111111111111111_1111100111100100_1111111101110001"; -- -0.023849520707147926
	pesos_i(8761) := b"0000000000000000_0000000000000000_0000100110001001_0001110000001100"; -- 0.037248375709981615
	pesos_i(8762) := b"1111111111111111_1111111111111111_1101101010000011_1001011110010101"; -- -0.1464295637090331
	pesos_i(8763) := b"1111111111111111_1111111111111111_1110111010001010_1000001111001001"; -- -0.06819893212231219
	pesos_i(8764) := b"0000000000000000_0000000000000000_0001100110100110_0111000001011000"; -- 0.10019590509379807
	pesos_i(8765) := b"1111111111111111_1111111111111111_1111011111010000_0111000100111101"; -- -0.03197567233755463
	pesos_i(8766) := b"1111111111111111_1111111111111111_1110101100100101_1110111101100011"; -- -0.08145240626109729
	pesos_i(8767) := b"0000000000000000_0000000000000000_0001010010111001_0001100111001001"; -- 0.08094941289269007
	pesos_i(8768) := b"0000000000000000_0000000000000000_0000101011100010_0010101111110010"; -- 0.04251360572223939
	pesos_i(8769) := b"0000000000000000_0000000000000000_0001001001011001_0000111011010001"; -- 0.07167141528750556
	pesos_i(8770) := b"1111111111111111_1111111111111111_1111010110110011_0010111101110000"; -- -0.04023459927454664
	pesos_i(8771) := b"1111111111111111_1111111111111111_1110110010111001_0100000100000010"; -- -0.07529824920995459
	pesos_i(8772) := b"0000000000000000_0000000000000000_0000001100101001_1001001101010100"; -- 0.012353141776341623
	pesos_i(8773) := b"0000000000000000_0000000000000000_0001100000110001_1101000101011011"; -- 0.0945101592627283
	pesos_i(8774) := b"1111111111111111_1111111111111111_1111111101100110_0101011001011011"; -- -0.002344706281034814
	pesos_i(8775) := b"0000000000000000_0000000000000000_0000111111011101_0101001101111100"; -- 0.061970918436696235
	pesos_i(8776) := b"0000000000000000_0000000000000000_0000101101001100_1001010101111110"; -- 0.04413732844059388
	pesos_i(8777) := b"0000000000000000_0000000000000000_0000000100101010_0011111101010111"; -- 0.004550894383597123
	pesos_i(8778) := b"0000000000000000_0000000000000000_0010011010100101_0001111001111011"; -- 0.1509570169741546
	pesos_i(8779) := b"0000000000000000_0000000000000000_0000101011111111_1010101111110110"; -- 0.042963740783661164
	pesos_i(8780) := b"0000000000000000_0000000000000000_0000111111011101_1011110101011001"; -- 0.061977228361141085
	pesos_i(8781) := b"0000000000000000_0000000000000000_0000000011001111_0101000111110101"; -- 0.003163454411562675
	pesos_i(8782) := b"1111111111111111_1111111111111111_1111111100101111_1010101101001111"; -- -0.0031788760910356436
	pesos_i(8783) := b"0000000000000000_0000000000000000_0000010000000110_1100110010000010"; -- 0.01572874234594076
	pesos_i(8784) := b"0000000000000000_0000000000000000_0001100000100101_0010010100111110"; -- 0.09431679497075343
	pesos_i(8785) := b"0000000000000000_0000000000000000_0001101101101001_0000111001101011"; -- 0.1070717822397927
	pesos_i(8786) := b"0000000000000000_0000000000000000_0000100011111111_1001111001000111"; -- 0.03515042516658382
	pesos_i(8787) := b"0000000000000000_0000000000000000_0001011111000001_1110100000010101"; -- 0.09280252955593071
	pesos_i(8788) := b"1111111111111111_1111111111111111_1110111111111000_1011010001011100"; -- -0.06261131997823526
	pesos_i(8789) := b"0000000000000000_0000000000000000_0001010100100001_0001100111100100"; -- 0.08253633315020759
	pesos_i(8790) := b"0000000000000000_0000000000000000_0000001100011101_0000100110000100"; -- 0.01216182204001044
	pesos_i(8791) := b"0000000000000000_0000000000000000_0001111110010000_0010101011111111"; -- 0.12329357845039128
	pesos_i(8792) := b"1111111111111111_1111111111111111_1110100011100010_1001001011111011"; -- -0.09029275299862664
	pesos_i(8793) := b"0000000000000000_0000000000000000_0010011110110111_0011101111101011"; -- 0.1551396797726496
	pesos_i(8794) := b"0000000000000000_0000000000000000_0000011011011101_1100001000111010"; -- 0.026821269222220917
	pesos_i(8795) := b"0000000000000000_0000000000000000_0000000110110000_1001011101111100"; -- 0.006600826053867503
	pesos_i(8796) := b"1111111111111111_1111111111111111_1110010000100101_1010011101000001"; -- -0.10880045580929024
	pesos_i(8797) := b"0000000000000000_0000000000000000_0000001101011110_1111001011100001"; -- 0.013167552800744017
	pesos_i(8798) := b"0000000000000000_0000000000000000_0000110111010010_1110010101001011"; -- 0.05399926262885781
	pesos_i(8799) := b"1111111111111111_1111111111111111_1110100011000100_1100011000011010"; -- -0.09074746946763634
	pesos_i(8800) := b"1111111111111111_1111111111111111_1110110010011011_0110011110100100"; -- -0.07575371021819519
	pesos_i(8801) := b"1111111111111111_1111111111111111_1111101001101110_1000110001001000"; -- -0.021750671726109387
	pesos_i(8802) := b"0000000000000000_0000000000000000_0001001110000101_0101111010110100"; -- 0.07625381378744873
	pesos_i(8803) := b"0000000000000000_0000000000000000_0010000100100001_1010101010101011"; -- 0.12941996272382017
	pesos_i(8804) := b"1111111111111111_1111111111111111_1111000111100110_0111011111110000"; -- -0.05507707966166151
	pesos_i(8805) := b"0000000000000000_0000000000000000_0001011110101010_1001010110111010"; -- 0.092446668496166
	pesos_i(8806) := b"0000000000000000_0000000000000000_0010001001001010_1001101010011110"; -- 0.13395086639236903
	pesos_i(8807) := b"1111111111111111_1111111111111111_1111000101010010_1001001111001001"; -- -0.05733372073006398
	pesos_i(8808) := b"1111111111111111_1111111111111111_1111010111001110_1110010010001111"; -- -0.0398118163953668
	pesos_i(8809) := b"1111111111111111_1111111111111111_1110101111110011_1001011111110011"; -- -0.07831430729454694
	pesos_i(8810) := b"1111111111111111_1111111111111111_1110011001000110_0110011000111000"; -- -0.10048829215342536
	pesos_i(8811) := b"0000000000000000_0000000000000000_0001010010100110_0000001110110011"; -- 0.08065817953626843
	pesos_i(8812) := b"1111111111111111_1111111111111111_1110011010101100_1001011101000000"; -- -0.09892897297343009
	pesos_i(8813) := b"1111111111111111_1111111111111111_1110000000001000_1011110101101010"; -- -0.12486663973780233
	pesos_i(8814) := b"1111111111111111_1111111111111111_1111000011000110_0000010101000110"; -- -0.05947844550527547
	pesos_i(8815) := b"1111111111111111_1111111111111111_1110011010100110_0110101111001101"; -- -0.0990231155142524
	pesos_i(8816) := b"0000000000000000_0000000000000000_0000100011100111_0000000110110111"; -- 0.034774882510444076
	pesos_i(8817) := b"1111111111111111_1111111111111111_1110101000010010_1001011101101001"; -- -0.08565381699956566
	pesos_i(8818) := b"0000000000000000_0000000000000000_0001111000110010_1011101000000110"; -- 0.11796152735648624
	pesos_i(8819) := b"1111111111111111_1111111111111111_1101100111100010_1011011011110100"; -- -0.148884358791678
	pesos_i(8820) := b"1111111111111111_1111111111111111_1110000011100001_0101001010110101"; -- -0.12156184283983949
	pesos_i(8821) := b"1111111111111111_1111111111111111_1101110110000011_0011001000101101"; -- -0.13471685798766586
	pesos_i(8822) := b"0000000000000000_0000000000000000_0000100100000011_0001110111000001"; -- 0.03520379972885446
	pesos_i(8823) := b"1111111111111111_1111111111111111_1110111001110101_0101110101110100"; -- -0.06852165145757176
	pesos_i(8824) := b"1111111111111111_1111111111111111_1110000110011000_0110010011000101"; -- -0.11876840762401504
	pesos_i(8825) := b"0000000000000000_0000000000000000_0010001100001100_0101010000001101"; -- 0.1369068652897772
	pesos_i(8826) := b"0000000000000000_0000000000000000_0010000001101000_0001011011110100"; -- 0.12658828227927355
	pesos_i(8827) := b"1111111111111111_1111111111111111_1110101110001111_0110001011110110"; -- -0.07984334460784763
	pesos_i(8828) := b"1111111111111111_1111111111111111_1110000010111010_1011011001011100"; -- -0.1221509957288362
	pesos_i(8829) := b"0000000000000000_0000000000000000_0001000101011000_1011011110001010"; -- 0.06775996323054502
	pesos_i(8830) := b"0000000000000000_0000000000000000_0010000111010010_0100111100111111"; -- 0.13211531922452494
	pesos_i(8831) := b"1111111111111111_1111111111111111_1110101011101101_0011001000111111"; -- -0.08231817216787451
	pesos_i(8832) := b"1111111111111111_1111111111111111_1111100111100111_1001110101010110"; -- -0.02380959166226377
	pesos_i(8833) := b"1111111111111111_1111111111111111_1110000001111000_0000011101010111"; -- -0.1231685077511884
	pesos_i(8834) := b"0000000000000000_0000000000000000_0001110000100100_0100100010111110"; -- 0.10992865208026395
	pesos_i(8835) := b"1111111111111111_1111111111111111_1111101001101100_1010011001001010"; -- -0.021779639098787273
	pesos_i(8836) := b"1111111111111111_1111111111111111_1101100010011001_1000101101111010"; -- -0.15390709181500395
	pesos_i(8837) := b"0000000000000000_0000000000000000_0000100000111001_0100011001101101"; -- 0.03212394861423274
	pesos_i(8838) := b"0000000000000000_0000000000000000_0001111111111000_0100100011010110"; -- 0.12488227110018578
	pesos_i(8839) := b"1111111111111111_1111111111111111_1101111000100001_0000110000100000"; -- -0.13230823718702414
	pesos_i(8840) := b"1111111111111111_1111111111111111_1101101111101011_1100001001111000"; -- -0.14093384337189258
	pesos_i(8841) := b"1111111111111111_1111111111111111_1101111001011010_0110010011001001"; -- -0.13143320179582194
	pesos_i(8842) := b"1111111111111111_1111111111111111_1110111011001001_0001100101011001"; -- -0.06724397261556835
	pesos_i(8843) := b"1111111111111111_1111111111111111_1111101000100001_1100111011011110"; -- -0.022921629691214845
	pesos_i(8844) := b"0000000000000000_0000000000000000_0000110100010100_1010010001111010"; -- 0.05109622935022674
	pesos_i(8845) := b"1111111111111111_1111111111111111_1110100100100110_0110100110101101"; -- -0.08925761732550609
	pesos_i(8846) := b"1111111111111111_1111111111111111_1111100010010111_1110011100100110"; -- -0.02893214534551192
	pesos_i(8847) := b"0000000000000000_0000000000000000_0010011010000010_1101011110000101"; -- 0.15043398850855505
	pesos_i(8848) := b"1111111111111111_1111111111111111_1110001111011000_1101111001011010"; -- -0.10997209830239255
	pesos_i(8849) := b"0000000000000000_0000000000000000_0001101111111100_0000100101100110"; -- 0.10931452509200458
	pesos_i(8850) := b"0000000000000000_0000000000000000_0001010010110100_0011110001010000"; -- 0.08087517686884486
	pesos_i(8851) := b"1111111111111111_1111111111111111_1111110110000011_1101100011010101"; -- -0.009706924544426492
	pesos_i(8852) := b"1111111111111111_1111111111111111_1101100100111111_1110111110010110"; -- -0.1513681658759671
	pesos_i(8853) := b"0000000000000000_0000000000000000_0000100111111100_0101001101010010"; -- 0.03900643119998646
	pesos_i(8854) := b"0000000000000000_0000000000000000_0010001100111110_1000010100000001"; -- 0.13767272265170538
	pesos_i(8855) := b"1111111111111111_1111111111111111_1111011000100100_0110001010100011"; -- -0.03850730434960002
	pesos_i(8856) := b"0000000000000000_0000000000000000_0000001011101011_1011001001100000"; -- 0.01140894733829416
	pesos_i(8857) := b"1111111111111111_1111111111111111_1101110100110000_0001001011010111"; -- -0.1359852052246442
	pesos_i(8858) := b"0000000000000000_0000000000000000_0001100000010111_1001010111100011"; -- 0.094109886090683
	pesos_i(8859) := b"1111111111111111_1111111111111111_1110111110011100_1000100001111101"; -- -0.06401774349270024
	pesos_i(8860) := b"1111111111111111_1111111111111111_1110011010001100_0110000110111010"; -- -0.09942044453740281
	pesos_i(8861) := b"0000000000000000_0000000000000000_0001001101110010_0111100100110010"; -- 0.0759654757149098
	pesos_i(8862) := b"1111111111111111_1111111111111111_1110100101000000_1110101111111001"; -- -0.08885312237246042
	pesos_i(8863) := b"1111111111111111_1111111111111111_1111100111101011_0001100110111001"; -- -0.02375640141334422
	pesos_i(8864) := b"0000000000000000_0000000000000000_0010011001110001_0011011101011111"; -- 0.1501650436442905
	pesos_i(8865) := b"0000000000000000_0000000000000000_0010010001100101_1010101010011001"; -- 0.14217630600564926
	pesos_i(8866) := b"1111111111111111_1111111111111111_1111000010011011_1010100111111011"; -- -0.06012475596597169
	pesos_i(8867) := b"1111111111111111_1111111111111111_1110011111111110_1000001010111001"; -- -0.09377272590212375
	pesos_i(8868) := b"1111111111111111_1111111111111111_1110001101000110_1011011011010110"; -- -0.11220223684983695
	pesos_i(8869) := b"0000000000000000_0000000000000000_0010010111010111_0010101111110101"; -- 0.1478145095983788
	pesos_i(8870) := b"0000000000000000_0000000000000000_0000101010010010_1100001101101111"; -- 0.04130193188369976
	pesos_i(8871) := b"0000000000000000_0000000000000000_0000101100011101_0101010100111100"; -- 0.043416335254828485
	pesos_i(8872) := b"0000000000000000_0000000000000000_0000001101011110_1011111100011100"; -- 0.013164467069503498
	pesos_i(8873) := b"0000000000000000_0000000000000000_0000010101111101_1000010001011001"; -- 0.021446487245490708
	pesos_i(8874) := b"1111111111111111_1111111111111111_1111100011000100_0000100011000101"; -- -0.0282587546758106
	pesos_i(8875) := b"0000000000000000_0000000000000000_0001011001010011_1000101110110011"; -- 0.08721230622190677
	pesos_i(8876) := b"1111111111111111_1111111111111111_1101110111010100_0011000110111001"; -- -0.1334809229310841
	pesos_i(8877) := b"0000000000000000_0000000000000000_0001100000101000_0101001100111011"; -- 0.094365312564293
	pesos_i(8878) := b"0000000000000000_0000000000000000_0001111111111010_0001110111011101"; -- 0.1249102271462693
	pesos_i(8879) := b"0000000000000000_0000000000000000_0001110011111110_1000100110101010"; -- 0.11325893777492947
	pesos_i(8880) := b"0000000000000000_0000000000000000_0000110111110000_1101001001110010"; -- 0.05445590291778909
	pesos_i(8881) := b"1111111111111111_1111111111111111_1110011000101010_0100001100111011"; -- -0.10091762359785009
	pesos_i(8882) := b"1111111111111111_1111111111111111_1110010011000001_1001110010001111"; -- -0.10642072207987109
	pesos_i(8883) := b"0000000000000000_0000000000000000_0001110100111101_1001001110110001"; -- 0.11422083932182327
	pesos_i(8884) := b"1111111111111111_1111111111111111_1111111110100101_0011100111010100"; -- -0.001385103028105613
	pesos_i(8885) := b"1111111111111111_1111111111111111_1110001001111101_1101010111011010"; -- -0.11526740476217306
	pesos_i(8886) := b"0000000000000000_0000000000000000_0010010111100011_1100111101111100"; -- 0.14800736217511912
	pesos_i(8887) := b"1111111111111111_1111111111111111_1111000010101101_0000111000110111"; -- -0.05985938230087455
	pesos_i(8888) := b"1111111111111111_1111111111111111_1111100011111010_0001111111111000"; -- -0.02743339735053059
	pesos_i(8889) := b"1111111111111111_1111111111111111_1110100011000011_0110100011110101"; -- -0.09076828031443251
	pesos_i(8890) := b"1111111111111111_1111111111111111_1110101101011110_1001011001100011"; -- -0.08058796018998433
	pesos_i(8891) := b"0000000000000000_0000000000000000_0000100110100010_0111011011000100"; -- 0.0376352527972418
	pesos_i(8892) := b"1111111111111111_1111111111111111_1110110010100000_1010101101110101"; -- -0.07567337421908588
	pesos_i(8893) := b"0000000000000000_0000000000000000_0000000011000011_0000011101111011"; -- 0.002975909768894484
	pesos_i(8894) := b"1111111111111111_1111111111111111_1110011011100100_0011110110001011"; -- -0.09807982777665367
	pesos_i(8895) := b"1111111111111111_1111111111111111_1110110010101101_1000101000001101"; -- -0.0754770009672284
	pesos_i(8896) := b"1111111111111111_1111111111111111_1110100011111101_0110010110110000"; -- -0.08988346521218692
	pesos_i(8897) := b"1111111111111111_1111111111111111_1110101000001010_1110011010111110"; -- -0.08577115885015885
	pesos_i(8898) := b"0000000000000000_0000000000000000_0000000000001111_0000110001100011"; -- 0.00022962021495453322
	pesos_i(8899) := b"0000000000000000_0000000000000000_0010001101101111_0101000001101011"; -- 0.13841726881402622
	pesos_i(8900) := b"1111111111111111_1111111111111111_1101110001110100_1000101001010000"; -- -0.13884673650375737
	pesos_i(8901) := b"0000000000000000_0000000000000000_0000000001011101_0101111001010011"; -- 0.0014246896507816938
	pesos_i(8902) := b"1111111111111111_1111111111111111_1110110001100101_1101011111101010"; -- -0.07657099283859423
	pesos_i(8903) := b"1111111111111111_1111111111111111_1110011001001100_0100001001110111"; -- -0.10039887050652582
	pesos_i(8904) := b"0000000000000000_0000000000000000_0000001001010011_0000110111010111"; -- 0.009079804357866508
	pesos_i(8905) := b"1111111111111111_1111111111111111_1101100000101010_0010000100100100"; -- -0.15560715543915976
	pesos_i(8906) := b"0000000000000000_0000000000000000_0001110111000110_0100110011101011"; -- 0.11630707481221952
	pesos_i(8907) := b"0000000000000000_0000000000000000_0010011110010001_1001111000101111"; -- 0.15456570287433516
	pesos_i(8908) := b"1111111111111111_1111111111111111_1111011010110010_1001011001000111"; -- -0.036337478265767255
	pesos_i(8909) := b"1111111111111111_1111111111111111_1111010110000110_0111111000001011"; -- -0.04091655956794229
	pesos_i(8910) := b"0000000000000000_0000000000000000_0001000111001001_0001100101101110"; -- 0.06947478225545993
	pesos_i(8911) := b"0000000000000000_0000000000000000_0001100100011110_1111110010001100"; -- 0.09812906671839265
	pesos_i(8912) := b"0000000000000000_0000000000000000_0001011100010010_0100000001011100"; -- 0.09012224442664851
	pesos_i(8913) := b"0000000000000000_0000000000000000_0000100011000011_1101101010010010"; -- 0.03423849176320965
	pesos_i(8914) := b"1111111111111111_1111111111111111_1110111101010110_1000001001100101"; -- -0.06508622201496567
	pesos_i(8915) := b"1111111111111111_1111111111111111_1110010101100100_0011010001111010"; -- -0.10393974327414399
	pesos_i(8916) := b"1111111111111111_1111111111111111_1111001101011110_0101011010111001"; -- -0.04934175480083722
	pesos_i(8917) := b"0000000000000000_0000000000000000_0001000110100110_0000110000011111"; -- 0.06893993149616467
	pesos_i(8918) := b"0000000000000000_0000000000000000_0000100100011011_0011000010010101"; -- 0.03557113302538997
	pesos_i(8919) := b"1111111111111111_1111111111111111_1110100111111010_0110111010101110"; -- -0.08602245575751356
	pesos_i(8920) := b"1111111111111111_1111111111111111_1101010110001001_1000100010111011"; -- -0.16587014619938636
	pesos_i(8921) := b"1111111111111111_1111111111111111_1111110011001101_0001001101100010"; -- -0.012495793027680571
	pesos_i(8922) := b"0000000000000000_0000000000000000_0001010010000100_0110100011010110"; -- 0.0801454088592467
	pesos_i(8923) := b"1111111111111111_1111111111111111_1111011001100011_1001101000110111"; -- -0.03754268789183892
	pesos_i(8924) := b"0000000000000000_0000000000000000_0001001111110110_0100101110011100"; -- 0.07797691885206848
	pesos_i(8925) := b"0000000000000000_0000000000000000_0010000101110010_0110000000000110"; -- 0.13065147533007182
	pesos_i(8926) := b"0000000000000000_0000000000000000_0000100100010100_1100101010110010"; -- 0.035473507433201976
	pesos_i(8927) := b"1111111111111111_1111111111111111_1111001100001000_1111010100111011"; -- -0.05064456278245279
	pesos_i(8928) := b"1111111111111111_1111111111111111_1111110101001111_1111011000001001"; -- -0.010498640712735449
	pesos_i(8929) := b"1111111111111111_1111111111111111_1111111000010101_1001100000110100"; -- -0.007482993440431639
	pesos_i(8930) := b"1111111111111111_1111111111111111_1110101000001101_0101011011101111"; -- -0.08573395416540364
	pesos_i(8931) := b"1111111111111111_1111111111111111_1111010111100110_0001111100010001"; -- -0.039457376875123705
	pesos_i(8932) := b"1111111111111111_1111111111111111_1110101101001100_1010000100000010"; -- -0.0808619852527711
	pesos_i(8933) := b"0000000000000000_0000000000000000_0001111000001010_1010101101111101"; -- 0.11735030927311557
	pesos_i(8934) := b"1111111111111111_1111111111111111_1111110011000001_1001011111000000"; -- -0.012671008749224662
	pesos_i(8935) := b"1111111111111111_1111111111111111_1110100011010101_1100100001100010"; -- -0.09048793408065954
	pesos_i(8936) := b"1111111111111111_1111111111111111_1111111110010101_1000101100001101"; -- -0.0016244024600597013
	pesos_i(8937) := b"0000000000000000_0000000000000000_0001011110100010_0001000000100101"; -- 0.09231663609568573
	pesos_i(8938) := b"1111111111111111_1111111111111111_1101110011100011_1011001011000101"; -- -0.1371505993889196
	pesos_i(8939) := b"1111111111111111_1111111111111111_1101110110011110_0011111110110001"; -- -0.13430406502262743
	pesos_i(8940) := b"1111111111111111_1111111111111111_1110001010110011_0100101010000111"; -- -0.11445173456286473
	pesos_i(8941) := b"0000000000000000_0000000000000000_0000111110000110_1100111010010100"; -- 0.06065074080694206
	pesos_i(8942) := b"1111111111111111_1111111111111111_1111000100110100_1111010110101001"; -- -0.057785650448099024
	pesos_i(8943) := b"0000000000000000_0000000000000000_0010101001100100_1111110100110011"; -- 0.16560347084886393
	pesos_i(8944) := b"1111111111111111_1111111111111111_1110000001110011_0011010001101110"; -- -0.1232421143160208
	pesos_i(8945) := b"0000000000000000_0000000000000000_0000101001110001_1101110011110111"; -- 0.040799913695355544
	pesos_i(8946) := b"1111111111111111_1111111111111111_1110111011100100_0000100010110010"; -- -0.06683297790528954
	pesos_i(8947) := b"1111111111111111_1111111111111111_1101111100110010_0010000110000000"; -- -0.1281413138945248
	pesos_i(8948) := b"0000000000000000_0000000000000000_0000100101011000_0000001001100111"; -- 0.036499166679970364
	pesos_i(8949) := b"1111111111111111_1111111111111111_1110100000110100_0000111111001110"; -- -0.09295560098115618
	pesos_i(8950) := b"1111111111111111_1111111111111111_1111110111100011_1100001001100010"; -- -0.008243418852343089
	pesos_i(8951) := b"1111111111111111_1111111111111111_1110111101110010_1001100110001010"; -- -0.06465759630543343
	pesos_i(8952) := b"1111111111111111_1111111111111111_1110100101010011_1010111000100101"; -- -0.08856689072223303
	pesos_i(8953) := b"1111111111111111_1111111111111111_1111101100100111_1101101011011101"; -- -0.018923111876179108
	pesos_i(8954) := b"1111111111111111_1111111111111111_1111101000100100_0010111000001101"; -- -0.02288543874729504
	pesos_i(8955) := b"0000000000000000_0000000000000000_0001111110111100_0000000110001001"; -- 0.12396249384750946
	pesos_i(8956) := b"1111111111111111_1111111111111111_1110011001000010_1011001010101100"; -- -0.10054477015958188
	pesos_i(8957) := b"1111111111111111_1111111111111111_1110011111011111_1100100011100001"; -- -0.09424156677075037
	pesos_i(8958) := b"1111111111111111_1111111111111111_1101100110101011_1001100111111101"; -- -0.14972531868609
	pesos_i(8959) := b"0000000000000000_0000000000000000_0000100101011011_1101110110101011"; -- 0.036558012291917893
	pesos_i(8960) := b"0000000000000000_0000000000000000_0000100100101110_0001011010000000"; -- 0.035859495499797125
	pesos_i(8961) := b"0000000000000000_0000000000000000_0010010001011011_0010010111101101"; -- 0.14201581046636894
	pesos_i(8962) := b"0000000000000000_0000000000000000_0000111010001111_0111001010110110"; -- 0.05687634420482133
	pesos_i(8963) := b"1111111111111111_1111111111111111_1110011111110110_0000100101101010"; -- -0.09390202672745866
	pesos_i(8964) := b"1111111111111111_1111111111111111_1110101100011000_0110011111111111"; -- -0.08165884051366767
	pesos_i(8965) := b"0000000000000000_0000000000000000_0001101110100001_1011011011000001"; -- 0.10793630813450514
	pesos_i(8966) := b"0000000000000000_0000000000000000_0001100000100100_0000001010111111"; -- 0.09429948005227076
	pesos_i(8967) := b"1111111111111111_1111111111111111_1101111110001000_0011111110001101"; -- -0.1268272667302254
	pesos_i(8968) := b"0000000000000000_0000000000000000_0010011000000110_1000110100100001"; -- 0.1485374646503044
	pesos_i(8969) := b"1111111111111111_1111111111111111_1111100101101001_1110100100011101"; -- -0.025727682570706793
	pesos_i(8970) := b"0000000000000000_0000000000000000_0001000101110100_0011100110100001"; -- 0.068179704568871
	pesos_i(8971) := b"0000000000000000_0000000000000000_0001000010001001_0110111101110010"; -- 0.06459709664626179
	pesos_i(8972) := b"0000000000000000_0000000000000000_0010100100100010_0100001001010111"; -- 0.16067900289130635
	pesos_i(8973) := b"1111111111111111_1111111111111111_1101101101111111_0000111100101011"; -- -0.14259247971438882
	pesos_i(8974) := b"0000000000000000_0000000000000000_0000011011011110_1011011011011001"; -- 0.026835849849406814
	pesos_i(8975) := b"1111111111111111_1111111111111111_1110100111000110_1011010111111001"; -- -0.08681166344436023
	pesos_i(8976) := b"1111111111111111_1111111111111111_1110001111110000_1000010011110110"; -- -0.10961121557351407
	pesos_i(8977) := b"0000000000000000_0000000000000000_0001111110110101_0100111011101100"; -- 0.12386029490265436
	pesos_i(8978) := b"0000000000000000_0000000000000000_0010010010011110_1011000011010100"; -- 0.14304642847384313
	pesos_i(8979) := b"1111111111111111_1111111111111111_1110000001101101_1011011110000000"; -- -0.12332585453335464
	pesos_i(8980) := b"1111111111111111_1111111111111111_1110110100001011_1111110010001101"; -- -0.07403585009260774
	pesos_i(8981) := b"0000000000000000_0000000000000000_0000010100111011_1110010000101001"; -- 0.020445118075905707
	pesos_i(8982) := b"1111111111111111_1111111111111111_1110100001010100_0001001111110101"; -- -0.09246707214351803
	pesos_i(8983) := b"1111111111111111_1111111111111111_1101111101110100_0010000010000110"; -- -0.1271342920034826
	pesos_i(8984) := b"0000000000000000_0000000000000000_0010001010110001_0000010010000101"; -- 0.1355135750467461
	pesos_i(8985) := b"0000000000000000_0000000000000000_0001000110011001_1100100011111011"; -- 0.06875282414592253
	pesos_i(8986) := b"0000000000000000_0000000000000000_0001001110100000_0101001010110000"; -- 0.07666508492365462
	pesos_i(8987) := b"1111111111111111_1111111111111111_1111101011110000_1110111110111101"; -- -0.01976110103997204
	pesos_i(8988) := b"0000000000000000_0000000000000000_0001011000010011_1010010101011101"; -- 0.08623727340631984
	pesos_i(8989) := b"0000000000000000_0000000000000000_0001011100011100_0001101001010000"; -- 0.09027256446990573
	pesos_i(8990) := b"0000000000000000_0000000000000000_0010011110011001_1111010000000011"; -- 0.15469288899567693
	pesos_i(8991) := b"0000000000000000_0000000000000000_0001001001111010_0100000011101111"; -- 0.07217794261823827
	pesos_i(8992) := b"1111111111111111_1111111111111111_1110100011111111_0101110101110011"; -- -0.0898534388102882
	pesos_i(8993) := b"0000000000000000_0000000000000000_0001110101001000_1110000101111111"; -- 0.11439332353750513
	pesos_i(8994) := b"0000000000000000_0000000000000000_0010001101010111_0100010000110011"; -- 0.1380503295518449
	pesos_i(8995) := b"0000000000000000_0000000000000000_0000100011111110_1010001001111101"; -- 0.035135417449995085
	pesos_i(8996) := b"0000000000000000_0000000000000000_0000011111101100_0000110100100010"; -- 0.03094560687911812
	pesos_i(8997) := b"0000000000000000_0000000000000000_0010001111011001_0001001000000101"; -- 0.14003098128496608
	pesos_i(8998) := b"1111111111111111_1111111111111111_1111000100100111_1010100000110000"; -- -0.057988632475563004
	pesos_i(8999) := b"1111111111111111_1111111111111111_1111010101010111_1110101001001011"; -- -0.04162727038893719
	pesos_i(9000) := b"1111111111111111_1111111111111111_1101100010010000_0101111010101010"; -- -0.15404709195887298
	pesos_i(9001) := b"0000000000000000_0000000000000000_0001001001111110_1100010111001001"; -- 0.07224689633762928
	pesos_i(9002) := b"0000000000000000_0000000000000000_0001100111111101_1100000001111111"; -- 0.10152819739376094
	pesos_i(9003) := b"0000000000000000_0000000000000000_0000101011111111_0001110010100111"; -- 0.04295519901653156
	pesos_i(9004) := b"0000000000000000_0000000000000000_0001101100111011_1101011110001001"; -- 0.10638186538189956
	pesos_i(9005) := b"0000000000000000_0000000000000000_0000001011101010_0000011101100100"; -- 0.011383497177235637
	pesos_i(9006) := b"0000000000000000_0000000000000000_0010010000110111_1010110101001010"; -- 0.14147456222291344
	pesos_i(9007) := b"0000000000000000_0000000000000000_0010000011101001_0001001011011100"; -- 0.1285564220267951
	pesos_i(9008) := b"0000000000000000_0000000000000000_0001100011001011_0110010011101110"; -- 0.09685355013712749
	pesos_i(9009) := b"1111111111111111_1111111111111111_1111110000101111_1110000011111101"; -- -0.01489442663438957
	pesos_i(9010) := b"1111111111111111_1111111111111111_1110000000001110_0110001000101001"; -- -0.12478052606053107
	pesos_i(9011) := b"1111111111111111_1111111111111111_1110110011100001_0000100001001000"; -- -0.07469127880778359
	pesos_i(9012) := b"1111111111111111_1111111111111111_1110001000000000_0101011111001000"; -- -0.11718226776454203
	pesos_i(9013) := b"0000000000000000_0000000000000000_0000101010111101_1111111110000001"; -- 0.04196164033593265
	pesos_i(9014) := b"0000000000000000_0000000000000000_0010011100011010_0101101010001010"; -- 0.1527458750007366
	pesos_i(9015) := b"1111111111111111_1111111111111111_1101110001100100_0000010001000111"; -- -0.13909886614586586
	pesos_i(9016) := b"1111111111111111_1111111111111111_1111100110010010_1110100000111111"; -- -0.02510212382282008
	pesos_i(9017) := b"0000000000000000_0000000000000000_0000000001010001_1001101100001111"; -- 0.001245204093054958
	pesos_i(9018) := b"1111111111111111_1111111111111111_1110000000010000_1011111101011111"; -- -0.12474445286426995
	pesos_i(9019) := b"0000000000000000_0000000000000000_0000011101000111_0100110101100111"; -- 0.028431737474167697
	pesos_i(9020) := b"0000000000000000_0000000000000000_0000110001010010_1110110100110101"; -- 0.04814035935289701
	pesos_i(9021) := b"1111111111111111_1111111111111111_1111100101000011_0001111100011101"; -- -0.026319556658448304
	pesos_i(9022) := b"0000000000000000_0000000000000000_0010000000000110_1110000110110010"; -- 0.12510500522905882
	pesos_i(9023) := b"1111111111111111_1111111111111111_1111010101010010_0000110001010110"; -- -0.04171679405985484
	pesos_i(9024) := b"0000000000000000_0000000000000000_0000111000001110_1000010011111101"; -- 0.05490904972829723
	pesos_i(9025) := b"1111111111111111_1111111111111111_1110110011001001_0100010101001100"; -- -0.07505385291048813
	pesos_i(9026) := b"0000000000000000_0000000000000000_0000010001010100_0011010110100010"; -- 0.016909935131412476
	pesos_i(9027) := b"1111111111111111_1111111111111111_1101100001100110_1001101001111011"; -- -0.1546843958073434
	pesos_i(9028) := b"1111111111111111_1111111111111111_1111101011110110_1000010001111110"; -- -0.01967594065148499
	pesos_i(9029) := b"1111111111111111_1111111111111111_1110100001100110_1101001001000011"; -- -0.0921810708909002
	pesos_i(9030) := b"0000000000000000_0000000000000000_0001001110111000_0110101011001111"; -- 0.07703273355064963
	pesos_i(9031) := b"1111111111111111_1111111111111111_1110101000000101_0110101010111111"; -- -0.08585484353618072
	pesos_i(9032) := b"0000000000000000_0000000000000000_0010010110000100_1110111000101101"; -- 0.14655960657854927
	pesos_i(9033) := b"1111111111111111_1111111111111111_1101110001010010_0101100100001000"; -- -0.13936847252480114
	pesos_i(9034) := b"1111111111111111_1111111111111111_1111000000011110_1111110101010011"; -- -0.062027137064974334
	pesos_i(9035) := b"0000000000000000_0000000000000000_0000010000011110_0111101010000110"; -- 0.016090066531365313
	pesos_i(9036) := b"1111111111111111_1111111111111111_1110111110010000_1011000110001101"; -- -0.06419840145279086
	pesos_i(9037) := b"1111111111111111_1111111111111111_1111001101111011_1010110010110000"; -- -0.048894126061298344
	pesos_i(9038) := b"1111111111111111_1111111111111111_1110100110011010_0001000111110001"; -- -0.08749282700461254
	pesos_i(9039) := b"1111111111111111_1111111111111111_1110011011110001_1011010010000111"; -- -0.09787437163019777
	pesos_i(9040) := b"0000000000000000_0000000000000000_0001001111001110_1111101011001110"; -- 0.07737700963608825
	pesos_i(9041) := b"1111111111111111_1111111111111111_1111100001111101_1011111011100000"; -- -0.02933127422598785
	pesos_i(9042) := b"1111111111111111_1111111111111111_1111000001100100_0010011001010111"; -- -0.06097183589337527
	pesos_i(9043) := b"0000000000000000_0000000000000000_0000000001001110_1000101101000010"; -- 0.0011984860603231552
	pesos_i(9044) := b"1111111111111111_1111111111111111_1101101110110111_1100000001011101"; -- -0.1417274259131067
	pesos_i(9045) := b"1111111111111111_1111111111111111_1110011000100111_0001010000011110"; -- -0.10096620820403113
	pesos_i(9046) := b"1111111111111111_1111111111111111_1101100001101000_0110100011001101"; -- -0.1546568392685829
	pesos_i(9047) := b"1111111111111111_1111111111111111_1110100110010001_1001001111001110"; -- -0.08762241568338489
	pesos_i(9048) := b"1111111111111111_1111111111111111_1111010111011100_1101011110011000"; -- -0.039598966086508244
	pesos_i(9049) := b"1111111111111111_1111111111111111_1101111101101110_0010010101010000"; -- -0.12722555926164644
	pesos_i(9050) := b"1111111111111111_1111111111111111_1111010111101100_0110010000111001"; -- -0.039361702065182545
	pesos_i(9051) := b"0000000000000000_0000000000000000_0001110010010000_0010101001111011"; -- 0.11157479775948705
	pesos_i(9052) := b"0000000000000000_0000000000000000_0010000010001110_1000010100110001"; -- 0.1271746869155487
	pesos_i(9053) := b"1111111111111111_1111111111111111_1110110100110011_0010110011001010"; -- -0.0734378821094029
	pesos_i(9054) := b"0000000000000000_0000000000000000_0000001011100101_1010001101011011"; -- 0.011316499511995903
	pesos_i(9055) := b"0000000000000000_0000000000000000_0000000100010110_0010000000011110"; -- 0.0042438577370422
	pesos_i(9056) := b"1111111111111111_1111111111111111_1111000001111101_1010010011000110"; -- -0.06058283006044882
	pesos_i(9057) := b"1111111111111111_1111111111111111_1110110111110001_0110111100001001"; -- -0.07053476369146668
	pesos_i(9058) := b"0000000000000000_0000000000000000_0000100100101101_0000101111100100"; -- 0.035843604348797395
	pesos_i(9059) := b"0000000000000000_0000000000000000_0000011101011111_0111111001100001"; -- 0.028800867839495925
	pesos_i(9060) := b"0000000000000000_0000000000000000_0000010110001101_1111010011011100"; -- 0.021697334040933075
	pesos_i(9061) := b"1111111111111111_1111111111111111_1111111100110001_1110011101101011"; -- -0.0031447758059640406
	pesos_i(9062) := b"0000000000000000_0000000000000000_0010000010011101_0110110111001011"; -- 0.1274021740635334
	pesos_i(9063) := b"0000000000000000_0000000000000000_0010010000000001_1100101011111100"; -- 0.14065235760338948
	pesos_i(9064) := b"1111111111111111_1111111111111111_1101011110111010_0001011000011101"; -- -0.15731679720553474
	pesos_i(9065) := b"1111111111111111_1111111111111111_1111011010110111_0001100011100111"; -- -0.03626865740545895
	pesos_i(9066) := b"0000000000000000_0000000000000000_0000110011111000_0011011001000111"; -- 0.050662414890516726
	pesos_i(9067) := b"0000000000000000_0000000000000000_0000110101111101_1111101101001110"; -- 0.05270357753988196
	pesos_i(9068) := b"1111111111111111_1111111111111111_1101100010100000_0001010011000010"; -- -0.15380735649652535
	pesos_i(9069) := b"1111111111111111_1111111111111111_1101110010100100_1010100111110011"; -- -0.1381124287651714
	pesos_i(9070) := b"1111111111111111_1111111111111111_1101110011100100_0100010011100000"; -- -0.13714189077571998
	pesos_i(9071) := b"1111111111111111_1111111111111111_1110101101011011_1010010101111000"; -- -0.08063283755605315
	pesos_i(9072) := b"1111111111111111_1111111111111111_1110100000011010_1100101010000010"; -- -0.09334120113328744
	pesos_i(9073) := b"1111111111111111_1111111111111111_1101110011010101_1101110110001001"; -- -0.13736167329948312
	pesos_i(9074) := b"0000000000000000_0000000000000000_0010000110110000_1000100011101001"; -- 0.13159995737170865
	pesos_i(9075) := b"1111111111111111_1111111111111111_1110111001001001_0001100100100100"; -- -0.06919710989770943
	pesos_i(9076) := b"0000000000000000_0000000000000000_0001111110000011_0000011101111110"; -- 0.12309309786485957
	pesos_i(9077) := b"0000000000000000_0000000000000000_0010100001100001_1101110111111100"; -- 0.1577433337241869
	pesos_i(9078) := b"0000000000000000_0000000000000000_0010000000010101_0000010001101010"; -- 0.125320697715443
	pesos_i(9079) := b"1111111111111111_1111111111111111_1111111001000000_0011110010011110"; -- -0.006832324399133642
	pesos_i(9080) := b"0000000000000000_0000000000000000_0001101000000101_0010000101101010"; -- 0.10164078564385422
	pesos_i(9081) := b"1111111111111111_1111111111111111_1111000001110000_1110110010111101"; -- -0.06077690488117958
	pesos_i(9082) := b"1111111111111111_1111111111111111_1111010010011010_0100011010000100"; -- -0.04452094343942537
	pesos_i(9083) := b"0000000000000000_0000000000000000_0000111101111111_1100000001111011"; -- 0.0605430888306552
	pesos_i(9084) := b"0000000000000000_0000000000000000_0001000001001001_1010010111110111"; -- 0.06362378397825919
	pesos_i(9085) := b"1111111111111111_1111111111111111_1110000110001101_1110101100100101"; -- -0.11892824509584568
	pesos_i(9086) := b"1111111111111111_1111111111111111_1111001111000100_0110100010010111"; -- -0.04778429331297493
	pesos_i(9087) := b"0000000000000000_0000000000000000_0010000101001000_1011110010010010"; -- 0.13001612250031305
	pesos_i(9088) := b"0000000000000000_0000000000000000_0000011010011011_1011010010110001"; -- 0.025813382459457444
	pesos_i(9089) := b"0000000000000000_0000000000000000_0000111111101010_1000101000010101"; -- 0.06217253704806673
	pesos_i(9090) := b"0000000000000000_0000000000000000_0000011010010001_0110011111011110"; -- 0.025656215480850557
	pesos_i(9091) := b"0000000000000000_0000000000000000_0001001100001111_0101100101100111"; -- 0.0744529606908687
	pesos_i(9092) := b"0000000000000000_0000000000000000_0010000010100001_0100100000101101"; -- 0.12746096697169215
	pesos_i(9093) := b"1111111111111111_1111111111111111_1111101010011101_1110011011011110"; -- -0.021028109250850212
	pesos_i(9094) := b"1111111111111111_1111111111111111_1111111110011010_1010101011001010"; -- -0.0015462166821449414
	pesos_i(9095) := b"0000000000000000_0000000000000000_0001000000010100_1111010100001001"; -- 0.06281978095923996
	pesos_i(9096) := b"1111111111111111_1111111111111111_1110011111110000_0100011111110001"; -- -0.09398985256534031
	pesos_i(9097) := b"1111111111111111_1111111111111111_1110011101000001_1010110001000100"; -- -0.0966541609633006
	pesos_i(9098) := b"0000000000000000_0000000000000000_0000111100010110_1111011010101001"; -- 0.05894414546787511
	pesos_i(9099) := b"0000000000000000_0000000000000000_0001110110100100_0100000101101100"; -- 0.1157875908307423
	pesos_i(9100) := b"0000000000000000_0000000000000000_0000000010001011_1011011101011010"; -- 0.002131900182815047
	pesos_i(9101) := b"0000000000000000_0000000000000000_0001011111110001_0001001100101101"; -- 0.09352226122161675
	pesos_i(9102) := b"0000000000000000_0000000000000000_0001001011101001_0011100111110101"; -- 0.07387125230500961
	pesos_i(9103) := b"1111111111111111_1111111111111111_1111011011001101_1001101010110011"; -- -0.035925227450204496
	pesos_i(9104) := b"1111111111111111_1111111111111111_1101111000101000_0001111110110000"; -- -0.13220025980064895
	pesos_i(9105) := b"1111111111111111_1111111111111111_1111001010010100_1101110011111110"; -- -0.05241602717145559
	pesos_i(9106) := b"1111111111111111_1111111111111111_1111110100000011_0110111010010001"; -- -0.011666383268938303
	pesos_i(9107) := b"0000000000000000_0000000000000000_0001110011111010_0110010101010011"; -- 0.11319573666931156
	pesos_i(9108) := b"0000000000000000_0000000000000000_0010000101010000_0111010001010100"; -- 0.1301338868904803
	pesos_i(9109) := b"1111111111111111_1111111111111111_1110100001000010_1001100100001000"; -- -0.09273379857065825
	pesos_i(9110) := b"0000000000000000_0000000000000000_0001011011010101_0010100011111000"; -- 0.08919006404200558
	pesos_i(9111) := b"1111111111111111_1111111111111111_1111111111001001_0111100101101111"; -- -0.0008319953028294345
	pesos_i(9112) := b"0000000000000000_0000000000000000_0001101100100110_1000100010111001"; -- 0.10605673320225242
	pesos_i(9113) := b"1111111111111111_1111111111111111_1110001100000100_1100010001101001"; -- -0.11320850783947566
	pesos_i(9114) := b"0000000000000000_0000000000000000_0000111100100101_1011101001101110"; -- 0.05916943734250261
	pesos_i(9115) := b"1111111111111111_1111111111111111_1110110111110100_1011000011001101"; -- -0.07048506733022807
	pesos_i(9116) := b"1111111111111111_1111111111111111_1110101011001000_1010011101011010"; -- -0.08287576720196063
	pesos_i(9117) := b"0000000000000000_0000000000000000_0000100000000011_1010110110100100"; -- 0.03130612618388024
	pesos_i(9118) := b"1111111111111111_1111111111111111_1110111000010010_0100100001010100"; -- -0.07003353074426294
	pesos_i(9119) := b"0000000000000000_0000000000000000_0010100110100101_1110010000000100"; -- 0.16268754110171696
	pesos_i(9120) := b"0000000000000000_0000000000000000_0000000001100101_0101110011000011"; -- 0.0015466667708685313
	pesos_i(9121) := b"1111111111111111_1111111111111111_1110101100111101_1001011100011011"; -- -0.08109145725177277
	pesos_i(9122) := b"1111111111111111_1111111111111111_1110100110001001_1101110101011111"; -- -0.0877401012315446
	pesos_i(9123) := b"1111111111111111_1111111111111111_1111111111001011_1100000001101011"; -- -0.0007972467827165118
	pesos_i(9124) := b"1111111111111111_1111111111111111_1111001100100111_1000001100100001"; -- -0.05017834128550467
	pesos_i(9125) := b"1111111111111111_1111111111111111_1111001101011011_0000111101010001"; -- -0.04939178731631905
	pesos_i(9126) := b"0000000000000000_0000000000000000_0000110111001100_0101110110101101"; -- 0.05389962638024617
	pesos_i(9127) := b"0000000000000000_0000000000000000_0010010011000001_0101101111100010"; -- 0.14357542304605742
	pesos_i(9128) := b"1111111111111111_1111111111111111_1101100011110111_1101101110110001"; -- -0.15246798458293587
	pesos_i(9129) := b"1111111111111111_1111111111111111_1111001101001000_0001110001001010"; -- -0.04968093102203732
	pesos_i(9130) := b"0000000000000000_0000000000000000_0010000010001110_1011100111001101"; -- 0.12717782267984312
	pesos_i(9131) := b"0000000000000000_0000000000000000_0010000000101111_1001111100011110"; -- 0.12572664719813756
	pesos_i(9132) := b"0000000000000000_0000000000000000_0001001000101011_0110111100000101"; -- 0.07097524527327767
	pesos_i(9133) := b"1111111111111111_1111111111111111_1111000010101001_0110010001000110"; -- -0.059915287982854636
	pesos_i(9134) := b"0000000000000000_0000000000000000_0010000111111111_0101001010011010"; -- 0.1328021645838286
	pesos_i(9135) := b"0000000000000000_0000000000000000_0000111011010101_1010010101100000"; -- 0.057947479268165625
	pesos_i(9136) := b"0000000000000000_0000000000000000_0001111011100111_1110001010111001"; -- 0.12072579394369985
	pesos_i(9137) := b"1111111111111111_1111111111111111_1110011101001110_1111001010110110"; -- -0.09645159766790802
	pesos_i(9138) := b"1111111111111111_1111111111111111_1111010010000111_0101101101111100"; -- -0.04480961061956801
	pesos_i(9139) := b"0000000000000000_0000000000000000_0000110000011000_0010100110101101"; -- 0.047243694916997564
	pesos_i(9140) := b"1111111111111111_1111111111111111_1111001000100011_0100001110111101"; -- -0.05414940491235493
	pesos_i(9141) := b"1111111111111111_1111111111111111_1110100100100111_0001101011101000"; -- -0.0892470534780309
	pesos_i(9142) := b"1111111111111111_1111111111111111_1111010001011110_0001110000111110"; -- -0.0454389904300259
	pesos_i(9143) := b"1111111111111111_1111111111111111_1111011101000010_0001110001001010"; -- -0.03414748369943658
	pesos_i(9144) := b"1111111111111111_1111111111111111_1110101101000011_1111101011010010"; -- -0.08099396110424918
	pesos_i(9145) := b"1111111111111111_1111111111111111_1110110110000110_1011111110100011"; -- -0.07216264971823552
	pesos_i(9146) := b"0000000000000000_0000000000000000_0010011010100101_0010011101001101"; -- 0.15095754272904316
	pesos_i(9147) := b"0000000000000000_0000000000000000_0000110000011001_1110000110001000"; -- 0.04726991235527561
	pesos_i(9148) := b"1111111111111111_1111111111111111_1110000011110100_0000110001111010"; -- -0.12127611183063915
	pesos_i(9149) := b"1111111111111111_1111111111111111_1111111010110001_0000111011000101"; -- -0.005110814007216783
	pesos_i(9150) := b"0000000000000000_0000000000000000_0000010111111100_1101011011100101"; -- 0.0233892734429693
	pesos_i(9151) := b"1111111111111111_1111111111111111_1111101101110010_1000000001001011"; -- -0.017784101098769097
	pesos_i(9152) := b"0000000000000000_0000000000000000_0010101001111100_0010000001100000"; -- 0.16595651956951735
	pesos_i(9153) := b"0000000000000000_0000000000000000_0000101101000101_0100100010001101"; -- 0.04402593073274579
	pesos_i(9154) := b"1111111111111111_1111111111111111_1110110000111011_0111110101000111"; -- -0.07721726428734256
	pesos_i(9155) := b"0000000000000000_0000000000000000_0000111011001111_1001111000010110"; -- 0.057855491879266904
	pesos_i(9156) := b"0000000000000000_0000000000000000_0000000101101000_0011001110100010"; -- 0.005496241609469214
	pesos_i(9157) := b"1111111111111111_1111111111111111_1110000101110100_0111101101000110"; -- -0.11931638277461454
	pesos_i(9158) := b"0000000000000000_0000000000000000_0010011011000111_0000111010111100"; -- 0.15147487736783743
	pesos_i(9159) := b"1111111111111111_1111111111111111_1110100100011111_1011100000110100"; -- -0.08935974827069344
	pesos_i(9160) := b"0000000000000000_0000000000000000_0010000010110011_0100000011001110"; -- 0.1277351859778856
	pesos_i(9161) := b"0000000000000000_0000000000000000_0000011010101000_0001111110011110"; -- 0.026002861208918614
	pesos_i(9162) := b"0000000000000000_0000000000000000_0000011011111010_1100110001111100"; -- 0.02726438556933013
	pesos_i(9163) := b"1111111111111111_1111111111111111_1111101001100100_1010011100110100"; -- -0.021901655076176786
	pesos_i(9164) := b"0000000000000000_0000000000000000_0000010000010101_0111100111010111"; -- 0.01595269668864482
	pesos_i(9165) := b"0000000000000000_0000000000000000_0000001111000100_1010010101000110"; -- 0.01471932379400344
	pesos_i(9166) := b"0000000000000000_0000000000000000_0010100011011010_1110101000101101"; -- 0.15959037389235456
	pesos_i(9167) := b"1111111111111111_1111111111111111_1101111110101100_1011101111110001"; -- -0.12627053611903555
	pesos_i(9168) := b"0000000000000000_0000000000000000_0000000000001011_1010001110110111"; -- 0.00017760496007616683
	pesos_i(9169) := b"0000000000000000_0000000000000000_0000100110011010_1010100011111001"; -- 0.03751617514797718
	pesos_i(9170) := b"0000000000000000_0000000000000000_0000001100010010_1101100111010010"; -- 0.012006391299352874
	pesos_i(9171) := b"1111111111111111_1111111111111111_1110001001100011_0000110011011001"; -- -0.1156761140024329
	pesos_i(9172) := b"1111111111111111_1111111111111111_1101101100101101_1111101110001100"; -- -0.1438296111769628
	pesos_i(9173) := b"0000000000000000_0000000000000000_0000100000001001_0000111101111101"; -- 0.03138825225108479
	pesos_i(9174) := b"1111111111111111_1111111111111111_1110101011011101_0111001001100010"; -- -0.08255848976651113
	pesos_i(9175) := b"0000000000000000_0000000000000000_0000000111011101_0111011000100110"; -- 0.007285484682918466
	pesos_i(9176) := b"1111111111111111_1111111111111111_1111111000110100_0110010101100100"; -- -0.007012999573128291
	pesos_i(9177) := b"1111111111111111_1111111111111111_1110000011000011_0000101101001101"; -- -0.12202386259441612
	pesos_i(9178) := b"0000000000000000_0000000000000000_0000001010100010_0011110010011001"; -- 0.010288035813474202
	pesos_i(9179) := b"0000000000000000_0000000000000000_0001010101111000_0100001101001001"; -- 0.08386631530016359
	pesos_i(9180) := b"0000000000000000_0000000000000000_0000011110001101_0011011101001111"; -- 0.029498535839362443
	pesos_i(9181) := b"1111111111111111_1111111111111111_1110101100000001_0111011011010101"; -- -0.08200890831271386
	pesos_i(9182) := b"1111111111111111_1111111111111111_1111011011110110_1110110010011000"; -- -0.03529473575653739
	pesos_i(9183) := b"1111111111111111_1111111111111111_1101111000111001_0000101000100011"; -- -0.13194214486498532
	pesos_i(9184) := b"0000000000000000_0000000000000000_0000110011000100_0110001111101011"; -- 0.04987167829920597
	pesos_i(9185) := b"1111111111111111_1111111111111111_1111000111010000_0000001110100111"; -- -0.05541970423455404
	pesos_i(9186) := b"0000000000000000_0000000000000000_0000011111010011_1111011100010111"; -- 0.03057808221722808
	pesos_i(9187) := b"1111111111111111_1111111111111111_1110110011010101_1110100011001001"; -- -0.07486100284003143
	pesos_i(9188) := b"1111111111111111_1111111111111111_1110111100011011_1111110010010001"; -- -0.06597920853519759
	pesos_i(9189) := b"0000000000000000_0000000000000000_0010001110000101_0111011011111010"; -- 0.13875526040179262
	pesos_i(9190) := b"0000000000000000_0000000000000000_0000100000101100_1100100010101000"; -- 0.031933346682520944
	pesos_i(9191) := b"1111111111111111_1111111111111111_1101011111000010_1011010000111001"; -- -0.15718530281868728
	pesos_i(9192) := b"1111111111111111_1111111111111111_1111110110010000_1001010010010100"; -- -0.009512628506499393
	pesos_i(9193) := b"1111111111111111_1111111111111111_1111100001101010_1111110111111001"; -- -0.029617430395278088
	pesos_i(9194) := b"1111111111111111_1111111111111111_1111100100110001_0010000100100001"; -- -0.02659409461350578
	pesos_i(9195) := b"0000000000000000_0000000000000000_0000011010000110_1101000001100110"; -- 0.025494599170887977
	pesos_i(9196) := b"0000000000000000_0000000000000000_0001010001001111_0010111110001100"; -- 0.07933327836466782
	pesos_i(9197) := b"1111111111111111_1111111111111111_1110110000001001_1010110110010010"; -- -0.0779773252898136
	pesos_i(9198) := b"1111111111111111_1111111111111111_1111010010010000_0100001111001110"; -- -0.04467369292796911
	pesos_i(9199) := b"1111111111111111_1111111111111111_1110101100001110_0100010010011011"; -- -0.08181353780945873
	pesos_i(9200) := b"1111111111111111_1111111111111111_1111100110110111_0111110010100001"; -- -0.02454396322298829
	pesos_i(9201) := b"1111111111111111_1111111111111111_1110100001011001_1000001101010010"; -- -0.09238414046772762
	pesos_i(9202) := b"1111111111111111_1111111111111111_1111110110111110_1001100000101100"; -- -0.008810509897296832
	pesos_i(9203) := b"0000000000000000_0000000000000000_0001111110110000_0011100010101001"; -- 0.1237826741254611
	pesos_i(9204) := b"1111111111111111_1111111111111111_1111001100001010_1110010011100000"; -- -0.05061502010699885
	pesos_i(9205) := b"0000000000000000_0000000000000000_0001110001001000_0010101110111100"; -- 0.11047623949203471
	pesos_i(9206) := b"0000000000000000_0000000000000000_0001010010000011_0000010101100110"; -- 0.08012422307580873
	pesos_i(9207) := b"0000000000000000_0000000000000000_0001011110111011_1100110101011000"; -- 0.09270938308077935
	pesos_i(9208) := b"0000000000000000_0000000000000000_0010010000110101_1001111110010000"; -- 0.1414432264577426
	pesos_i(9209) := b"0000000000000000_0000000000000000_0000000010111101_1100000001111111"; -- 0.0028953849069552956
	pesos_i(9210) := b"0000000000000000_0000000000000000_0000010011100101_1010011101110001"; -- 0.019129242964190427
	pesos_i(9211) := b"0000000000000000_0000000000000000_0001110001010000_1001100101111001"; -- 0.11060485070333183
	pesos_i(9212) := b"1111111111111111_1111111111111111_1101011111011001_0111101010110010"; -- -0.1568377795381608
	pesos_i(9213) := b"0000000000000000_0000000000000000_0001100000101101_0101001111101100"; -- 0.09444164773496111
	pesos_i(9214) := b"1111111111111111_1111111111111111_1110011111011101_0000111111100001"; -- -0.09428311114932872
	pesos_i(9215) := b"0000000000000000_0000000000000000_0001011111000000_0110110100110100"; -- 0.09277994657953191
	pesos_i(9216) := b"1111111111111111_1111111111111111_1110101000011010_1101100001110111"; -- -0.08552786906552366
	pesos_i(9217) := b"0000000000000000_0000000000000000_0010000111110100_1001110100100111"; -- 0.13263876146555711
	pesos_i(9218) := b"1111111111111111_1111111111111111_1101110110000011_0001110000111011"; -- -0.13471816585639634
	pesos_i(9219) := b"0000000000000000_0000000000000000_0000001011001101_1100010010001111"; -- 0.010952267605737358
	pesos_i(9220) := b"1111111111111111_1111111111111111_1101011000001000_1101000011100111"; -- -0.1639279780504608
	pesos_i(9221) := b"0000000000000000_0000000000000000_0010001111100100_1100001001101011"; -- 0.1402093422062245
	pesos_i(9222) := b"1111111111111111_1111111111111111_1101101110011001_0100001101101000"; -- -0.14219263748121444
	pesos_i(9223) := b"1111111111111111_1111111111111111_1101110100101100_1110111100011101"; -- -0.13603311094212572
	pesos_i(9224) := b"1111111111111111_1111111111111111_1111011100010110_0110100111111100"; -- -0.0348142394992219
	pesos_i(9225) := b"0000000000000000_0000000000000000_0001110100010000_0011001000010011"; -- 0.11352837535128428
	pesos_i(9226) := b"0000000000000000_0000000000000000_0010000111010101_1001100010100101"; -- 0.13216547038502205
	pesos_i(9227) := b"1111111111111111_1111111111111111_1101111111001010_1001001001001011"; -- -0.12581525480286254
	pesos_i(9228) := b"0000000000000000_0000000000000000_0001010010010100_1110111111100010"; -- 0.08039759899201754
	pesos_i(9229) := b"1111111111111111_1111111111111111_1110100110001111_1111000011110011"; -- -0.08764738149941673
	pesos_i(9230) := b"0000000000000000_0000000000000000_0001010010110110_0100101110011110"; -- 0.08090660676319186
	pesos_i(9231) := b"1111111111111111_1111111111111111_1111000100101110_0001111100100110"; -- -0.057889988997561606
	pesos_i(9232) := b"0000000000000000_0000000000000000_0000110100110010_1011101100000110"; -- 0.05155533682873476
	pesos_i(9233) := b"1111111111111111_1111111111111111_1111000101101111_0100000110011011"; -- -0.0568961139595572
	pesos_i(9234) := b"0000000000000000_0000000000000000_0000001111001111_1110110111110111"; -- 0.014891503121198716
	pesos_i(9235) := b"1111111111111111_1111111111111111_1111100100100101_1000000001000001"; -- -0.0267715303894008
	pesos_i(9236) := b"1111111111111111_1111111111111111_1110000100100001_1010010100111111"; -- -0.12058036057039338
	pesos_i(9237) := b"1111111111111111_1111111111111111_1111010011011000_0010000110110001"; -- -0.04357709331433433
	pesos_i(9238) := b"1111111111111111_1111111111111111_1111011000001001_1000011010001100"; -- -0.038917151273894675
	pesos_i(9239) := b"0000000000000000_0000000000000000_0000000011100001_0110101010111011"; -- 0.003439589214235284
	pesos_i(9240) := b"0000000000000000_0000000000000000_0001001111000111_1101110100010100"; -- 0.07726842640755253
	pesos_i(9241) := b"1111111111111111_1111111111111111_1110110110000010_0110001010111100"; -- -0.07222922230586366
	pesos_i(9242) := b"0000000000000000_0000000000000000_0001001010011110_0101000110110011"; -- 0.0727282582321481
	pesos_i(9243) := b"1111111111111111_1111111111111111_1101101101100011_0101010011011010"; -- -0.14301557241979665
	pesos_i(9244) := b"0000000000000000_0000000000000000_0000000000110001_0100110111110011"; -- 0.0007523268649503045
	pesos_i(9245) := b"1111111111111111_1111111111111111_1111001101011011_1001110010011101"; -- -0.049383365377970584
	pesos_i(9246) := b"0000000000000000_0000000000000000_0010001011000011_1010011100010101"; -- 0.1357979226401014
	pesos_i(9247) := b"1111111111111111_1111111111111111_1111010101101100_0011111001111010"; -- -0.04131707694308269
	pesos_i(9248) := b"1111111111111111_1111111111111111_1110010110110011_0010111011001100"; -- -0.10273463737885619
	pesos_i(9249) := b"0000000000000000_0000000000000000_0001110100100000_1001011101110101"; -- 0.113778558693557
	pesos_i(9250) := b"0000000000000000_0000000000000000_0001011100111111_1110001100101111"; -- 0.09081859480675876
	pesos_i(9251) := b"0000000000000000_0000000000000000_0001011101101110_1000111111100111"; -- 0.09153079392866793
	pesos_i(9252) := b"0000000000000000_0000000000000000_0001101010101101_0011001101011001"; -- 0.10420533116821586
	pesos_i(9253) := b"1111111111111111_1111111111111111_1110101010111011_1010011101111111"; -- -0.08307412285649499
	pesos_i(9254) := b"1111111111111111_1111111111111111_1111100010101100_0010100001000111"; -- -0.028623087642290206
	pesos_i(9255) := b"1111111111111111_1111111111111111_1110000111101000_1110111111001001"; -- -0.11753941863117759
	pesos_i(9256) := b"1111111111111111_1111111111111111_1111111100001110_1001001011100101"; -- -0.0036838713883723304
	pesos_i(9257) := b"0000000000000000_0000000000000000_0000000111011001_0001110100000110"; -- 0.007219137045357265
	pesos_i(9258) := b"1111111111111111_1111111111111111_1111111110000100_0011001100101110"; -- -0.0018890392104385398
	pesos_i(9259) := b"0000000000000000_0000000000000000_0001101011111001_0010001111000110"; -- 0.10536407076078624
	pesos_i(9260) := b"0000000000000000_0000000000000000_0010001011101110_0111111001000001"; -- 0.13645161712808881
	pesos_i(9261) := b"0000000000000000_0000000000000000_0010010001101100_0100101110111100"; -- 0.14227746328981675
	pesos_i(9262) := b"0000000000000000_0000000000000000_0000001010100110_1001110101110001"; -- 0.010354843185732413
	pesos_i(9263) := b"0000000000000000_0000000000000000_0000110001001001_0110110101110001"; -- 0.04799541479229559
	pesos_i(9264) := b"0000000000000000_0000000000000000_0000111100001101_1110100101110111"; -- 0.05880602983496808
	pesos_i(9265) := b"1111111111111111_1111111111111111_1111011101010110_0010000100011011"; -- -0.03384202101040827
	pesos_i(9266) := b"1111111111111111_1111111111111111_1110010010011111_1100011010110011"; -- -0.10693700916444697
	pesos_i(9267) := b"0000000000000000_0000000000000000_0010001010000000_1011000100011100"; -- 0.13477618161367755
	pesos_i(9268) := b"0000000000000000_0000000000000000_0010000111001001_1110011111011010"; -- 0.13198708613383864
	pesos_i(9269) := b"1111111111111111_1111111111111111_1110111000011000_1100110101100101"; -- -0.06993404661746061
	pesos_i(9270) := b"1111111111111111_1111111111111111_1111111100011100_1000000010011011"; -- -0.003471338323621328
	pesos_i(9271) := b"0000000000000000_0000000000000000_0001100100010110_0101011001111010"; -- 0.0979970976589115
	pesos_i(9272) := b"1111111111111111_1111111111111111_1101111101110010_0000010010111011"; -- -0.1271664660060757
	pesos_i(9273) := b"0000000000000000_0000000000000000_0001100101100011_0001110001101110"; -- 0.09916856476173896
	pesos_i(9274) := b"0000000000000000_0000000000000000_0000101100101010_0101001010001001"; -- 0.043614538650919764
	pesos_i(9275) := b"0000000000000000_0000000000000000_0001000011010011_0100000100011111"; -- 0.06572348596104832
	pesos_i(9276) := b"1111111111111111_1111111111111111_1111110111111000_0111000110010011"; -- -0.007927800711897262
	pesos_i(9277) := b"0000000000000000_0000000000000000_0000110000001101_1000011101011011"; -- 0.04708143203382195
	pesos_i(9278) := b"1111111111111111_1111111111111111_1111111000001001_1001010101001101"; -- -0.007666271925600766
	pesos_i(9279) := b"1111111111111111_1111111111111111_1110001100101011_1111000100001000"; -- -0.11261075555219757
	pesos_i(9280) := b"0000000000000000_0000000000000000_0010001000101100_1111110101100100"; -- 0.1334989900808685
	pesos_i(9281) := b"0000000000000000_0000000000000000_0000101011011111_0001011010011111"; -- 0.042466558356344275
	pesos_i(9282) := b"1111111111111111_1111111111111111_1111000001101010_1001100000100110"; -- -0.06087349969687161
	pesos_i(9283) := b"0000000000000000_0000000000000000_0000000110101010_1110111101110011"; -- 0.006514516485816648
	pesos_i(9284) := b"0000000000000000_0000000000000000_0000000001101111_1111101001000010"; -- 0.001708642111185156
	pesos_i(9285) := b"1111111111111111_1111111111111111_1110101100110000_1101001111011010"; -- -0.08128620075947608
	pesos_i(9286) := b"0000000000000000_0000000000000000_0000001011011100_1111010011111010"; -- 0.011184035236459958
	pesos_i(9287) := b"1111111111111111_1111111111111111_1111001010110000_0100011110000000"; -- -0.05199769141563205
	pesos_i(9288) := b"1111111111111111_1111111111111111_1110100111100010_0001101001110010"; -- -0.0863936873915094
	pesos_i(9289) := b"0000000000000000_0000000000000000_0001000001001100_1000111000001101"; -- 0.06366813491543952
	pesos_i(9290) := b"0000000000000000_0000000000000000_0001101000010001_0100010100110100"; -- 0.10182602419272702
	pesos_i(9291) := b"0000000000000000_0000000000000000_0001011111101110_0010111011110111"; -- 0.09347814119659566
	pesos_i(9292) := b"1111111111111111_1111111111111111_1111011001010101_1110010111011000"; -- -0.03775180317663518
	pesos_i(9293) := b"0000000000000000_0000000000000000_0000100010100100_0111011111111100"; -- 0.03375959303747701
	pesos_i(9294) := b"1111111111111111_1111111111111111_1111000000000000_1001101001000111"; -- -0.06249080434912423
	pesos_i(9295) := b"1111111111111111_1111111111111111_1111010101111111_0010100101110001"; -- -0.041028413605003776
	pesos_i(9296) := b"1111111111111111_1111111111111111_1110011110011000_0110010010110110"; -- -0.09533091121337474
	pesos_i(9297) := b"0000000000000000_0000000000000000_0000100110111101_1011111100011111"; -- 0.03805155288775413
	pesos_i(9298) := b"1111111111111111_1111111111111111_1110000100000000_1010110101000111"; -- -0.12108342196021264
	pesos_i(9299) := b"1111111111111111_1111111111111111_1110011110010110_1011101110100110"; -- -0.09535624682734123
	pesos_i(9300) := b"1111111111111111_1111111111111111_1110101000110001_1111011101001001"; -- -0.08517507999886928
	pesos_i(9301) := b"1111111111111111_1111111111111111_1110001100010010_0010011100101100"; -- -0.11300425693690806
	pesos_i(9302) := b"1111111111111111_1111111111111111_1110001000011111_0111011110101101"; -- -0.11670734434656066
	pesos_i(9303) := b"0000000000000000_0000000000000000_0001000110111100_1111111101110000"; -- 0.06929012767350776
	pesos_i(9304) := b"0000000000000000_0000000000000000_0001010010101001_0110000101111001"; -- 0.08070954527066525
	pesos_i(9305) := b"1111111111111111_1111111111111111_1101101101111001_0111001000000111"; -- -0.1426781400557369
	pesos_i(9306) := b"1111111111111111_1111111111111111_1110111110100100_0111101000101111"; -- -0.06389652593952397
	pesos_i(9307) := b"0000000000000000_0000000000000000_0001101111110001_0100101011011111"; -- 0.10915058089275712
	pesos_i(9308) := b"0000000000000000_0000000000000000_0001111001100111_0101010110000111"; -- 0.11876425305532133
	pesos_i(9309) := b"0000000000000000_0000000000000000_0001111010000001_0011101011010100"; -- 0.11915939027109995
	pesos_i(9310) := b"0000000000000000_0000000000000000_0000111111000010_1010110001001011"; -- 0.061564224571738484
	pesos_i(9311) := b"1111111111111111_1111111111111111_1110011100111010_0000010011111101"; -- -0.09677094287524224
	pesos_i(9312) := b"0000000000000000_0000000000000000_0001101111001010_0001100001011100"; -- 0.10855247739406473
	pesos_i(9313) := b"1111111111111111_1111111111111111_1110011111001010_0011111101101000"; -- -0.09457019540846075
	pesos_i(9314) := b"0000000000000000_0000000000000000_0001100010000111_1110011000101100"; -- 0.09582365573720052
	pesos_i(9315) := b"1111111111111111_1111111111111111_1111001111010101_1001000011010010"; -- -0.04752249598377387
	pesos_i(9316) := b"0000000000000000_0000000000000000_0010010011101010_1001001100001010"; -- 0.14420432084205986
	pesos_i(9317) := b"1111111111111111_1111111111111111_1110001011100000_0110100001000100"; -- -0.11376331643020052
	pesos_i(9318) := b"1111111111111111_1111111111111111_1110100101101110_0100001010101110"; -- -0.08816130875899214
	pesos_i(9319) := b"1111111111111111_1111111111111111_1111000101010111_1010011110010110"; -- -0.057256246406928106
	pesos_i(9320) := b"1111111111111111_1111111111111111_1110011111110110_0010111100010101"; -- -0.0938997814948181
	pesos_i(9321) := b"0000000000000000_0000000000000000_0000111100110000_1000001000001111"; -- 0.05933392398471727
	pesos_i(9322) := b"1111111111111111_1111111111111111_1111110001101111_1000110011011000"; -- -0.013922879500381829
	pesos_i(9323) := b"0000000000000000_0000000000000000_0001000100010101_0111110110011101"; -- 0.06673417168187666
	pesos_i(9324) := b"1111111111111111_1111111111111111_1110101011111110_0000001111000001"; -- -0.08206154376427692
	pesos_i(9325) := b"1111111111111111_1111111111111111_1110100001110001_1110111011000000"; -- -0.09201152628665486
	pesos_i(9326) := b"1111111111111111_1111111111111111_1110010100011011_0001101100110101"; -- -0.10505514102857692
	pesos_i(9327) := b"1111111111111111_1111111111111111_1111001101110111_1011010110111100"; -- -0.04895462194701989
	pesos_i(9328) := b"0000000000000000_0000000000000000_0000110000001101_0101000010101000"; -- 0.04707817169192413
	pesos_i(9329) := b"0000000000000000_0000000000000000_0001011101000011_1110011011001011"; -- 0.0908798452519109
	pesos_i(9330) := b"1111111111111111_1111111111111111_1110010010111010_1011011010111110"; -- -0.1065259728394298
	pesos_i(9331) := b"0000000000000000_0000000000000000_0001101111011011_1101100000110010"; -- 0.10882331098149874
	pesos_i(9332) := b"0000000000000000_0000000000000000_0001000000110000_0001111100001111"; -- 0.06323427315628008
	pesos_i(9333) := b"1111111111111111_1111111111111111_1101101010011100_1010101111000010"; -- -0.1460468912413962
	pesos_i(9334) := b"1111111111111111_1111111111111111_1111011000011001_0011100001101110"; -- -0.03867766669724635
	pesos_i(9335) := b"0000000000000000_0000000000000000_0001001000111011_1100001011000011"; -- 0.07122437727350285
	pesos_i(9336) := b"1111111111111111_1111111111111111_1110001001100101_0110110001011111"; -- -0.11563990280763663
	pesos_i(9337) := b"0000000000000000_0000000000000000_0001100100111001_1110011101011000"; -- 0.09853979009370326
	pesos_i(9338) := b"1111111111111111_1111111111111111_1110010111001110_1011111000100110"; -- -0.10231410580124996
	pesos_i(9339) := b"0000000000000000_0000000000000000_0000010001101001_0000111000010101"; -- 0.017228012122214774
	pesos_i(9340) := b"1111111111111111_1111111111111111_1111111101000111_1001101100111101"; -- -0.002813622941455177
	pesos_i(9341) := b"0000000000000000_0000000000000000_0000101011000010_0000101000101100"; -- 0.0420233113986068
	pesos_i(9342) := b"1111111111111111_1111111111111111_1111010000101011_0111111111001011"; -- -0.04621125510320409
	pesos_i(9343) := b"0000000000000000_0000000000000000_0001011011011001_0101010110111100"; -- 0.08925376734507441
	pesos_i(9344) := b"1111111111111111_1111111111111111_1111000010011110_1001110011101101"; -- -0.06007975770893293
	pesos_i(9345) := b"1111111111111111_1111111111111111_1111000010011111_1010010110001110"; -- -0.06006398481378493
	pesos_i(9346) := b"0000000000000000_0000000000000000_0001100011010100_1110011101100000"; -- 0.09699865440237754
	pesos_i(9347) := b"1111111111111111_1111111111111111_1110101011011111_1010000111100001"; -- -0.08252514124745688
	pesos_i(9348) := b"1111111111111111_1111111111111111_1111000000101100_1000110101010011"; -- -0.061820189716951794
	pesos_i(9349) := b"0000000000000000_0000000000000000_0010101001000110_0010011111010011"; -- 0.16513298894726958
	pesos_i(9350) := b"0000000000000000_0000000000000000_0001110000011011_1011101111111011"; -- 0.10979819183440112
	pesos_i(9351) := b"1111111111111111_1111111111111111_1101111000000110_0001000000000011"; -- -0.13271999284747857
	pesos_i(9352) := b"0000000000000000_0000000000000000_0001011011110100_0000010100101100"; -- 0.089660952715521
	pesos_i(9353) := b"1111111111111111_1111111111111111_1110001110111010_1100100010001110"; -- -0.11043116132335924
	pesos_i(9354) := b"0000000000000000_0000000000000000_0000111011011111_0110000011111110"; -- 0.05809599110674222
	pesos_i(9355) := b"0000000000000000_0000000000000000_0000010100000101_0101100101100101"; -- 0.01961287217444475
	pesos_i(9356) := b"1111111111111111_1111111111111111_1111001010100100_0110101001110101"; -- -0.05217871330340597
	pesos_i(9357) := b"0000000000000000_0000000000000000_0010011011100101_1101110111000100"; -- 0.15194498092702804
	pesos_i(9358) := b"1111111111111111_1111111111111111_1110111010111110_1101100000000011"; -- -0.0674004547399329
	pesos_i(9359) := b"0000000000000000_0000000000000000_0001101011011100_1100110101101100"; -- 0.10493167779392333
	pesos_i(9360) := b"1111111111111111_1111111111111111_1111110101111001_0110011110101000"; -- -0.00986625801867228
	pesos_i(9361) := b"1111111111111111_1111111111111111_1111010001001000_1000110111110110"; -- -0.04576790570362712
	pesos_i(9362) := b"0000000000000000_0000000000000000_0001100101100010_0000001100000110"; -- 0.099151791471969
	pesos_i(9363) := b"0000000000000000_0000000000000000_0001011100001011_1001001101101100"; -- 0.09002038360460443
	pesos_i(9364) := b"0000000000000000_0000000000000000_0001001101110101_0010001100000110"; -- 0.07600611577917175
	pesos_i(9365) := b"0000000000000000_0000000000000000_0001010010101010_0000010100000111"; -- 0.0807192937453899
	pesos_i(9366) := b"1111111111111111_1111111111111111_1111101101110110_0010110110000000"; -- -0.017728000805547994
	pesos_i(9367) := b"0000000000000000_0000000000000000_0010010011101100_0001101111110011"; -- 0.14422774016466455
	pesos_i(9368) := b"1111111111111111_1111111111111111_1110100001111011_1100100111101101"; -- -0.09186113316594273
	pesos_i(9369) := b"1111111111111111_1111111111111111_1111011000110001_0010000001110101"; -- -0.038312884801081304
	pesos_i(9370) := b"0000000000000000_0000000000000000_0001101100100110_0100111101011101"; -- 0.10605331437737109
	pesos_i(9371) := b"1111111111111111_1111111111111111_1110111011001011_0101011110111001"; -- -0.06720973714160675
	pesos_i(9372) := b"1111111111111111_1111111111111111_1101101000110011_1011001000010001"; -- -0.147648688248433
	pesos_i(9373) := b"0000000000000000_0000000000000000_0001100010110010_0111011111101101"; -- 0.09647321266915705
	pesos_i(9374) := b"1111111111111111_1111111111111111_1111110010100111_0001011110101010"; -- -0.013075371806882717
	pesos_i(9375) := b"0000000000000000_0000000000000000_0010000001011100_0101010110100101"; -- 0.12640891349207498
	pesos_i(9376) := b"0000000000000000_0000000000000000_0000001110111010_0001001010000000"; -- 0.014557987411361734
	pesos_i(9377) := b"1111111111111111_1111111111111111_1111111001001111_0000011000100001"; -- -0.006606690446654932
	pesos_i(9378) := b"1111111111111111_1111111111111111_1110000110010110_0111011010101010"; -- -0.11879785871929506
	pesos_i(9379) := b"0000000000000000_0000000000000000_0000100011001101_0111011111100010"; -- 0.03438519734112952
	pesos_i(9380) := b"0000000000000000_0000000000000000_0000100000110101_1010011010001001"; -- 0.03206864199960313
	pesos_i(9381) := b"1111111111111111_1111111111111111_1101100101000100_1011001001100110"; -- -0.15129551906450636
	pesos_i(9382) := b"1111111111111111_1111111111111111_1110101101101101_0010100011010111"; -- -0.0803656078544124
	pesos_i(9383) := b"1111111111111111_1111111111111111_1111010000100101_1110010100101000"; -- -0.046296766021307674
	pesos_i(9384) := b"1111111111111111_1111111111111111_1110100000101110_1001111100010110"; -- -0.09303861334965854
	pesos_i(9385) := b"1111111111111111_1111111111111111_1111100001010111_1001100010010011"; -- -0.029913391233830734
	pesos_i(9386) := b"0000000000000000_0000000000000000_0001010011011000_0000100111101010"; -- 0.08142148943907442
	pesos_i(9387) := b"0000000000000000_0000000000000000_0001011101110000_1001010101110000"; -- 0.09156164159816813
	pesos_i(9388) := b"1111111111111111_1111111111111111_1111110011010001_1010011111000010"; -- -0.012425913952825262
	pesos_i(9389) := b"0000000000000000_0000000000000000_0000110100101110_0100000100011111"; -- 0.051487035769699464
	pesos_i(9390) := b"1111111111111111_1111111111111111_1111000111011001_1100000011101001"; -- -0.05527109454125063
	pesos_i(9391) := b"0000000000000000_0000000000000000_0000001100110100_0010000011110010"; -- 0.012514170709300996
	pesos_i(9392) := b"0000000000000000_0000000000000000_0001101101100100_0111011001100011"; -- 0.10700168540012611
	pesos_i(9393) := b"0000000000000000_0000000000000000_0001101111001100_0101101101001011"; -- 0.10858698456992041
	pesos_i(9394) := b"1111111111111111_1111111111111111_1110100100110001_1000110100001010"; -- -0.08908766275202024
	pesos_i(9395) := b"1111111111111111_1111111111111111_1101111000000110_1100011111001111"; -- -0.1327090378524571
	pesos_i(9396) := b"1111111111111111_1111111111111111_1110110111111010_0111110011101101"; -- -0.07039660655830356
	pesos_i(9397) := b"1111111111111111_1111111111111111_1110100010111000_1010110011000001"; -- -0.09093208596451766
	pesos_i(9398) := b"0000000000000000_0000000000000000_0000011101100001_0100010011100001"; -- 0.02882795807454146
	pesos_i(9399) := b"0000000000000000_0000000000000000_0010100001010110_0000100001111100"; -- 0.15756276156969823
	pesos_i(9400) := b"1111111111111111_1111111111111111_1111111111011110_1001010001010101"; -- -0.0005099576535838782
	pesos_i(9401) := b"1111111111111111_1111111111111111_1111000111111000_0101010010010001"; -- -0.05480452979820174
	pesos_i(9402) := b"1111111111111111_1111111111111111_1101110011011001_0100110001010010"; -- -0.13730929380806556
	pesos_i(9403) := b"1111111111111111_1111111111111111_1110100111101011_0000010101100100"; -- -0.08625761333490937
	pesos_i(9404) := b"1111111111111111_1111111111111111_1111010100000111_1010001010011000"; -- -0.04285224718848723
	pesos_i(9405) := b"1111111111111111_1111111111111111_1111000010110101_1100100100100111"; -- -0.0597261695692517
	pesos_i(9406) := b"0000000000000000_0000000000000000_0000001011010110_1000011011001111"; -- 0.01108591605614389
	pesos_i(9407) := b"0000000000000000_0000000000000000_0010001011101110_0001100000010010"; -- 0.13644552648482206
	pesos_i(9408) := b"1111111111111111_1111111111111111_1111000010100110_0100001101001011"; -- -0.05996303006990167
	pesos_i(9409) := b"1111111111111111_1111111111111111_1111100110101010_1111100010010100"; -- -0.024734939489408466
	pesos_i(9410) := b"1111111111111111_1111111111111111_1110110010110010_1100001001001001"; -- -0.07539735529102981
	pesos_i(9411) := b"1111111111111111_1111111111111111_1111100001111000_1111111111010111"; -- -0.029403696127278327
	pesos_i(9412) := b"1111111111111111_1111111111111111_1111100101100110_0101010010010011"; -- -0.025782312556547095
	pesos_i(9413) := b"1111111111111111_1111111111111111_1111000101100100_0000010111000010"; -- -0.05706752786084948
	pesos_i(9414) := b"0000000000000000_0000000000000000_0001000110110111_1110111100011111"; -- 0.06921286101525374
	pesos_i(9415) := b"0000000000000000_0000000000000000_0001011111000111_1011101001110010"; -- 0.09289136210834598
	pesos_i(9416) := b"1111111111111111_1111111111111111_1111000100001001_1101100011000100"; -- -0.058443500751163106
	pesos_i(9417) := b"0000000000000000_0000000000000000_0001111001011000_0001101101111110"; -- 0.1185319121791468
	pesos_i(9418) := b"0000000000000000_0000000000000000_0000000010101110_1011110011011011"; -- 0.0026662860402911466
	pesos_i(9419) := b"0000000000000000_0000000000000000_0001010010010000_0011100101111111"; -- 0.08032569275141467
	pesos_i(9420) := b"0000000000000000_0000000000000000_0010001000110000_1011101101000100"; -- 0.13355608383408138
	pesos_i(9421) := b"0000000000000000_0000000000000000_0001110011001101_0100001100010110"; -- 0.11250705043859854
	pesos_i(9422) := b"0000000000000000_0000000000000000_0001110011101101_0100101100000010"; -- 0.11299580378796838
	pesos_i(9423) := b"0000000000000000_0000000000000000_0010000111110111_0101101101111011"; -- 0.13268062354953963
	pesos_i(9424) := b"1111111111111111_1111111111111111_1101111101011110_1010100010100001"; -- -0.12746187280820612
	pesos_i(9425) := b"1111111111111111_1111111111111111_1101110010000000_0011010110010101"; -- -0.13866868116594339
	pesos_i(9426) := b"1111111111111111_1111111111111111_1111010010111000_1111001011000010"; -- -0.044052913430367234
	pesos_i(9427) := b"1111111111111111_1111111111111111_1111110001110101_0011101111001001"; -- -0.013836158104448215
	pesos_i(9428) := b"0000000000000000_0000000000000000_0000011111100000_0010111111101010"; -- 0.030764574654317905
	pesos_i(9429) := b"1111111111111111_1111111111111111_1110101000101111_1111111001010001"; -- -0.08520517855299532
	pesos_i(9430) := b"0000000000000000_0000000000000000_0000010100010111_1011101001000010"; -- 0.01989330392689041
	pesos_i(9431) := b"1111111111111111_1111111111111111_1111111100110111_1001010100110001"; -- -0.0030581240176435
	pesos_i(9432) := b"0000000000000000_0000000000000000_0000010101101111_1100101000101100"; -- 0.021237025863091227
	pesos_i(9433) := b"1111111111111111_1111111111111111_1111101000000111_0110100010111100"; -- -0.02332444582840463
	pesos_i(9434) := b"0000000000000000_0000000000000000_0010100101010100_1011010000100111"; -- 0.161448726108641
	pesos_i(9435) := b"1111111111111111_1111111111111111_1111100100011100_0101011000100000"; -- -0.0269113704202712
	pesos_i(9436) := b"1111111111111111_1111111111111111_1111000100110111_0010010110110100"; -- -0.05775226939779824
	pesos_i(9437) := b"1111111111111111_1111111111111111_1110000000010110_0001011101101100"; -- -0.12466291065997692
	pesos_i(9438) := b"1111111111111111_1111111111111111_1101110000010111_0001011000110011"; -- -0.1402727247584431
	pesos_i(9439) := b"1111111111111111_1111111111111111_1110110001100011_1111111110010000"; -- -0.07659914714797667
	pesos_i(9440) := b"1111111111111111_1111111111111111_1111001011001101_1010010100110000"; -- -0.05154960222179417
	pesos_i(9441) := b"1111111111111111_1111111111111111_1101110011101001_0110110100110110"; -- -0.13706319262008818
	pesos_i(9442) := b"0000000000000000_0000000000000000_0000011011001100_0110000101001010"; -- 0.026556091749442515
	pesos_i(9443) := b"0000000000000000_0000000000000000_0001101111001110_0110001100000111"; -- 0.10861796296741999
	pesos_i(9444) := b"0000000000000000_0000000000000000_0000100000110111_0111100111000101"; -- 0.032096491356258444
	pesos_i(9445) := b"1111111111111111_1111111111111111_1110110000101111_0100100010101001"; -- -0.0774035060499225
	pesos_i(9446) := b"1111111111111111_1111111111111111_1111101101100011_1011100000110101"; -- -0.018009650222837483
	pesos_i(9447) := b"0000000000000000_0000000000000000_0000010010110101_1110011110100000"; -- 0.018400646734266567
	pesos_i(9448) := b"0000000000000000_0000000000000000_0001001010100101_1110010110000000"; -- 0.0728438793984836
	pesos_i(9449) := b"1111111111111111_1111111111111111_1110101010010010_0101010000001110"; -- -0.08370470674741097
	pesos_i(9450) := b"0000000000000000_0000000000000000_0010001000001010_1010011011001110"; -- 0.1329750302069923
	pesos_i(9451) := b"1111111111111111_1111111111111111_1110100110111110_0001111010110011"; -- -0.08694275026038761
	pesos_i(9452) := b"0000000000000000_0000000000000000_0001100001101100_0100101101111000"; -- 0.0954024474263763
	pesos_i(9453) := b"1111111111111111_1111111111111111_1110101111011100_1101011000000000"; -- -0.07866156105644193
	pesos_i(9454) := b"0000000000000000_0000000000000000_0000011111100010_0000010101100010"; -- 0.030792557267523973
	pesos_i(9455) := b"0000000000000000_0000000000000000_0000111100000011_1000010111001101"; -- 0.05864750147362216
	pesos_i(9456) := b"1111111111111111_1111111111111111_1111110001100101_0010101110000101"; -- -0.014081268344693816
	pesos_i(9457) := b"0000000000000000_0000000000000000_0000011100000100_1011000001010001"; -- 0.027415294521985448
	pesos_i(9458) := b"0000000000000000_0000000000000000_0000100001100011_0001011101101001"; -- 0.032762015504172105
	pesos_i(9459) := b"0000000000000000_0000000000000000_0001101111101011_1111100101111100"; -- 0.10906943589401319
	pesos_i(9460) := b"1111111111111111_1111111111111111_1110110101111001_1010001010010000"; -- -0.07236274700908815
	pesos_i(9461) := b"1111111111111111_1111111111111111_1110010101111101_0110011010101100"; -- -0.10355528156370682
	pesos_i(9462) := b"1111111111111111_1111111111111111_1101101100100100_1111011111000001"; -- -0.14396716631260215
	pesos_i(9463) := b"1111111111111111_1111111111111111_1111010000100001_1001011000100100"; -- -0.04636251090810955
	pesos_i(9464) := b"1111111111111111_1111111111111111_1110000101011101_1101010111101010"; -- -0.11966193226323568
	pesos_i(9465) := b"0000000000000000_0000000000000000_0000110100110000_0001010111100010"; -- 0.051514976276361785
	pesos_i(9466) := b"0000000000000000_0000000000000000_0000111110101010_0110000111101111"; -- 0.06119358134166755
	pesos_i(9467) := b"1111111111111111_1111111111111111_1110011111101100_1011001110010011"; -- -0.09404447229173134
	pesos_i(9468) := b"0000000000000000_0000000000000000_0000101011000011_0110110111111110"; -- 0.04204451989832828
	pesos_i(9469) := b"1111111111111111_1111111111111111_1111000101101000_0001110100100000"; -- -0.05700510003938203
	pesos_i(9470) := b"1111111111111111_1111111111111111_1110111111110101_0100101001111000"; -- -0.06266340802732234
	pesos_i(9471) := b"0000000000000000_0000000000000000_0001101100001101_0011011011100011"; -- 0.10567038571474147
	pesos_i(9472) := b"1111111111111111_1111111111111111_1110100010111011_1111111001111111"; -- -0.09088143735093987
	pesos_i(9473) := b"1111111111111111_1111111111111111_1111110000010100_0010010110001010"; -- -0.01531758664585097
	pesos_i(9474) := b"1111111111111111_1111111111111111_1101111010011110_0101111010000001"; -- -0.13039597843565925
	pesos_i(9475) := b"0000000000000000_0000000000000000_0000101101101110_0000001011010000"; -- 0.04464738435575233
	pesos_i(9476) := b"1111111111111111_1111111111111111_1111101000010110_0000000101110100"; -- -0.02310172007051638
	pesos_i(9477) := b"1111111111111111_1111111111111111_1101111101111111_0111111101010011"; -- -0.1269607946783124
	pesos_i(9478) := b"1111111111111111_1111111111111111_1111111001000100_0110111101101110"; -- -0.006768260551288201
	pesos_i(9479) := b"1111111111111111_1111111111111111_1110110101011111_1011100100010111"; -- -0.07275813273664195
	pesos_i(9480) := b"0000000000000000_0000000000000000_0001110101101000_1011000010101110"; -- 0.11487869499313827
	pesos_i(9481) := b"1111111111111111_1111111111111111_1111110110000101_0101101101000110"; -- -0.009683890754265359
	pesos_i(9482) := b"0000000000000000_0000000000000000_0001010001001001_1010000011101100"; -- 0.07924848321594292
	pesos_i(9483) := b"0000000000000000_0000000000000000_0001111010100011_0000110100010000"; -- 0.11967546119168024
	pesos_i(9484) := b"0000000000000000_0000000000000000_0001100011100100_1001111101111011"; -- 0.09723850957336441
	pesos_i(9485) := b"0000000000000000_0000000000000000_0001100000011010_1001011111111101"; -- 0.09415578771732798
	pesos_i(9486) := b"1111111111111111_1111111111111111_1101111000100010_0000110111100001"; -- -0.1322928739630522
	pesos_i(9487) := b"1111111111111111_1111111111111111_1110111100010000_0110001001011100"; -- -0.06615624676475769
	pesos_i(9488) := b"1111111111111111_1111111111111111_1111011110111001_0111101001010011"; -- -0.03232608302256627
	pesos_i(9489) := b"1111111111111111_1111111111111111_1110010011100101_1110100100100010"; -- -0.1058668414874286
	pesos_i(9490) := b"1111111111111111_1111111111111111_1110010000000100_1011111000010111"; -- -0.10930263456287821
	pesos_i(9491) := b"0000000000000000_0000000000000000_0000100010110111_0111000001000011"; -- 0.03404904972850652
	pesos_i(9492) := b"1111111111111111_1111111111111111_1101110011000010_0011111011100101"; -- -0.13766104611760518
	pesos_i(9493) := b"1111111111111111_1111111111111111_1111100100110010_1010100001000101"; -- -0.026570780832058025
	pesos_i(9494) := b"1111111111111111_1111111111111111_1101101101000010_1011011000001110"; -- -0.14351331860122676
	pesos_i(9495) := b"1111111111111111_1111111111111111_1110100111001010_0101111000000001"; -- -0.08675587157797068
	pesos_i(9496) := b"1111111111111111_1111111111111111_1101010110011110_1010011001010111"; -- -0.16554794671681253
	pesos_i(9497) := b"1111111111111111_1111111111111111_1111100110001011_1100100011111111"; -- -0.02521079807517392
	pesos_i(9498) := b"0000000000000000_0000000000000000_0010000100010100_0111001001010100"; -- 0.12921824024893855
	pesos_i(9499) := b"1111111111111111_1111111111111111_1111100011000000_0111000110001011"; -- -0.02831354492394731
	pesos_i(9500) := b"0000000000000000_0000000000000000_0001101011011000_0111000110110001"; -- 0.10486517499419616
	pesos_i(9501) := b"0000000000000000_0000000000000000_0000101010100001_0111011011111010"; -- 0.04152625659804057
	pesos_i(9502) := b"0000000000000000_0000000000000000_0000111000000110_1001000011001010"; -- 0.05478768282424649
	pesos_i(9503) := b"1111111111111111_1111111111111111_1111101010010100_1110010101111001"; -- -0.02116552157991216
	pesos_i(9504) := b"0000000000000000_0000000000000000_0010000100100001_0111000011111101"; -- 0.12941652474569232
	pesos_i(9505) := b"1111111111111111_1111111111111111_1111010100000100_0100011110001001"; -- -0.04290345097629714
	pesos_i(9506) := b"1111111111111111_1111111111111111_1110101110110100_1011101000110001"; -- -0.07927357002348963
	pesos_i(9507) := b"1111111111111111_1111111111111111_1110000010011101_0110101101111000"; -- -0.12259796454197774
	pesos_i(9508) := b"0000000000000000_0000000000000000_0000011010000010_0001001010010100"; -- 0.025422250003759177
	pesos_i(9509) := b"1111111111111111_1111111111111111_1110000011001111_1111111001010001"; -- -0.1218262721336549
	pesos_i(9510) := b"1111111111111111_1111111111111111_1110110010110001_0110011000100011"; -- -0.07541810647932544
	pesos_i(9511) := b"1111111111111111_1111111111111111_1111010010010100_0101011010101101"; -- -0.04461153285647374
	pesos_i(9512) := b"0000000000000000_0000000000000000_0010000011000110_0000111101100101"; -- 0.12802215788000185
	pesos_i(9513) := b"0000000000000000_0000000000000000_0001000100100000_0101011101001010"; -- 0.06689973418816429
	pesos_i(9514) := b"0000000000000000_0000000000000000_0000010010000011_1110110100001110"; -- 0.017638030906984438
	pesos_i(9515) := b"1111111111111111_1111111111111111_1111010010000000_1100101010110000"; -- -0.044909793982495026
	pesos_i(9516) := b"1111111111111111_1111111111111111_1110011011011101_1001100111110101"; -- -0.09818113106150685
	pesos_i(9517) := b"1111111111111111_1111111111111111_1101110111011010_1111110011001111"; -- -0.13337726545418627
	pesos_i(9518) := b"1111111111111111_1111111111111111_1101110110101100_1000010000011100"; -- -0.13408636385263384
	pesos_i(9519) := b"0000000000000000_0000000000000000_0001001011011010_1010101011100010"; -- 0.07364910139201233
	pesos_i(9520) := b"0000000000000000_0000000000000000_0010010100010110_1000101101010101"; -- 0.14487524827922524
	pesos_i(9521) := b"0000000000000000_0000000000000000_0010000110110111_1011001010100110"; -- 0.1317092566906862
	pesos_i(9522) := b"1111111111111111_1111111111111111_1110001011010100_0110111011111001"; -- -0.11394602222469873
	pesos_i(9523) := b"1111111111111111_1111111111111111_1111100110111000_1001100000100111"; -- -0.02452706376467631
	pesos_i(9524) := b"1111111111111111_1111111111111111_1111010010110101_0111010010001101"; -- -0.04410621221235436
	pesos_i(9525) := b"0000000000000000_0000000000000000_0000011111010110_1101011101111111"; -- 0.03062197535429244
	pesos_i(9526) := b"0000000000000000_0000000000000000_0001111100001101_1001111100110111"; -- 0.12130160410193738
	pesos_i(9527) := b"0000000000000000_0000000000000000_0010000110101110_1000110101000111"; -- 0.13156970012299082
	pesos_i(9528) := b"1111111111111111_1111111111111111_1111101010110011_0000010100100111"; -- -0.020705869563019594
	pesos_i(9529) := b"0000000000000000_0000000000000000_0000011101011101_1000100000011111"; -- 0.028770930826465733
	pesos_i(9530) := b"0000000000000000_0000000000000000_0001010010001000_1001011110110010"; -- 0.08020923701881866
	pesos_i(9531) := b"1111111111111111_1111111111111111_1101111010110011_0000010110001110"; -- -0.13008084560270222
	pesos_i(9532) := b"1111111111111111_1111111111111111_1111111010000110_1110011111000101"; -- -0.005754007775172294
	pesos_i(9533) := b"0000000000000000_0000000000000000_0001111011101101_0011010110100000"; -- 0.12080702919958021
	pesos_i(9534) := b"1111111111111111_1111111111111111_1111110111010111_0110110011010000"; -- -0.008431624515613906
	pesos_i(9535) := b"0000000000000000_0000000000000000_0000100110000111_1010101101010000"; -- 0.0372263975819118
	pesos_i(9536) := b"0000000000000000_0000000000000000_0000001001001010_0110111001011010"; -- 0.008948227964799767
	pesos_i(9537) := b"0000000000000000_0000000000000000_0001111100101010_0000100100010110"; -- 0.12173516076338985
	pesos_i(9538) := b"1111111111111111_1111111111111111_1111101010011011_0100000100110110"; -- -0.021068500816066076
	pesos_i(9539) := b"1111111111111111_1111111111111111_1110000110000111_0001011011111110"; -- -0.11903244299320498
	pesos_i(9540) := b"0000000000000000_0000000000000000_0000010011000001_1101000111010111"; -- 0.018582453824239075
	pesos_i(9541) := b"1111111111111111_1111111111111111_1110011000111111_1000001000011011"; -- -0.1005934413948841
	pesos_i(9542) := b"1111111111111111_1111111111111111_1110111001010101_0010111010001101"; -- -0.06901272833243659
	pesos_i(9543) := b"0000000000000000_0000000000000000_0001110011100101_1100010010010010"; -- 0.11288097930077365
	pesos_i(9544) := b"0000000000000000_0000000000000000_0000001110000000_1110011111101000"; -- 0.013685697580032609
	pesos_i(9545) := b"1111111111111111_1111111111111111_1111110110001101_0010101110111000"; -- -0.009564654844398198
	pesos_i(9546) := b"0000000000000000_0000000000000000_0001101001100100_1111100000000000"; -- 0.10310316086682912
	pesos_i(9547) := b"0000000000000000_0000000000000000_0000001010101101_1011010001001000"; -- 0.010463016138327452
	pesos_i(9548) := b"0000000000000000_0000000000000000_0000010010101011_1010011010001010"; -- 0.018244179356056142
	pesos_i(9549) := b"0000000000000000_0000000000000000_0000000000001011_0110010111100100"; -- 0.00017391972913662768
	pesos_i(9550) := b"0000000000000000_0000000000000000_0010001110101111_1010110111110100"; -- 0.13939940639928797
	pesos_i(9551) := b"0000000000000000_0000000000000000_0001101100000011_0110010001010000"; -- 0.10552050552106637
	pesos_i(9552) := b"1111111111111111_1111111111111111_1110000101011111_0001111101100000"; -- -0.11964229486081818
	pesos_i(9553) := b"0000000000000000_0000000000000000_0000101101011111_0111011101111011"; -- 0.04442545652635068
	pesos_i(9554) := b"1111111111111111_1111111111111111_1111101100001000_1010000111011010"; -- -0.019399532588702716
	pesos_i(9555) := b"0000000000000000_0000000000000000_0001101111010110_1011000001011110"; -- 0.10874464316367108
	pesos_i(9556) := b"1111111111111111_1111111111111111_1111001100101000_1110011000010011"; -- -0.05015718503359846
	pesos_i(9557) := b"1111111111111111_1111111111111111_1101101011010100_1011011000011111"; -- -0.14519178148426615
	pesos_i(9558) := b"0000000000000000_0000000000000000_0001101100100001_0100100000111011"; -- 0.10597659523515812
	pesos_i(9559) := b"0000000000000000_0000000000000000_0000010111011110_1001010010110100"; -- 0.022927564566022633
	pesos_i(9560) := b"1111111111111111_1111111111111111_1111111110111001_0010000010011101"; -- -0.0010814300155056766
	pesos_i(9561) := b"1111111111111111_1111111111111111_1110101110100010_0000101101010000"; -- -0.07955865178966555
	pesos_i(9562) := b"1111111111111111_1111111111111111_1111011010111010_0110010100111010"; -- -0.03621833164337747
	pesos_i(9563) := b"1111111111111111_1111111111111111_1111100111110011_1000000111100011"; -- -0.023628122509280976
	pesos_i(9564) := b"0000000000000000_0000000000000000_0000001001011011_0101100010001000"; -- 0.009206326585430857
	pesos_i(9565) := b"1111111111111111_1111111111111111_1101110001001000_0001001001101010"; -- -0.13952526963375983
	pesos_i(9566) := b"0000000000000000_0000000000000000_0010000111110101_1001101001111001"; -- 0.1326538606596843
	pesos_i(9567) := b"1111111111111111_1111111111111111_1110110001001110_1001100111001111"; -- -0.07692564665044681
	pesos_i(9568) := b"0000000000000000_0000000000000000_0000000100111100_0000011011110000"; -- 0.004822190805177755
	pesos_i(9569) := b"0000000000000000_0000000000000000_0000000001011001_0101000000110110"; -- 0.001362813067188789
	pesos_i(9570) := b"0000000000000000_0000000000000000_0000010100010111_1010001001010010"; -- 0.01989187713323095
	pesos_i(9571) := b"0000000000000000_0000000000000000_0000010010010010_0010110111101011"; -- 0.017855520240189427
	pesos_i(9572) := b"0000000000000000_0000000000000000_0000100100011010_0100101101110000"; -- 0.03555747495522952
	pesos_i(9573) := b"1111111111111111_1111111111111111_1111001010001101_0110111110010100"; -- -0.052529360260714315
	pesos_i(9574) := b"1111111111111111_1111111111111111_1101111011100110_1100111000011011"; -- -0.12929069358585354
	pesos_i(9575) := b"1111111111111111_1111111111111111_1111101101001111_0010101000110101"; -- -0.018323289845999003
	pesos_i(9576) := b"0000000000000000_0000000000000000_0000100111111101_1001101011111110"; -- 0.03902596190734697
	pesos_i(9577) := b"0000000000000000_0000000000000000_0001100010101101_0100011001011110"; -- 0.09639396477471388
	pesos_i(9578) := b"0000000000000000_0000000000000000_0010000110111100_1100101101111000"; -- 0.13178702997450867
	pesos_i(9579) := b"0000000000000000_0000000000000000_0001110000111100_0000110001010011"; -- 0.11029126192721925
	pesos_i(9580) := b"1111111111111111_1111111111111111_1111100000101001_1010110001000010"; -- -0.030614122248201932
	pesos_i(9581) := b"0000000000000000_0000000000000000_0000011010001101_1010011100011110"; -- 0.02559895012085262
	pesos_i(9582) := b"0000000000000000_0000000000000000_0000110100000010_1011001011001100"; -- 0.050822424636073546
	pesos_i(9583) := b"1111111111111111_1111111111111111_1111100000101011_0000001000001101"; -- -0.030593749765508733
	pesos_i(9584) := b"1111111111111111_1111111111111111_1101110100100110_1111111110101101"; -- -0.1361236765875426
	pesos_i(9585) := b"1111111111111111_1111111111111111_1110011010000110_1100100101001011"; -- -0.09950582436562662
	pesos_i(9586) := b"1111111111111111_1111111111111111_1111000011101001_1000010010101010"; -- -0.0589367946454048
	pesos_i(9587) := b"1111111111111111_1111111111111111_1111100010100011_0001110110111101"; -- -0.028761044764424964
	pesos_i(9588) := b"1111111111111111_1111111111111111_1110101111001000_0011110000001100"; -- -0.07897591316160862
	pesos_i(9589) := b"1111111111111111_1111111111111111_1110101100010111_0000001000110001"; -- -0.08168016731088162
	pesos_i(9590) := b"1111111111111111_1111111111111111_1111111000111000_1001010111101100"; -- -0.0069490717448337175
	pesos_i(9591) := b"0000000000000000_0000000000000000_0001111110101110_0011001001000111"; -- 0.12375177610435603
	pesos_i(9592) := b"1111111111111111_1111111111111111_1111101101100010_1101010100101110"; -- -0.01802318209259646
	pesos_i(9593) := b"1111111111111111_1111111111111111_1111111111110011_0010011110001011"; -- -0.0001960072634708341
	pesos_i(9594) := b"1111111111111111_1111111111111111_1110110001110011_0011001100001010"; -- -0.07636719699946128
	pesos_i(9595) := b"0000000000000000_0000000000000000_0001110110001101_0111111001100000"; -- 0.11544027189545389
	pesos_i(9596) := b"0000000000000000_0000000000000000_0001011101111101_0000111001100111"; -- 0.09175195700401241
	pesos_i(9597) := b"0000000000000000_0000000000000000_0001101101101010_1101100110101101"; -- 0.10709915614894978
	pesos_i(9598) := b"1111111111111111_1111111111111111_1110110100110111_0010011110001110"; -- -0.07337715888259501
	pesos_i(9599) := b"1111111111111111_1111111111111111_1111011011110101_1110100100010101"; -- -0.03531020383587673
	pesos_i(9600) := b"1111111111111111_1111111111111111_1111000011100101_0011000111100101"; -- -0.05900276333231558
	pesos_i(9601) := b"0000000000000000_0000000000000000_0000100110110100_1010000101100111"; -- 0.0379124524705775
	pesos_i(9602) := b"1111111111111111_1111111111111111_1111000000111011_1100111010010011"; -- -0.06158741870839053
	pesos_i(9603) := b"0000000000000000_0000000000000000_0000011001111000_1101000110100010"; -- 0.025281049757138557
	pesos_i(9604) := b"0000000000000000_0000000000000000_0001000111110011_1111000000101111"; -- 0.07012845181870855
	pesos_i(9605) := b"1111111111111111_1111111111111111_1111010011110011_0101011110010011"; -- -0.04316189449335993
	pesos_i(9606) := b"1111111111111111_1111111111111111_1111001101111111_1000001001000100"; -- -0.04883561926381223
	pesos_i(9607) := b"1111111111111111_1111111111111111_1110010100110011_1101011001111001"; -- -0.10467776828965028
	pesos_i(9608) := b"1111111111111111_1111111111111111_1101100110100000_1011101000101100"; -- -0.14989124713358126
	pesos_i(9609) := b"0000000000000000_0000000000000000_0010101001101110_0101111000100001"; -- 0.1657465772822901
	pesos_i(9610) := b"1111111111111111_1111111111111111_1111010001011001_0001000110000100"; -- -0.04551592382142579
	pesos_i(9611) := b"0000000000000000_0000000000000000_0000101101100100_0100111010101000"; -- 0.044499317112868884
	pesos_i(9612) := b"1111111111111111_1111111111111111_1101111100010011_0100100000110100"; -- -0.12861202936194693
	pesos_i(9613) := b"0000000000000000_0000000000000000_0000100111111100_1001100000011010"; -- 0.03901053072332577
	pesos_i(9614) := b"1111111111111111_1111111111111111_1101110101101000_1101110000111100"; -- -0.13511870884905225
	pesos_i(9615) := b"0000000000000000_0000000000000000_0001111110010001_0000110001010000"; -- 0.1233070083768355
	pesos_i(9616) := b"1111111111111111_1111111111111111_1111100111011001_1011101100011001"; -- -0.024021440966867934
	pesos_i(9617) := b"1111111111111111_1111111111111111_1111001110100110_0010110111011111"; -- -0.04824555698653998
	pesos_i(9618) := b"1111111111111111_1111111111111111_1111000010010011_0011011000000101"; -- -0.06025373810445648
	pesos_i(9619) := b"0000000000000000_0000000000000000_0000010000011101_0111011000000100"; -- 0.016074539193831477
	pesos_i(9620) := b"0000000000000000_0000000000000000_0000101000110001_1111110000100001"; -- 0.039825208680991306
	pesos_i(9621) := b"1111111111111111_1111111111111111_1110001100000101_0101101001001111"; -- -0.11319957330682917
	pesos_i(9622) := b"1111111111111111_1111111111111111_1110001101111010_1000110111100100"; -- -0.11141122036212678
	pesos_i(9623) := b"1111111111111111_1111111111111111_1110001000101100_1010111100000010"; -- -0.11650568194984885
	pesos_i(9624) := b"0000000000000000_0000000000000000_0001011110111011_0011111101101000"; -- 0.09270092284943111
	pesos_i(9625) := b"0000000000000000_0000000000000000_0001101001101100_0010111110101101"; -- 0.10321329083107927
	pesos_i(9626) := b"0000000000000000_0000000000000000_0000010010010000_1110010100111000"; -- 0.01783592818862567
	pesos_i(9627) := b"1111111111111111_1111111111111111_1110111101111101_0011110000111111"; -- -0.06449531037927714
	pesos_i(9628) := b"0000000000000000_0000000000000000_0000100010000101_0110101011011100"; -- 0.03328578817092573
	pesos_i(9629) := b"0000000000000000_0000000000000000_0001100011011110_1110110101110100"; -- 0.09715160451452427
	pesos_i(9630) := b"0000000000000000_0000000000000000_0001110011110000_1000111011111110"; -- 0.11304563232629039
	pesos_i(9631) := b"1111111111111111_1111111111111111_1111101100101000_1100001101000111"; -- -0.018909258933968696
	pesos_i(9632) := b"1111111111111111_1111111111111111_1111100011010000_1101101011100011"; -- -0.02806312524780631
	pesos_i(9633) := b"1111111111111111_1111111111111111_1110000100100111_1000010111101111"; -- -0.12049067417069356
	pesos_i(9634) := b"0000000000000000_0000000000000000_0000001111110011_0110011011010110"; -- 0.015432765326770344
	pesos_i(9635) := b"1111111111111111_1111111111111111_1111100010100101_0110011100111001"; -- -0.028726147277824354
	pesos_i(9636) := b"1111111111111111_1111111111111111_1111100000100110_1111100011110110"; -- -0.030655326785925585
	pesos_i(9637) := b"1111111111111111_1111111111111111_1110000010001100_1001101100100010"; -- -0.12285452295064268
	pesos_i(9638) := b"0000000000000000_0000000000000000_0010100101100001_1101100111011010"; -- 0.16164933741275014
	pesos_i(9639) := b"0000000000000000_0000000000000000_0000101101100011_1000111000011010"; -- 0.044487840021945606
	pesos_i(9640) := b"0000000000000000_0000000000000000_0010010000010100_1000001010100101"; -- 0.14093796286899685
	pesos_i(9641) := b"0000000000000000_0000000000000000_0000110011011010_1000110001010111"; -- 0.05020978087342282
	pesos_i(9642) := b"1111111111111111_1111111111111111_1111110111100010_0101110011010110"; -- -0.008264730275878165
	pesos_i(9643) := b"0000000000000000_0000000000000000_0000010100101110_0001110000100001"; -- 0.020234831013825495
	pesos_i(9644) := b"1111111111111111_1111111111111111_1101011100110100_1000111100100100"; -- -0.1593542612094539
	pesos_i(9645) := b"0000000000000000_0000000000000000_0010100101110111_0110011111000011"; -- 0.16197823051920504
	pesos_i(9646) := b"1111111111111111_1111111111111111_1110001111010100_0011101000001100"; -- -0.11004292674286235
	pesos_i(9647) := b"1111111111111111_1111111111111111_1111100111001111_0101000101011100"; -- -0.02418033133085012
	pesos_i(9648) := b"0000000000000000_0000000000000000_0000101010101100_0100011000011110"; -- 0.04169119113129277
	pesos_i(9649) := b"1111111111111111_1111111111111111_1110001011110000_1000100010001110"; -- -0.11351725121506907
	pesos_i(9650) := b"1111111111111111_1111111111111111_1101110101000111_0110001111010101"; -- -0.13562942557321195
	pesos_i(9651) := b"1111111111111111_1111111111111111_1101111110101010_1110001001001101"; -- -0.1262987672121579
	pesos_i(9652) := b"1111111111111111_1111111111111111_1111111110010001_0111110110111011"; -- -0.0016862314645361123
	pesos_i(9653) := b"0000000000000000_0000000000000000_0000111010101111_0101010010000000"; -- 0.05736282476902807
	pesos_i(9654) := b"1111111111111111_1111111111111111_1110100100101010_0011101111011111"; -- -0.08919931233081091
	pesos_i(9655) := b"1111111111111111_1111111111111111_1110010100111101_0001011011010010"; -- -0.10453660360267154
	pesos_i(9656) := b"1111111111111111_1111111111111111_1101110111011001_1100100001011011"; -- -0.1333956505755722
	pesos_i(9657) := b"1111111111111111_1111111111111111_1111001100000100_1001001110101001"; -- -0.05071141356781332
	pesos_i(9658) := b"1111111111111111_1111111111111111_1110110111011110_0101100101100000"; -- -0.07082597157497394
	pesos_i(9659) := b"1111111111111111_1111111111111111_1111101010101010_1011010001100010"; -- -0.020832754163642844
	pesos_i(9660) := b"1111111111111111_1111111111111111_1111000010000101_1101111100000001"; -- -0.06045728893240172
	pesos_i(9661) := b"0000000000000000_0000000000000000_0001111000111000_0010101111111010"; -- 0.11804461344417022
	pesos_i(9662) := b"1111111111111111_1111111111111111_1111010011111000_1010000110011101"; -- -0.04308118729583441
	pesos_i(9663) := b"1111111111111111_1111111111111111_1101111100110011_0001001111110001"; -- -0.12812686310117627
	pesos_i(9664) := b"0000000000000000_0000000000000000_0001010010111001_1111000100110011"; -- 0.080962252575826
	pesos_i(9665) := b"1111111111111111_1111111111111111_1110110111001111_1000100000010101"; -- -0.0710520695613315
	pesos_i(9666) := b"0000000000000000_0000000000000000_0001010010111100_1110110011111011"; -- 0.08100777750530178
	pesos_i(9667) := b"0000000000000000_0000000000000000_0000110000101111_0101100100011011"; -- 0.04759747419191107
	pesos_i(9668) := b"1111111111111111_1111111111111111_1110110000000010_0001110000001010"; -- -0.07809281108229903
	pesos_i(9669) := b"1111111111111111_1111111111111111_1111111111001101_0011111101010011"; -- -0.0007744238734922761
	pesos_i(9670) := b"1111111111111111_1111111111111111_1110101010010101_1101011101010000"; -- -0.08365110673806608
	pesos_i(9671) := b"1111111111111111_1111111111111111_1111101010000110_1101110110000000"; -- -0.02137961972891259
	pesos_i(9672) := b"1111111111111111_1111111111111111_1110100000001000_0010001000100001"; -- -0.09362589551270792
	pesos_i(9673) := b"1111111111111111_1111111111111111_1110101000010110_1010100110111101"; -- -0.08559168951788697
	pesos_i(9674) := b"0000000000000000_0000000000000000_0000000001011111_0100111001010110"; -- 0.0014542540321818335
	pesos_i(9675) := b"0000000000000000_0000000000000000_0001011000001010_0100001100111001"; -- 0.08609409467074998
	pesos_i(9676) := b"0000000000000000_0000000000000000_0001001100010111_1010010110111010"; -- 0.0745795801874995
	pesos_i(9677) := b"0000000000000000_0000000000000000_0010100001110000_0010001101100011"; -- 0.1579610936353199
	pesos_i(9678) := b"0000000000000000_0000000000000000_0000011000011011_0100000111101111"; -- 0.023853417143723722
	pesos_i(9679) := b"1111111111111111_1111111111111111_1110101000000100_0111011010011000"; -- -0.08586939606316431
	pesos_i(9680) := b"1111111111111111_1111111111111111_1110011111100000_1111011101100100"; -- -0.09422353571208991
	pesos_i(9681) := b"1111111111111111_1111111111111111_1110000011101011_1010011110011110"; -- -0.1214041937707705
	pesos_i(9682) := b"1111111111111111_1111111111111111_1111010010101110_1001111100011101"; -- -0.04421048687986764
	pesos_i(9683) := b"1111111111111111_1111111111111111_1110100100000100_0100100000000011"; -- -0.08977842267512878
	pesos_i(9684) := b"1111111111111111_1111111111111111_1110000111011101_0110110000100110"; -- -0.11771511144571475
	pesos_i(9685) := b"0000000000000000_0000000000000000_0001110011001111_0000100010010101"; -- 0.11253408084532712
	pesos_i(9686) := b"0000000000000000_0000000000000000_0001000100001111_0000110101111110"; -- 0.0666359360301598
	pesos_i(9687) := b"1111111111111111_1111111111111111_1101111111101011_0011011100001110"; -- -0.12531715304187954
	pesos_i(9688) := b"1111111111111111_1111111111111111_1111000000011000_1100110111001000"; -- -0.06212152357581714
	pesos_i(9689) := b"1111111111111111_1111111111111111_1110000000110101_0010001001010110"; -- -0.12418923753651323
	pesos_i(9690) := b"1111111111111111_1111111111111111_1110010011110010_0110100100010001"; -- -0.10567611049946213
	pesos_i(9691) := b"0000000000000000_0000000000000000_0001000011111110_0000011101101100"; -- 0.0663761746952123
	pesos_i(9692) := b"0000000000000000_0000000000000000_0000101001111000_0010100001011001"; -- 0.040895959641877595
	pesos_i(9693) := b"0000000000000000_0000000000000000_0000010111001000_1000001101010010"; -- 0.022590835166567232
	pesos_i(9694) := b"1111111111111111_1111111111111111_1110001110111010_0110011110001111"; -- -0.11043694274813304
	pesos_i(9695) := b"1111111111111111_1111111111111111_1111100000111101_0011011110001101"; -- -0.030315902718301715
	pesos_i(9696) := b"1111111111111111_1111111111111111_1111100111000010_0001001100011000"; -- -0.02438240691932951
	pesos_i(9697) := b"0000000000000000_0000000000000000_0010100010000000_0101100101100111"; -- 0.15820845385110668
	pesos_i(9698) := b"1111111111111111_1111111111111111_1101111101111101_1101010101011011"; -- -0.12698618447470983
	pesos_i(9699) := b"0000000000000000_0000000000000000_0001110101100100_0101100011010001"; -- 0.11481242278245285
	pesos_i(9700) := b"0000000000000000_0000000000000000_0000100100111001_0111000011010110"; -- 0.03603272647713148
	pesos_i(9701) := b"0000000000000000_0000000000000000_0001001101011110_0101111010001111"; -- 0.0756587122324768
	pesos_i(9702) := b"1111111111111111_1111111111111111_1110000110000101_1010110101101100"; -- -0.11905399427331557
	pesos_i(9703) := b"0000000000000000_0000000000000000_0000111110110101_0100100100000101"; -- 0.06135994304809858
	pesos_i(9704) := b"0000000000000000_0000000000000000_0000001010111011_1001010000100000"; -- 0.010674722465629883
	pesos_i(9705) := b"1111111111111111_1111111111111111_1110100110110000_1001101010100110"; -- -0.08714898538712136
	pesos_i(9706) := b"1111111111111111_1111111111111111_1110111011110001_0100000000100111"; -- -0.06663130810033267
	pesos_i(9707) := b"0000000000000000_0000000000000000_0001010010001000_0000101001010011"; -- 0.0802008106240852
	pesos_i(9708) := b"0000000000000000_0000000000000000_0010101111110010_0100110011000010"; -- 0.17166595203400017
	pesos_i(9709) := b"0000000000000000_0000000000000000_0000111111110101_0001111000001000"; -- 0.062333943351086246
	pesos_i(9710) := b"1111111111111111_1111111111111111_1111001110110110_0011010100011010"; -- -0.04800098521443868
	pesos_i(9711) := b"0000000000000000_0000000000000000_0010010101100000_0111100110111010"; -- 0.14600334926437555
	pesos_i(9712) := b"0000000000000000_0000000000000000_0010000010011100_0000111111101110"; -- 0.12738132048092468
	pesos_i(9713) := b"0000000000000000_0000000000000000_0000101101000010_0100001111100111"; -- 0.043979877399757734
	pesos_i(9714) := b"1111111111111111_1111111111111111_1111010110011101_0000011111110010"; -- -0.040572646429324205
	pesos_i(9715) := b"1111111111111111_1111111111111111_1101110010110111_1100100010010001"; -- -0.1378206869617527
	pesos_i(9716) := b"1111111111111111_1111111111111111_1110111100100101_0110011100010100"; -- -0.06583553084604096
	pesos_i(9717) := b"0000000000000000_0000000000000000_0000111001000011_1100010110110010"; -- 0.05572162243757744
	pesos_i(9718) := b"0000000000000000_0000000000000000_0000001101011011_0100011110110100"; -- 0.013111573732904402
	pesos_i(9719) := b"1111111111111111_1111111111111111_1110010100001100_1111001001100010"; -- -0.10527119740391062
	pesos_i(9720) := b"0000000000000000_0000000000000000_0000000100100000_0010001011010010"; -- 0.004396606814380236
	pesos_i(9721) := b"1111111111111111_1111111111111111_1110011000111011_1101011111100111"; -- -0.1006493627653393
	pesos_i(9722) := b"0000000000000000_0000000000000000_0000100000001010_1001001001101100"; -- 0.03141131533788239
	pesos_i(9723) := b"1111111111111111_1111111111111111_1111101110111110_1100111010110100"; -- -0.01661975960212108
	pesos_i(9724) := b"1111111111111111_1111111111111111_1110110001000001_0101001001011001"; -- -0.07712827044731764
	pesos_i(9725) := b"1111111111111111_1111111111111111_1101100110011001_0101111101010101"; -- -0.1500034730773076
	pesos_i(9726) := b"1111111111111111_1111111111111111_1111000110110010_0101100011001010"; -- -0.05587239322271731
	pesos_i(9727) := b"0000000000000000_0000000000000000_0010010111011011_0110000000011001"; -- 0.147878652577702
	pesos_i(9728) := b"1111111111111111_1111111111111111_1111011011100101_0010101110010111"; -- -0.03556563909048937
	pesos_i(9729) := b"1111111111111111_1111111111111111_1110111101001011_1001101010010111"; -- -0.06525262652617841
	pesos_i(9730) := b"0000000000000000_0000000000000000_0000111010011011_1000110100010101"; -- 0.05706102140253223
	pesos_i(9731) := b"1111111111111111_1111111111111111_1110111110111100_1101101100100110"; -- -0.06352453540177888
	pesos_i(9732) := b"0000000000000000_0000000000000000_0001110111111011_1110000110000010"; -- 0.11712464728112187
	pesos_i(9733) := b"1111111111111111_1111111111111111_1110110011000000_1110111110001000"; -- -0.07518103527633474
	pesos_i(9734) := b"0000000000000000_0000000000000000_0001101101001101_1000110100110100"; -- 0.10665209308640268
	pesos_i(9735) := b"1111111111111111_1111111111111111_1110110101111010_0011000001011111"; -- -0.0723542946127136
	pesos_i(9736) := b"0000000000000000_0000000000000000_0001000001100110_0101010011111100"; -- 0.06406146197086289
	pesos_i(9737) := b"0000000000000000_0000000000000000_0000001101111100_1100010011011010"; -- 0.013622573200753926
	pesos_i(9738) := b"1111111111111111_1111111111111111_1111101110011110_0110101111100001"; -- -0.0171139312771181
	pesos_i(9739) := b"0000000000000000_0000000000000000_0001110101101011_1001110101001001"; -- 0.11492331542446167
	pesos_i(9740) := b"1111111111111111_1111111111111111_1111101011011101_1010000110011000"; -- -0.02005567594378631
	pesos_i(9741) := b"0000000000000000_0000000000000000_0000110100101101_0111001100010110"; -- 0.051474755254518646
	pesos_i(9742) := b"0000000000000000_0000000000000000_0000000000111000_0001110010000100"; -- 0.0008561917552934495
	pesos_i(9743) := b"0000000000000000_0000000000000000_0010010010111010_1000101110110000"; -- 0.1434714606966244
	pesos_i(9744) := b"1111111111111111_1111111111111111_1101101111000011_1011001111101100"; -- -0.1415450619427984
	pesos_i(9745) := b"0000000000000000_0000000000000000_0001110000001011_0000011100101000"; -- 0.10954327320387737
	pesos_i(9746) := b"1111111111111111_1111111111111111_1110100010101010_1100011010001101"; -- -0.09114417119563531
	pesos_i(9747) := b"1111111111111111_1111111111111111_1101111000000010_1110010000001100"; -- -0.13276838986961195
	pesos_i(9748) := b"1111111111111111_1111111111111111_1111101000001101_1010011101111110"; -- -0.02322915235012643
	pesos_i(9749) := b"1111111111111111_1111111111111111_1110010101001100_1000100001011100"; -- -0.1043009542828617
	pesos_i(9750) := b"0000000000000000_0000000000000000_0000001001101100_0101000110001000"; -- 0.009465308971520606
	pesos_i(9751) := b"1111111111111111_1111111111111111_1111011010011000_0101100101111111"; -- -0.036737829652031914
	pesos_i(9752) := b"1111111111111111_1111111111111111_1101011101110110_1010000000010100"; -- -0.15834617157759442
	pesos_i(9753) := b"1111111111111111_1111111111111111_1110000011110011_1110011010000011"; -- -0.12127837460251865
	pesos_i(9754) := b"0000000000000000_0000000000000000_0001110110010101_0000110100100001"; -- 0.11555559214521982
	pesos_i(9755) := b"1111111111111111_1111111111111111_1111110010100011_0111010010001011"; -- -0.013130870902448443
	pesos_i(9756) := b"1111111111111111_1111111111111111_1101101100110011_0000110111101111"; -- -0.14375222120962017
	pesos_i(9757) := b"0000000000000000_0000000000000000_0010000110101011_1111001110011101"; -- 0.13153002337766165
	pesos_i(9758) := b"0000000000000000_0000000000000000_0001101110110110_1010011010110110"; -- 0.10825578642158104
	pesos_i(9759) := b"0000000000000000_0000000000000000_0000010101100011_1011001011110001"; -- 0.021052535918195593
	pesos_i(9760) := b"0000000000000000_0000000000000000_0000101000011010_1101101101111000"; -- 0.03947230982722151
	pesos_i(9761) := b"0000000000000000_0000000000000000_0001101100110001_1001001011110110"; -- 0.10622519018798755
	pesos_i(9762) := b"0000000000000000_0000000000000000_0000011110000010_0111111110111010"; -- 0.029335005670264678
	pesos_i(9763) := b"1111111111111111_1111111111111111_1111101111000001_1110111010100001"; -- -0.016572080276837674
	pesos_i(9764) := b"1111111111111111_1111111111111111_1111111001100101_0111100100110010"; -- -0.0062641385511439844
	pesos_i(9765) := b"1111111111111111_1111111111111111_1110101000010000_0110011110010101"; -- -0.0856871854138016
	pesos_i(9766) := b"1111111111111111_1111111111111111_1111110000001111_0001111001001110"; -- -0.015394311847278297
	pesos_i(9767) := b"1111111111111111_1111111111111111_1111110010011011_0110110100011101"; -- -0.013253384140908072
	pesos_i(9768) := b"1111111111111111_1111111111111111_1110101001100011_1000101110111011"; -- -0.0844185514070143
	pesos_i(9769) := b"1111111111111111_1111111111111111_1111110001000111_1011101110101101"; -- -0.014530439606229817
	pesos_i(9770) := b"1111111111111111_1111111111111111_1110110000001000_0100100001101101"; -- -0.07799861279576506
	pesos_i(9771) := b"0000000000000000_0000000000000000_0001000100101111_1110000100010001"; -- 0.06713682800467738
	pesos_i(9772) := b"0000000000000000_0000000000000000_0000110111010100_0110010010100010"; -- 0.05402211153832462
	pesos_i(9773) := b"0000000000000000_0000000000000000_0001011101111001_0000100110100101"; -- 0.09169063834548405
	pesos_i(9774) := b"0000000000000000_0000000000000000_0000000101000110_1011010100000001"; -- 0.0049851539179231776
	pesos_i(9775) := b"1111111111111111_1111111111111111_1111001100101110_0000101100111011"; -- -0.05007867622781316
	pesos_i(9776) := b"0000000000000000_0000000000000000_0001001010110000_0000101011011001"; -- 0.07299869355103311
	pesos_i(9777) := b"1111111111111111_1111111111111111_1111001000100110_1011001011110010"; -- -0.05409699996312669
	pesos_i(9778) := b"1111111111111111_1111111111111111_1111000110001000_0111001010000000"; -- -0.05651172994090011
	pesos_i(9779) := b"1111111111111111_1111111111111111_1111001100001010_0100110100101101"; -- -0.050624062063002226
	pesos_i(9780) := b"1111111111111111_1111111111111111_1111111001110100_0000101001101011"; -- -0.006041859603834058
	pesos_i(9781) := b"0000000000000000_0000000000000000_0010000010011001_1100000100001100"; -- 0.12734610113099556
	pesos_i(9782) := b"0000000000000000_0000000000000000_0001111010111001_0100001010011110"; -- 0.12001434655488512
	pesos_i(9783) := b"0000000000000000_0000000000000000_0001100001001110_1110110111000110"; -- 0.09495435803820428
	pesos_i(9784) := b"1111111111111111_1111111111111111_1111011110010001_1100110010010110"; -- -0.032931531398583104
	pesos_i(9785) := b"1111111111111111_1111111111111111_1101111010111110_1101010000110010"; -- -0.12990068225480725
	pesos_i(9786) := b"0000000000000000_0000000000000000_0000100011011000_1101111100111101"; -- 0.034559204371249645
	pesos_i(9787) := b"0000000000000000_0000000000000000_0010010100011100_0000111000011010"; -- 0.144959336712867
	pesos_i(9788) := b"0000000000000000_0000000000000000_0010011010010111_0010111011010001"; -- 0.1507443677084624
	pesos_i(9789) := b"1111111111111111_1111111111111111_1111010111100100_1001110011101110"; -- -0.039480392254980144
	pesos_i(9790) := b"0000000000000000_0000000000000000_0001101100001010_1111011011010000"; -- 0.10563604907193222
	pesos_i(9791) := b"1111111111111111_1111111111111111_1110010000001011_0010010010000010"; -- -0.10920497722198325
	pesos_i(9792) := b"1111111111111111_1111111111111111_1111111100000001_0010100101100101"; -- -0.0038885239147357785
	pesos_i(9793) := b"0000000000000000_0000000000000000_0001101111000111_0111010010110001"; -- 0.10851220438100222
	pesos_i(9794) := b"0000000000000000_0000000000000000_0000011110101110_1000010101100100"; -- 0.030006730037595165
	pesos_i(9795) := b"1111111111111111_1111111111111111_1110010010010101_0101100010100100"; -- -0.10709615703796808
	pesos_i(9796) := b"0000000000000000_0000000000000000_0000000001010100_1111110000010100"; -- 0.0012967633464598695
	pesos_i(9797) := b"0000000000000000_0000000000000000_0001111111110011_0010011110101100"; -- 0.12480400045408514
	pesos_i(9798) := b"0000000000000000_0000000000000000_0001111101010001_1011110111110110"; -- 0.12234103447408395
	pesos_i(9799) := b"0000000000000000_0000000000000000_0000111111111010_0000010101110111"; -- 0.062408772911607326
	pesos_i(9800) := b"1111111111111111_1111111111111111_1101110001111001_1011010111010011"; -- -0.13876784895473593
	pesos_i(9801) := b"0000000000000000_0000000000000000_0000101000011001_1100100001001011"; -- 0.03945590822467205
	pesos_i(9802) := b"0000000000000000_0000000000000000_0010010100101010_0111100110110110"; -- 0.14517937375515658
	pesos_i(9803) := b"1111111111111111_1111111111111111_1110101111100100_1111100001101000"; -- -0.07853743985148197
	pesos_i(9804) := b"0000000000000000_0000000000000000_0001100100110010_1111101110011111"; -- 0.0984341871381674
	pesos_i(9805) := b"0000000000000000_0000000000000000_0010011010111000_0100001111100101"; -- 0.15124916413176234
	pesos_i(9806) := b"1111111111111111_1111111111111111_1111111101101001_1001100010001101"; -- -0.0022949844481313995
	pesos_i(9807) := b"0000000000000000_0000000000000000_0000011100101111_0000001011100111"; -- 0.028061085988089544
	pesos_i(9808) := b"0000000000000000_0000000000000000_0010100000110010_1100111101101100"; -- 0.15702530283063604
	pesos_i(9809) := b"1111111111111111_1111111111111111_1111100000011111_0101100011011100"; -- -0.030771681141024795
	pesos_i(9810) := b"1111111111111111_1111111111111111_1101111000100100_0110111000101111"; -- -0.13225661607485006
	pesos_i(9811) := b"1111111111111111_1111111111111111_1111111111011000_1001010001110001"; -- -0.000601503719100417
	pesos_i(9812) := b"1111111111111111_1111111111111111_1110111000100101_0001110110011011"; -- -0.06974616023410614
	pesos_i(9813) := b"1111111111111111_1111111111111111_1110100010110110_0110011111110010"; -- -0.09096670487394615
	pesos_i(9814) := b"0000000000000000_0000000000000000_0000010010100101_1100010110110111"; -- 0.018154485024966006
	pesos_i(9815) := b"1111111111111111_1111111111111111_1101111000111001_0001100000111001"; -- -0.13194130534217827
	pesos_i(9816) := b"1111111111111111_1111111111111111_1111010101100101_0011000101010010"; -- -0.04142467250902391
	pesos_i(9817) := b"1111111111111111_1111111111111111_1110101011100101_1001111001101110"; -- -0.08243379426935597
	pesos_i(9818) := b"1111111111111111_1111111111111111_1110010001010011_0010010100100111"; -- -0.10810630608296792
	pesos_i(9819) := b"0000000000000000_0000000000000000_0001011111100100_1001111110100011"; -- 0.09333226899883897
	pesos_i(9820) := b"1111111111111111_1111111111111111_1101111101101100_1010101010010001"; -- -0.127248134221477
	pesos_i(9821) := b"0000000000000000_0000000000000000_0000010100101111_1000001011010011"; -- 0.020256210764521394
	pesos_i(9822) := b"1111111111111111_1111111111111111_1111010000000010_0101101110001010"; -- -0.046839026165422674
	pesos_i(9823) := b"0000000000000000_0000000000000000_0010010100011010_0101100010110000"; -- 0.14493326469000392
	pesos_i(9824) := b"0000000000000000_0000000000000000_0001010001101100_0011001111011011"; -- 0.07977604003562545
	pesos_i(9825) := b"1111111111111111_1111111111111111_1111101111011111_1111001110101011"; -- -0.016114016296601353
	pesos_i(9826) := b"1111111111111111_1111111111111111_1111010111011110_1011110010110010"; -- -0.03957005180968402
	pesos_i(9827) := b"1111111111111111_1111111111111111_1111011100001001_1010000010010111"; -- -0.03500934890055677
	pesos_i(9828) := b"1111111111111111_1111111111111111_1111011011101101_0011101111001100"; -- -0.03544260278659616
	pesos_i(9829) := b"1111111111111111_1111111111111111_1110001111000011_1101100111101011"; -- -0.11029279730569357
	pesos_i(9830) := b"0000000000000000_0000000000000000_0001001010110000_0111000010111001"; -- 0.07300476560894195
	pesos_i(9831) := b"1111111111111111_1111111111111111_1110101001101110_1101011001000001"; -- -0.08424626277534382
	pesos_i(9832) := b"1111111111111111_1111111111111111_1111101101101100_0010100011101100"; -- -0.017880861553747046
	pesos_i(9833) := b"1111111111111111_1111111111111111_1110101011100101_0101001001011000"; -- -0.08243832928094967
	pesos_i(9834) := b"1111111111111111_1111111111111111_1101101101000111_0111011001111010"; -- -0.14344081428629163
	pesos_i(9835) := b"1111111111111111_1111111111111111_1101111111010110_0001011010101010"; -- -0.12563951831253758
	pesos_i(9836) := b"0000000000000000_0000000000000000_0010000100000111_0110100010011010"; -- 0.12901929616983387
	pesos_i(9837) := b"1111111111111111_1111111111111111_1101111000010101_1000100100100100"; -- -0.13248389130763621
	pesos_i(9838) := b"0000000000000000_0000000000000000_0001111100011010_0101110001100000"; -- 0.12149598455642781
	pesos_i(9839) := b"1111111111111111_1111111111111111_1101011111001001_0001100100110110"; -- -0.15708773060452796
	pesos_i(9840) := b"1111111111111111_1111111111111111_1111001000111111_0011000110000110"; -- -0.05372324441425913
	pesos_i(9841) := b"0000000000000000_0000000000000000_0001110001111001_0011000111110010"; -- 0.11122429042408129
	pesos_i(9842) := b"1111111111111111_1111111111111111_1111110011100011_0100100010010010"; -- -0.012156929334119293
	pesos_i(9843) := b"1111111111111111_1111111111111111_1111111001010010_1110100101011011"; -- -0.0065473701593796755
	pesos_i(9844) := b"1111111111111111_1111111111111111_1111101100111000_0001100100001011"; -- -0.018675265221906986
	pesos_i(9845) := b"0000000000000000_0000000000000000_0000111101011101_1111011110101111"; -- 0.06002758051153093
	pesos_i(9846) := b"0000000000000000_0000000000000000_0001000010101101_1101101100110000"; -- 0.06515283503637187
	pesos_i(9847) := b"1111111111111111_1111111111111111_1110111011011101_1101000001101100"; -- -0.06692788480463394
	pesos_i(9848) := b"0000000000000000_0000000000000000_0010001111000111_0000110010110011"; -- 0.13975600599531643
	pesos_i(9849) := b"0000000000000000_0000000000000000_0001011111000110_0110000100010011"; -- 0.09287077628642215
	pesos_i(9850) := b"0000000000000000_0000000000000000_0001000011100111_0010011100111010"; -- 0.0660271184197595
	pesos_i(9851) := b"1111111111111111_1111111111111111_1101110010010011_0111101001101001"; -- -0.13837466188547698
	pesos_i(9852) := b"1111111111111111_1111111111111111_1110000111010111_0000110100001010"; -- -0.11781233319422424
	pesos_i(9853) := b"0000000000000000_0000000000000000_0010001001101010_0000101101010100"; -- 0.1344306069019866
	pesos_i(9854) := b"1111111111111111_1111111111111111_1111000111010001_1000100101111101"; -- -0.055396468138092604
	pesos_i(9855) := b"0000000000000000_0000000000000000_0010000100110011_0010001000100110"; -- 0.12968648362353707
	pesos_i(9856) := b"1111111111111111_1111111111111111_1101111011111001_1000100100101000"; -- -0.12900488638186283
	pesos_i(9857) := b"1111111111111111_1111111111111111_1111010110101110_1111001010000110"; -- -0.040299265285236516
	pesos_i(9858) := b"0000000000000000_0000000000000000_0001110110100001_0111100100110010"; -- 0.11574513879753547
	pesos_i(9859) := b"1111111111111111_1111111111111111_1110000011110101_0011010010100100"; -- -0.12125845911512434
	pesos_i(9860) := b"0000000000000000_0000000000000000_0001000011110101_0011000100000001"; -- 0.06624132421277255
	pesos_i(9861) := b"0000000000000000_0000000000000000_0000101001100010_0100111111010000"; -- 0.04056261850533836
	pesos_i(9862) := b"1111111111111111_1111111111111111_1110100000011000_0101100110100010"; -- -0.09337844659881107
	pesos_i(9863) := b"0000000000000000_0000000000000000_0001010000100100_0110100001101011"; -- 0.07868054021384949
	pesos_i(9864) := b"0000000000000000_0000000000000000_0000110100110111_1000110000001001"; -- 0.05162883014694132
	pesos_i(9865) := b"1111111111111111_1111111111111111_1110100110000100_1110011110101001"; -- -0.08781578181264182
	pesos_i(9866) := b"0000000000000000_0000000000000000_0001011001110110_1000101111000111"; -- 0.0877463684619783
	pesos_i(9867) := b"0000000000000000_0000000000000000_0000010111111011_1101101011110001"; -- 0.023374255949915757
	pesos_i(9868) := b"0000000000000000_0000000000000000_0010000101001010_0110001011011011"; -- 0.1300412925445317
	pesos_i(9869) := b"1111111111111111_1111111111111111_1101100111001011_0110100110100001"; -- -0.14923991989615223
	pesos_i(9870) := b"1111111111111111_1111111111111111_1111001010101111_1101011010011000"; -- -0.052004421074726144
	pesos_i(9871) := b"1111111111111111_1111111111111111_1110010100101100_0100011000111111"; -- -0.10479317640234193
	pesos_i(9872) := b"1111111111111111_1111111111111111_1111000000100010_1001011011001010"; -- -0.06197221352385383
	pesos_i(9873) := b"1111111111111111_1111111111111111_1110010111010010_1001000001110010"; -- -0.1022557946036411
	pesos_i(9874) := b"1111111111111111_1111111111111111_1110010101011110_1010111000001100"; -- -0.10402404973550669
	pesos_i(9875) := b"0000000000000000_0000000000000000_0001101110000010_1110101100111010"; -- 0.1074664132555736
	pesos_i(9876) := b"1111111111111111_1111111111111111_1101111101111000_1100100000010110"; -- -0.12706326919022243
	pesos_i(9877) := b"1111111111111111_1111111111111111_1110001111111000_0001110010011001"; -- -0.10949536583881098
	pesos_i(9878) := b"0000000000000000_0000000000000000_0000000010111101_0111111111010010"; -- 0.002891529774049275
	pesos_i(9879) := b"0000000000000000_0000000000000000_0000110101001100_0101101000111101"; -- 0.05194629661609103
	pesos_i(9880) := b"1111111111111111_1111111111111111_1111011101011001_1111011000101101"; -- -0.03378354463735455
	pesos_i(9881) := b"0000000000000000_0000000000000000_0001000001001111_1001101111100100"; -- 0.06371473622341718
	pesos_i(9882) := b"1111111111111111_1111111111111111_1111000100011100_1011001101000000"; -- -0.05815581979699994
	pesos_i(9883) := b"0000000000000000_0000000000000000_0010011000011011_1110011000011111"; -- 0.14886320353333718
	pesos_i(9884) := b"0000000000000000_0000000000000000_0000000011010111_0111000100001001"; -- 0.003287377028971019
	pesos_i(9885) := b"1111111111111111_1111111111111111_1110010000000000_1010000101000011"; -- -0.10936538795026814
	pesos_i(9886) := b"1111111111111111_1111111111111111_1101111010100001_0001001000110010"; -- -0.13035475044410286
	pesos_i(9887) := b"0000000000000000_0000000000000000_0000011110100000_1000101110000011"; -- 0.029793471907951678
	pesos_i(9888) := b"1111111111111111_1111111111111111_1111101101110111_1010011001111110"; -- -0.017705530349551264
	pesos_i(9889) := b"0000000000000000_0000000000000000_0000101000011110_0111000110110101"; -- 0.03952704124024105
	pesos_i(9890) := b"0000000000000000_0000000000000000_0000100101111010_0101001100011001"; -- 0.03702277534687352
	pesos_i(9891) := b"1111111111111111_1111111111111111_1111011110001001_1011110100110011"; -- -0.03305451876079684
	pesos_i(9892) := b"1111111111111111_1111111111111111_1111010111010110_1011110010101100"; -- -0.039692123479321786
	pesos_i(9893) := b"1111111111111111_1111111111111111_1111101111101010_0000001110100101"; -- -0.01596047608278101
	pesos_i(9894) := b"0000000000000000_0000000000000000_0010001110110110_0011110111001100"; -- 0.139499533006972
	pesos_i(9895) := b"1111111111111111_1111111111111111_1111111011111111_1100001100110100"; -- -0.003909873755527204
	pesos_i(9896) := b"1111111111111111_1111111111111111_1111110110011111_0011001001011111"; -- -0.009289600280880866
	pesos_i(9897) := b"0000000000000000_0000000000000000_0001001111001110_1001100111000101"; -- 0.07737122591529018
	pesos_i(9898) := b"0000000000000000_0000000000000000_0000101110010110_1101110100100101"; -- 0.0452707495796043
	pesos_i(9899) := b"1111111111111111_1111111111111111_1110110101000001_0110101110100001"; -- -0.07322051342058689
	pesos_i(9900) := b"1111111111111111_1111111111111111_1110010000100010_0101111010100011"; -- -0.10885056041107406
	pesos_i(9901) := b"1111111111111111_1111111111111111_1110011000110001_0111101110000111"; -- -0.10080745641662162
	pesos_i(9902) := b"0000000000000000_0000000000000000_0001100000110011_0101110100000111"; -- 0.09453374317297748
	pesos_i(9903) := b"0000000000000000_0000000000000000_0000001111001011_0100010100101101"; -- 0.01482040735467918
	pesos_i(9904) := b"0000000000000000_0000000000000000_0000000100101101_0101011111100111"; -- 0.004598134888204851
	pesos_i(9905) := b"1111111111111111_1111111111111111_1110001100011011_0010001101100111"; -- -0.11286715264878362
	pesos_i(9906) := b"1111111111111111_1111111111111111_1111100101000011_0011110001000000"; -- -0.026317820032324992
	pesos_i(9907) := b"0000000000000000_0000000000000000_0010001101010010_1111101110011001"; -- 0.13798496714095046
	pesos_i(9908) := b"0000000000000000_0000000000000000_0001100110000111_0101001011111100"; -- 0.09972113280374666
	pesos_i(9909) := b"1111111111111111_1111111111111111_1110101101110100_1100100001111111"; -- -0.08024927991831973
	pesos_i(9910) := b"0000000000000000_0000000000000000_0000111101110101_0011101011010101"; -- 0.06038253494656542
	pesos_i(9911) := b"0000000000000000_0000000000000000_0010000100001001_0010101101110001"; -- 0.12904616842685354
	pesos_i(9912) := b"0000000000000000_0000000000000000_0010010000000010_1001101110000100"; -- 0.1406647869157831
	pesos_i(9913) := b"0000000000000000_0000000000000000_0000011011000101_1110100111000001"; -- 0.026457414312870586
	pesos_i(9914) := b"0000000000000000_0000000000000000_0001010001100111_0010000110011010"; -- 0.07969865797726915
	pesos_i(9915) := b"1111111111111111_1111111111111111_1111110010111101_0101100100001001"; -- -0.012735781948517108
	pesos_i(9916) := b"1111111111111111_1111111111111111_1111110101000100_0011101110111110"; -- -0.010677591501643597
	pesos_i(9917) := b"1111111111111111_1111111111111111_1110101011100001_1111000000111011"; -- -0.08248995354503441
	pesos_i(9918) := b"1111111111111111_1111111111111111_1111100011110111_1110100000111110"; -- -0.027467236476544237
	pesos_i(9919) := b"0000000000000000_0000000000000000_0000001100010100_0111110001011101"; -- 0.012031338325599017
	pesos_i(9920) := b"1111111111111111_1111111111111111_1111000110010010_1110100110010010"; -- -0.056352044833069145
	pesos_i(9921) := b"0000000000000000_0000000000000000_0010000000000100_1111110001011010"; -- 0.1250760763685069
	pesos_i(9922) := b"0000000000000000_0000000000000000_0000001011110010_0100110100110111"; -- 0.01150972925543021
	pesos_i(9923) := b"1111111111111111_1111111111111111_1110101011101001_0000001110000000"; -- -0.08238199364390361
	pesos_i(9924) := b"0000000000000000_0000000000000000_0000011111001000_0000000011100100"; -- 0.030395560978848695
	pesos_i(9925) := b"1111111111111111_1111111111111111_1101111100101110_1011110101000000"; -- -0.12819306555493326
	pesos_i(9926) := b"1111111111111111_1111111111111111_1111100100001010_1001110011010000"; -- -0.027181815352118065
	pesos_i(9927) := b"1111111111111111_1111111111111111_1110100000001100_1100110010110000"; -- -0.09355469427917205
	pesos_i(9928) := b"0000000000000000_0000000000000000_0010011010100101_0001010000010000"; -- 0.1509563960962762
	pesos_i(9929) := b"0000000000000000_0000000000000000_0010011011101111_1110101110100101"; -- 0.15209839612221682
	pesos_i(9930) := b"0000000000000000_0000000000000000_0000001101100111_0111001001001011"; -- 0.013297217679771102
	pesos_i(9931) := b"0000000000000000_0000000000000000_0001111010010001_1100000001111101"; -- 0.11941149771631791
	pesos_i(9932) := b"0000000000000000_0000000000000000_0001000001111100_0000111100100001"; -- 0.06439299150468956
	pesos_i(9933) := b"1111111111111111_1111111111111111_1111000110000100_0110001011101001"; -- -0.05657369425404386
	pesos_i(9934) := b"0000000000000000_0000000000000000_0000100101110011_0001111010011100"; -- 0.036912835238690656
	pesos_i(9935) := b"0000000000000000_0000000000000000_0001100110010111_1100001011010011"; -- 0.09997193968889995
	pesos_i(9936) := b"0000000000000000_0000000000000000_0000001011011110_1110110100001010"; -- 0.0112140797288709
	pesos_i(9937) := b"0000000000000000_0000000000000000_0000100011101100_1110001101010011"; -- 0.034864623837833314
	pesos_i(9938) := b"1111111111111111_1111111111111111_1110011000010011_0000111010010010"; -- -0.10127171444614419
	pesos_i(9939) := b"1111111111111111_1111111111111111_1111000101100010_1011000010111110"; -- -0.057087853935911356
	pesos_i(9940) := b"1111111111111111_1111111111111111_1111100110111111_1110011010100110"; -- -0.024415573617427987
	pesos_i(9941) := b"1111111111111111_1111111111111111_1101110011011111_0010011000001001"; -- -0.13722002291638707
	pesos_i(9942) := b"0000000000000000_0000000000000000_0001010001000011_1110010101011000"; -- 0.07916100879216023
	pesos_i(9943) := b"1111111111111111_1111111111111111_1101111100101000_1010110010110000"; -- -0.1282856055705156
	pesos_i(9944) := b"1111111111111111_1111111111111111_1111010011010110_0011001001100100"; -- -0.0436066156798831
	pesos_i(9945) := b"1111111111111111_1111111111111111_1110010011010011_1010101100101001"; -- -0.10614519354307095
	pesos_i(9946) := b"0000000000000000_0000000000000000_0001001011001100_1011100001000110"; -- 0.0734362765841745
	pesos_i(9947) := b"1111111111111111_1111111111111111_1101111001110000_1100111100010101"; -- -0.13109117261299996
	pesos_i(9948) := b"0000000000000000_0000000000000000_0000011001011101_1110111100001110"; -- 0.02487081622416034
	pesos_i(9949) := b"1111111111111111_1111111111111111_1111010110000001_0101011000110001"; -- -0.04099522870093094
	pesos_i(9950) := b"0000000000000000_0000000000000000_0010100110001000_1101000001111000"; -- 0.1622438710153152
	pesos_i(9951) := b"1111111111111111_1111111111111111_1111011111010011_1100111001110011"; -- -0.03192434012269976
	pesos_i(9952) := b"0000000000000000_0000000000000000_0000000111110101_0000000110110110"; -- 0.00764475535729927
	pesos_i(9953) := b"0000000000000000_0000000000000000_0000010111011010_1101110101001110"; -- 0.02287085669804134
	pesos_i(9954) := b"0000000000000000_0000000000000000_0001101100111111_1001001110101100"; -- 0.10643885560227669
	pesos_i(9955) := b"1111111111111111_1111111111111111_1101101111101010_0110010100111011"; -- -0.14095465958958914
	pesos_i(9956) := b"0000000000000000_0000000000000000_0000011101011010_0111001100001011"; -- 0.028723898115782055
	pesos_i(9957) := b"0000000000000000_0000000000000000_0000011111110000_0110100010000001"; -- 0.031012088259646214
	pesos_i(9958) := b"1111111111111111_1111111111111111_1110010011011011_0001100110111001"; -- -0.10603179211761937
	pesos_i(9959) := b"1111111111111111_1111111111111111_1101111011000100_0010101111011011"; -- -0.1298191633972329
	pesos_i(9960) := b"0000000000000000_0000000000000000_0000011100001010_0100111101010010"; -- 0.027501065851277356
	pesos_i(9961) := b"1111111111111111_1111111111111111_1110111101110001_1010110111101001"; -- -0.06467164093207699
	pesos_i(9962) := b"1111111111111111_1111111111111111_1111110100100011_0000110101110011"; -- -0.011183890649210585
	pesos_i(9963) := b"1111111111111111_1111111111111111_1111001110000100_0010011011000010"; -- -0.04876477980867764
	pesos_i(9964) := b"0000000000000000_0000000000000000_0000110101011101_1101001101111101"; -- 0.052212923056520436
	pesos_i(9965) := b"1111111111111111_1111111111111111_1101101011101010_1110110110010110"; -- -0.14485278214358685
	pesos_i(9966) := b"0000000000000000_0000000000000000_0001110101010100_1101100010111000"; -- 0.11457590568144174
	pesos_i(9967) := b"0000000000000000_0000000000000000_0000111101000001_1001111011111011"; -- 0.05959504737065934
	pesos_i(9968) := b"0000000000000000_0000000000000000_0000101001101011_0100011100101010"; -- 0.04069943209253918
	pesos_i(9969) := b"0000000000000000_0000000000000000_0000001011001011_0001101001111000"; -- 0.010911611767927968
	pesos_i(9970) := b"0000000000000000_0000000000000000_0001000111011110_0110000110010110"; -- 0.06979951774407375
	pesos_i(9971) := b"1111111111111111_1111111111111111_1110100100000011_0111011110111000"; -- -0.08979083783150572
	pesos_i(9972) := b"0000000000000000_0000000000000000_0001001011011000_1010010011111000"; -- 0.07361823143019927
	pesos_i(9973) := b"0000000000000000_0000000000000000_0001101101001111_0100111001110111"; -- 0.10667887119506272
	pesos_i(9974) := b"1111111111111111_1111111111111111_1111111000101010_0100001000111111"; -- -0.0071676822356448455
	pesos_i(9975) := b"0000000000000000_0000000000000000_0010001110001110_1111000101111000"; -- 0.13889989059994587
	pesos_i(9976) := b"0000000000000000_0000000000000000_0000111100111010_0101000000010101"; -- 0.059483532978718404
	pesos_i(9977) := b"1111111111111111_1111111111111111_1110001111111010_0000010010010010"; -- -0.10946628022176395
	pesos_i(9978) := b"1111111111111111_1111111111111111_1111011101100101_0100101111011011"; -- -0.033610590935725417
	pesos_i(9979) := b"1111111111111111_1111111111111111_1101111000011111_1110000000001101"; -- -0.13232612307208555
	pesos_i(9980) := b"1111111111111111_1111111111111111_1111101101010001_1110011011101110"; -- -0.018281523569873514
	pesos_i(9981) := b"1111111111111111_1111111111111111_1110011110111001_0000000011010001"; -- -0.09483332537579514
	pesos_i(9982) := b"1111111111111111_1111111111111111_1111100000000111_1011010000111011"; -- -0.031132445963799108
	pesos_i(9983) := b"1111111111111111_1111111111111111_1110110001011111_0000000001000111"; -- -0.07667539856507176
	pesos_i(9984) := b"0000000000000000_0000000000000000_0001010100101110_0010111100001100"; -- 0.08273595844295761
	pesos_i(9985) := b"0000000000000000_0000000000000000_0001001011100001_1010101011100111"; -- 0.073755914025424
	pesos_i(9986) := b"1111111111111111_1111111111111111_1110001011110100_0010010111111101"; -- -0.1134620911969403
	pesos_i(9987) := b"0000000000000000_0000000000000000_0001000100100001_0011111001110110"; -- 0.06691351297721443
	pesos_i(9988) := b"0000000000000000_0000000000000000_0000100000100100_1111111001001111"; -- 0.031814474337785614
	pesos_i(9989) := b"0000000000000000_0000000000000000_0000101110101010_0111101100001010"; -- 0.045570077936949456
	pesos_i(9990) := b"0000000000000000_0000000000000000_0000011011011000_1101000011101101"; -- 0.02674585137004118
	pesos_i(9991) := b"0000000000000000_0000000000000000_0000011001101010_0111100011011110"; -- 0.025062135935039753
	pesos_i(9992) := b"1111111111111111_1111111111111111_1110010111010101_0011011010110010"; -- -0.10221536791613516
	pesos_i(9993) := b"1111111111111111_1111111111111111_1111000011010011_0000000111101000"; -- -0.05928028184170206
	pesos_i(9994) := b"0000000000000000_0000000000000000_0000011100001101_0100111100010111"; -- 0.02754682834541211
	pesos_i(9995) := b"1111111111111111_1111111111111111_1111100001110001_0100011011011000"; -- -0.029521534266544826
	pesos_i(9996) := b"1111111111111111_1111111111111111_1101100101111111_1000010000101011"; -- -0.1503980058967484
	pesos_i(9997) := b"0000000000000000_0000000000000000_0000010110111111_1110010100101001"; -- 0.02245933765347281
	pesos_i(9998) := b"0000000000000000_0000000000000000_0000001100110110_0000010010011100"; -- 0.012542999397620463
	pesos_i(9999) := b"0000000000000000_0000000000000000_0001011110111011_0001101011100100"; -- 0.0926987464676537
	pesos_i(10000) := b"1111111111111111_1111111111111111_1101111010011110_0010010000000101"; -- -0.1303994644571403
	pesos_i(10001) := b"0000000000000000_0000000000000000_0001010110100100_1110001101110100"; -- 0.08454724862573007
	pesos_i(10002) := b"1111111111111111_1111111111111111_1111000011100111_1000101001010110"; -- -0.058966974185526946
	pesos_i(10003) := b"1111111111111111_1111111111111111_1111010100110100_1001100001011111"; -- -0.042166211003132927
	pesos_i(10004) := b"0000000000000000_0000000000000000_0001100010101100_1110010010010000"; -- 0.09638813519746033
	pesos_i(10005) := b"0000000000000000_0000000000000000_0000110010001101_1110001100101001"; -- 0.04904002907585035
	pesos_i(10006) := b"0000000000000000_0000000000000000_0000100111010100_1101011000000000"; -- 0.03840386865291662
	pesos_i(10007) := b"1111111111111111_1111111111111111_1111100000110110_0110000010100011"; -- -0.030420265416019013
	pesos_i(10008) := b"1111111111111111_1111111111111111_1110010111010001_1110101010110001"; -- -0.10226567438053229
	pesos_i(10009) := b"1111111111111111_1111111111111111_1111001110010110_0000000101011010"; -- -0.04849235101895415
	pesos_i(10010) := b"0000000000000000_0000000000000000_0001110111000001_0001000001000000"; -- 0.11622716496679052
	pesos_i(10011) := b"0000000000000000_0000000000000000_0001111001111101_1001101011010101"; -- 0.11910407727053544
	pesos_i(10012) := b"1111111111111111_1111111111111111_1111001001011010_1110001000011101"; -- -0.0533007315822104
	pesos_i(10013) := b"1111111111111111_1111111111111111_1110111100101101_1011110000111111"; -- -0.06570838423338267
	pesos_i(10014) := b"0000000000000000_0000000000000000_0000100000011001_0011111111100100"; -- 0.0316352780092118
	pesos_i(10015) := b"1111111111111111_1111111111111111_1110111100101000_1011011110100011"; -- -0.06578495279263809
	pesos_i(10016) := b"1111111111111111_1111111111111111_1111010010100001_0111110011010101"; -- -0.0444108944244534
	pesos_i(10017) := b"1111111111111111_1111111111111111_1101101000101110_1111000010110111"; -- -0.147721247990696
	pesos_i(10018) := b"0000000000000000_0000000000000000_0000100111111001_1110011001010101"; -- 0.038969417289275235
	pesos_i(10019) := b"1111111111111111_1111111111111111_1110100101100101_0011110000111010"; -- -0.08829902246015969
	pesos_i(10020) := b"1111111111111111_1111111111111111_1111001010011100_0110110001010101"; -- -0.05230067188358211
	pesos_i(10021) := b"1111111111111111_1111111111111111_1110011110110001_1110101101101110"; -- -0.09494141169684002
	pesos_i(10022) := b"1111111111111111_1111111111111111_1101100010001011_0101111010010111"; -- -0.15412339034665076
	pesos_i(10023) := b"1111111111111111_1111111111111111_1111110001011110_1000101111011100"; -- -0.014182337598851348
	pesos_i(10024) := b"1111111111111111_1111111111111111_1111000000001010_1100111010010001"; -- -0.062335099765244956
	pesos_i(10025) := b"1111111111111111_1111111111111111_1101111110011011_0011100001001110"; -- -0.12653778173458818
	pesos_i(10026) := b"1111111111111111_1111111111111111_1111111101111000_1110000100110100"; -- -0.0020617722230784376
	pesos_i(10027) := b"0000000000000000_0000000000000000_0000010110101100_1011101010111101"; -- 0.022166892078274006
	pesos_i(10028) := b"0000000000000000_0000000000000000_0001110110001000_0011110101110001"; -- 0.11536010758534467
	pesos_i(10029) := b"1111111111111111_1111111111111111_1110001011011100_1010011000110101"; -- -0.11382065957989733
	pesos_i(10030) := b"1111111111111111_1111111111111111_1110110000100101_1010000001101000"; -- -0.07755086393653919
	pesos_i(10031) := b"1111111111111111_1111111111111111_1111101010001101_0010111111011011"; -- -0.021283158383478062
	pesos_i(10032) := b"0000000000000000_0000000000000000_0001011011100000_0110110100101111"; -- 0.0893619764913007
	pesos_i(10033) := b"1111111111111111_1111111111111111_1110010110010101_0001111010011101"; -- -0.10319336572167666
	pesos_i(10034) := b"0000000000000000_0000000000000000_0001010000001110_1100011010001110"; -- 0.07835045781595368
	pesos_i(10035) := b"1111111111111111_1111111111111111_1101101100000100_1111101010011101"; -- -0.1444552771871298
	pesos_i(10036) := b"0000000000000000_0000000000000000_0001010100111110_1011001101111001"; -- 0.08298799239443494
	pesos_i(10037) := b"1111111111111111_1111111111111111_1101110011100000_1110001010101010"; -- -0.13719352092022832
	pesos_i(10038) := b"0000000000000000_0000000000000000_0001110001000101_1100011011011000"; -- 0.11043970850497518
	pesos_i(10039) := b"1111111111111111_1111111111111111_1111011000000000_0011111100001100"; -- -0.039058742157947204
	pesos_i(10040) := b"0000000000000000_0000000000000000_0000111000100111_0110011001111000"; -- 0.05528870029542353
	pesos_i(10041) := b"1111111111111111_1111111111111111_1111001110111011_1001100011101001"; -- -0.04791874236114215
	pesos_i(10042) := b"1111111111111111_1111111111111111_1110101001000000_0100001001001110"; -- -0.08495698537858457
	pesos_i(10043) := b"0000000000000000_0000000000000000_0001101011000001_1000100111001101"; -- 0.10451565982923301
	pesos_i(10044) := b"1111111111111111_1111111111111111_1110011100011010_1110101101010110"; -- -0.0972454944354227
	pesos_i(10045) := b"1111111111111111_1111111111111111_1111010000100000_1000000111010110"; -- -0.04637897996618142
	pesos_i(10046) := b"0000000000000000_0000000000000000_0001100111101111_1100001110010111"; -- 0.10131475861585074
	pesos_i(10047) := b"1111111111111111_1111111111111111_1101111100011001_0010110001001101"; -- -0.1285221397028117
	pesos_i(10048) := b"1111111111111111_1111111111111111_1111101101011111_1001011100101010"; -- -0.018072654993092838
	pesos_i(10049) := b"0000000000000000_0000000000000000_0001100100101100_1011100011101110"; -- 0.09833865936873565
	pesos_i(10050) := b"0000000000000000_0000000000000000_0000000110100100_1011101001011000"; -- 0.0064197984280182155
	pesos_i(10051) := b"0000000000000000_0000000000000000_0001111010111111_1010011000111011"; -- 0.12011183687630278
	pesos_i(10052) := b"0000000000000000_0000000000000000_0000110101110010_0100000100111100"; -- 0.052524640327267995
	pesos_i(10053) := b"0000000000000000_0000000000000000_0000101001111111_1100011010100001"; -- 0.041012205384136705
	pesos_i(10054) := b"1111111111111111_1111111111111111_1111110111010101_0011111010110100"; -- -0.008464890525510015
	pesos_i(10055) := b"0000000000000000_0000000000000000_0001001110011000_1111111110011011"; -- 0.07655332120759645
	pesos_i(10056) := b"0000000000000000_0000000000000000_0001100111111010_0001101010110100"; -- 0.1014725388652139
	pesos_i(10057) := b"1111111111111111_1111111111111111_1110100001010101_1000010111000000"; -- -0.0924450308016149
	pesos_i(10058) := b"0000000000000000_0000000000000000_0001110100001110_1101000011001010"; -- 0.11350731793096866
	pesos_i(10059) := b"0000000000000000_0000000000000000_0001110101000111_1101100100101000"; -- 0.11437756744051142
	pesos_i(10060) := b"0000000000000000_0000000000000000_0001110111000011_0100001011111010"; -- 0.1162607060692297
	pesos_i(10061) := b"0000000000000000_0000000000000000_0000100110111001_1111010111000110"; -- 0.03799377524800891
	pesos_i(10062) := b"1111111111111111_1111111111111111_1110001101111101_1001111110001100"; -- -0.1113643917320969
	pesos_i(10063) := b"0000000000000000_0000000000000000_0000110100110000_0101000110011000"; -- 0.051518535150755475
	pesos_i(10064) := b"1111111111111111_1111111111111111_1110111011001011_1011101101101011"; -- -0.0672037948289844
	pesos_i(10065) := b"1111111111111111_1111111111111111_1110000011101100_1101110010010001"; -- -0.1213857790160364
	pesos_i(10066) := b"0000000000000000_0000000000000000_0000010100110001_0111110010001111"; -- 0.02028635483541521
	pesos_i(10067) := b"0000000000000000_0000000000000000_0000100100111111_1000010000010100"; -- 0.036125426225596904
	pesos_i(10068) := b"0000000000000000_0000000000000000_0000010100001111_0001001010011000"; -- 0.01976124020912215
	pesos_i(10069) := b"1111111111111111_1111111111111111_1110100010011000_1001000110110100"; -- -0.09142197948833586
	pesos_i(10070) := b"0000000000000000_0000000000000000_0001101000101100_0001111001010000"; -- 0.10223569347382437
	pesos_i(10071) := b"1111111111111111_1111111111111111_1110010101111111_0011001111100010"; -- -0.10352779121679052
	pesos_i(10072) := b"1111111111111111_1111111111111111_1110111111110000_0101010110011100"; -- -0.06273903779420535
	pesos_i(10073) := b"1111111111111111_1111111111111111_1110011111001100_0101111101100111"; -- -0.0945377705727815
	pesos_i(10074) := b"1111111111111111_1111111111111111_1111101100110111_1111111011101101"; -- -0.018676821738423187
	pesos_i(10075) := b"1111111111111111_1111111111111111_1111111001100001_0011100100000110"; -- -0.006328998489903544
	pesos_i(10076) := b"0000000000000000_0000000000000000_0000110101000010_0010010101111011"; -- 0.05179056414027904
	pesos_i(10077) := b"1111111111111111_1111111111111111_1111010111111000_0010001000110000"; -- -0.03918253255210425
	pesos_i(10078) := b"0000000000000000_0000000000000000_0000100001111101_0000111001111101"; -- 0.03315821229304021
	pesos_i(10079) := b"0000000000000000_0000000000000000_0000110010001010_1101110100001000"; -- 0.04899388745113983
	pesos_i(10080) := b"1111111111111111_1111111111111111_1111010100001011_0101111000000101"; -- -0.04279529925607389
	pesos_i(10081) := b"0000000000000000_0000000000000000_0010000000110101_0000110110000100"; -- 0.12580952137525922
	pesos_i(10082) := b"1111111111111111_1111111111111111_1111000101100001_1000110101000101"; -- -0.057105227154232774
	pesos_i(10083) := b"0000000000000000_0000000000000000_0001010010010010_0000010110110101"; -- 0.08035312338516266
	pesos_i(10084) := b"1111111111111111_1111111111111111_1111100000011111_0001100101000010"; -- -0.030775472024956098
	pesos_i(10085) := b"1111111111111111_1111111111111111_1110010100100101_0001000100111101"; -- -0.10490314740285786
	pesos_i(10086) := b"0000000000000000_0000000000000000_0001110101010101_0001100110011111"; -- 0.114579774296092
	pesos_i(10087) := b"1111111111111111_1111111111111111_1111110000001001_0110010010101010"; -- -0.015481670805653141
	pesos_i(10088) := b"1111111111111111_1111111111111111_1110110100100101_1000000000010110"; -- -0.07364654029778019
	pesos_i(10089) := b"1111111111111111_1111111111111111_1110001101111001_0111011110111011"; -- -0.11142779995475666
	pesos_i(10090) := b"0000000000000000_0000000000000000_0000011111010000_0101101001000011"; -- 0.030522958057378348
	pesos_i(10091) := b"1111111111111111_1111111111111111_1101111101111010_0000111010110110"; -- -0.1270438007851956
	pesos_i(10092) := b"1111111111111111_1111111111111111_1111111001000010_1010100011111101"; -- -0.006795347367323704
	pesos_i(10093) := b"0000000000000000_0000000000000000_0000101101000011_0011110011011011"; -- 0.04399471624076969
	pesos_i(10094) := b"0000000000000000_0000000000000000_0010000110001010_0101111111010111"; -- 0.13101767534962974
	pesos_i(10095) := b"1111111111111111_1111111111111111_1110000111000010_0010010101011111"; -- -0.11813131733593345
	pesos_i(10096) := b"0000000000000000_0000000000000000_0010010100011011_0111001100001100"; -- 0.14495009459905756
	pesos_i(10097) := b"1111111111111111_1111111111111111_1110000010100101_0111110111001111"; -- -0.1224748009607064
	pesos_i(10098) := b"1111111111111111_1111111111111111_1110100100110000_0010000011100111"; -- -0.0891093670338037
	pesos_i(10099) := b"0000000000000000_0000000000000000_0001000101110101_0100111011010000"; -- 0.06819622585388929
	pesos_i(10100) := b"0000000000000000_0000000000000000_0001001100101011_1101101000001111"; -- 0.0748878753073859
	pesos_i(10101) := b"1111111111111111_1111111111111111_1110000111110100_0100011011011000"; -- -0.1173663829583723
	pesos_i(10102) := b"0000000000000000_0000000000000000_0001010101000100_0110011011000001"; -- 0.08307497234192855
	pesos_i(10103) := b"0000000000000000_0000000000000000_0001111100111011_1001110110010100"; -- 0.12200341103593201
	pesos_i(10104) := b"1111111111111111_1111111111111111_1111010101011011_1010101101000111"; -- -0.041569991322191344
	pesos_i(10105) := b"1111111111111111_1111111111111111_1111011001001000_1010110011110111"; -- -0.03795355775347465
	pesos_i(10106) := b"1111111111111111_1111111111111111_1111011100001001_1110101100000101"; -- -0.03500491269193643
	pesos_i(10107) := b"1111111111111111_1111111111111111_1110000111010101_1011001001110010"; -- -0.11783299167328697
	pesos_i(10108) := b"0000000000000000_0000000000000000_0001111011001011_0110101010001100"; -- 0.1202913848302228
	pesos_i(10109) := b"1111111111111111_1111111111111111_1111111101100001_0010111010110111"; -- -0.002423363115388354
	pesos_i(10110) := b"1111111111111111_1111111111111111_1111100101100110_0000111000000000"; -- -0.02578651894283288
	pesos_i(10111) := b"1111111111111111_1111111111111111_1101101101110101_1000010010100011"; -- -0.14273806599001257
	pesos_i(10112) := b"0000000000000000_0000000000000000_0010001100000100_1100100000111000"; -- 0.13679171906187132
	pesos_i(10113) := b"1111111111111111_1111111111111111_1110110011100010_1011011101110011"; -- -0.07466557915921086
	pesos_i(10114) := b"0000000000000000_0000000000000000_0010000011001011_0101011111101111"; -- 0.1281027754463096
	pesos_i(10115) := b"1111111111111111_1111111111111111_1101110101111100_1000111010101101"; -- -0.13481815597721064
	pesos_i(10116) := b"1111111111111111_1111111111111111_1110001001110100_0000001011110111"; -- -0.1154173038616128
	pesos_i(10117) := b"0000000000000000_0000000000000000_0001110010111111_1111000001011110"; -- 0.11230375561120019
	pesos_i(10118) := b"1111111111111111_1111111111111111_1110010010010001_1100000111111000"; -- -0.10715091420105982
	pesos_i(10119) := b"1111111111111111_1111111111111111_1110010011101011_0001100110111000"; -- -0.10578765152812457
	pesos_i(10120) := b"0000000000000000_0000000000000000_0001010000100100_0000001011110111"; -- 0.07867449310436817
	pesos_i(10121) := b"0000000000000000_0000000000000000_0000110000011011_0011100011101011"; -- 0.047290379841830925
	pesos_i(10122) := b"0000000000000000_0000000000000000_0001100100101000_0110111111011001"; -- 0.09827326817081763
	pesos_i(10123) := b"1111111111111111_1111111111111111_1110000101001000_1111100100111000"; -- -0.1199802626944165
	pesos_i(10124) := b"0000000000000000_0000000000000000_0000011010110000_1001100111000111"; -- 0.02613221264111803
	pesos_i(10125) := b"0000000000000000_0000000000000000_0001110100001010_0001000110000101"; -- 0.11343488209394616
	pesos_i(10126) := b"0000000000000000_0000000000000000_0000001011011001_0010110001100011"; -- 0.011126302956147293
	pesos_i(10127) := b"1111111111111111_1111111111111111_1110010010001110_1100111110010101"; -- -0.10719587904774822
	pesos_i(10128) := b"1111111111111111_1111111111111111_1110001000110000_0010010001011110"; -- -0.11645291041741147
	pesos_i(10129) := b"1111111111111111_1111111111111111_1111001001010000_0010101111010001"; -- -0.05346418525163612
	pesos_i(10130) := b"1111111111111111_1111111111111111_1101011110101011_0010100011000100"; -- -0.1575445671401011
	pesos_i(10131) := b"1111111111111111_1111111111111111_1110010000110010_0100100000011101"; -- -0.10860776227819155
	pesos_i(10132) := b"1111111111111111_1111111111111111_1110110100001100_1011110111111110"; -- -0.07402432006137076
	pesos_i(10133) := b"0000000000000000_0000000000000000_0001001100011010_1110001001101000"; -- 0.07462897343809204
	pesos_i(10134) := b"0000000000000000_0000000000000000_0001111110101010_0000010111001111"; -- 0.12368809037047114
	pesos_i(10135) := b"1111111111111111_1111111111111111_1101111001110000_0100011101110010"; -- -0.1310992570837014
	pesos_i(10136) := b"0000000000000000_0000000000000000_0000001011011010_0111110101010111"; -- 0.011146386754477914
	pesos_i(10137) := b"0000000000000000_0000000000000000_0000111000110101_1100011010011110"; -- 0.05550805423952506
	pesos_i(10138) := b"0000000000000000_0000000000000000_0001001000000101_0010101110010001"; -- 0.07039139069052582
	pesos_i(10139) := b"1111111111111111_1111111111111111_1110001000100010_0001110000100110"; -- -0.11666702339811662
	pesos_i(10140) := b"1111111111111111_1111111111111111_1101111010010101_0001100000011011"; -- -0.1305375036272219
	pesos_i(10141) := b"0000000000000000_0000000000000000_0000011001010110_0111011011001011"; -- 0.024756836471026594
	pesos_i(10142) := b"1111111111111111_1111111111111111_1101101001100011_1111111110110011"; -- -0.14691163907792426
	pesos_i(10143) := b"1111111111111111_1111111111111111_1110011000111001_0111011110001001"; -- -0.10068562412010928
	pesos_i(10144) := b"0000000000000000_0000000000000000_0010001010000010_0010001110110010"; -- 0.13479827027403915
	pesos_i(10145) := b"1111111111111111_1111111111111111_1111010001000000_0000101101000000"; -- -0.045897766933140356
	pesos_i(10146) := b"0000000000000000_0000000000000000_0010011011000101_1010011011010101"; -- 0.15145342534983205
	pesos_i(10147) := b"0000000000000000_0000000000000000_0000001110110011_1111000100011101"; -- 0.014464444737189747
	pesos_i(10148) := b"1111111111111111_1111111111111111_1110001011111011_1110010100111011"; -- -0.11334388082736405
	pesos_i(10149) := b"1111111111111111_1111111111111111_1111001100000000_0100000101101101"; -- -0.050777350268518186
	pesos_i(10150) := b"0000000000000000_0000000000000000_0010010001100011_1101111110001110"; -- 0.14214894495809455
	pesos_i(10151) := b"1111111111111111_1111111111111111_1110011111111000_0100011011000100"; -- -0.09386785240206394
	pesos_i(10152) := b"1111111111111111_1111111111111111_1101111000101110_1010011100100101"; -- -0.1321006331763478
	pesos_i(10153) := b"1111111111111111_1111111111111111_1110001001001011_0011110000000111"; -- -0.11603951292881695
	pesos_i(10154) := b"0000000000000000_0000000000000000_0001000000010101_0011111011000110"; -- 0.06282417614329609
	pesos_i(10155) := b"0000000000000000_0000000000000000_0000101111110001_1011011010011110"; -- 0.046657002888485406
	pesos_i(10156) := b"0000000000000000_0000000000000000_0010001011001000_0001100111101110"; -- 0.135865803341249
	pesos_i(10157) := b"0000000000000000_0000000000000000_0000010101100111_0110001111101100"; -- 0.021108861111026493
	pesos_i(10158) := b"0000000000000000_0000000000000000_0000110101011110_1001100000001011"; -- 0.05222463864946935
	pesos_i(10159) := b"1111111111111111_1111111111111111_1111011011101101_1111001111000111"; -- -0.03543163680837683
	pesos_i(10160) := b"0000000000000000_0000000000000000_0001110100100101_1001010010001001"; -- 0.11385467852629923
	pesos_i(10161) := b"0000000000000000_0000000000000000_0000111011110110_1111000011101001"; -- 0.05845552139676199
	pesos_i(10162) := b"1111111111111111_1111111111111111_1111001110100011_0000011100010000"; -- -0.04829364640424564
	pesos_i(10163) := b"1111111111111111_1111111111111111_1110011110001110_1000111011001001"; -- -0.09548099129906049
	pesos_i(10164) := b"1111111111111111_1111111111111111_1111110111111011_0010001110101001"; -- -0.007886668529371992
	pesos_i(10165) := b"1111111111111111_1111111111111111_1111100110011100_0101010001001000"; -- -0.024958355356435227
	pesos_i(10166) := b"1111111111111111_1111111111111111_1111100011001000_0101011111000101"; -- -0.028193010775890995
	pesos_i(10167) := b"1111111111111111_1111111111111111_1111001101011101_0100000110000100"; -- -0.049358277624687294
	pesos_i(10168) := b"1111111111111111_1111111111111111_1110000110001101_1010110011011011"; -- -0.11893195763840882
	pesos_i(10169) := b"1111111111111111_1111111111111111_1110111110111101_1011001011110110"; -- -0.0635116719789188
	pesos_i(10170) := b"1111111111111111_1111111111111111_1101111010110001_0101111101101010"; -- -0.13010600715546403
	pesos_i(10171) := b"0000000000000000_0000000000000000_0001011100100010_0110011110110100"; -- 0.09036873003184306
	pesos_i(10172) := b"0000000000000000_0000000000000000_0001000000011000_0101000110101001"; -- 0.06287107828893072
	pesos_i(10173) := b"0000000000000000_0000000000000000_0000101111111100_1111000011101101"; -- 0.046828325179981124
	pesos_i(10174) := b"1111111111111111_1111111111111111_1110111001010001_1010100100111001"; -- -0.06906645170682216
	pesos_i(10175) := b"1111111111111111_1111111111111111_1110100010110111_1010110111100001"; -- -0.09094727752706683
	pesos_i(10176) := b"1111111111111111_1111111111111111_1111110111011101_1000010101101101"; -- -0.008338604761544181
	pesos_i(10177) := b"1111111111111111_1111111111111111_1110110100000100_0010011101000011"; -- -0.07415537467244879
	pesos_i(10178) := b"0000000000000000_0000000000000000_0000011111101100_1111110001101001"; -- 0.03095986894871456
	pesos_i(10179) := b"1111111111111111_1111111111111111_1110000000001001_0000111000010010"; -- -0.12486183228672462
	pesos_i(10180) := b"0000000000000000_0000000000000000_0001000101000101_0100100011101100"; -- 0.06746345300208313
	pesos_i(10181) := b"1111111111111111_1111111111111111_1111001001111010_0101001011011011"; -- -0.05282098921098243
	pesos_i(10182) := b"1111111111111111_1111111111111111_1101100101010011_0011011010000110"; -- -0.15107402067966538
	pesos_i(10183) := b"1111111111111111_1111111111111111_1110001111000110_1101011011000100"; -- -0.11024720877164103
	pesos_i(10184) := b"0000000000000000_0000000000000000_0001001011110111_1001100001010101"; -- 0.07409050052975713
	pesos_i(10185) := b"1111111111111111_1111111111111111_1101111100111011_0100010010011110"; -- -0.12800189144840898
	pesos_i(10186) := b"0000000000000000_0000000000000000_0000110100110000_0000011110011011"; -- 0.05151412527565952
	pesos_i(10187) := b"0000000000000000_0000000000000000_0000101011000010_1100101101000010"; -- 0.04203482023290936
	pesos_i(10188) := b"1111111111111111_1111111111111111_1110001000000100_1111000101000010"; -- -0.1171120847010968
	pesos_i(10189) := b"0000000000000000_0000000000000000_0000110010011110_1000001001001010"; -- 0.04929365458976693
	pesos_i(10190) := b"0000000000000000_0000000000000000_0001111101100101_1001101101111001"; -- 0.12264415453736424
	pesos_i(10191) := b"0000000000000000_0000000000000000_0010000010100111_0010101110101101"; -- 0.12755082101706594
	pesos_i(10192) := b"1111111111111111_1111111111111111_1101101110010001_1101100001010010"; -- -0.14230583186161944
	pesos_i(10193) := b"1111111111111111_1111111111111111_1110010010100101_0101000111110101"; -- -0.10685241471333816
	pesos_i(10194) := b"1111111111111111_1111111111111111_1110001110000100_0111000111101101"; -- -0.11126029924422014
	pesos_i(10195) := b"0000000000000000_0000000000000000_0010100010110100_0111111001101010"; -- 0.15900411679575704
	pesos_i(10196) := b"1111111111111111_1111111111111111_1110101100110001_0111101001111100"; -- -0.08127626873286603
	pesos_i(10197) := b"1111111111111111_1111111111111111_1110000010100011_0001111110010111"; -- -0.12251093448902448
	pesos_i(10198) := b"0000000000000000_0000000000000000_0001000111101000_1101111001001010"; -- 0.06995953851854957
	pesos_i(10199) := b"0000000000000000_0000000000000000_0010001001111000_1110000110101110"; -- 0.13465700626868457
	pesos_i(10200) := b"0000000000000000_0000000000000000_0001000100111111_0101010010000001"; -- 0.06737259043739137
	pesos_i(10201) := b"0000000000000000_0000000000000000_0001110100001110_0001000000110011"; -- 0.11349583854517525
	pesos_i(10202) := b"1111111111111111_1111111111111111_1111110110111001_1000101111010000"; -- -0.008887540574021146
	pesos_i(10203) := b"0000000000000000_0000000000000000_0001100011111110_0100000101100111"; -- 0.097629630632663
	pesos_i(10204) := b"1111111111111111_1111111111111111_1110110100000100_1010010100100010"; -- -0.07414787209302831
	pesos_i(10205) := b"0000000000000000_0000000000000000_0001000111011010_0111000110101000"; -- 0.0697394403853286
	pesos_i(10206) := b"1111111111111111_1111111111111111_1110110011011010_1000010010010001"; -- -0.07479068231696019
	pesos_i(10207) := b"1111111111111111_1111111111111111_1111111001000011_1001110010011100"; -- -0.006780826395256093
	pesos_i(10208) := b"1111111111111111_1111111111111111_1110100111101000_1011110110111010"; -- -0.08629240238286799
	pesos_i(10209) := b"0000000000000000_0000000000000000_0010001010010001_0010011011011010"; -- 0.1350273401132366
	pesos_i(10210) := b"1111111111111111_1111111111111111_1101111000100000_0011111000100000"; -- -0.1323205157712264
	pesos_i(10211) := b"1111111111111111_1111111111111111_1110011111000101_0010000101100101"; -- -0.09464827813820689
	pesos_i(10212) := b"0000000000000000_0000000000000000_0000110010101100_0010001000000111"; -- 0.04950153979460236
	pesos_i(10213) := b"1111111111111111_1111111111111111_1110001001011011_0000110001101110"; -- -0.11579820940210288
	pesos_i(10214) := b"1111111111111111_1111111111111111_1110101010111011_0000000010101111"; -- -0.08308406571037419
	pesos_i(10215) := b"1111111111111111_1111111111111111_1111111110100001_1100111100101110"; -- -0.0014372360817457405
	pesos_i(10216) := b"0000000000000000_0000000000000000_0001011100011000_1000000010110101"; -- 0.09021763253797854
	pesos_i(10217) := b"1111111111111111_1111111111111111_1111011100111111_0011100000111111"; -- -0.034191593858792536
	pesos_i(10218) := b"1111111111111111_1111111111111111_1111001111010110_0101001010100011"; -- -0.04751094351565566
	pesos_i(10219) := b"0000000000000000_0000000000000000_0001000111110101_0011111011010010"; -- 0.07014839775698187
	pesos_i(10220) := b"1111111111111111_1111111111111111_1110111101110101_0110000111001010"; -- -0.06461514311246326
	pesos_i(10221) := b"0000000000000000_0000000000000000_0001111100100110_1011110000100001"; -- 0.12168479738679176
	pesos_i(10222) := b"1111111111111111_1111111111111111_1110101110110110_0101011011110011"; -- -0.0792489678951277
	pesos_i(10223) := b"0000000000000000_0000000000000000_0001011100001100_0010111000011011"; -- 0.09002960345364844
	pesos_i(10224) := b"0000000000000000_0000000000000000_0001101010100110_0101101000000000"; -- 0.10410082333318517
	pesos_i(10225) := b"0000000000000000_0000000000000000_0001110110000101_0011110110011110"; -- 0.11531434151674212
	pesos_i(10226) := b"1111111111111111_1111111111111111_1111110001000001_0110001000000001"; -- -0.014627337276905596
	pesos_i(10227) := b"1111111111111111_1111111111111111_1111100100110010_1111010010001000"; -- -0.026566235382255877
	pesos_i(10228) := b"0000000000000000_0000000000000000_0010000000100101_1001100101000001"; -- 0.12557370991545674
	pesos_i(10229) := b"0000000000000000_0000000000000000_0000000100011101_1001110010100001"; -- 0.004358090787951393
	pesos_i(10230) := b"0000000000000000_0000000000000000_0000000111111100_0101000111001010"; -- 0.007756339779239665
	pesos_i(10231) := b"1111111111111111_1111111111111111_1111111101011011_1101111010110101"; -- -0.002504425709508137
	pesos_i(10232) := b"1111111111111111_1111111111111111_1111101011100000_0101010111110100"; -- -0.020014408057734967
	pesos_i(10233) := b"0000000000000000_0000000000000000_0000101111111111_0010011001010010"; -- 0.046862025393661716
	pesos_i(10234) := b"0000000000000000_0000000000000000_0000010101101101_1100000101110000"; -- 0.0212059877627251
	pesos_i(10235) := b"1111111111111111_1111111111111111_1101110111111110_0110010101001001"; -- -0.1328369805998394
	pesos_i(10236) := b"1111111111111111_1111111111111111_1101111000011101_0011100101000100"; -- -0.13236658186102945
	pesos_i(10237) := b"1111111111111111_1111111111111111_1111011010001000_1100101011011110"; -- -0.036975212932920144
	pesos_i(10238) := b"1111111111111111_1111111111111111_1101111001111010_0101001100010011"; -- -0.1309459762125572
	pesos_i(10239) := b"1111111111111111_1111111111111111_1110100010001100_0100011010101011"; -- -0.09160955737191155
	pesos_i(10240) := b"1111111111111111_1111111111111111_1110100011000101_0010010011111011"; -- -0.09074181445121769
	pesos_i(10241) := b"1111111111111111_1111111111111111_1110101010011010_1101100000111011"; -- -0.0835747581279464
	pesos_i(10242) := b"0000000000000000_0000000000000000_0000011010000000_0011110101111100"; -- 0.02539428967990135
	pesos_i(10243) := b"1111111111111111_1111111111111111_1110011001010111_0011000011100001"; -- -0.10023207184949236
	pesos_i(10244) := b"0000000000000000_0000000000000000_0001110010111100_1000110111111000"; -- 0.11225211444689291
	pesos_i(10245) := b"0000000000000000_0000000000000000_0010000100101110_0110100001111101"; -- 0.12961438219517374
	pesos_i(10246) := b"0000000000000000_0000000000000000_0001100101010111_1100111000110100"; -- 0.09899605523262921
	pesos_i(10247) := b"1111111111111111_1111111111111111_1101110100001111_1110100011001100"; -- -0.13647599244839773
	pesos_i(10248) := b"0000000000000000_0000000000000000_0001111000000000_0101101000111100"; -- 0.11719287843410608
	pesos_i(10249) := b"0000000000000000_0000000000000000_0001001101100101_1000011001100111"; -- 0.07576789874217203
	pesos_i(10250) := b"1111111111111111_1111111111111111_1111010101010101_1110001101110011"; -- -0.04165819595109916
	pesos_i(10251) := b"1111111111111111_1111111111111111_1101111011111001_0010110011000001"; -- -0.12901039397271064
	pesos_i(10252) := b"1111111111111111_1111111111111111_1110111110011001_1001001111100101"; -- -0.06406284000507206
	pesos_i(10253) := b"1111111111111111_1111111111111111_1111000001110110_1100001001000101"; -- -0.06068788349466381
	pesos_i(10254) := b"0000000000000000_0000000000000000_0010001111000101_1011110001001001"; -- 0.13973595415392484
	pesos_i(10255) := b"1111111111111111_1111111111111111_1110101111010100_0111111111111111"; -- -0.07878875753181833
	pesos_i(10256) := b"1111111111111111_1111111111111111_1110111111100000_1011010111000111"; -- -0.06297744639027442
	pesos_i(10257) := b"1111111111111111_1111111111111111_1110110110100011_1001110101000100"; -- -0.07172219362273792
	pesos_i(10258) := b"1111111111111111_1111111111111111_1110111000110010_1000010101100111"; -- -0.06954160904351177
	pesos_i(10259) := b"0000000000000000_0000000000000000_0010010110100011_0000101001101001"; -- 0.14701905319719757
	pesos_i(10260) := b"1111111111111111_1111111111111111_1110001111110101_1011000010110110"; -- -0.10953231397203034
	pesos_i(10261) := b"0000000000000000_0000000000000000_0000110010000011_0111110001101111"; -- 0.048881318073602124
	pesos_i(10262) := b"0000000000000000_0000000000000000_0010010000110011_0100100011100000"; -- 0.14140754187692006
	pesos_i(10263) := b"1111111111111111_1111111111111111_1110101110001110_1100111100111100"; -- -0.07985214971230334
	pesos_i(10264) := b"1111111111111111_1111111111111111_1111011011111000_0000111111001001"; -- -0.035277379355001644
	pesos_i(10265) := b"1111111111111111_1111111111111111_1110111000111101_0010100001100011"; -- -0.0693793065884543
	pesos_i(10266) := b"1111111111111111_1111111111111111_1110110000111000_1110100111000011"; -- -0.07725657443148261
	pesos_i(10267) := b"0000000000000000_0000000000000000_0000110010101101_0110011001000110"; -- 0.04952086655494011
	pesos_i(10268) := b"1111111111111111_1111111111111111_1111110111001111_1001000110010100"; -- -0.008551503639714098
	pesos_i(10269) := b"1111111111111111_1111111111111111_1111001110110000_1110111101101101"; -- -0.04808143213012021
	pesos_i(10270) := b"1111111111111111_1111111111111111_1110001110010100_0100101100100111"; -- -0.11101846985496036
	pesos_i(10271) := b"1111111111111111_1111111111111111_1110100000011111_1011011011001011"; -- -0.09326608231393077
	pesos_i(10272) := b"1111111111111111_1111111111111111_1111101010010101_0101001000111101"; -- -0.021159038707089187
	pesos_i(10273) := b"1111111111111111_1111111111111111_1101110011011011_1111010110101011"; -- -0.13726868231819866
	pesos_i(10274) := b"0000000000000000_0000000000000000_0010000111110100_0010110000101110"; -- 0.13263202773231555
	pesos_i(10275) := b"1111111111111111_1111111111111111_1110011010001001_1111101001011011"; -- -0.09945712348084376
	pesos_i(10276) := b"0000000000000000_0000000000000000_0001000110000001_1000000010111110"; -- 0.06838230733445853
	pesos_i(10277) := b"0000000000000000_0000000000000000_0000000101011101_0011000100101101"; -- 0.005328248427913129
	pesos_i(10278) := b"0000000000000000_0000000000000000_0001010000100101_0001110100111001"; -- 0.0786913169066551
	pesos_i(10279) := b"1111111111111111_1111111111111111_1110101010111000_0101110000001001"; -- -0.08312439708546482
	pesos_i(10280) := b"1111111111111111_1111111111111111_1101101001111100_1110111000000001"; -- -0.14653122410745215
	pesos_i(10281) := b"1111111111111111_1111111111111111_1110011111111100_1100101100101011"; -- -0.09379892550183937
	pesos_i(10282) := b"0000000000000000_0000000000000000_0000100011011101_0010000100101011"; -- 0.03462416927158455
	pesos_i(10283) := b"0000000000000000_0000000000000000_0001000011101011_1011101011111110"; -- 0.06609696101149358
	pesos_i(10284) := b"0000000000000000_0000000000000000_0001100001000010_1011001111100100"; -- 0.09476780230505402
	pesos_i(10285) := b"0000000000000000_0000000000000000_0000011111110000_1011110101101110"; -- 0.031017150236856847
	pesos_i(10286) := b"1111111111111111_1111111111111111_1110100111110100_1011100011011101"; -- -0.08610958674641225
	pesos_i(10287) := b"0000000000000000_0000000000000000_0010011011100000_1101010100110100"; -- 0.15186817662812888
	pesos_i(10288) := b"0000000000000000_0000000000000000_0000010000100100_0001001101101011"; -- 0.016175473747159032
	pesos_i(10289) := b"1111111111111111_1111111111111111_1111100011011011_0101001111000110"; -- -0.027903331912704707
	pesos_i(10290) := b"1111111111111111_1111111111111111_1110011110010101_0000100010011110"; -- -0.09538217672765001
	pesos_i(10291) := b"0000000000000000_0000000000000000_0000100000110001_0101111100000101"; -- 0.03200334420844333
	pesos_i(10292) := b"0000000000000000_0000000000000000_0000000001110100_0011100100111001"; -- 0.0017734303204209793
	pesos_i(10293) := b"1111111111111111_1111111111111111_1110011110011010_1010100000000001"; -- -0.09529638268310116
	pesos_i(10294) := b"1111111111111111_1111111111111111_1111111010010000_1000010001000101"; -- -0.005607350591424544
	pesos_i(10295) := b"1111111111111111_1111111111111111_1111111100100001_0111110101001101"; -- -0.0033952413652600473
	pesos_i(10296) := b"1111111111111111_1111111111111111_1110110011101010_1000110010110101"; -- -0.07454605666524955
	pesos_i(10297) := b"0000000000000000_0000000000000000_0000110100111111_0111110001100011"; -- 0.05174996780671566
	pesos_i(10298) := b"1111111111111111_1111111111111111_1101111101100100_1000001100001101"; -- -0.1273725599051427
	pesos_i(10299) := b"0000000000000000_0000000000000000_0010000110110111_0101101101010001"; -- 0.13170405126794563
	pesos_i(10300) := b"0000000000000000_0000000000000000_0000101101110101_1110000000100010"; -- 0.04476738769265689
	pesos_i(10301) := b"1111111111111111_1111111111111111_1101101001101110_0100001110000110"; -- -0.1467550085376702
	pesos_i(10302) := b"0000000000000000_0000000000000000_0000011100110110_1011100001010011"; -- 0.02817871112118577
	pesos_i(10303) := b"0000000000000000_0000000000000000_0001011001001010_0010010001000101"; -- 0.08706881231588869
	pesos_i(10304) := b"1111111111111111_1111111111111111_1110001001101110_0000011010010110"; -- -0.11550864065612737
	pesos_i(10305) := b"0000000000000000_0000000000000000_0000011001110100_0100010101110010"; -- 0.02521165884552783
	pesos_i(10306) := b"0000000000000000_0000000000000000_0000011100001010_0011011110101011"; -- 0.027499656018128985
	pesos_i(10307) := b"1111111111111111_1111111111111111_1111111010000010_1100010110100110"; -- -0.005817076581222583
	pesos_i(10308) := b"0000000000000000_0000000000000000_0001100010000011_0000011001011110"; -- 0.09574928092759454
	pesos_i(10309) := b"0000000000000000_0000000000000000_0000110010110001_1011010011011100"; -- 0.049586585656445095
	pesos_i(10310) := b"0000000000000000_0000000000000000_0001011101000000_0111111111000000"; -- 0.09082792700174602
	pesos_i(10311) := b"0000000000000000_0000000000000000_0010001101111000_1110110110100101"; -- 0.1385639693373769
	pesos_i(10312) := b"0000000000000000_0000000000000000_0001110000001001_0011110010111101"; -- 0.10951594948515964
	pesos_i(10313) := b"0000000000000000_0000000000000000_0000001111011101_1101001110010110"; -- 0.015103553958814351
	pesos_i(10314) := b"1111111111111111_1111111111111111_1110000010100011_0100100011101001"; -- -0.12250847166208431
	pesos_i(10315) := b"0000000000000000_0000000000000000_0000000001100111_0110001100011000"; -- 0.0015775618294676971
	pesos_i(10316) := b"0000000000000000_0000000000000000_0000010010110110_0110111001101001"; -- 0.01840868065359279
	pesos_i(10317) := b"0000000000000000_0000000000000000_0010001111000010_0011011010011100"; -- 0.1396822101106634
	pesos_i(10318) := b"1111111111111111_1111111111111111_1111001110100100_0000110111111101"; -- -0.04827797488463437
	pesos_i(10319) := b"1111111111111111_1111111111111111_1110111000010010_0110010000100111"; -- -0.07003187213776914
	pesos_i(10320) := b"0000000000000000_0000000000000000_0001100001111100_1100100000111111"; -- 0.09565402546082019
	pesos_i(10321) := b"1111111111111111_1111111111111111_1111000100011111_1111000111101110"; -- -0.05810630746696703
	pesos_i(10322) := b"0000000000000000_0000000000000000_0001110011000111_1100101111100011"; -- 0.11242365162340451
	pesos_i(10323) := b"1111111111111111_1111111111111111_1110011111001100_0111111000000110"; -- -0.0945359454404838
	pesos_i(10324) := b"1111111111111111_1111111111111111_1110011111000101_1011111101010001"; -- -0.09463886514673191
	pesos_i(10325) := b"1111111111111111_1111111111111111_1110110110111010_0000010000101001"; -- -0.07138036730295938
	pesos_i(10326) := b"1111111111111111_1111111111111111_1110010101010101_0111010100110101"; -- -0.10416476687553154
	pesos_i(10327) := b"1111111111111111_1111111111111111_1110101111000000_0000001111010011"; -- -0.07910133454174546
	pesos_i(10328) := b"0000000000000000_0000000000000000_0000110101001111_1101010001100000"; -- 0.05199935297869617
	pesos_i(10329) := b"0000000000000000_0000000000000000_0001011000111110_1111111011110001"; -- 0.08689874061926872
	pesos_i(10330) := b"0000000000000000_0000000000000000_0001010010011011_0011000000001001"; -- 0.08049297547305322
	pesos_i(10331) := b"1111111111111111_1111111111111111_1111010000011100_0100110110110001"; -- -0.04644312310213157
	pesos_i(10332) := b"1111111111111111_1111111111111111_1111111000011100_1100000110110101"; -- -0.0073737080900994996
	pesos_i(10333) := b"1111111111111111_1111111111111111_1110011010111000_0011000011100000"; -- -0.09875196969860876
	pesos_i(10334) := b"1111111111111111_1111111111111111_1110011111010110_0111110110001101"; -- -0.09438338577744099
	pesos_i(10335) := b"1111111111111111_1111111111111111_1110010101100100_0011100101101100"; -- -0.1039394485303361
	pesos_i(10336) := b"1111111111111111_1111111111111111_1111001001011010_1101001001010110"; -- -0.053301672045696934
	pesos_i(10337) := b"1111111111111111_1111111111111111_1101110110000101_1110000011011011"; -- -0.13467592871886755
	pesos_i(10338) := b"1111111111111111_1111111111111111_1110010111001011_0101100000010001"; -- -0.10236596674094353
	pesos_i(10339) := b"0000000000000000_0000000000000000_0001111000111101_1111100010010111"; -- 0.11813310313467972
	pesos_i(10340) := b"1111111111111111_1111111111111111_1110011101110001_1010100010111010"; -- -0.09592194994472468
	pesos_i(10341) := b"1111111111111111_1111111111111111_1110110111011100_1010001001000010"; -- -0.07085214512742602
	pesos_i(10342) := b"1111111111111111_1111111111111111_1101010111001110_0010000011010110"; -- -0.16482348238523825
	pesos_i(10343) := b"0000000000000000_0000000000000000_0010000000001110_1100010100011100"; -- 0.12522537165446662
	pesos_i(10344) := b"0000000000000000_0000000000000000_0001110111100100_1001001010101001"; -- 0.11676899554198636
	pesos_i(10345) := b"1111111111111111_1111111111111111_1110101111010101_1010010101010111"; -- -0.07877127288880152
	pesos_i(10346) := b"0000000000000000_0000000000000000_0000011001000001_0001101000001101"; -- 0.02443087396864296
	pesos_i(10347) := b"0000000000000000_0000000000000000_0000000000110100_1110100001010011"; -- 0.0008073046738914432
	pesos_i(10348) := b"1111111111111111_1111111111111111_1111111000011001_0000000001010010"; -- -0.007431011067893805
	pesos_i(10349) := b"1111111111111111_1111111111111111_1111100110111001_1110101000111111"; -- -0.024506911976459295
	pesos_i(10350) := b"0000000000000000_0000000000000000_0000011101101100_1011001100100111"; -- 0.02900237752085819
	pesos_i(10351) := b"1111111111111111_1111111111111111_1111101110000011_0010010101110101"; -- -0.017530115990778607
	pesos_i(10352) := b"1111111111111111_1111111111111111_1110010111011011_0100010100110001"; -- -0.10212295115056909
	pesos_i(10353) := b"0000000000000000_0000000000000000_0001100001010111_0100000101111101"; -- 0.0950814180295062
	pesos_i(10354) := b"0000000000000000_0000000000000000_0001001011101101_1000110001010111"; -- 0.07393719792716276
	pesos_i(10355) := b"0000000000000000_0000000000000000_0001010011001010_0010010100111101"; -- 0.08120949504049906
	pesos_i(10356) := b"0000000000000000_0000000000000000_0010001000011011_1110000010111110"; -- 0.133237883011646
	pesos_i(10357) := b"0000000000000000_0000000000000000_0000100010111000_0100010010001010"; -- 0.034061702508636674
	pesos_i(10358) := b"1111111111111111_1111111111111111_1111010110111011_1001000100101101"; -- -0.040106703328917914
	pesos_i(10359) := b"1111111111111111_1111111111111111_1111001110000010_1110000011011000"; -- -0.04878420558988646
	pesos_i(10360) := b"0000000000000000_0000000000000000_0010001000100000_1101011011011110"; -- 0.13331358839977453
	pesos_i(10361) := b"1111111111111111_1111111111111111_1111000101111001_0110011010000111"; -- -0.05674132549490622
	pesos_i(10362) := b"1111111111111111_1111111111111111_1110101110000001_0110111001100001"; -- -0.08005628717728117
	pesos_i(10363) := b"0000000000000000_0000000000000000_0010011100111001_0100110100011010"; -- 0.15321809658823596
	pesos_i(10364) := b"1111111111111111_1111111111111111_1101110000010111_1101010111110010"; -- -0.14026129560502837
	pesos_i(10365) := b"1111111111111111_1111111111111111_1110100100110110_1010101110100001"; -- -0.08900954560695472
	pesos_i(10366) := b"0000000000000000_0000000000000000_0010001100101010_0001010111110010"; -- 0.13736092728635038
	pesos_i(10367) := b"0000000000000000_0000000000000000_0001110001101101_1111000101001101"; -- 0.1110525905783149
	pesos_i(10368) := b"1111111111111111_1111111111111111_1111100000110010_1110010101000011"; -- -0.030473395508616875
	pesos_i(10369) := b"0000000000000000_0000000000000000_0000010010110111_1000010001101110"; -- 0.018425251878569523
	pesos_i(10370) := b"0000000000000000_0000000000000000_0010001111101001_1001001111000111"; -- 0.14028285617923064
	pesos_i(10371) := b"1111111111111111_1111111111111111_1110000111101010_0001001000101110"; -- -0.1175221096979339
	pesos_i(10372) := b"0000000000000000_0000000000000000_0001010001101011_1101010100111101"; -- 0.07977040048879752
	pesos_i(10373) := b"1111111111111111_1111111111111111_1110100001000111_1110110000011010"; -- -0.09265255322831913
	pesos_i(10374) := b"1111111111111111_1111111111111111_1101110011111110_1100011011100001"; -- -0.13673741347764426
	pesos_i(10375) := b"0000000000000000_0000000000000000_0010011001011010_1111001010100110"; -- 0.14982525397976484
	pesos_i(10376) := b"1111111111111111_1111111111111111_1101111001101100_1101001011001100"; -- -0.1311519864226595
	pesos_i(10377) := b"1111111111111111_1111111111111111_1110110101110011_1110100101111001"; -- -0.07245007311810318
	pesos_i(10378) := b"0000000000000000_0000000000000000_0010010110001001_1001110101011010"; -- 0.1466310830013624
	pesos_i(10379) := b"0000000000000000_0000000000000000_0001101100110101_0000111001000101"; -- 0.10627831634368824
	pesos_i(10380) := b"1111111111111111_1111111111111111_1111011100010001_1001100111101101"; -- -0.034887675880008726
	pesos_i(10381) := b"1111111111111111_1111111111111111_1110001010010110_1100000000110110"; -- -0.11488722494433208
	pesos_i(10382) := b"0000000000000000_0000000000000000_0001001011001010_1010111101100000"; -- 0.07340522860359587
	pesos_i(10383) := b"1111111111111111_1111111111111111_1110010100010111_0010000100011100"; -- -0.10511582439398638
	pesos_i(10384) := b"1111111111111111_1111111111111111_1101111111001110_1110000101011000"; -- -0.12574950794805118
	pesos_i(10385) := b"0000000000000000_0000000000000000_0000010010111000_1000100001111001"; -- 0.018440751558702746
	pesos_i(10386) := b"0000000000000000_0000000000000000_0000110100111010_1111010001101001"; -- 0.05168082768686271
	pesos_i(10387) := b"0000000000000000_0000000000000000_0000011100000101_1000100100101011"; -- 0.02742821989718983
	pesos_i(10388) := b"0000000000000000_0000000000000000_0010001110101111_1101010110111101"; -- 0.13940177783784946
	pesos_i(10389) := b"1111111111111111_1111111111111111_1111111110100101_0001100011010001"; -- -0.0013870707191897486
	pesos_i(10390) := b"1111111111111111_1111111111111111_1101111011110000_1100110011100011"; -- -0.1291381784436599
	pesos_i(10391) := b"0000000000000000_0000000000000000_0000011010000111_0100001000111110"; -- 0.02550138479191768
	pesos_i(10392) := b"1111111111111111_1111111111111111_1111111011010000_1001111100100101"; -- -0.00462918611740233
	pesos_i(10393) := b"1111111111111111_1111111111111111_1111001010101001_0110011011100110"; -- -0.052102631481719376
	pesos_i(10394) := b"1111111111111111_1111111111111111_1111001111111011_0100110010100101"; -- -0.0469467256778342
	pesos_i(10395) := b"1111111111111111_1111111111111111_1110110000100101_0100100000001101"; -- -0.07755613014934785
	pesos_i(10396) := b"0000000000000000_0000000000000000_0000001000000001_0111100001101100"; -- 0.00783493638605492
	pesos_i(10397) := b"1111111111111111_1111111111111111_1101110110001001_1011010101100110"; -- -0.13461748369381446
	pesos_i(10398) := b"0000000000000000_0000000000000000_0001011100011001_0101111011100110"; -- 0.09023087617131441
	pesos_i(10399) := b"1111111111111111_1111111111111111_1110101001001111_1001000010110110"; -- -0.08472343032400048
	pesos_i(10400) := b"0000000000000000_0000000000000000_0010000111000111_1010001001100000"; -- 0.1319524273726303
	pesos_i(10401) := b"1111111111111111_1111111111111111_1111111000111110_0011100010000101"; -- -0.0068630862370601614
	pesos_i(10402) := b"1111111111111111_1111111111111111_1111101000010000_0011101000000011"; -- -0.023189901548553306
	pesos_i(10403) := b"1111111111111111_1111111111111111_1111001010101100_1011011111011001"; -- -0.05205203017951587
	pesos_i(10404) := b"1111111111111111_1111111111111111_1110101001010101_1000001110101110"; -- -0.08463265422767494
	pesos_i(10405) := b"1111111111111111_1111111111111111_1110111111000011_1100111100110101"; -- -0.06341843553212154
	pesos_i(10406) := b"1111111111111111_1111111111111111_1110110100000101_0010000110100000"; -- -0.0741404518784479
	pesos_i(10407) := b"0000000000000000_0000000000000000_0001111000100001_1101000111111011"; -- 0.1177035557719998
	pesos_i(10408) := b"1111111111111111_1111111111111111_1111111011110011_0001001001100110"; -- -0.004103517556049377
	pesos_i(10409) := b"1111111111111111_1111111111111111_1111010101010000_1001001001000011"; -- -0.04173932890323581
	pesos_i(10410) := b"1111111111111111_1111111111111111_1110001110011100_0110111111010000"; -- -0.11089421425469864
	pesos_i(10411) := b"1111111111111111_1111111111111111_1110011010000010_1111101000100011"; -- -0.09956394807854124
	pesos_i(10412) := b"0000000000000000_0000000000000000_0000110101001001_1010101100101110"; -- 0.05190534463478377
	pesos_i(10413) := b"1111111111111111_1111111111111111_1111100001101100_1110101011111111"; -- -0.0295880439757568
	pesos_i(10414) := b"0000000000000000_0000000000000000_0010100001110100_1000001101111011"; -- 0.15802785640939518
	pesos_i(10415) := b"1111111111111111_1111111111111111_1110000100011101_0100111101001011"; -- -0.12064651878088008
	pesos_i(10416) := b"1111111111111111_1111111111111111_1111000010100110_1000110001001111"; -- -0.05995867792463435
	pesos_i(10417) := b"1111111111111111_1111111111111111_1111001011110011_1101001001011111"; -- -0.050967075123059084
	pesos_i(10418) := b"0000000000000000_0000000000000000_0010000110010110_1110101110001100"; -- 0.13120910813959646
	pesos_i(10419) := b"0000000000000000_0000000000000000_0000001110010100_1100011100101101"; -- 0.013988922695217945
	pesos_i(10420) := b"0000000000000000_0000000000000000_0001001000011101_1000011011001110"; -- 0.07076303982315124
	pesos_i(10421) := b"1111111111111111_1111111111111111_1111000110000101_0101111010001110"; -- -0.05655869520732592
	pesos_i(10422) := b"0000000000000000_0000000000000000_0000111111011111_0010010011011101"; -- 0.06199865709679268
	pesos_i(10423) := b"1111111111111111_1111111111111111_1110011011000101_1010111111100000"; -- -0.09854603558503641
	pesos_i(10424) := b"0000000000000000_0000000000000000_0001011110100100_0111011111110111"; -- 0.09235334190365092
	pesos_i(10425) := b"1111111111111111_1111111111111111_1111011100000001_0001000110000011"; -- -0.035139947374517456
	pesos_i(10426) := b"1111111111111111_1111111111111111_1110100100111111_1001111010001111"; -- -0.08887299551255545
	pesos_i(10427) := b"0000000000000000_0000000000000000_0001000101101010_1000110110001100"; -- 0.06803211856429846
	pesos_i(10428) := b"0000000000000000_0000000000000000_0010001010000001_0100110110110011"; -- 0.13478551503611572
	pesos_i(10429) := b"1111111111111111_1111111111111111_1110101011010101_1010010001001111"; -- -0.0826775843875035
	pesos_i(10430) := b"0000000000000000_0000000000000000_0001110101001010_0010001001011011"; -- 0.1144124481563249
	pesos_i(10431) := b"1111111111111111_1111111111111111_1101111010011010_0100100101000001"; -- -0.13045828031884868
	pesos_i(10432) := b"0000000000000000_0000000000000000_0010001101101011_0001111000110000"; -- 0.13835323965202667
	pesos_i(10433) := b"1111111111111111_1111111111111111_1110001011001110_0011101001100011"; -- -0.11404070928466005
	pesos_i(10434) := b"1111111111111111_1111111111111111_1110001111111101_0001001001001110"; -- -0.10941968524661648
	pesos_i(10435) := b"0000000000000000_0000000000000000_0001100011010011_0101110110100100"; -- 0.09697518579801319
	pesos_i(10436) := b"0000000000000000_0000000000000000_0001111101101000_0101100111101011"; -- 0.12268602366505066
	pesos_i(10437) := b"0000000000000000_0000000000000000_0000110001110101_1001100010011010"; -- 0.04866937406826598
	pesos_i(10438) := b"1111111111111111_1111111111111111_1111101100001011_0000000011001011"; -- -0.019363356068519976
	pesos_i(10439) := b"0000000000000000_0000000000000000_0010001111111011_0011110100101101"; -- 0.14055235248772824
	pesos_i(10440) := b"0000000000000000_0000000000000000_0000001001010011_1010000011111010"; -- 0.009088574411777784
	pesos_i(10441) := b"1111111111111111_1111111111111111_1101110001000100_1010000001001010"; -- -0.13957784837844917
	pesos_i(10442) := b"1111111111111111_1111111111111111_1111101000101011_0010100001101110"; -- -0.022778962257685966
	pesos_i(10443) := b"1111111111111111_1111111111111111_1111101011100100_0011100010001111"; -- -0.01995512501536011
	pesos_i(10444) := b"1111111111111111_1111111111111111_1111011110010010_1011110101001001"; -- -0.03291718455975436
	pesos_i(10445) := b"0000000000000000_0000000000000000_0001101001110111_1111000010100110"; -- 0.10339263970707369
	pesos_i(10446) := b"0000000000000000_0000000000000000_0000101011101001_0001110111100110"; -- 0.04261957997382327
	pesos_i(10447) := b"0000000000000000_0000000000000000_0000100011010101_1011111010011111"; -- 0.03451148390830584
	pesos_i(10448) := b"0000000000000000_0000000000000000_0000110001110110_0110100111000101"; -- 0.04868184149541042
	pesos_i(10449) := b"1111111111111111_1111111111111111_1101110010001110_1100110111010100"; -- -0.13844598365107302
	pesos_i(10450) := b"1111111111111111_1111111111111111_1101110011000100_0011010110101000"; -- -0.13763107913409212
	pesos_i(10451) := b"0000000000000000_0000000000000000_0010110001101011_1111010100001100"; -- 0.17352229642149364
	pesos_i(10452) := b"1111111111111111_1111111111111111_1110001010101001_0011001000000011"; -- -0.11460578371743164
	pesos_i(10453) := b"1111111111111111_1111111111111111_1110101000011011_1001100011001011"; -- -0.08551640542010533
	pesos_i(10454) := b"0000000000000000_0000000000000000_0010001100001010_1010100101010011"; -- 0.136881430343154
	pesos_i(10455) := b"1111111111111111_1111111111111111_1110010101011001_1010001100010001"; -- -0.10410099830306492
	pesos_i(10456) := b"1111111111111111_1111111111111111_1101111010111000_1101111001101010"; -- -0.12999162595968622
	pesos_i(10457) := b"0000000000000000_0000000000000000_0010100110001001_0010010001011010"; -- 0.16224887076689673
	pesos_i(10458) := b"1111111111111111_1111111111111111_1101100101101100_1011001100001110"; -- -0.15068512837603143
	pesos_i(10459) := b"0000000000000000_0000000000000000_0001010011011001_1001110110011011"; -- 0.08144555133733843
	pesos_i(10460) := b"1111111111111111_1111111111111111_1111001000110011_1000111100110011"; -- -0.05390076632183977
	pesos_i(10461) := b"1111111111111111_1111111111111111_1110100000110000_1111111101011010"; -- -0.09300235806854695
	pesos_i(10462) := b"1111111111111111_1111111111111111_1110111010101001_1100110010010000"; -- -0.06772157166918019
	pesos_i(10463) := b"1111111111111111_1111111111111111_1110101000110001_1100011000110011"; -- -0.08517800572434558
	pesos_i(10464) := b"1111111111111111_1111111111111111_1101011000011001_1111011101110000"; -- -0.1636662818878831
	pesos_i(10465) := b"0000000000000000_0000000000000000_0000110100100010_1000010100010010"; -- 0.05130798040501392
	pesos_i(10466) := b"1111111111111111_1111111111111111_1110011101001100_0000000101110001"; -- -0.0964964960159494
	pesos_i(10467) := b"1111111111111111_1111111111111111_1110010101100010_1000011001001110"; -- -0.10396538349824667
	pesos_i(10468) := b"0000000000000000_0000000000000000_0001100000010010_1110100111010100"; -- 0.09403859542634095
	pesos_i(10469) := b"1111111111111111_1111111111111111_1101110101011110_1100110011110010"; -- -0.1352722081133454
	pesos_i(10470) := b"0000000000000000_0000000000000000_0000010001010111_1011110010111101"; -- 0.016963764361585056
	pesos_i(10471) := b"0000000000000000_0000000000000000_0010010000100001_0010010000101100"; -- 0.1411306959835984
	pesos_i(10472) := b"1111111111111111_1111111111111111_1111110000100110_0100110001110110"; -- -0.015040608487264916
	pesos_i(10473) := b"0000000000000000_0000000000000000_0000111110111001_1110101111001111"; -- 0.0614306813337166
	pesos_i(10474) := b"1111111111111111_1111111111111111_1110001000111110_0001111010101100"; -- -0.11623962686695302
	pesos_i(10475) := b"1111111111111111_1111111111111111_1101111110110011_0100111000001101"; -- -0.1261702746506438
	pesos_i(10476) := b"1111111111111111_1111111111111111_1111010110110110_1111010010111010"; -- -0.04017706364865918
	pesos_i(10477) := b"0000000000000000_0000000000000000_0001001110101010_1101100001001100"; -- 0.07682563646147406
	pesos_i(10478) := b"1111111111111111_1111111111111111_1111110111011010_0001101101001110"; -- -0.008390706417509688
	pesos_i(10479) := b"0000000000000000_0000000000000000_0000101101010000_0001100110111110"; -- 0.044190987449446134
	pesos_i(10480) := b"1111111111111111_1111111111111111_1110110110100010_1110001011111000"; -- -0.07173329779489766
	pesos_i(10481) := b"1111111111111111_1111111111111111_1111010001110101_0000011100011011"; -- -0.04508929820098684
	pesos_i(10482) := b"1111111111111111_1111111111111111_1110100011101010_0111111011111111"; -- -0.0901718737532067
	pesos_i(10483) := b"0000000000000000_0000000000000000_0000010101010001_0100011000100011"; -- 0.02077139239087659
	pesos_i(10484) := b"0000000000000000_0000000000000000_0000000010011001_1111001111110110"; -- 0.0023491358982847977
	pesos_i(10485) := b"1111111111111111_1111111111111111_1110110100000011_0100100111110100"; -- -0.07416856579540114
	pesos_i(10486) := b"1111111111111111_1111111111111111_1111010001000001_0110101011000010"; -- -0.045876815555915815
	pesos_i(10487) := b"0000000000000000_0000000000000000_0000100110101001_0011001010100100"; -- 0.03773800377003124
	pesos_i(10488) := b"0000000000000000_0000000000000000_0000000110011111_0100100100100101"; -- 0.006336757244020643
	pesos_i(10489) := b"0000000000000000_0000000000000000_0001101001001111_1110100000111110"; -- 0.10278178715391835
	pesos_i(10490) := b"1111111111111111_1111111111111111_1110100000010111_1111000100100110"; -- -0.0933846743288089
	pesos_i(10491) := b"1111111111111111_1111111111111111_1111000110111000_0011110111001110"; -- -0.055782448895011445
	pesos_i(10492) := b"0000000000000000_0000000000000000_0001001110001101_1111101101110010"; -- 0.07638522659628695
	pesos_i(10493) := b"1111111111111111_1111111111111111_1111010101110100_0011101110111001"; -- -0.041195170624468175
	pesos_i(10494) := b"1111111111111111_1111111111111111_1110111100101000_1100100101100111"; -- -0.06578389394055084
	pesos_i(10495) := b"0000000000000000_0000000000000000_0010000110100011_1101110000111111"; -- 0.13140656032844208
	pesos_i(10496) := b"1111111111111111_1111111111111111_1101111011100001_1110100000110110"; -- -0.12936543154155325
	pesos_i(10497) := b"1111111111111111_1111111111111111_1101100111010111_1111111110101000"; -- -0.14904787193642036
	pesos_i(10498) := b"0000000000000000_0000000000000000_0000001100010010_1000100000001000"; -- 0.012001516289588864
	pesos_i(10499) := b"1111111111111111_1111111111111111_1110001101110110_1100011110000010"; -- -0.11146882138164087
	pesos_i(10500) := b"0000000000000000_0000000000000000_0000100100011100_1101010001001001"; -- 0.035596149368980805
	pesos_i(10501) := b"1111111111111111_1111111111111111_1111001010100100_1000110000101000"; -- -0.05217670470541154
	pesos_i(10502) := b"0000000000000000_0000000000000000_0001000010011001_0100000000100011"; -- 0.06483841746111439
	pesos_i(10503) := b"1111111111111111_1111111111111111_1110010010110111_0101001101100000"; -- -0.10657767212984062
	pesos_i(10504) := b"1111111111111111_1111111111111111_1111001100000110_0010101100000101"; -- -0.050687133110860566
	pesos_i(10505) := b"0000000000000000_0000000000000000_0000110001111011_0101000011111110"; -- 0.04875665850947585
	pesos_i(10506) := b"1111111111111111_1111111111111111_1110110011101010_0100010010110110"; -- -0.07455034780269476
	pesos_i(10507) := b"1111111111111111_1111111111111111_1110010111111000_0101000101000011"; -- -0.10167972675211188
	pesos_i(10508) := b"1111111111111111_1111111111111111_1111101000101010_1001100111000000"; -- -0.022787466698125668
	pesos_i(10509) := b"0000000000000000_0000000000000000_0001111101101101_1100000111100100"; -- 0.12276851483263918
	pesos_i(10510) := b"1111111111111111_1111111111111111_1110001001101011_1000011111010000"; -- -0.11554671452746283
	pesos_i(10511) := b"0000000000000000_0000000000000000_0000101000000100_0010010101000100"; -- 0.03912575646650114
	pesos_i(10512) := b"1111111111111111_1111111111111111_1110011100011110_1010001101001010"; -- -0.09718875353275078
	pesos_i(10513) := b"1111111111111111_1111111111111111_1111100000101100_1101010011000101"; -- -0.03056593113516779
	pesos_i(10514) := b"1111111111111111_1111111111111111_1110001000111110_0100001110000011"; -- -0.11623743103302744
	pesos_i(10515) := b"0000000000000000_0000000000000000_0001000100111100_0110001001100100"; -- 0.06732764181364587
	pesos_i(10516) := b"0000000000000000_0000000000000000_0000111011101000_1011010001111100"; -- 0.05823829666279737
	pesos_i(10517) := b"0000000000000000_0000000000000000_0001111011000100_1011100001110110"; -- 0.12018921740276552
	pesos_i(10518) := b"1111111111111111_1111111111111111_1110110110111110_0110101110001100"; -- -0.07131316975903294
	pesos_i(10519) := b"0000000000000000_0000000000000000_0010001110110000_0100010010101001"; -- 0.1394083892572539
	pesos_i(10520) := b"1111111111111111_1111111111111111_1111001110111000_0101011110000111"; -- -0.04796841574145235
	pesos_i(10521) := b"0000000000000000_0000000000000000_0001110010111111_1000000010010111"; -- 0.11229709322013573
	pesos_i(10522) := b"0000000000000000_0000000000000000_0001000000001011_1100011011001101"; -- 0.06267969611018692
	pesos_i(10523) := b"0000000000000000_0000000000000000_0001110000100110_1001111101011000"; -- 0.10996433159917778
	pesos_i(10524) := b"0000000000000000_0000000000000000_0000111101000010_1010011100100000"; -- 0.059610791539477986
	pesos_i(10525) := b"0000000000000000_0000000000000000_0001011101011100_1111011101000111"; -- 0.09126229752302327
	pesos_i(10526) := b"0000000000000000_0000000000000000_0010010100101110_0000100010011000"; -- 0.1452336664714709
	pesos_i(10527) := b"1111111111111111_1111111111111111_1111010100011010_1111111011000111"; -- -0.04255683566025123
	pesos_i(10528) := b"0000000000000000_0000000000000000_0001110010010011_1001001001011101"; -- 0.11162676601013806
	pesos_i(10529) := b"0000000000000000_0000000000000000_0000111010111110_0010111011011011"; -- 0.057589462726593
	pesos_i(10530) := b"1111111111111111_1111111111111111_1110000001011100_1000001101110001"; -- -0.12358835688272164
	pesos_i(10531) := b"0000000000000000_0000000000000000_0001001100111011_1100010110001010"; -- 0.07513079290550712
	pesos_i(10532) := b"0000000000000000_0000000000000000_0001110100011001_0011010001010111"; -- 0.11366583952656911
	pesos_i(10533) := b"0000000000000000_0000000000000000_0010010000011100_0000110010001000"; -- 0.14105299312583716
	pesos_i(10534) := b"1111111111111111_1111111111111111_1111110101111110_0101111011101110"; -- -0.009790484352903134
	pesos_i(10535) := b"1111111111111111_1111111111111111_1111101001100101_1000011001110101"; -- -0.021888348001555463
	pesos_i(10536) := b"0000000000000000_0000000000000000_0010001100111010_0001101001111010"; -- 0.13760533786085574
	pesos_i(10537) := b"0000000000000000_0000000000000000_0000011101110011_1011111100111010"; -- 0.029109908682851814
	pesos_i(10538) := b"1111111111111111_1111111111111111_1110010011101011_1100101011100011"; -- -0.1057770915008142
	pesos_i(10539) := b"1111111111111111_1111111111111111_1110111000110110_1100001100100111"; -- -0.06947689351369794
	pesos_i(10540) := b"0000000000000000_0000000000000000_0000011100100001_1010101010111100"; -- 0.02785746668112928
	pesos_i(10541) := b"0000000000000000_0000000000000000_0000100000100100_0110110000011010"; -- 0.031805759862228916
	pesos_i(10542) := b"1111111111111111_1111111111111111_1110101001101010_1010101011000011"; -- -0.08430989007146468
	pesos_i(10543) := b"0000000000000000_0000000000000000_0001110111011100_0110101100010010"; -- 0.11664456557283945
	pesos_i(10544) := b"1111111111111111_1111111111111111_1110100011110001_0010011111001000"; -- -0.09007026076016164
	pesos_i(10545) := b"1111111111111111_1111111111111111_1111110011010110_1011000111011100"; -- -0.012349018007645735
	pesos_i(10546) := b"0000000000000000_0000000000000000_0000111011101001_1000111011111001"; -- 0.05825131957865026
	pesos_i(10547) := b"0000000000000000_0000000000000000_0001100100101011_1000000011111110"; -- 0.09832006649519999
	pesos_i(10548) := b"0000000000000000_0000000000000000_0000111010111100_0001110001000110"; -- 0.057557837580807625
	pesos_i(10549) := b"1111111111111111_1111111111111111_1110011100001011_1111011111011101"; -- -0.09747362962969315
	pesos_i(10550) := b"0000000000000000_0000000000000000_0000111100111101_0100110011111100"; -- 0.059529124643862404
	pesos_i(10551) := b"0000000000000000_0000000000000000_0000111001010001_1111001000011101"; -- 0.05593789306526151
	pesos_i(10552) := b"1111111111111111_1111111111111111_1110001000000010_0101011101001100"; -- -0.11715177923294108
	pesos_i(10553) := b"0000000000000000_0000000000000000_0000110111110010_1100011000111110"; -- 0.054485693154241545
	pesos_i(10554) := b"1111111111111111_1111111111111111_1110111000111100_0000100000101100"; -- -0.06939648550923064
	pesos_i(10555) := b"0000000000000000_0000000000000000_0000011011010000_1010101000011000"; -- 0.026621466586116117
	pesos_i(10556) := b"1111111111111111_1111111111111111_1111101001011001_1110100000100010"; -- -0.02206563158888493
	pesos_i(10557) := b"0000000000000000_0000000000000000_0000011010001110_0000101110000101"; -- 0.02560493471773185
	pesos_i(10558) := b"1111111111111111_1111111111111111_1110111000111100_0000011100111001"; -- -0.06939654220926855
	pesos_i(10559) := b"0000000000000000_0000000000000000_0000011110010001_1001101011001000"; -- 0.029565500022844176
	pesos_i(10560) := b"1111111111111111_1111111111111111_1111011111101010_1000011010101011"; -- -0.031577666520321755
	pesos_i(10561) := b"0000000000000000_0000000000000000_0001001000000110_1101011001111111"; -- 0.07041683760891634
	pesos_i(10562) := b"1111111111111111_1111111111111111_1110000110111101_0000100100101100"; -- -0.11820929220277289
	pesos_i(10563) := b"0000000000000000_0000000000000000_0001011110101100_0100110110101111"; -- 0.09247289200464243
	pesos_i(10564) := b"1111111111111111_1111111111111111_1110011110000010_1011011110110010"; -- -0.09566165833382081
	pesos_i(10565) := b"1111111111111111_1111111111111111_1110000011000101_1010111001000011"; -- -0.12198363168270246
	pesos_i(10566) := b"1111111111111111_1111111111111111_1111111111110101_0000110001011001"; -- -0.00016711072650813796
	pesos_i(10567) := b"0000000000000000_0000000000000000_0001101000001010_0110101011110000"; -- 0.10172146176963519
	pesos_i(10568) := b"1111111111111111_1111111111111111_1111010101111110_1101100000001101"; -- -0.041033264833948827
	pesos_i(10569) := b"0000000000000000_0000000000000000_0001001010100100_1100111110100101"; -- 0.07282731790777178
	pesos_i(10570) := b"1111111111111111_1111111111111111_1111001000000101_0100110110011100"; -- -0.05460658025603774
	pesos_i(10571) := b"1111111111111111_1111111111111111_1110110000101111_1100000001110001"; -- -0.07739636644321443
	pesos_i(10572) := b"1111111111111111_1111111111111111_1101101111000111_0000001001101101"; -- -0.14149460629498475
	pesos_i(10573) := b"0000000000000000_0000000000000000_0000010101000101_0010000101110110"; -- 0.02058610092917464
	pesos_i(10574) := b"0000000000000000_0000000000000000_0001101101001101_0100110000001111"; -- 0.10664821029050868
	pesos_i(10575) := b"0000000000000000_0000000000000000_0000000110000101_1100010111110110"; -- 0.0059474683151967385
	pesos_i(10576) := b"0000000000000000_0000000000000000_0010000011101110_1111100000010010"; -- 0.12864637797542852
	pesos_i(10577) := b"1111111111111111_1111111111111111_1110000101101011_1011101110110011"; -- -0.11944987185051155
	pesos_i(10578) := b"0000000000000000_0000000000000000_0010000110100110_1001000011010011"; -- 0.13144784110121777
	pesos_i(10579) := b"0000000000000000_0000000000000000_0001110010001010_1001111111010010"; -- 0.11149023885151102
	pesos_i(10580) := b"1111111111111111_1111111111111111_1101111101001010_0110010111101010"; -- -0.12777102506414953
	pesos_i(10581) := b"0000000000000000_0000000000000000_0001011111100110_1001101111111100"; -- 0.0933625689454531
	pesos_i(10582) := b"0000000000000000_0000000000000000_0001111010110110_1010111111111101"; -- 0.11997508931424229
	pesos_i(10583) := b"1111111111111111_1111111111111111_1110010100111110_0001101110010001"; -- -0.10452106203618271
	pesos_i(10584) := b"1111111111111111_1111111111111111_1111000010111111_0000101110110110"; -- -0.059584873310155974
	pesos_i(10585) := b"0000000000000000_0000000000000000_0001110001001001_0000101110110001"; -- 0.11048958853078804
	pesos_i(10586) := b"1111111111111111_1111111111111111_1110100111010000_1000010000111100"; -- -0.08666203998065047
	pesos_i(10587) := b"1111111111111111_1111111111111111_1110010001100001_0010011000010100"; -- -0.10789262793379098
	pesos_i(10588) := b"0000000000000000_0000000000000000_0000000001001110_0001100111100001"; -- 0.0011917280608176042
	pesos_i(10589) := b"1111111111111111_1111111111111111_1101111100000000_0001111011000001"; -- -0.12890441687856272
	pesos_i(10590) := b"1111111111111111_1111111111111111_1110000001000101_1101101010011100"; -- -0.1239341133218609
	pesos_i(10591) := b"0000000000000000_0000000000000000_0001101011001011_0000001100100001"; -- 0.10466022075979424
	pesos_i(10592) := b"1111111111111111_1111111111111111_1111100011001011_0010110100101010"; -- -0.028149773778570458
	pesos_i(10593) := b"1111111111111111_1111111111111111_1101110001001000_0110101100011111"; -- -0.13951998224099255
	pesos_i(10594) := b"1111111111111111_1111111111111111_1110110010111101_1000101011101000"; -- -0.0752328094790333
	pesos_i(10595) := b"1111111111111111_1111111111111111_1111001010111000_0001010111000101"; -- -0.05187858521729022
	pesos_i(10596) := b"0000000000000000_0000000000000000_0001110100001111_0010000110100101"; -- 0.11351213713045576
	pesos_i(10597) := b"0000000000000000_0000000000000000_0000010011101000_1111100111110000"; -- 0.01917993651528307
	pesos_i(10598) := b"0000000000000000_0000000000000000_0000001000001100_1100110101111000"; -- 0.008007852300595933
	pesos_i(10599) := b"1111111111111111_1111111111111111_1110000001001010_1110100111100111"; -- -0.12385690802885961
	pesos_i(10600) := b"1111111111111111_1111111111111111_1110001100110101_1100010000111110"; -- -0.11246083730043126
	pesos_i(10601) := b"1111111111111111_1111111111111111_1101101110101110_1100100010011000"; -- -0.14186426447911324
	pesos_i(10602) := b"0000000000000000_0000000000000000_0000010110010000_0100100001111000"; -- 0.021732835115989356
	pesos_i(10603) := b"0000000000000000_0000000000000000_0001101000000011_1100010100010101"; -- 0.10162002347117036
	pesos_i(10604) := b"0000000000000000_0000000000000000_0001100100111101_1010010001001011"; -- 0.09859682876506531
	pesos_i(10605) := b"1111111111111111_1111111111111111_1110000001010000_1100010111100110"; -- -0.12376750128753769
	pesos_i(10606) := b"0000000000000000_0000000000000000_0000111111001001_1101101010111000"; -- 0.061673803154232106
	pesos_i(10607) := b"0000000000000000_0000000000000000_0000010100010101_1111111000100011"; -- 0.01986683220953719
	pesos_i(10608) := b"0000000000000000_0000000000000000_0000100111100001_0111000100101110"; -- 0.03859622364117185
	pesos_i(10609) := b"0000000000000000_0000000000000000_0001111101000101_0001001111110000"; -- 0.12214779488234231
	pesos_i(10610) := b"1111111111111111_1111111111111111_1110111110100100_0101000111001100"; -- -0.06389893317184947
	pesos_i(10611) := b"1111111111111111_1111111111111111_1110101011011110_0011100011101110"; -- -0.08254665552990911
	pesos_i(10612) := b"0000000000000000_0000000000000000_0001000011010110_0100011001011101"; -- 0.06576957483517056
	pesos_i(10613) := b"0000000000000000_0000000000000000_0010010010000100_0001100101010100"; -- 0.1426406698910446
	pesos_i(10614) := b"1111111111111111_1111111111111111_1101100101100100_0001111101100111"; -- -0.15081599937443405
	pesos_i(10615) := b"1111111111111111_1111111111111111_1110101111101001_0111110110110011"; -- -0.07846845990991552
	pesos_i(10616) := b"1111111111111111_1111111111111111_1110000000000100_0110010110000100"; -- -0.12493291407289661
	pesos_i(10617) := b"0000000000000000_0000000000000000_0001000101001111_0100100110010011"; -- 0.06761607978821763
	pesos_i(10618) := b"1111111111111111_1111111111111111_1101110100101010_1100101110101110"; -- -0.13606574058052096
	pesos_i(10619) := b"1111111111111111_1111111111111111_1111011101010010_1010011110011001"; -- -0.033895039678777675
	pesos_i(10620) := b"1111111111111111_1111111111111111_1110001111111000_0100001100101101"; -- -0.10949306637717258
	pesos_i(10621) := b"0000000000000000_0000000000000000_0000110101100100_0101100101000110"; -- 0.0523124499631486
	pesos_i(10622) := b"0000000000000000_0000000000000000_0001101101111110_1000010100011011"; -- 0.10739929109195197
	pesos_i(10623) := b"0000000000000000_0000000000000000_0001010101111111_0011101101011011"; -- 0.08397265417220241
	pesos_i(10624) := b"1111111111111111_1111111111111111_1111001001110011_1101000111110100"; -- -0.052920225124565914
	pesos_i(10625) := b"0000000000000000_0000000000000000_0001100000111101_1111011100100011"; -- 0.09469551663954344
	pesos_i(10626) := b"1111111111111111_1111111111111111_1101101110101011_1010011010101101"; -- -0.14191206244893234
	pesos_i(10627) := b"1111111111111111_1111111111111111_1111101110000011_0011110010101011"; -- -0.017528732544045286
	pesos_i(10628) := b"0000000000000000_0000000000000000_0000111001100101_0000011110000100"; -- 0.0562290856839228
	pesos_i(10629) := b"1111111111111111_1111111111111111_1110101111010000_0011000101111000"; -- -0.07885447320314654
	pesos_i(10630) := b"1111111111111111_1111111111111111_1111001000010011_0001100001000000"; -- -0.05439613769518013
	pesos_i(10631) := b"1111111111111111_1111111111111111_1111010011110111_1100001011111100"; -- -0.04309445701239702
	pesos_i(10632) := b"0000000000000000_0000000000000000_0000100001110001_0010001011000011"; -- 0.03297631514004005
	pesos_i(10633) := b"0000000000000000_0000000000000000_0001101100111010_0110011101011100"; -- 0.10635992054996965
	pesos_i(10634) := b"1111111111111111_1111111111111111_1110111010111101_1101000001101001"; -- -0.06741616674375274
	pesos_i(10635) := b"0000000000000000_0000000000000000_0000111101010110_0100010011100010"; -- 0.059910111542194396
	pesos_i(10636) := b"1111111111111111_1111111111111111_1111111001110001_1110001000110010"; -- -0.00607477455324078
	pesos_i(10637) := b"1111111111111111_1111111111111111_1111011011100100_1110010111010000"; -- -0.03556979829676585
	pesos_i(10638) := b"0000000000000000_0000000000000000_0001001100001111_0001011010110011"; -- 0.07444898484809466
	pesos_i(10639) := b"1111111111111111_1111111111111111_1110100000011111_1111010010000010"; -- -0.09326240367269488
	pesos_i(10640) := b"1111111111111111_1111111111111111_1110010011011100_1000000000000001"; -- -0.10601043689516432
	pesos_i(10641) := b"0000000000000000_0000000000000000_0000000100010111_1111110010011010"; -- 0.004272258483491794
	pesos_i(10642) := b"0000000000000000_0000000000000000_0000110010111111_0111111111100101"; -- 0.04979705173248331
	pesos_i(10643) := b"0000000000000000_0000000000000000_0001110111010011_0101001110110111"; -- 0.11650584428410417
	pesos_i(10644) := b"0000000000000000_0000000000000000_0010011101100011_1100110011010100"; -- 0.15386657885978156
	pesos_i(10645) := b"0000000000000000_0000000000000000_0001001001001111_0111110000001010"; -- 0.07152533773253762
	pesos_i(10646) := b"1111111111111111_1111111111111111_1111010011110101_1001000101011010"; -- -0.043127933049544084
	pesos_i(10647) := b"1111111111111111_1111111111111111_1110111111110101_0000000001101111"; -- -0.06266782094324932
	pesos_i(10648) := b"1111111111111111_1111111111111111_1101010110011001_1000011001011110"; -- -0.165626146463201
	pesos_i(10649) := b"1111111111111111_1111111111111111_1110101111011100_0000011010000001"; -- -0.07867392883130896
	pesos_i(10650) := b"0000000000000000_0000000000000000_0000110100010110_1010011001010101"; -- 0.051126857418381084
	pesos_i(10651) := b"1111111111111111_1111111111111111_1110101011110111_0111000110101100"; -- -0.08216180374697295
	pesos_i(10652) := b"0000000000000000_0000000000000000_0000111010110000_1011011011110111"; -- 0.05738395248167342
	pesos_i(10653) := b"1111111111111111_1111111111111111_1110010001110011_0011010000111011"; -- -0.10761712607794363
	pesos_i(10654) := b"1111111111111111_1111111111111111_1110110100011100_0000000011001000"; -- -0.07379145722556797
	pesos_i(10655) := b"0000000000000000_0000000000000000_0000001001001001_1110000101111000"; -- 0.008939830557139681
	pesos_i(10656) := b"1111111111111111_1111111111111111_1101111111000100_1110010001111100"; -- -0.1259019086386315
	pesos_i(10657) := b"0000000000000000_0000000000000000_0000010111000000_1101100010100000"; -- 0.02247384928206115
	pesos_i(10658) := b"1111111111111111_1111111111111111_1111011110101000_0011010010101000"; -- -0.03258963486412373
	pesos_i(10659) := b"1111111111111111_1111111111111111_1110010100110111_1100000100010101"; -- -0.10461800801515461
	pesos_i(10660) := b"1111111111111111_1111111111111111_1110110110001010_1000101111010111"; -- -0.0721047021093229
	pesos_i(10661) := b"0000000000000000_0000000000000000_0000101101111101_1000000001011001"; -- 0.04488374880124964
	pesos_i(10662) := b"1111111111111111_1111111111111111_1110101011011111_0001001110110111"; -- -0.08253361503756529
	pesos_i(10663) := b"0000000000000000_0000000000000000_0001010110101010_0111111001110101"; -- 0.08463278167190884
	pesos_i(10664) := b"0000000000000000_0000000000000000_0001101010100110_0110101111001100"; -- 0.10410188428765839
	pesos_i(10665) := b"1111111111111111_1111111111111111_1111101110001100_1010010110101011"; -- -0.017385144934881885
	pesos_i(10666) := b"1111111111111111_1111111111111111_1111101101001100_0101100111101011"; -- -0.018366222430071716
	pesos_i(10667) := b"1111111111111111_1111111111111111_1110110000100001_1101000011101000"; -- -0.07760900810308304
	pesos_i(10668) := b"1111111111111111_1111111111111111_1101101111001100_1011011000100001"; -- -0.14140760130993954
	pesos_i(10669) := b"0000000000000000_0000000000000000_0001101101000001_0110000100011011"; -- 0.10646635924847503
	pesos_i(10670) := b"1111111111111111_1111111111111111_1101111001101011_1001011010101000"; -- -0.13117082972727795
	pesos_i(10671) := b"0000000000000000_0000000000000000_0010010010010111_1011010110010010"; -- 0.1429398996148673
	pesos_i(10672) := b"0000000000000000_0000000000000000_0001111110101100_1100101100111011"; -- 0.12373037523194287
	pesos_i(10673) := b"0000000000000000_0000000000000000_0000111101011100_1010011000000110"; -- 0.060007454404940035
	pesos_i(10674) := b"0000000000000000_0000000000000000_0000010100101011_1010001110101100"; -- 0.02019713352999486
	pesos_i(10675) := b"1111111111111111_1111111111111111_1111001111101111_0000011100111001"; -- -0.04713396900500516
	pesos_i(10676) := b"0000000000000000_0000000000000000_0010011010111010_0000011110011011"; -- 0.15127608802667936
	pesos_i(10677) := b"0000000000000000_0000000000000000_0001011111110011_1011111111000110"; -- 0.09356306634549662
	pesos_i(10678) := b"1111111111111111_1111111111111111_1111111100110101_0110100111011101"; -- -0.0030912241333889237
	pesos_i(10679) := b"0000000000000000_0000000000000000_0000001101011011_0101000000010100"; -- 0.013112072718509726
	pesos_i(10680) := b"1111111111111111_1111111111111111_1111100001100001_1111111000001000"; -- -0.029754756046661026
	pesos_i(10681) := b"0000000000000000_0000000000000000_0000110001011111_1100011111100011"; -- 0.048336499201156964
	pesos_i(10682) := b"1111111111111111_1111111111111111_1110001110100010_1100100000110110"; -- -0.1107973925821102
	pesos_i(10683) := b"1111111111111111_1111111111111111_1111101000100101_0101001110000110"; -- -0.022867946311330403
	pesos_i(10684) := b"0000000000000000_0000000000000000_0001001110011100_0100011111111001"; -- 0.07660341094622337
	pesos_i(10685) := b"0000000000000000_0000000000000000_0001001010001110_1100111100111110"; -- 0.07249160067890542
	pesos_i(10686) := b"1111111111111111_1111111111111111_1110100010000010_0111001110011010"; -- -0.09175946713077184
	pesos_i(10687) := b"0000000000000000_0000000000000000_0010000001101101_0101100000000010"; -- 0.12666845377750025
	pesos_i(10688) := b"0000000000000000_0000000000000000_0010001011100000_1011011110101000"; -- 0.13624141558704508
	pesos_i(10689) := b"1111111111111111_1111111111111111_1110100011111110_0011101010011110"; -- -0.08987077380442153
	pesos_i(10690) := b"1111111111111111_1111111111111111_1110100111000101_0101000000010010"; -- -0.08683299608647971
	pesos_i(10691) := b"0000000000000000_0000000000000000_0001111101111001_0111001101110111"; -- 0.1229469456716226
	pesos_i(10692) := b"1111111111111111_1111111111111111_1111101011100000_1111101010000111"; -- -0.020004598648770466
	pesos_i(10693) := b"1111111111111111_1111111111111111_1111000100000101_0010000010111111"; -- -0.058515504301088185
	pesos_i(10694) := b"0000000000000000_0000000000000000_0001000111010110_0110000100111011"; -- 0.06967742628791378
	pesos_i(10695) := b"1111111111111111_1111111111111111_1110110111111010_1110010000000000"; -- -0.0703904628732472
	pesos_i(10696) := b"0000000000000000_0000000000000000_0000011111110100_1100101011111001"; -- 0.031078992547781892
	pesos_i(10697) := b"0000000000000000_0000000000000000_0001001001011111_1100000000110011"; -- 0.07177354083094294
	pesos_i(10698) := b"0000000000000000_0000000000000000_0000101110111110_1001111000001011"; -- 0.04587733992860337
	pesos_i(10699) := b"1111111111111111_1111111111111111_1110111001010001_1001110101110111"; -- -0.06906715239501643
	pesos_i(10700) := b"0000000000000000_0000000000000000_0000011110100001_1010100000001111"; -- 0.02981043208134434
	pesos_i(10701) := b"0000000000000000_0000000000000000_0000011010110011_0000111001011010"; -- 0.026169678760592074
	pesos_i(10702) := b"0000000000000000_0000000000000000_0001101000001010_1001100011011100"; -- 0.10172419912025517
	pesos_i(10703) := b"1111111111111111_1111111111111111_1110100011010110_1010110010111011"; -- -0.09047432364818586
	pesos_i(10704) := b"1111111111111111_1111111111111111_1110000011111011_0000100000000000"; -- -0.12116956699240085
	pesos_i(10705) := b"0000000000000000_0000000000000000_0000000000111101_0101011010110001"; -- 0.0009359533189172272
	pesos_i(10706) := b"0000000000000000_0000000000000000_0000110001001010_1000010000111111"; -- 0.048012032964867536
	pesos_i(10707) := b"1111111111111111_1111111111111111_1110011100101010_1001110001101010"; -- -0.09700605787754309
	pesos_i(10708) := b"0000000000000000_0000000000000000_0000010001001011_0010000110111101"; -- 0.016771420065902716
	pesos_i(10709) := b"0000000000000000_0000000000000000_0010000100101010_1001001000000000"; -- 0.12955582149958525
	pesos_i(10710) := b"1111111111111111_1111111111111111_1110100111011011_1101010011100101"; -- -0.08648938574215197
	pesos_i(10711) := b"1111111111111111_1111111111111111_1110110110111010_0100111101001110"; -- -0.07137588823438382
	pesos_i(10712) := b"0000000000000000_0000000000000000_0000000000101001_1110101011000110"; -- 0.0006396038425380066
	pesos_i(10713) := b"1111111111111111_1111111111111111_1111110101101010_1001100101110011"; -- -0.01009217213945785
	pesos_i(10714) := b"1111111111111111_1111111111111111_1111001101101101_0100111101010000"; -- -0.04911331469102535
	pesos_i(10715) := b"1111111111111111_1111111111111111_1111001100011101_0001010111001101"; -- -0.050337445767545896
	pesos_i(10716) := b"0000000000000000_0000000000000000_0000110000111011_0001010110000001"; -- 0.04777655022081647
	pesos_i(10717) := b"0000000000000000_0000000000000000_0000100110000101_0111001001001110"; -- 0.037192481980996464
	pesos_i(10718) := b"0000000000000000_0000000000000000_0001110101011001_0101101111000110"; -- 0.11464475227281021
	pesos_i(10719) := b"0000000000000000_0000000000000000_0000010101000000_1011010101101001"; -- 0.020518625365840138
	pesos_i(10720) := b"0000000000000000_0000000000000000_0001110011000111_1001000110001100"; -- 0.11242017425141157
	pesos_i(10721) := b"1111111111111111_1111111111111111_1101110001011111_0001010000111100"; -- -0.13917420890020488
	pesos_i(10722) := b"0000000000000000_0000000000000000_0001101011000100_0101001011101001"; -- 0.10455816442604733
	pesos_i(10723) := b"0000000000000000_0000000000000000_0000101111000011_0000101010100110"; -- 0.045944848547291535
	pesos_i(10724) := b"1111111111111111_1111111111111111_1101101100101010_1010111010001110"; -- -0.14387997659802976
	pesos_i(10725) := b"0000000000000000_0000000000000000_0000011000100001_1011011010001011"; -- 0.02395192038124776
	pesos_i(10726) := b"0000000000000000_0000000000000000_0001011000101101_1010111101010011"; -- 0.08663459570319548
	pesos_i(10727) := b"1111111111111111_1111111111111111_1111100110010001_0111001111010010"; -- -0.025124322160044035
	pesos_i(10728) := b"1111111111111111_1111111111111111_1111110001101010_1001111111000010"; -- -0.01399804606249182
	pesos_i(10729) := b"1111111111111111_1111111111111111_1110100101100001_1111110000010011"; -- -0.0883486225556934
	pesos_i(10730) := b"1111111111111111_1111111111111111_1101101111010100_1100111010101100"; -- -0.14128406810865546
	pesos_i(10731) := b"0000000000000000_0000000000000000_0001111101101101_0101010011001001"; -- 0.12276201165831288
	pesos_i(10732) := b"1111111111111111_1111111111111111_1110001001111001_1011010110101110"; -- -0.1153303576217255
	pesos_i(10733) := b"1111111111111111_1111111111111111_1111101101010110_0010001011011110"; -- -0.01821691594842443
	pesos_i(10734) := b"0000000000000000_0000000000000000_0000100111111010_1011110101011000"; -- 0.03898223313640291
	pesos_i(10735) := b"0000000000000000_0000000000000000_0010001000101100_1011101111011100"; -- 0.13349508396412013
	pesos_i(10736) := b"0000000000000000_0000000000000000_0001000010001001_0100010001001110"; -- 0.0645945253555751
	pesos_i(10737) := b"1111111111111111_1111111111111111_1111010000111000_1100111000101000"; -- -0.046008220006348445
	pesos_i(10738) := b"0000000000000000_0000000000000000_0010011000001011_0111100011010101"; -- 0.14861254880017347
	pesos_i(10739) := b"0000000000000000_0000000000000000_0000111000110111_0011001011111111"; -- 0.05552977294042287
	pesos_i(10740) := b"0000000000000000_0000000000000000_0000111101000001_1100001010110100"; -- 0.05959717650606503
	pesos_i(10741) := b"1111111111111111_1111111111111111_1110111001110111_0010011011000010"; -- -0.06849439395256984
	pesos_i(10742) := b"1111111111111111_1111111111111111_1110100110101101_1100011000010101"; -- -0.08719217278003687
	pesos_i(10743) := b"1111111111111111_1111111111111111_1111110111001011_0011111110011101"; -- -0.00861742411777842
	pesos_i(10744) := b"1111111111111111_1111111111111111_1110101110010110_0100011100001110"; -- -0.07973819640217707
	pesos_i(10745) := b"1111111111111111_1111111111111111_1101110100101001_0110101101100010"; -- -0.13608673919535447
	pesos_i(10746) := b"0000000000000000_0000000000000000_0010000111011010_0001110000011111"; -- 0.1322343420802213
	pesos_i(10747) := b"0000000000000000_0000000000000000_0001000000101000_1010101100001100"; -- 0.06312054676513171
	pesos_i(10748) := b"1111111111111111_1111111111111111_1110100111100010_0010111001101010"; -- -0.08639249724502863
	pesos_i(10749) := b"0000000000000000_0000000000000000_0001110100110001_1111111000001100"; -- 0.11404407295728468
	pesos_i(10750) := b"1111111111111111_1111111111111111_1110100011101000_0101011100100010"; -- -0.09020476748108185
	pesos_i(10751) := b"0000000000000000_0000000000000000_0010000001010011_1101010111000110"; -- 0.12627922127646402
	pesos_i(10752) := b"1111111111111111_1111111111111111_1111010101110000_1000001110100100"; -- -0.041251919245791246
	pesos_i(10753) := b"1111111111111111_1111111111111111_1110011010000110_1101110000000010"; -- -0.09950470869185007
	pesos_i(10754) := b"0000000000000000_0000000000000000_0000010011110000_0010010001110010"; -- 0.019289281781268604
	pesos_i(10755) := b"0000000000000000_0000000000000000_0000011100001011_1100101110011001"; -- 0.027523732030656327
	pesos_i(10756) := b"1111111111111111_1111111111111111_1110011000111111_0010010111001100"; -- -0.10059894338705182
	pesos_i(10757) := b"1111111111111111_1111111111111111_1111110111110000_1110101001100000"; -- -0.008042670687832102
	pesos_i(10758) := b"0000000000000000_0000000000000000_0001111111010111_0110000100110101"; -- 0.12438018365392023
	pesos_i(10759) := b"0000000000000000_0000000000000000_0000010111000101_0111000100101011"; -- 0.022543976865848483
	pesos_i(10760) := b"0000000000000000_0000000000000000_0001000110001010_0001001110000101"; -- 0.0685131264447273
	pesos_i(10761) := b"1111111111111111_1111111111111111_1110101001110001_1101111011101101"; -- -0.08419996948878723
	pesos_i(10762) := b"1111111111111111_1111111111111111_1111111101011110_0110011010111101"; -- -0.00246580009808589
	pesos_i(10763) := b"0000000000000000_0000000000000000_0000100010110000_0111110100001100"; -- 0.033943000246083196
	pesos_i(10764) := b"1111111111111111_1111111111111111_1110110000101100_0000010000010011"; -- -0.07745337048524595
	pesos_i(10765) := b"0000000000000000_0000000000000000_0010011010100101_0110101010001000"; -- 0.15096154990336905
	pesos_i(10766) := b"0000000000000000_0000000000000000_0001100110100010_0010101010100101"; -- 0.10013071554132802
	pesos_i(10767) := b"1111111111111111_1111111111111111_1111000100100110_0001001001011101"; -- -0.05801282147984718
	pesos_i(10768) := b"1111111111111111_1111111111111111_1111101001101111_0110000011100000"; -- -0.02173800013623859
	pesos_i(10769) := b"1111111111111111_1111111111111111_1111000011110010_1011100011000101"; -- -0.058796359959736415
	pesos_i(10770) := b"1111111111111111_1111111111111111_1110110111001000_0111010001000011"; -- -0.07116006242047587
	pesos_i(10771) := b"1111111111111111_1111111111111111_1111011000111111_0010110111110011"; -- -0.03809845761801259
	pesos_i(10772) := b"1111111111111111_1111111111111111_1111011100011100_0111010111001110"; -- -0.03472198220104337
	pesos_i(10773) := b"0000000000000000_0000000000000000_0001001110000001_1011110101001001"; -- 0.0761984161271994
	pesos_i(10774) := b"1111111111111111_1111111111111111_1111100010001011_0010000010011011"; -- -0.029127084815561026
	pesos_i(10775) := b"0000000000000000_0000000000000000_0000000110111010_1110001100000110"; -- 0.006757916514007742
	pesos_i(10776) := b"0000000000000000_0000000000000000_0000000001001111_1001000011001000"; -- 0.0012140739950552784
	pesos_i(10777) := b"0000000000000000_0000000000000000_0001000011110010_0111111011001111"; -- 0.06620018541724149
	pesos_i(10778) := b"1111111111111111_1111111111111111_1110010011100111_1111111000101100"; -- -0.10583506993739263
	pesos_i(10779) := b"0000000000000000_0000000000000000_0000101101001110_0100000111101100"; -- 0.044162864903293374
	pesos_i(10780) := b"1111111111111111_1111111111111111_1101110110100001_0100100000101010"; -- -0.1342577835486511
	pesos_i(10781) := b"1111111111111111_1111111111111111_1111001011001100_0001010111100111"; -- -0.05157340150346528
	pesos_i(10782) := b"1111111111111111_1111111111111111_1111100000010111_1000110110000000"; -- -0.030890613703903985
	pesos_i(10783) := b"0000000000000000_0000000000000000_0000011101110101_0010011010101010"; -- 0.029131332946105152
	pesos_i(10784) := b"1111111111111111_1111111111111111_1101100010110010_1010100110100110"; -- -0.1535238236999643
	pesos_i(10785) := b"0000000000000000_0000000000000000_0001011100111000_1100001101111101"; -- 0.09070989408081064
	pesos_i(10786) := b"0000000000000000_0000000000000000_0001011010000100_0001000010100100"; -- 0.0879526520387923
	pesos_i(10787) := b"0000000000000000_0000000000000000_0001110110110101_1111100111100101"; -- 0.11605798560796236
	pesos_i(10788) := b"1111111111111111_1111111111111111_1110100011000000_1100010110110110"; -- -0.09080852808489706
	pesos_i(10789) := b"0000000000000000_0000000000000000_0001111110000011_0001000000101111"; -- 0.12309361600863322
	pesos_i(10790) := b"0000000000000000_0000000000000000_0001001001010101_0110101111000101"; -- 0.07161592060219021
	pesos_i(10791) := b"1111111111111111_1111111111111111_1111101010011000_0010010010100111"; -- -0.021115979402326394
	pesos_i(10792) := b"0000000000000000_0000000000000000_0000010111100011_1101000111111001"; -- 0.02300751050269919
	pesos_i(10793) := b"0000000000000000_0000000000000000_0000011000100001_0011110111000000"; -- 0.02394472053166291
	pesos_i(10794) := b"0000000000000000_0000000000000000_0001000101001010_1001111111011100"; -- 0.06754492882930543
	pesos_i(10795) := b"0000000000000000_0000000000000000_0001011010011110_1101100110010101"; -- 0.08836135761894563
	pesos_i(10796) := b"1111111111111111_1111111111111111_1101110001111011_0101000101001010"; -- -0.1387433236794765
	pesos_i(10797) := b"1111111111111111_1111111111111111_1110011001111011_0111110110011111"; -- -0.09967818133544425
	pesos_i(10798) := b"1111111111111111_1111111111111111_1110010001110010_1011000000100101"; -- -0.10762499891376677
	pesos_i(10799) := b"1111111111111111_1111111111111111_1111001010101001_0111101001101010"; -- -0.05210146828458525
	pesos_i(10800) := b"1111111111111111_1111111111111111_1101110101000111_0110110100010000"; -- -0.13562887537221016
	pesos_i(10801) := b"1111111111111111_1111111111111111_1111100100011010_1110100000000101"; -- -0.02693319214826066
	pesos_i(10802) := b"1111111111111111_1111111111111111_1110010111110011_1000101101000011"; -- -0.10175256363607352
	pesos_i(10803) := b"1111111111111111_1111111111111111_1110100111110010_1101010000100000"; -- -0.08613847945923675
	pesos_i(10804) := b"1111111111111111_1111111111111111_1101111000110011_0111100100101100"; -- -0.13202707943742492
	pesos_i(10805) := b"0000000000000000_0000000000000000_0000011110010111_1100010000111001"; -- 0.02965952284657463
	pesos_i(10806) := b"0000000000000000_0000000000000000_0001001100111110_1111111001001001"; -- 0.07517995149506998
	pesos_i(10807) := b"0000000000000000_0000000000000000_0010000010000110_0000111111110101"; -- 0.12704562888686424
	pesos_i(10808) := b"0000000000000000_0000000000000000_0001010001011100_1000111010011010"; -- 0.07953730821660006
	pesos_i(10809) := b"1111111111111111_1111111111111111_1111011111001110_1010101010010011"; -- -0.032002772484691376
	pesos_i(10810) := b"1111111111111111_1111111111111111_1110101010101010_0011100001101111"; -- -0.08334014209521566
	pesos_i(10811) := b"0000000000000000_0000000000000000_0001110110000001_0100111100010000"; -- 0.115254346334716
	pesos_i(10812) := b"0000000000000000_0000000000000000_0000100010011111_1101110110101010"; -- 0.03368935968260007
	pesos_i(10813) := b"0000000000000000_0000000000000000_0000011111100001_0110010110111111"; -- 0.030783041993941388
	pesos_i(10814) := b"0000000000000000_0000000000000000_0010010011001001_1001111011011010"; -- 0.14370148484465037
	pesos_i(10815) := b"1111111111111111_1111111111111111_1110111011111001_0111000000101001"; -- -0.06650637627392397
	pesos_i(10816) := b"0000000000000000_0000000000000000_0000011100001011_0011011100001010"; -- 0.027514877175135132
	pesos_i(10817) := b"0000000000000000_0000000000000000_0000000001111101_1111111011000100"; -- 0.0019225339635029035
	pesos_i(10818) := b"0000000000000000_0000000000000000_0001011001100110_0101100010010111"; -- 0.08749917684332185
	pesos_i(10819) := b"0000000000000000_0000000000000000_0000001011111101_1110110111000100"; -- 0.01168714548248018
	pesos_i(10820) := b"1111111111111111_1111111111111111_1111100011101011_1000110111101110"; -- -0.027655724984763267
	pesos_i(10821) := b"1111111111111111_1111111111111111_1110100100110011_1101000011110101"; -- -0.08905309684747488
	pesos_i(10822) := b"0000000000000000_0000000000000000_0001100000110011_1011001111001001"; -- 0.09453891419702849
	pesos_i(10823) := b"0000000000000000_0000000000000000_0001101010101001_1001000110110001"; -- 0.10414991932673247
	pesos_i(10824) := b"0000000000000000_0000000000000000_0001101011100101_1101001111010110"; -- 0.10506938920733218
	pesos_i(10825) := b"1111111111111111_1111111111111111_1101110110001101_1011010001101111"; -- -0.1345565059726293
	pesos_i(10826) := b"1111111111111111_1111111111111111_1101110001000011_1010111011101000"; -- -0.13959223598817372
	pesos_i(10827) := b"0000000000000000_0000000000000000_0001101010110001_0101011100001101"; -- 0.10426849421609843
	pesos_i(10828) := b"1111111111111111_1111111111111111_1111000100001101_1111100000010101"; -- -0.05838059900996215
	pesos_i(10829) := b"0000000000000000_0000000000000000_0001110110011000_0000110000011111"; -- 0.115601308373748
	pesos_i(10830) := b"0000000000000000_0000000000000000_0010011000111000_1110010100110110"; -- 0.1493056541758676
	pesos_i(10831) := b"0000000000000000_0000000000000000_0010010100110101_0111010010011100"; -- 0.14534691633305505
	pesos_i(10832) := b"0000000000000000_0000000000000000_0000010010010111_0000110101011000"; -- 0.017929872424774403
	pesos_i(10833) := b"1111111111111111_1111111111111111_1110111110001111_0011110010111100"; -- -0.06422062316468514
	pesos_i(10834) := b"1111111111111111_1111111111111111_1111100000101111_0010110110010001"; -- -0.03053012083554069
	pesos_i(10835) := b"0000000000000000_0000000000000000_0000101010011110_0100101101010010"; -- 0.041477878063728525
	pesos_i(10836) := b"0000000000000000_0000000000000000_0010011001100000_1111100011011110"; -- 0.14991717739784186
	pesos_i(10837) := b"0000000000000000_0000000000000000_0000101010001000_1001110001000110"; -- 0.0411470099379689
	pesos_i(10838) := b"1111111111111111_1111111111111111_1110111011100010_1111111101001011"; -- -0.06684879696111413
	pesos_i(10839) := b"0000000000000000_0000000000000000_0000110001000101_1110100000100110"; -- 0.04794169357308713
	pesos_i(10840) := b"1111111111111111_1111111111111111_1110110001011011_1010001000111011"; -- -0.07672678051718362
	pesos_i(10841) := b"1111111111111111_1111111111111111_1111000101110001_1111111000101001"; -- -0.05685435767236472
	pesos_i(10842) := b"0000000000000000_0000000000000000_0000010101011100_1000110010101000"; -- 0.020943442417360125
	pesos_i(10843) := b"1111111111111111_1111111111111111_1110001000101111_0010011001011101"; -- -0.11646805032060308
	pesos_i(10844) := b"0000000000000000_0000000000000000_0001101101111000_0010101101011110"; -- 0.10730238952566128
	pesos_i(10845) := b"0000000000000000_0000000000000000_0000101001100001_0111010000100111"; -- 0.04054952566390847
	pesos_i(10846) := b"0000000000000000_0000000000000000_0010001010110000_1011100010111101"; -- 0.13550905804032592
	pesos_i(10847) := b"1111111111111111_1111111111111111_1111111000100010_0000011010000100"; -- -0.0072933127622527155
	pesos_i(10848) := b"1111111111111111_1111111111111111_1101110101001001_0100110001010100"; -- -0.1356003087763796
	pesos_i(10849) := b"0000000000000000_0000000000000000_0000010011011101_0100101101100111"; -- 0.019001686655304054
	pesos_i(10850) := b"1111111111111111_1111111111111111_1101101100011001_0001010100010111"; -- -0.14414852322366692
	pesos_i(10851) := b"0000000000000000_0000000000000000_0001110000001000_0111000111010100"; -- 0.10950385503972074
	pesos_i(10852) := b"1111111111111111_1111111111111111_1111100111011010_1000101100111001"; -- -0.02400903558466085
	pesos_i(10853) := b"1111111111111111_1111111111111111_1101110001111111_0100000101100111"; -- -0.13868323544827263
	pesos_i(10854) := b"1111111111111111_1111111111111111_1110001100100001_0101111111101000"; -- -0.11277199345172256
	pesos_i(10855) := b"0000000000000000_0000000000000000_0001010000010110_1010001100101000"; -- 0.07847041820206999
	pesos_i(10856) := b"0000000000000000_0000000000000000_0000111101000101_0000111111010001"; -- 0.0596475491114249
	pesos_i(10857) := b"0000000000000000_0000000000000000_0000011001100000_0100100101001000"; -- 0.024906711660621073
	pesos_i(10858) := b"1111111111111111_1111111111111111_1111001010010100_0111101101110101"; -- -0.05242184054307123
	pesos_i(10859) := b"1111111111111111_1111111111111111_1111111101011011_0110010111001001"; -- -0.0025116332459163494
	pesos_i(10860) := b"1111111111111111_1111111111111111_1111100100011011_1101111111001000"; -- -0.026918424206355526
	pesos_i(10861) := b"1111111111111111_1111111111111111_1101100011011101_1000010011001100"; -- -0.15286989221465563
	pesos_i(10862) := b"1111111111111111_1111111111111111_1101101010101101_0100110011111110"; -- -0.1457931403703188
	pesos_i(10863) := b"1111111111111111_1111111111111111_1101110000010001_0001100100100000"; -- -0.1403641029591504
	pesos_i(10864) := b"0000000000000000_0000000000000000_0001010101001110_1001011111110111"; -- 0.08323049332892976
	pesos_i(10865) := b"0000000000000000_0000000000000000_0001101100101101_0000000110001010"; -- 0.10615548719617278
	pesos_i(10866) := b"0000000000000000_0000000000000000_0001001011101001_1010011100011111"; -- 0.07387775909578781
	pesos_i(10867) := b"0000000000000000_0000000000000000_0000011001010111_0111001010010010"; -- 0.024771843534234804
	pesos_i(10868) := b"0000000000000000_0000000000000000_0010001000101100_1110000100010110"; -- 0.13349730291794754
	pesos_i(10869) := b"1111111111111111_1111111111111111_1111011001011110_1010011110000110"; -- -0.03761818876441584
	pesos_i(10870) := b"0000000000000000_0000000000000000_0010001111000111_0010100111111011"; -- 0.13975775123965684
	pesos_i(10871) := b"0000000000000000_0000000000000000_0010001110111001_0010111011000100"; -- 0.13954441332024448
	pesos_i(10872) := b"0000000000000000_0000000000000000_0010010100101010_0000111010001100"; -- 0.145172986260145
	pesos_i(10873) := b"1111111111111111_1111111111111111_1110111111111010_0010111011001111"; -- -0.06258876263302748
	pesos_i(10874) := b"0000000000000000_0000000000000000_0000011110000110_0011011101011010"; -- 0.02939172686423331
	pesos_i(10875) := b"1111111111111111_1111111111111111_1101110010110101_0001101011101111"; -- -0.1378615537088178
	pesos_i(10876) := b"0000000000000000_0000000000000000_0000000011110101_1010100111100010"; -- 0.0037485290422707308
	pesos_i(10877) := b"1111111111111111_1111111111111111_1110101001000111_1001101001001011"; -- -0.0848449293476282
	pesos_i(10878) := b"0000000000000000_0000000000000000_0010100010011110_0100110101100100"; -- 0.15866550147522573
	pesos_i(10879) := b"0000000000000000_0000000000000000_0000010010100011_0111101100100100"; -- 0.018119522481368448
	pesos_i(10880) := b"1111111111111111_1111111111111111_1110011100100000_1010100100000101"; -- -0.09715789442434764
	pesos_i(10881) := b"0000000000000000_0000000000000000_0000110000011100_0011000111011000"; -- 0.0473052169971772
	pesos_i(10882) := b"1111111111111111_1111111111111111_1111100111000001_0101111000110010"; -- -0.02439318931915455
	pesos_i(10883) := b"0000000000000000_0000000000000000_0010001010000001_1111110111011100"; -- 0.13479601496765267
	pesos_i(10884) := b"0000000000000000_0000000000000000_0000111101111111_0111011010101111"; -- 0.06053869023725002
	pesos_i(10885) := b"0000000000000000_0000000000000000_0000011001110101_0100100110111101"; -- 0.02522717354408463
	pesos_i(10886) := b"0000000000000000_0000000000000000_0000001111100111_1100100011010110"; -- 0.015255501013388935
	pesos_i(10887) := b"1111111111111111_1111111111111111_1110000011001001_0100100101001001"; -- -0.12192861532602935
	pesos_i(10888) := b"0000000000000000_0000000000000000_0000000000101011_1001011011000001"; -- 0.0006651135381996635
	pesos_i(10889) := b"0000000000000000_0000000000000000_0001011011011111_1100001011001111"; -- 0.08935182136655373
	pesos_i(10890) := b"1111111111111111_1111111111111111_1111111110100110_1011111101000001"; -- -0.0013618914381480442
	pesos_i(10891) := b"0000000000000000_0000000000000000_0000010111110100_0011100111110000"; -- 0.023257847786187412
	pesos_i(10892) := b"0000000000000000_0000000000000000_0010000100100111_0111000000111111"; -- 0.12950803306611172
	pesos_i(10893) := b"0000000000000000_0000000000000000_0001100110100011_1000001000011011"; -- 0.10015118753938917
	pesos_i(10894) := b"0000000000000000_0000000000000000_0001111100110101_1100101001101110"; -- 0.1219145316027123
	pesos_i(10895) := b"0000000000000000_0000000000000000_0000110111011111_1000111111011111"; -- 0.05419253525563764
	pesos_i(10896) := b"1111111111111111_1111111111111111_1110110101011000_1011110000110011"; -- -0.07286475900518596
	pesos_i(10897) := b"0000000000000000_0000000000000000_0000100000011101_1100011000101111"; -- 0.031704317658353735
	pesos_i(10898) := b"0000000000000000_0000000000000000_0001110101011111_0101110011111010"; -- 0.11473637685351962
	pesos_i(10899) := b"0000000000000000_0000000000000000_0000111101110001_1110000100011001"; -- 0.06033140996151119
	pesos_i(10900) := b"0000000000000000_0000000000000000_0010001001100001_1100011011000101"; -- 0.13430445018471224
	pesos_i(10901) := b"1111111111111111_1111111111111111_1111110001100110_0101100100100101"; -- -0.01406329010857199
	pesos_i(10902) := b"1111111111111111_1111111111111111_1111111101010111_0001010100001101"; -- -0.0025774805827307487
	pesos_i(10903) := b"0000000000000000_0000000000000000_0000000101111100_0111011111010011"; -- 0.005805481876439094
	pesos_i(10904) := b"1111111111111111_1111111111111111_1111001110000011_0101101111000110"; -- -0.048776878580489944
	pesos_i(10905) := b"0000000000000000_0000000000000000_0001101100101110_0110010001010001"; -- 0.1061766336681077
	pesos_i(10906) := b"1111111111111111_1111111111111111_1111100011010101_0111001011110010"; -- -0.027993026748042237
	pesos_i(10907) := b"0000000000000000_0000000000000000_0001100100001000_1011100110101001"; -- 0.09778938659197418
	pesos_i(10908) := b"1111111111111111_1111111111111111_1101100101101000_1011000011001111"; -- -0.15074629727286942
	pesos_i(10909) := b"0000000000000000_0000000000000000_0000101010001100_1010001101100111"; -- 0.04120847008308157
	pesos_i(10910) := b"1111111111111111_1111111111111111_1110001000010111_1001000010111000"; -- -0.11682792196204125
	pesos_i(10911) := b"1111111111111111_1111111111111111_1110010000011010_1001010001010000"; -- -0.10896943137798033
	pesos_i(10912) := b"0000000000000000_0000000000000000_0000100111110010_0001100010101001"; -- 0.038850346842230994
	pesos_i(10913) := b"0000000000000000_0000000000000000_0000111011001011_0001111010111101"; -- 0.057786866433719136
	pesos_i(10914) := b"1111111111111111_1111111111111111_1110100011111100_1001011011011011"; -- -0.08989579341982074
	pesos_i(10915) := b"0000000000000000_0000000000000000_0000111011011110_1111100010001111"; -- 0.058089766305241604
	pesos_i(10916) := b"0000000000000000_0000000000000000_0001000010001011_0101011010110100"; -- 0.06462613957122693
	pesos_i(10917) := b"0000000000000000_0000000000000000_0000000111110100_0111010110110001"; -- 0.007636409447988868
	pesos_i(10918) := b"1111111111111111_1111111111111111_1111011110011001_0110101011000101"; -- -0.03281529128910168
	pesos_i(10919) := b"0000000000000000_0000000000000000_0000101111000100_1101111000110101"; -- 0.04597271717407108
	pesos_i(10920) := b"0000000000000000_0000000000000000_0001100110000011_1100000001101010"; -- 0.09966662005835629
	pesos_i(10921) := b"0000000000000000_0000000000000000_0001000001001101_1111110101010010"; -- 0.0636900257940076
	pesos_i(10922) := b"1111111111111111_1111111111111111_1111110010010110_1111001111101011"; -- -0.013321642984782953
	pesos_i(10923) := b"1111111111111111_1111111111111111_1110111010101111_0011001001111101"; -- -0.06763920259710123
	pesos_i(10924) := b"1111111111111111_1111111111111111_1101100011111111_0010100011100001"; -- -0.15235657229228652
	pesos_i(10925) := b"1111111111111111_1111111111111111_1111111101110010_1110000101000010"; -- -0.0021533216150385857
	pesos_i(10926) := b"0000000000000000_0000000000000000_0000001110011010_0110010100101111"; -- 0.014074634544760059
	pesos_i(10927) := b"0000000000000000_0000000000000000_0000101100100101_1100000010000100"; -- 0.043544799929341536
	pesos_i(10928) := b"0000000000000000_0000000000000000_0010011100111001_1100111111111010"; -- 0.1532258973359785
	pesos_i(10929) := b"0000000000000000_0000000000000000_0001100110000011_1011110001100001"; -- 0.09966637968324671
	pesos_i(10930) := b"1111111111111111_1111111111111111_1110111111001011_1010011101111000"; -- -0.06329873384248104
	pesos_i(10931) := b"1111111111111111_1111111111111111_1110001001111111_1011010011000011"; -- -0.11523885963007587
	pesos_i(10932) := b"1111111111111111_1111111111111111_1111000110001111_1110110011101001"; -- -0.05639762216253304
	pesos_i(10933) := b"0000000000000000_0000000000000000_0001101100011101_1101100101010001"; -- 0.10592420789234465
	pesos_i(10934) := b"0000000000000000_0000000000000000_0000011010001010_0100011000000100"; -- 0.025547386118146234
	pesos_i(10935) := b"0000000000000000_0000000000000000_0010001100111101_0111011110010001"; -- 0.1376566627313395
	pesos_i(10936) := b"1111111111111111_1111111111111111_1101101100010110_0111101000110001"; -- -0.1441882734844682
	pesos_i(10937) := b"0000000000000000_0000000000000000_0001001011100000_0010011110000000"; -- 0.07373282315027171
	pesos_i(10938) := b"1111111111111111_1111111111111111_1101111101011010_1001000000000010"; -- -0.12752437553692073
	pesos_i(10939) := b"0000000000000000_0000000000000000_0000001111111011_1110010101100100"; -- 0.015562378818828278
	pesos_i(10940) := b"1111111111111111_1111111111111111_1111110100000011_1110010010101101"; -- -0.01165934346396602
	pesos_i(10941) := b"0000000000000000_0000000000000000_0000011110011111_1011011010100001"; -- 0.029780783066943442
	pesos_i(10942) := b"1111111111111111_1111111111111111_1111111011001010_1111100110101110"; -- -0.004715342454104653
	pesos_i(10943) := b"1111111111111111_1111111111111111_1110001111100111_0111100000001011"; -- -0.10974931465288451
	pesos_i(10944) := b"1111111111111111_1111111111111111_1110011101011111_0010110111110010"; -- -0.09620392638647757
	pesos_i(10945) := b"1111111111111111_1111111111111111_1111011001100100_1100000000100011"; -- -0.0375251689379344
	pesos_i(10946) := b"1111111111111111_1111111111111111_1110111010001100_1100000111110011"; -- -0.06816470918406334
	pesos_i(10947) := b"1111111111111111_1111111111111111_1110011111001111_1110110011111000"; -- -0.09448355625375422
	pesos_i(10948) := b"1111111111111111_1111111111111111_1110011111000100_0111011100101101"; -- -0.09465842392165
	pesos_i(10949) := b"1111111111111111_1111111111111111_1111111010100100_1101001110001010"; -- -0.005297449958320058
	pesos_i(10950) := b"0000000000000000_0000000000000000_0001010011110011_0010100010001100"; -- 0.0818353024547863
	pesos_i(10951) := b"0000000000000000_0000000000000000_0001011111000110_1010001000010010"; -- 0.09287465026918762
	pesos_i(10952) := b"1111111111111111_1111111111111111_1110110101001001_0000111101011101"; -- -0.07310394259726632
	pesos_i(10953) := b"1111111111111111_1111111111111111_1101111101100111_0100100010010000"; -- -0.12733026955805288
	pesos_i(10954) := b"0000000000000000_0000000000000000_0001010110011011_1000011001110111"; -- 0.08440437708907879
	pesos_i(10955) := b"0000000000000000_0000000000000000_0000010011101110_1110011100100111"; -- 0.01927036945402095
	pesos_i(10956) := b"0000000000000000_0000000000000000_0000110000011100_1110000110001000"; -- 0.047315688726105795
	pesos_i(10957) := b"0000000000000000_0000000000000000_0000001010100010_1101001000011001"; -- 0.010296946598727234
	pesos_i(10958) := b"0000000000000000_0000000000000000_0000101001001111_0111110111011010"; -- 0.040275445626025176
	pesos_i(10959) := b"1111111111111111_1111111111111111_1101110111100001_1101011001110000"; -- -0.13327274108597323
	pesos_i(10960) := b"1111111111111111_1111111111111111_1111010111001000_1100001010010001"; -- -0.03990539521963355
	pesos_i(10961) := b"0000000000000000_0000000000000000_0000010111001100_1110010100100110"; -- 0.022657701251065625
	pesos_i(10962) := b"0000000000000000_0000000000000000_0000001111011001_0100011111100101"; -- 0.015034192532186097
	pesos_i(10963) := b"0000000000000000_0000000000000000_0000110110001010_1001100111101100"; -- 0.05289613732509157
	pesos_i(10964) := b"1111111111111111_1111111111111111_1111010111110100_1101011100100001"; -- -0.039232782676032654
	pesos_i(10965) := b"1111111111111111_1111111111111111_1111011101101110_0011001011001110"; -- -0.033474754984998724
	pesos_i(10966) := b"0000000000000000_0000000000000000_0000011101011100_0001100000011111"; -- 0.028748996240839687
	pesos_i(10967) := b"1111111111111111_1111111111111111_1110011001000110_0100100011111101"; -- -0.10049003440245369
	pesos_i(10968) := b"0000000000000000_0000000000000000_0001000010111110_0110010111010110"; -- 0.06540523974432705
	pesos_i(10969) := b"1111111111111111_1111111111111111_1111010000001000_1011110010000111"; -- -0.04674169263850438
	pesos_i(10970) := b"1111111111111111_1111111111111111_1111100100100001_0010101000001110"; -- -0.026837703237402397
	pesos_i(10971) := b"1111111111111111_1111111111111111_1101100111111100_1011100101100001"; -- -0.1484874857308535
	pesos_i(10972) := b"0000000000000000_0000000000000000_0010000111011101_0001001000100111"; -- 0.1322795242852478
	pesos_i(10973) := b"0000000000000000_0000000000000000_0000001010110000_0010011100000010"; -- 0.010500371988874067
	pesos_i(10974) := b"0000000000000000_0000000000000000_0000101011111001_1011000001100101"; -- 0.04287245232294306
	pesos_i(10975) := b"0000000000000000_0000000000000000_0001111110001111_1010000011001001"; -- 0.12328534036852819
	pesos_i(10976) := b"0000000000000000_0000000000000000_0001100011110010_1110011000001011"; -- 0.09745633848385311
	pesos_i(10977) := b"0000000000000000_0000000000000000_0010100101111011_1110101101000010"; -- 0.16204710358397262
	pesos_i(10978) := b"1111111111111111_1111111111111111_1110001011100100_0001110100001011"; -- -0.11370676500071336
	pesos_i(10979) := b"1111111111111111_1111111111111111_1111101110000001_0010000111100000"; -- -0.017560847162175396
	pesos_i(10980) := b"0000000000000000_0000000000000000_0001010101100110_1110001111001010"; -- 0.08360122386264449
	pesos_i(10981) := b"0000000000000000_0000000000000000_0001100111011101_1011110000110011"; -- 0.10103965990130885
	pesos_i(10982) := b"0000000000000000_0000000000000000_0001101011100000_0100110111001001"; -- 0.10498510513601188
	pesos_i(10983) := b"0000000000000000_0000000000000000_0001100010010010_1011011011111101"; -- 0.09598869016412985
	pesos_i(10984) := b"1111111111111111_1111111111111111_1110011011000000_0001011011000000"; -- -0.0986314564519521
	pesos_i(10985) := b"1111111111111111_1111111111111111_1111000001000000_0001010000011011"; -- -0.061522239064806444
	pesos_i(10986) := b"1111111111111111_1111111111111111_1110111111011010_1001110101101000"; -- -0.06307045183865886
	pesos_i(10987) := b"1111111111111111_1111111111111111_1110111011111101_0110111101111100"; -- -0.06644538146098573
	pesos_i(10988) := b"0000000000000000_0000000000000000_0001101011111100_0101111011010101"; -- 0.10541336727725159
	pesos_i(10989) := b"1111111111111111_1111111111111111_1110010110010110_0001011011011101"; -- -0.1031785688189226
	pesos_i(10990) := b"0000000000000000_0000000000000000_0000000000001110_1101110100001100"; -- 0.00022679856249254867
	pesos_i(10991) := b"0000000000000000_0000000000000000_0010000100001001_0100100010000111"; -- 0.12904790200137617
	pesos_i(10992) := b"1111111111111111_1111111111111111_1110010110101111_1111110111111101"; -- -0.1027833230136168
	pesos_i(10993) := b"0000000000000000_0000000000000000_0001110001001111_0111011111111101"; -- 0.1105875962165683
	pesos_i(10994) := b"1111111111111111_1111111111111111_1110010110100101_0110101001110001"; -- -0.10294470534331894
	pesos_i(10995) := b"0000000000000000_0000000000000000_0010011010001011_0111111000000110"; -- 0.150565983362315
	pesos_i(10996) := b"0000000000000000_0000000000000000_0001100110101010_0110110100101010"; -- 0.10025675093660244
	pesos_i(10997) := b"1111111111111111_1111111111111111_1101011101011100_0100101110010101"; -- -0.15874793631599687
	pesos_i(10998) := b"0000000000000000_0000000000000000_0001101001011010_1010000011011101"; -- 0.10294537919125574
	pesos_i(10999) := b"1111111111111111_1111111111111111_1111010011011001_1100010011110001"; -- -0.04355210417721763
	pesos_i(11000) := b"0000000000000000_0000000000000000_0001001001001001_0110101111110100"; -- 0.07143282611361439
	pesos_i(11001) := b"1111111111111111_1111111111111111_1110111000010100_0011000100001000"; -- -0.07000440172885215
	pesos_i(11002) := b"1111111111111111_1111111111111111_1101110011010111_1101010100011010"; -- -0.13733165854943896
	pesos_i(11003) := b"0000000000000000_0000000000000000_0000100111100011_0000100110100010"; -- 0.03862056922279122
	pesos_i(11004) := b"1111111111111111_1111111111111111_1110100000010010_0110011001100001"; -- -0.093469239536214
	pesos_i(11005) := b"1111111111111111_1111111111111111_1111100101001010_0101101111010101"; -- -0.0262091260050166
	pesos_i(11006) := b"0000000000000000_0000000000000000_0000110100011111_1010001000000000"; -- 0.05126392848347696
	pesos_i(11007) := b"0000000000000000_0000000000000000_0001111011101011_0011110110001011"; -- 0.12077698366272262
	pesos_i(11008) := b"0000000000000000_0000000000000000_0000011011010101_0011100010001011"; -- 0.02669099228632705
	pesos_i(11009) := b"0000000000000000_0000000000000000_0000000110000111_0111011001100001"; -- 0.005973242483249506
	pesos_i(11010) := b"1111111111111111_1111111111111111_1110000100111100_0010001100100011"; -- -0.12017612845606555
	pesos_i(11011) := b"0000000000000000_0000000000000000_0001101001000101_1111001001110110"; -- 0.10262980823673759
	pesos_i(11012) := b"1111111111111111_1111111111111111_1110101011010110_0001100101111000"; -- -0.08267060106719804
	pesos_i(11013) := b"1111111111111111_1111111111111111_1111001101001011_0000011010001011"; -- -0.049636450776731664
	pesos_i(11014) := b"1111111111111111_1111111111111111_1101110001001010_0010101010101010"; -- -0.13949330666974416
	pesos_i(11015) := b"1111111111111111_1111111111111111_1110111011110011_1101110010111001"; -- -0.06659145819024803
	pesos_i(11016) := b"1111111111111111_1111111111111111_1111100100001000_0000000110011011"; -- -0.027221583936408986
	pesos_i(11017) := b"0000000000000000_0000000000000000_0001010100100111_1000000000010100"; -- 0.08263397673792013
	pesos_i(11018) := b"0000000000000000_0000000000000000_0000000010110000_1010101011010010"; -- 0.002695728633398245
	pesos_i(11019) := b"0000000000000000_0000000000000000_0001011001111011_0110001100110011"; -- 0.08782024368490958
	pesos_i(11020) := b"0000000000000000_0000000000000000_0000010111011010_0100011001111101"; -- 0.022861867553872428
	pesos_i(11021) := b"1111111111111111_1111111111111111_1110001101000111_0010010011110001"; -- -0.11219567401876455
	pesos_i(11022) := b"1111111111111111_1111111111111111_1110001100011010_1000100101110110"; -- -0.11287632820767271
	pesos_i(11023) := b"1111111111111111_1111111111111111_1101111010101100_0001101011110000"; -- -0.13018638269748337
	pesos_i(11024) := b"1111111111111111_1111111111111111_1110011000000110_0000100010101011"; -- -0.10147043064581203
	pesos_i(11025) := b"1111111111111111_1111111111111111_1111100010101010_1111111111000011"; -- -0.028640761162279392
	pesos_i(11026) := b"0000000000000000_0000000000000000_0010000111011010_0100010111001000"; -- 0.13223682537295234
	pesos_i(11027) := b"0000000000000000_0000000000000000_0000101010100011_0100001110001000"; -- 0.04155370780041357
	pesos_i(11028) := b"1111111111111111_1111111111111111_1110100110001100_1010001011111111"; -- -0.08769780424588952
	pesos_i(11029) := b"1111111111111111_1111111111111111_1110000111000101_0010100001101101"; -- -0.11808535909523268
	pesos_i(11030) := b"0000000000000000_0000000000000000_0000000101011011_0000101011110011"; -- 0.005295452453330768
	pesos_i(11031) := b"1111111111111111_1111111111111111_1111101000101011_0111001011100011"; -- -0.022774524278264544
	pesos_i(11032) := b"1111111111111111_1111111111111111_1110100100100100_1100000011110010"; -- -0.08928293327027646
	pesos_i(11033) := b"0000000000000000_0000000000000000_0001111001000110_0111110110001011"; -- 0.1182630982532132
	pesos_i(11034) := b"1111111111111111_1111111111111111_1110001010010110_0111111111010010"; -- -0.11489106296960586
	pesos_i(11035) := b"0000000000000000_0000000000000000_0001001110011100_1000011010001110"; -- 0.07660714122103453
	pesos_i(11036) := b"1111111111111111_1111111111111111_1101100110111000_0101100111011011"; -- -0.14953077701381537
	pesos_i(11037) := b"0000000000000000_0000000000000000_0001111111010101_1100110000010111"; -- 0.124356036691215
	pesos_i(11038) := b"1111111111111111_1111111111111111_1111000011011011_0110010100110000"; -- -0.0591522939941763
	pesos_i(11039) := b"0000000000000000_0000000000000000_0001110011111101_0010101101111011"; -- 0.113238065227577
	pesos_i(11040) := b"1111111111111111_1111111111111111_1111100001110100_1101101101110110"; -- -0.029466899657963553
	pesos_i(11041) := b"0000000000000000_0000000000000000_0010000111111000_1111101101010110"; -- 0.13270541041762526
	pesos_i(11042) := b"0000000000000000_0000000000000000_0000111011010101_0011100111101010"; -- 0.05794107407967334
	pesos_i(11043) := b"0000000000000000_0000000000000000_0001100010100010_1101010000100111"; -- 0.09623456920772194
	pesos_i(11044) := b"1111111111111111_1111111111111111_1110111010001110_1110000111101001"; -- -0.06813228676366534
	pesos_i(11045) := b"1111111111111111_1111111111111111_1110101010111111_1011001100101100"; -- -0.08301239170613113
	pesos_i(11046) := b"0000000000000000_0000000000000000_0001110101101101_0011111001111011"; -- 0.1149481820800195
	pesos_i(11047) := b"1111111111111111_1111111111111111_1110110100001101_0110110001100011"; -- -0.0740139254979677
	pesos_i(11048) := b"1111111111111111_1111111111111111_1101101001011001_1100010100110111"; -- -0.1470677128590122
	pesos_i(11049) := b"0000000000000000_0000000000000000_0000011011010111_1101100001101111"; -- 0.026731040188300727
	pesos_i(11050) := b"1111111111111111_1111111111111111_1111001101011010_0111001101101111"; -- -0.049401078554801116
	pesos_i(11051) := b"1111111111111111_1111111111111111_1111010111110011_0010111101100011"; -- -0.03925803971215746
	pesos_i(11052) := b"0000000000000000_0000000000000000_0000101010000010_0100100101010100"; -- 0.04105051326016448
	pesos_i(11053) := b"0000000000000000_0000000000000000_0001001110000101_0011111001101000"; -- 0.07625188870195455
	pesos_i(11054) := b"0000000000000000_0000000000000000_0001101000100000_0001000100000010"; -- 0.10205179506495834
	pesos_i(11055) := b"1111111111111111_1111111111111111_1110110101001011_1110100100100000"; -- -0.07306044554175205
	pesos_i(11056) := b"0000000000000000_0000000000000000_0010011110010011_0010000001001110"; -- 0.1545887174505049
	pesos_i(11057) := b"1111111111111111_1111111111111111_1110101100000111_1111010101111101"; -- -0.0819098061821715
	pesos_i(11058) := b"0000000000000000_0000000000000000_0010000100101000_1011101000110101"; -- 0.129527700310245
	pesos_i(11059) := b"1111111111111111_1111111111111111_1101110110100101_0110000111111001"; -- -0.13419521016881017
	pesos_i(11060) := b"0000000000000000_0000000000000000_0000110101111001_1010010010101101"; -- 0.052637378918634216
	pesos_i(11061) := b"1111111111111111_1111111111111111_1101110100010011_1111001111110111"; -- -0.1364142915388535
	pesos_i(11062) := b"1111111111111111_1111111111111111_1110010000001111_1111001010100011"; -- -0.10913165592121556
	pesos_i(11063) := b"0000000000000000_0000000000000000_0001011000100100_0101001101000100"; -- 0.08649177942802652
	pesos_i(11064) := b"1111111111111111_1111111111111111_1111010010110110_0011000011100100"; -- -0.04409498639222297
	pesos_i(11065) := b"1111111111111111_1111111111111111_1110111111010110_0010001110000101"; -- -0.06313875209519752
	pesos_i(11066) := b"1111111111111111_1111111111111111_1101110110001011_1101010001001111"; -- -0.13458512372641102
	pesos_i(11067) := b"1111111111111111_1111111111111111_1110000011011100_1101000100100101"; -- -0.12163060034038903
	pesos_i(11068) := b"0000000000000000_0000000000000000_0001111011110100_0010101110011110"; -- 0.12091324438608375
	pesos_i(11069) := b"0000000000000000_0000000000000000_0000000001101001_1000111000110101"; -- 0.0016106490178728439
	pesos_i(11070) := b"1111111111111111_1111111111111111_1111000100001001_0110010010000110"; -- -0.0584504292273791
	pesos_i(11071) := b"1111111111111111_1111111111111111_1111111110001010_1011001110100011"; -- -0.0017898299813379269
	pesos_i(11072) := b"0000000000000000_0000000000000000_0010001001100000_0010000110011101"; -- 0.13427934727095983
	pesos_i(11073) := b"0000000000000000_0000000000000000_0001111101100000_1100010000101001"; -- 0.12257028587345721
	pesos_i(11074) := b"0000000000000000_0000000000000000_0010011000100100_1010110101111010"; -- 0.14899715642840347
	pesos_i(11075) := b"0000000000000000_0000000000000000_0010011001111011_1100010111110011"; -- 0.1503261296928655
	pesos_i(11076) := b"0000000000000000_0000000000000000_0000100111110001_1100100000000010"; -- 0.03884553951063846
	pesos_i(11077) := b"0000000000000000_0000000000000000_0010000000111111_1110110011111101"; -- 0.12597542932907269
	pesos_i(11078) := b"1111111111111111_1111111111111111_1111011100111101_0101000011010001"; -- -0.034220646781366784
	pesos_i(11079) := b"0000000000000000_0000000000000000_0000010101000110_0101101011010011"; -- 0.020604778794823524
	pesos_i(11080) := b"0000000000000000_0000000000000000_0001110010110001_1011100110010100"; -- 0.11208686704521591
	pesos_i(11081) := b"1111111111111111_1111111111111111_1111010000000011_0110011001000000"; -- -0.04682312912012221
	pesos_i(11082) := b"0000000000000000_0000000000000000_0010010111100000_1010101010111100"; -- 0.14795939529563634
	pesos_i(11083) := b"0000000000000000_0000000000000000_0001000010111011_0001010000101110"; -- 0.06535459640213612
	pesos_i(11084) := b"1111111111111111_1111111111111111_1110100100100100_0101010000000001"; -- -0.08928942663247814
	pesos_i(11085) := b"0000000000000000_0000000000000000_0000110001010111_0010011111100001"; -- 0.048204891532133136
	pesos_i(11086) := b"1111111111111111_1111111111111111_1110010001100010_0101010010010100"; -- -0.10787459744326293
	pesos_i(11087) := b"1111111111111111_1111111111111111_1111010010000011_0101011100101100"; -- -0.04487090274861013
	pesos_i(11088) := b"0000000000000000_0000000000000000_0000101110001010_1011010000101011"; -- 0.04508520176632782
	pesos_i(11089) := b"1111111111111111_1111111111111111_1101110111101001_1111101000101101"; -- -0.1331485405026621
	pesos_i(11090) := b"1111111111111111_1111111111111111_1111010011111001_1111010111010011"; -- -0.04306090933155247
	pesos_i(11091) := b"1111111111111111_1111111111111111_1110100011111000_1001111110011110"; -- -0.08995630642171216
	pesos_i(11092) := b"1111111111111111_1111111111111111_1110111101001010_0101011100111101"; -- -0.06527189968706669
	pesos_i(11093) := b"1111111111111111_1111111111111111_1110011111111101_0010111010101011"; -- -0.09379299468074505
	pesos_i(11094) := b"0000000000000000_0000000000000000_0000011111111010_1101100001101110"; -- 0.031171347589980764
	pesos_i(11095) := b"0000000000000000_0000000000000000_0000010000000110_1101110011001010"; -- 0.015729712736835866
	pesos_i(11096) := b"0000000000000000_0000000000000000_0001000011001011_1100111111011110"; -- 0.06560992413677955
	pesos_i(11097) := b"1111111111111111_1111111111111111_1101110111000111_0011101000010010"; -- -0.13367878971117922
	pesos_i(11098) := b"1111111111111111_1111111111111111_1111010011000011_0010101001011110"; -- -0.04389701093955177
	pesos_i(11099) := b"1111111111111111_1111111111111111_1110100110000111_1001010011011011"; -- -0.08777494101260704
	pesos_i(11100) := b"0000000000000000_0000000000000000_0000010111011110_0101010100010001"; -- 0.022923771471175147
	pesos_i(11101) := b"0000000000000000_0000000000000000_0001110110001100_0100100100100010"; -- 0.11542183953369699
	pesos_i(11102) := b"0000000000000000_0000000000000000_0010011101110101_0110010100100100"; -- 0.15413505682624754
	pesos_i(11103) := b"1111111111111111_1111111111111111_1110100100010001_0000101010001001"; -- -0.08958372274824439
	pesos_i(11104) := b"1111111111111111_1111111111111111_1111100101110100_1011010101101110"; -- -0.025562916389893442
	pesos_i(11105) := b"1111111111111111_1111111111111111_1111101001001110_1000011010010011"; -- -0.022239293172923096
	pesos_i(11106) := b"0000000000000000_0000000000000000_0001010111001010_1111010001011111"; -- 0.08512809103541517
	pesos_i(11107) := b"1111111111111111_1111111111111111_1111000111011110_0111110101010010"; -- -0.055198829217029656
	pesos_i(11108) := b"1111111111111111_1111111111111111_1101111101110000_1111011101110101"; -- -0.12718251599612454
	pesos_i(11109) := b"0000000000000000_0000000000000000_0001111000111011_1111111001011001"; -- 0.11810292893503656
	pesos_i(11110) := b"1111111111111111_1111111111111111_1111100111110101_0001100111010111"; -- -0.02360380640000881
	pesos_i(11111) := b"1111111111111111_1111111111111111_1101100110011001_1010110011100001"; -- -0.14999885091425316
	pesos_i(11112) := b"1111111111111111_1111111111111111_1110011110101110_1111100110100001"; -- -0.09498634157564896
	pesos_i(11113) := b"1111111111111111_1111111111111111_1110001010011100_1110011101011000"; -- -0.1147933398297013
	pesos_i(11114) := b"0000000000000000_0000000000000000_0000100011110000_0011011100101000"; -- 0.034915397052899734
	pesos_i(11115) := b"0000000000000000_0000000000000000_0000001011110111_1011111010111111"; -- 0.011592790226923286
	pesos_i(11116) := b"0000000000000000_0000000000000000_0000000111101111_0100101101101011"; -- 0.007557595737239113
	pesos_i(11117) := b"0000000000000000_0000000000000000_0001101111100101_1111100001101111"; -- 0.10897782046358478
	pesos_i(11118) := b"1111111111111111_1111111111111111_1110100011101100_1011010111011110"; -- -0.09013808561146862
	pesos_i(11119) := b"1111111111111111_1111111111111111_1111011011111000_0111000011010010"; -- -0.03527159562810193
	pesos_i(11120) := b"1111111111111111_1111111111111111_1110111100111010_1011000010001000"; -- -0.06551071806723081
	pesos_i(11121) := b"0000000000000000_0000000000000000_0000000011001110_0110101011011110"; -- 0.003149680278095163
	pesos_i(11122) := b"1111111111111111_1111111111111111_1111010110000101_0111110000100001"; -- -0.04093193230418446
	pesos_i(11123) := b"0000000000000000_0000000000000000_0001110010010111_1101001010001111"; -- 0.11169162749662934
	pesos_i(11124) := b"0000000000000000_0000000000000000_0001101100111011_0001011000100011"; -- 0.10637033805594455
	pesos_i(11125) := b"1111111111111111_1111111111111111_1101011001111011_0101111111101001"; -- -0.1621799522290395
	pesos_i(11126) := b"1111111111111111_1111111111111111_1111011000001111_1001000000010101"; -- -0.0388250303158738
	pesos_i(11127) := b"1111111111111111_1111111111111111_1101110000100001_0101011100111111"; -- -0.1401162596091857
	pesos_i(11128) := b"1111111111111111_1111111111111111_1111110110111110_1110001010011101"; -- -0.008806072821913894
	pesos_i(11129) := b"0000000000000000_0000000000000000_0001001010100001_0111110101110011"; -- 0.07277664229892228
	pesos_i(11130) := b"0000000000000000_0000000000000000_0000001001110010_1101110010111110"; -- 0.009565159128557163
	pesos_i(11131) := b"1111111111111111_1111111111111111_1111010100100001_1000111011000100"; -- -0.0424567003505572
	pesos_i(11132) := b"1111111111111111_1111111111111111_1111100111111000_1110101000100110"; -- -0.023545613970466096
	pesos_i(11133) := b"0000000000000000_0000000000000000_0000100110010010_1110001111010110"; -- 0.037397613398015596
	pesos_i(11134) := b"1111111111111111_1111111111111111_1101110111011110_1111101101110000"; -- -0.13331631197689442
	pesos_i(11135) := b"0000000000000000_0000000000000000_0000010100000010_1010101110010011"; -- 0.019571994148677795
	pesos_i(11136) := b"1111111111111111_1111111111111111_1111011001010010_0100100100111001"; -- -0.03780691495610903
	pesos_i(11137) := b"0000000000000000_0000000000000000_0001110010100011_0101101010011100"; -- 0.11186758343059625
	pesos_i(11138) := b"1111111111111111_1111111111111111_1111100001001000_0000111000010110"; -- -0.03015052752180693
	pesos_i(11139) := b"1111111111111111_1111111111111111_1111110000010000_0000110001101001"; -- -0.015380119721588903
	pesos_i(11140) := b"0000000000000000_0000000000000000_0001001110001010_1100000010101011"; -- 0.07633594681335641
	pesos_i(11141) := b"1111111111111111_1111111111111111_1110110011101010_0000010011100010"; -- -0.0745541522308202
	pesos_i(11142) := b"1111111111111111_1111111111111111_1110110000111100_1010001010001010"; -- -0.07719978446814059
	pesos_i(11143) := b"0000000000000000_0000000000000000_0000000101100010_1110010111011010"; -- 0.005415311543292428
	pesos_i(11144) := b"0000000000000000_0000000000000000_0001011001110110_1011101110101101"; -- 0.08774922338465646
	pesos_i(11145) := b"1111111111111111_1111111111111111_1111011010111010_0110100111000000"; -- -0.036218062088490835
	pesos_i(11146) := b"1111111111111111_1111111111111111_1110101010100010_1001010111101101"; -- -0.08345663985926974
	pesos_i(11147) := b"1111111111111111_1111111111111111_1111100111000000_1100001101011001"; -- -0.024402418862675586
	pesos_i(11148) := b"0000000000000000_0000000000000000_0000110011001111_1010000011000001"; -- 0.05004315113062282
	pesos_i(11149) := b"1111111111111111_1111111111111111_1110010001010111_1101000100110101"; -- -0.10803501564786792
	pesos_i(11150) := b"0000000000000000_0000000000000000_0000011011011101_1001001110111101"; -- 0.02681849828465706
	pesos_i(11151) := b"0000000000000000_0000000000000000_0000111111010011_0000011110001010"; -- 0.061813803875691326
	pesos_i(11152) := b"1111111111111111_1111111111111111_1111100001101111_0001110110000101"; -- -0.029554514826984075
	pesos_i(11153) := b"0000000000000000_0000000000000000_0001010011101101_1001011110101111"; -- 0.0817503740491811
	pesos_i(11154) := b"0000000000000000_0000000000000000_0001011101111101_1011001001001000"; -- 0.09176172509986825
	pesos_i(11155) := b"0000000000000000_0000000000000000_0001100111100110_0001101011001000"; -- 0.10116736779702422
	pesos_i(11156) := b"1111111111111111_1111111111111111_1110010001110001_1100010010010000"; -- -0.10763904072084228
	pesos_i(11157) := b"1111111111111111_1111111111111111_1110000100110100_0100101100101100"; -- -0.12029581228605746
	pesos_i(11158) := b"1111111111111111_1111111111111111_1101011111101000_1110000100001110"; -- -0.1566027965411552
	pesos_i(11159) := b"1111111111111111_1111111111111111_1110000010101111_0001010011011111"; -- -0.12232846790766025
	pesos_i(11160) := b"1111111111111111_1111111111111111_1111011100000111_1011110000010010"; -- -0.03503822861929648
	pesos_i(11161) := b"1111111111111111_1111111111111111_1110100111111101_1100001101110000"; -- -0.08597162734818413
	pesos_i(11162) := b"1111111111111111_1111111111111111_1110000101001101_1101110010101110"; -- -0.11990566966246356
	pesos_i(11163) := b"0000000000000000_0000000000000000_0001100010100100_0000110110010000"; -- 0.09625324979169939
	pesos_i(11164) := b"1111111111111111_1111111111111111_1111001011110100_1110010000101010"; -- -0.050950755929259094
	pesos_i(11165) := b"0000000000000000_0000000000000000_0000101110111001_0101010010110010"; -- 0.045796674214206
	pesos_i(11166) := b"1111111111111111_1111111111111111_1101101101000001_1111101010010010"; -- -0.14352449357346478
	pesos_i(11167) := b"1111111111111111_1111111111111111_1110001000011011_1111001100101010"; -- -0.11676101889663416
	pesos_i(11168) := b"1111111111111111_1111111111111111_1111111110001111_0001001010100001"; -- -0.0017231328932685974
	pesos_i(11169) := b"1111111111111111_1111111111111111_1111101101111100_0011101010011110"; -- -0.017635666349989594
	pesos_i(11170) := b"0000000000000000_0000000000000000_0010010110001101_1100010010111100"; -- 0.14669446554347088
	pesos_i(11171) := b"1111111111111111_1111111111111111_1110110111110010_0000100100000010"; -- -0.07052558623061417
	pesos_i(11172) := b"0000000000000000_0000000000000000_0001011001100101_0000110111100001"; -- 0.08747946485536746
	pesos_i(11173) := b"1111111111111111_1111111111111111_1111111100101111_0010110111010000"; -- -0.0031863563001595665
	pesos_i(11174) := b"1111111111111111_1111111111111111_1101100000111100_1111100100010111"; -- -0.15531962584116263
	pesos_i(11175) := b"1111111111111111_1111111111111111_1110111111101011_1110101101001010"; -- -0.06280641028751091
	pesos_i(11176) := b"1111111111111111_1111111111111111_1101110100010001_1111010100001100"; -- -0.13644474454601277
	pesos_i(11177) := b"1111111111111111_1111111111111111_1111111110111101_1001110111011001"; -- -0.0010129304488874391
	pesos_i(11178) := b"0000000000000000_0000000000000000_0010001000111100_0000100100001001"; -- 0.13372856592620613
	pesos_i(11179) := b"0000000000000000_0000000000000000_0001100110100100_0110001111101110"; -- 0.10016464763861148
	pesos_i(11180) := b"0000000000000000_0000000000000000_0010001111110000_0001011111101011"; -- 0.14038228495615443
	pesos_i(11181) := b"0000000000000000_0000000000000000_0010001011011111_1110111000110111"; -- 0.13622940857976645
	pesos_i(11182) := b"0000000000000000_0000000000000000_0010001010010001_1100001101011110"; -- 0.13503666912808326
	pesos_i(11183) := b"0000000000000000_0000000000000000_0000100111011101_1101011100101000"; -- 0.038541266686032895
	pesos_i(11184) := b"1111111111111111_1111111111111111_1111111001010000_1010001100100010"; -- -0.006582073372582996
	pesos_i(11185) := b"1111111111111111_1111111111111111_1110001001001001_1010011010101111"; -- -0.11606367336326102
	pesos_i(11186) := b"1111111111111111_1111111111111111_1101111100001010_0000010011110101"; -- -0.12875336668815304
	pesos_i(11187) := b"0000000000000000_0000000000000000_0001100100100101_0100100100100010"; -- 0.09822518421590666
	pesos_i(11188) := b"0000000000000000_0000000000000000_0001101000010101_1000100111000000"; -- 0.10189114500945472
	pesos_i(11189) := b"0000000000000000_0000000000000000_0001100001110000_0110100001100011"; -- 0.09546520628994516
	pesos_i(11190) := b"1111111111111111_1111111111111111_1110010010010100_1111000110101011"; -- -0.10710229479468199
	pesos_i(11191) := b"1111111111111111_1111111111111111_1110100100111101_1111001110000011"; -- -0.08889844948350763
	pesos_i(11192) := b"0000000000000000_0000000000000000_0001111100000010_1011100001001001"; -- 0.12113525175761349
	pesos_i(11193) := b"0000000000000000_0000000000000000_0000010111111010_0111100111000110"; -- 0.023353205625387008
	pesos_i(11194) := b"1111111111111111_1111111111111111_1111011011000110_0000011001000001"; -- -0.03604088704939094
	pesos_i(11195) := b"0000000000000000_0000000000000000_0001100110010110_0011100101011110"; -- 0.09994848768669777
	pesos_i(11196) := b"0000000000000000_0000000000000000_0010011001101111_1100101111000101"; -- 0.15014337116830134
	pesos_i(11197) := b"1111111111111111_1111111111111111_1111010101110001_1110111100111000"; -- -0.04123024828917828
	pesos_i(11198) := b"1111111111111111_1111111111111111_1111100110001100_0101000111011000"; -- -0.02520264129504782
	pesos_i(11199) := b"0000000000000000_0000000000000000_0001011000100010_1111101110111100"; -- 0.08647130328579647
	pesos_i(11200) := b"0000000000000000_0000000000000000_0001000100001001_1011101000010110"; -- 0.06655467073903051
	pesos_i(11201) := b"0000000000000000_0000000000000000_0001100101011010_0111110110001011"; -- 0.09903702400456092
	pesos_i(11202) := b"1111111111111111_1111111111111111_1101111110001011_1010000100111001"; -- -0.1267756687237188
	pesos_i(11203) := b"0000000000000000_0000000000000000_0001001101010110_0100100100011011"; -- 0.0755353633743606
	pesos_i(11204) := b"0000000000000000_0000000000000000_0010001010101011_1011101000101010"; -- 0.13543284906419523
	pesos_i(11205) := b"0000000000000000_0000000000000000_0000010011001110_1011010110111000"; -- 0.018779141723140803
	pesos_i(11206) := b"0000000000000000_0000000000000000_0001110011101110_1010111010011100"; -- 0.11301699923993828
	pesos_i(11207) := b"1111111111111111_1111111111111111_1101101111010001_1110011101111010"; -- -0.14132836608861124
	pesos_i(11208) := b"1111111111111111_1111111111111111_1111010100010111_1100101101001010"; -- -0.042605680948367704
	pesos_i(11209) := b"1111111111111111_1111111111111111_1111110011011101_0110000111001101"; -- -0.012246978160418536
	pesos_i(11210) := b"0000000000000000_0000000000000000_0000011000001011_0100010001111011"; -- 0.023609428336527332
	pesos_i(11211) := b"1111111111111111_1111111111111111_1111000011001011_1010010110100001"; -- -0.05939259359359699
	pesos_i(11212) := b"0000000000000000_0000000000000000_0001101111111001_1111110001000101"; -- 0.10928322494284146
	pesos_i(11213) := b"0000000000000000_0000000000000000_0000000001110110_1001111111011011"; -- 0.001810065198757129
	pesos_i(11214) := b"1111111111111111_1111111111111111_1111101110010100_0001001001101101"; -- -0.017271851028219168
	pesos_i(11215) := b"1111111111111111_1111111111111111_1111110011111011_0101111100111001"; -- -0.011789368309847755
	pesos_i(11216) := b"0000000000000000_0000000000000000_0001010001111100_1010000010101001"; -- 0.08002666602079311
	pesos_i(11217) := b"0000000000000000_0000000000000000_0010000101100001_1100110110100001"; -- 0.13039860897918434
	pesos_i(11218) := b"1111111111111111_1111111111111111_1110011100101111_1001110011100001"; -- -0.09692973625070786
	pesos_i(11219) := b"1111111111111111_1111111111111111_1110000111101000_0010010100111011"; -- -0.11755149181065214
	pesos_i(11220) := b"0000000000000000_0000000000000000_0001010001000011_1001101010001101"; -- 0.07915655079433603
	pesos_i(11221) := b"0000000000000000_0000000000000000_0001011100111110_0110010110101011"; -- 0.0907958546932274
	pesos_i(11222) := b"1111111111111111_1111111111111111_1111001101000101_0111001110100101"; -- -0.049721500578405214
	pesos_i(11223) := b"1111111111111111_1111111111111111_1101101100000110_0100001011111011"; -- -0.14443570484867807
	pesos_i(11224) := b"0000000000000000_0000000000000000_0001011010010101_0100110100010111"; -- 0.08821565442705662
	pesos_i(11225) := b"1111111111111111_1111111111111111_1101110101100011_0111010111001111"; -- -0.1352011078992043
	pesos_i(11226) := b"1111111111111111_1111111111111111_1110101100010100_0111111101111111"; -- -0.08171847480104363
	pesos_i(11227) := b"0000000000000000_0000000000000000_0001100001110010_0100110111101100"; -- 0.09549414649211099
	pesos_i(11228) := b"1111111111111111_1111111111111111_1111001100111100_1010010110100101"; -- -0.04985584948776029
	pesos_i(11229) := b"0000000000000000_0000000000000000_0010010000011111_1100111110111010"; -- 0.14111040403312045
	pesos_i(11230) := b"0000000000000000_0000000000000000_0001100111011110_0110011111101010"; -- 0.1010498948943745
	pesos_i(11231) := b"1111111111111111_1111111111111111_1110010010001111_1011000000001000"; -- -0.10718250098040816
	pesos_i(11232) := b"1111111111111111_1111111111111111_1111111100010111_0010011101001010"; -- -0.0035529560790707048
	pesos_i(11233) := b"1111111111111111_1111111111111111_1110101001011000_0111001111001001"; -- -0.0845878252863863
	pesos_i(11234) := b"1111111111111111_1111111111111111_1101111110100111_1000000001011000"; -- -0.12635038241425836
	pesos_i(11235) := b"1111111111111111_1111111111111111_1111101100100010_1010111000000110"; -- -0.01900207856031929
	pesos_i(11236) := b"1111111111111111_1111111111111111_1110011010011010_1110010101110001"; -- -0.09919897078675675
	pesos_i(11237) := b"1111111111111111_1111111111111111_1101110101101011_1000000000101100"; -- -0.13507842002497006
	pesos_i(11238) := b"1111111111111111_1111111111111111_1111110111101010_1001010010110101"; -- -0.008139329815978858
	pesos_i(11239) := b"1111111111111111_1111111111111111_1111100101010011_1100001000100111"; -- -0.02606569822567523
	pesos_i(11240) := b"1111111111111111_1111111111111111_1111101010101100_1001010010101100"; -- -0.02080412663462683
	pesos_i(11241) := b"0000000000000000_0000000000000000_0001100010111001_0010011101001110"; -- 0.09657521878615748
	pesos_i(11242) := b"0000000000000000_0000000000000000_0010000001011101_0000100101100101"; -- 0.12641962745291718
	pesos_i(11243) := b"0000000000000000_0000000000000000_0000101001111001_0001101101110010"; -- 0.04091044943193033
	pesos_i(11244) := b"0000000000000000_0000000000000000_0010001001011011_1100011011011011"; -- 0.13421290248085174
	pesos_i(11245) := b"1111111111111111_1111111111111111_1101101101000101_0101001111001100"; -- -0.14347339895327202
	pesos_i(11246) := b"1111111111111111_1111111111111111_1111000111101110_0111100100110010"; -- -0.05495493445894333
	pesos_i(11247) := b"0000000000000000_0000000000000000_0000100110000111_1100111010110010"; -- 0.03722850654890168
	pesos_i(11248) := b"0000000000000000_0000000000000000_0010010111010001_0100010010111101"; -- 0.14772443393428927
	pesos_i(11249) := b"1111111111111111_1111111111111111_1110101000000111_1101011110111001"; -- -0.0858178305104676
	pesos_i(11250) := b"0000000000000000_0000000000000000_0000011010111001_0001011100101111"; -- 0.026261757825724423
	pesos_i(11251) := b"0000000000000000_0000000000000000_0001001000001011_1100001110011110"; -- 0.07049200633751175
	pesos_i(11252) := b"0000000000000000_0000000000000000_0010011010100000_0101000110110010"; -- 0.15088377556519567
	pesos_i(11253) := b"1111111111111111_1111111111111111_1110111000111000_1111011011101000"; -- -0.06944329097437955
	pesos_i(11254) := b"1111111111111111_1111111111111111_1111010000101001_1101100010000011"; -- -0.046236484657212695
	pesos_i(11255) := b"1111111111111111_1111111111111111_1111100001011001_0000110000100011"; -- -0.029891244292697478
	pesos_i(11256) := b"0000000000000000_0000000000000000_0000101010000000_1001000010010110"; -- 0.04102424297107534
	pesos_i(11257) := b"1111111111111111_1111111111111111_1110000111101000_1100001101010000"; -- -0.11754206935240816
	pesos_i(11258) := b"1111111111111111_1111111111111111_1111001111011101_0111100010111101"; -- -0.04740186107573618
	pesos_i(11259) := b"0000000000000000_0000000000000000_0000111001100101_1111001110000011"; -- 0.056243152103027175
	pesos_i(11260) := b"0000000000000000_0000000000000000_0001110101010101_1001101110011011"; -- 0.11458752185886466
	pesos_i(11261) := b"0000000000000000_0000000000000000_0000100110111000_0001010100111110"; -- 0.037965133230009177
	pesos_i(11262) := b"0000000000000000_0000000000000000_0000011110000101_1000010111100111"; -- 0.029381150083738566
	pesos_i(11263) := b"0000000000000000_0000000000000000_0010000100011011_0100111101011001"; -- 0.12932296670202634
	pesos_i(11264) := b"1111111111111111_1111111111111111_1111001111010010_1011001101111100"; -- -0.04756620624174536
	pesos_i(11265) := b"1111111111111111_1111111111111111_1110101100111001_0101110001100000"; -- -0.081155993122813
	pesos_i(11266) := b"0000000000000000_0000000000000000_0010100001000001_1001100000111101"; -- 0.15725089531752534
	pesos_i(11267) := b"1111111111111111_1111111111111111_1110100101010110_0101000001101010"; -- -0.08852670098025761
	pesos_i(11268) := b"1111111111111111_1111111111111111_1110110010001010_0010011111011001"; -- -0.07601691198840199
	pesos_i(11269) := b"1111111111111111_1111111111111111_1110100110100010_1111010100101000"; -- -0.087357213733007
	pesos_i(11270) := b"1111111111111111_1111111111111111_1111100100111101_0101011110100001"; -- -0.026407740700128725
	pesos_i(11271) := b"1111111111111111_1111111111111111_1111101111111111_0101001110111101"; -- -0.015635267701238922
	pesos_i(11272) := b"1111111111111111_1111111111111111_1110111100011110_0001000111010010"; -- -0.06594742421987965
	pesos_i(11273) := b"0000000000000000_0000000000000000_0001000011101100_1111010011001110"; -- 0.0661156656445138
	pesos_i(11274) := b"0000000000000000_0000000000000000_0010010101101000_1101001010001010"; -- 0.14613071316107046
	pesos_i(11275) := b"1111111111111111_1111111111111111_1110000110111101_0000110110101010"; -- -0.1182090244672103
	pesos_i(11276) := b"0000000000000000_0000000000000000_0000101011001010_1111011000101111"; -- 0.042159449178989866
	pesos_i(11277) := b"0000000000000000_0000000000000000_0001110111111000_1100111101011000"; -- 0.11707778827858555
	pesos_i(11278) := b"1111111111111111_1111111111111111_1111000111101001_0111001001100001"; -- -0.05503163465390027
	pesos_i(11279) := b"0000000000000000_0000000000000000_0000111100001111_0101010100010110"; -- 0.058827703432956825
	pesos_i(11280) := b"1111111111111111_1111111111111111_1110100110000010_1011010001010011"; -- -0.08784935936548781
	pesos_i(11281) := b"1111111111111111_1111111111111111_1110100100000111_0111000001100111"; -- -0.08973023875362564
	pesos_i(11282) := b"0000000000000000_0000000000000000_0000011010000001_0111000101000100"; -- 0.025412634843703572
	pesos_i(11283) := b"0000000000000000_0000000000000000_0001101000001110_0000100100000011"; -- 0.10177666028476194
	pesos_i(11284) := b"1111111111111111_1111111111111111_1111100111011101_0011100000110000"; -- -0.023968208503195514
	pesos_i(11285) := b"1111111111111111_1111111111111111_1111011000000001_0111110101101111"; -- -0.0390397648572539
	pesos_i(11286) := b"1111111111111111_1111111111111111_1110101100100010_0111100101101000"; -- -0.0815052147531937
	pesos_i(11287) := b"1111111111111111_1111111111111111_1111001000000100_1101001000001110"; -- -0.05461394458449526
	pesos_i(11288) := b"1111111111111111_1111111111111111_1111010101010110_0110100101110011"; -- -0.04165020881543062
	pesos_i(11289) := b"0000000000000000_0000000000000000_0001001010110000_0111101000101111"; -- 0.07300532956933117
	pesos_i(11290) := b"1111111111111111_1111111111111111_1110000111011100_0010011110101101"; -- -0.1177344515494689
	pesos_i(11291) := b"0000000000000000_0000000000000000_0001100111101111_1111000011000110"; -- 0.10131745169526213
	pesos_i(11292) := b"1111111111111111_1111111111111111_1111100000010010_1111101110101111"; -- -0.03096034030528741
	pesos_i(11293) := b"1111111111111111_1111111111111111_1110111101100011_0111100010000111"; -- -0.06488844595673776
	pesos_i(11294) := b"0000000000000000_0000000000000000_0010001111110100_0010111110000100"; -- 0.14044472667048347
	pesos_i(11295) := b"0000000000000000_0000000000000000_0001101110101111_1010101000110010"; -- 0.1081491824010594
	pesos_i(11296) := b"0000000000000000_0000000000000000_0000111000110111_1110111011010000"; -- 0.05554096780440017
	pesos_i(11297) := b"0000000000000000_0000000000000000_0010000110111011_0101001010111100"; -- 0.13176457497111654
	pesos_i(11298) := b"0000000000000000_0000000000000000_0000010101110101_0010000011110011"; -- 0.021318492289043083
	pesos_i(11299) := b"1111111111111111_1111111111111111_1111101011011001_0101011010101111"; -- -0.020121176025655278
	pesos_i(11300) := b"0000000000000000_0000000000000000_0001010100010011_0011110001111000"; -- 0.08232477132124351
	pesos_i(11301) := b"1111111111111111_1111111111111111_1111111000111110_1100100110011111"; -- -0.006854437620895178
	pesos_i(11302) := b"0000000000000000_0000000000000000_0010010001101110_1000010000011001"; -- 0.14231134032084802
	pesos_i(11303) := b"0000000000000000_0000000000000000_0010001100110100_1111100001001011"; -- 0.13752700645845134
	pesos_i(11304) := b"1111111111111111_1111111111111111_1110111101100101_1101111000010011"; -- -0.06485187560488716
	pesos_i(11305) := b"1111111111111111_1111111111111111_1111111010111011_0110110000011000"; -- -0.004952663513784551
	pesos_i(11306) := b"1111111111111111_1111111111111111_1101101000100010_1010000111010001"; -- -0.1479090562581368
	pesos_i(11307) := b"1111111111111111_1111111111111111_1110010010101001_0100100001010100"; -- -0.10679195366649828
	pesos_i(11308) := b"0000000000000000_0000000000000000_0010001001011000_0110010100101011"; -- 0.1341613036016565
	pesos_i(11309) := b"0000000000000000_0000000000000000_0000001000001111_1011011100100011"; -- 0.0080522977380175
	pesos_i(11310) := b"1111111111111111_1111111111111111_1111010111001011_1010100110101000"; -- -0.03986110341874427
	pesos_i(11311) := b"0000000000000000_0000000000000000_0001101011101000_1111001010010001"; -- 0.10511699712965071
	pesos_i(11312) := b"0000000000000000_0000000000000000_0000110101001010_1101001110111111"; -- 0.05192302143239162
	pesos_i(11313) := b"1111111111111111_1111111111111111_1101100101000100_0000111000100111"; -- -0.15130530874141707
	pesos_i(11314) := b"0000000000000000_0000000000000000_0000101000100011_1000101111101011"; -- 0.03960489731818187
	pesos_i(11315) := b"1111111111111111_1111111111111111_1110110101011000_0011000111001110"; -- -0.07287300799727076
	pesos_i(11316) := b"1111111111111111_1111111111111111_1111101010000000_1101010011011010"; -- -0.0214716880538944
	pesos_i(11317) := b"0000000000000000_0000000000000000_0010011010010001_0010010100111001"; -- 0.15065224305226035
	pesos_i(11318) := b"0000000000000000_0000000000000000_0001011111110111_1101001010111100"; -- 0.09362523153799372
	pesos_i(11319) := b"0000000000000000_0000000000000000_0001000010011001_1101101111100011"; -- 0.06484770106433481
	pesos_i(11320) := b"0000000000000000_0000000000000000_0010001100001001_0010110111010010"; -- 0.13685881027485852
	pesos_i(11321) := b"0000000000000000_0000000000000000_0001011001101111_1010001110100000"; -- 0.08764097849532801
	pesos_i(11322) := b"1111111111111111_1111111111111111_1110110110010011_1000111001011000"; -- -0.07196722376679009
	pesos_i(11323) := b"1111111111111111_1111111111111111_1111111101110000_1110110101100000"; -- -0.0021831170024678524
	pesos_i(11324) := b"1111111111111111_1111111111111111_1101100010110110_0001111000101010"; -- -0.15347110258717897
	pesos_i(11325) := b"0000000000000000_0000000000000000_0000010111110100_0011011101100000"; -- 0.023257695050441063
	pesos_i(11326) := b"1111111111111111_1111111111111111_1110001000010011_0011010000010000"; -- -0.11689447991776358
	pesos_i(11327) := b"0000000000000000_0000000000000000_0000011001001110_0110101001100110"; -- 0.024634027488612355
	pesos_i(11328) := b"0000000000000000_0000000000000000_0001000011101110_1001000110111010"; -- 0.06614027767244905
	pesos_i(11329) := b"1111111111111111_1111111111111111_1111001101101100_1110000110110010"; -- -0.04911984840684735
	pesos_i(11330) := b"1111111111111111_1111111111111111_1110001111100000_1110010111111010"; -- -0.10984957356011615
	pesos_i(11331) := b"0000000000000000_0000000000000000_0000111011100010_1011011010110001"; -- 0.058146875688045316
	pesos_i(11332) := b"0000000000000000_0000000000000000_0000110100111110_1010000010110110"; -- 0.051736874055909314
	pesos_i(11333) := b"1111111111111111_1111111111111111_1110101010011110_0000110100011110"; -- -0.08352582944781968
	pesos_i(11334) := b"1111111111111111_1111111111111111_1110100001101101_1110111010100101"; -- -0.09207256773455225
	pesos_i(11335) := b"1111111111111111_1111111111111111_1111001110110010_0010000110000001"; -- -0.04806318850666139
	pesos_i(11336) := b"1111111111111111_1111111111111111_1111111000010001_0101010010000011"; -- -0.007548063261565219
	pesos_i(11337) := b"1111111111111111_1111111111111111_1111001110000001_0100100101001011"; -- -0.04880849758244988
	pesos_i(11338) := b"1111111111111111_1111111111111111_1111010011111111_0111100011101000"; -- -0.04297680211275975
	pesos_i(11339) := b"0000000000000000_0000000000000000_0001111010011010_0011011110010000"; -- 0.11954066528630708
	pesos_i(11340) := b"1111111111111111_1111111111111111_1111000110010000_0111111110000011"; -- -0.056388884126069766
	pesos_i(11341) := b"1111111111111111_1111111111111111_1111000001111000_1010111100111110"; -- -0.06065849998423273
	pesos_i(11342) := b"1111111111111111_1111111111111111_1110101001100011_0000111011110110"; -- -0.08442598819270562
	pesos_i(11343) := b"1111111111111111_1111111111111111_1101110111000001_0010111011001010"; -- -0.13377101494499147
	pesos_i(11344) := b"1111111111111111_1111111111111111_1101100101101100_0010101101110110"; -- -0.15069321019956625
	pesos_i(11345) := b"0000000000000000_0000000000000000_0001110010011101_1111001010011111"; -- 0.11178509131379662
	pesos_i(11346) := b"1111111111111111_1111111111111111_1111111010111100_0010100001111100"; -- -0.004941434699935817
	pesos_i(11347) := b"0000000000000000_0000000000000000_0000010101111010_0100000001101100"; -- 0.02139666200239558
	pesos_i(11348) := b"1111111111111111_1111111111111111_1111000000101111_1101100100000010"; -- -0.06176990230960993
	pesos_i(11349) := b"0000000000000000_0000000000000000_0001011110110010_1011100111110000"; -- 0.09257089729251039
	pesos_i(11350) := b"0000000000000000_0000000000000000_0001011101001101_0101110101011101"; -- 0.09102424163890874
	pesos_i(11351) := b"0000000000000000_0000000000000000_0001011111110100_1111011000100010"; -- 0.09358156515031428
	pesos_i(11352) := b"1111111111111111_1111111111111111_1111100110101011_0001110101101110"; -- -0.02473274291875584
	pesos_i(11353) := b"0000000000000000_0000000000000000_0001010100011000_0111011001011101"; -- 0.08240451584046371
	pesos_i(11354) := b"1111111111111111_1111111111111111_1111010100001000_0101100101110011"; -- -0.04284134801293299
	pesos_i(11355) := b"0000000000000000_0000000000000000_0010001100100001_1000111110101000"; -- 0.137230852657546
	pesos_i(11356) := b"0000000000000000_0000000000000000_0010001000101011_1111110100111101"; -- 0.13348372200440184
	pesos_i(11357) := b"0000000000000000_0000000000000000_0001111110111101_0101010010000101"; -- 0.12398269887627972
	pesos_i(11358) := b"0000000000000000_0000000000000000_0010010110111000_0010100111111111"; -- 0.14734137030270342
	pesos_i(11359) := b"1111111111111111_1111111111111111_1110110011111010_0001110011000110"; -- -0.07430858776884809
	pesos_i(11360) := b"1111111111111111_1111111111111111_1111101100100000_0000101100000110"; -- -0.019042311787969488
	pesos_i(11361) := b"1111111111111111_1111111111111111_1110000100011011_0111001010010000"; -- -0.12067493425692166
	pesos_i(11362) := b"1111111111111111_1111111111111111_1111010111010101_0010100111101101"; -- -0.03971612886263404
	pesos_i(11363) := b"1111111111111111_1111111111111111_1110111001111110_1010100011100000"; -- -0.06837982693204217
	pesos_i(11364) := b"0000000000000000_0000000000000000_0000111110011110_0001100100100111"; -- 0.06100613789072385
	pesos_i(11365) := b"0000000000000000_0000000000000000_0001000000001100_0110011011101010"; -- 0.06268923960768943
	pesos_i(11366) := b"1111111111111111_1111111111111111_1110001011000001_0000011100111001"; -- -0.11424212318362234
	pesos_i(11367) := b"1111111111111111_1111111111111111_1110110101011010_0011011110000001"; -- -0.07284215067199842
	pesos_i(11368) := b"1111111111111111_1111111111111111_1111011001001110_0100111010010100"; -- -0.03786763078051212
	pesos_i(11369) := b"1111111111111111_1111111111111111_1101110100000011_0111001011001010"; -- -0.1366661317797146
	pesos_i(11370) := b"1111111111111111_1111111111111111_1110110011100101_0100110101011000"; -- -0.07462612729449376
	pesos_i(11371) := b"0000000000000000_0000000000000000_0001111101110001_0011011000100011"; -- 0.12282121993092195
	pesos_i(11372) := b"0000000000000000_0000000000000000_0001111100001000_0101011011111110"; -- 0.12122100536990602
	pesos_i(11373) := b"0000000000000000_0000000000000000_0000101010101000_0100010100101100"; -- 0.04163009963823397
	pesos_i(11374) := b"1111111111111111_1111111111111111_1101100100010010_0000111001001001"; -- -0.15206824037052577
	pesos_i(11375) := b"1111111111111111_1111111111111111_1111110001010100_0010001011000000"; -- -0.014341190436206559
	pesos_i(11376) := b"1111111111111111_1111111111111111_1110000111110011_0111011011101110"; -- -0.11737877541671309
	pesos_i(11377) := b"0000000000000000_0000000000000000_0010000100011111_1011110110011011"; -- 0.12939057389004127
	pesos_i(11378) := b"1111111111111111_1111111111111111_1111110110101110_1111011010100001"; -- -0.009049020460490206
	pesos_i(11379) := b"1111111111111111_1111111111111111_1111111110100101_1000011010001101"; -- -0.0013805298760992048
	pesos_i(11380) := b"0000000000000000_0000000000000000_0000110000101111_0001101000010011"; -- 0.047593717274278614
	pesos_i(11381) := b"0000000000000000_0000000000000000_0001110001010111_0101101001001000"; -- 0.11070789590821267
	pesos_i(11382) := b"1111111111111111_1111111111111111_1110000010101101_0000111010111001"; -- -0.12235935201853228
	pesos_i(11383) := b"0000000000000000_0000000000000000_0000000111100101_1111100110111100"; -- 0.00741539805191141
	pesos_i(11384) := b"0000000000000000_0000000000000000_0000010011010100_1110011010110101"; -- 0.018873614496398187
	pesos_i(11385) := b"1111111111111111_1111111111111111_1101110011101010_0100000101111110"; -- -0.13705053975726386
	pesos_i(11386) := b"0000000000000000_0000000000000000_0010011100111001_1011111000011000"; -- 0.15322483141216123
	pesos_i(11387) := b"1111111111111111_1111111111111111_1110010001001100_0111101011001000"; -- -0.10820801364325083
	pesos_i(11388) := b"1111111111111111_1111111111111111_1110100101101001_0110011100000010"; -- -0.0882354375027896
	pesos_i(11389) := b"0000000000000000_0000000000000000_0010010111110111_1001101111011101"; -- 0.14830946102950765
	pesos_i(11390) := b"0000000000000000_0000000000000000_0000110110001100_0000100100001000"; -- 0.05291801887113542
	pesos_i(11391) := b"0000000000000000_0000000000000000_0001111110010000_0101000010100110"; -- 0.12329582266713536
	pesos_i(11392) := b"1111111111111111_1111111111111111_1101001001110000_1111110011101001"; -- -0.17796344095745142
	pesos_i(11393) := b"1111111111111111_1111111111111111_1110111100001011_0111101001100100"; -- -0.06623110834099963
	pesos_i(11394) := b"0000000000000000_0000000000000000_0000111101010010_0110010111100111"; -- 0.05985104451740266
	pesos_i(11395) := b"1111111111111111_1111111111111111_1111110100110001_0010000110001010"; -- -0.010969070149872742
	pesos_i(11396) := b"0000000000000000_0000000000000000_0010001000001000_1010101100100010"; -- 0.13294477065122992
	pesos_i(11397) := b"1111111111111111_1111111111111111_1110100101100001_0110000001010100"; -- -0.08835790585612563
	pesos_i(11398) := b"0000000000000000_0000000000000000_0001101101011011_1110001111000111"; -- 0.10687087642804487
	pesos_i(11399) := b"0000000000000000_0000000000000000_0001111010111111_1100100001000010"; -- 0.12011386489356216
	pesos_i(11400) := b"1111111111111111_1111111111111111_1111111010100010_0011101011010101"; -- -0.005337069457603108
	pesos_i(11401) := b"0000000000000000_0000000000000000_0001011001101010_0101000111001001"; -- 0.08755980642861465
	pesos_i(11402) := b"0000000000000000_0000000000000000_0010100010110011_1011101100010101"; -- 0.1589924742534382
	pesos_i(11403) := b"0000000000000000_0000000000000000_0000100011111100_0101101001001000"; -- 0.03510059600238609
	pesos_i(11404) := b"0000000000000000_0000000000000000_0001001010011000_0100100010100110"; -- 0.07263616602636523
	pesos_i(11405) := b"1111111111111111_1111111111111111_1110011111010000_0110110101001101"; -- -0.09447590702505544
	pesos_i(11406) := b"0000000000000000_0000000000000000_0000000001010101_1110100111001011"; -- 0.001310932245961803
	pesos_i(11407) := b"0000000000000000_0000000000000000_0001101011111001_1100000111010110"; -- 0.10537349197325828
	pesos_i(11408) := b"1111111111111111_1111111111111111_1111010010101011_0011110111110100"; -- -0.044262054334169826
	pesos_i(11409) := b"1111111111111111_1111111111111111_1101101011100001_0111101000111011"; -- -0.14499698695791488
	pesos_i(11410) := b"0000000000000000_0000000000000000_0000111110011000_0000100111101000"; -- 0.06091367642344859
	pesos_i(11411) := b"0000000000000000_0000000000000000_0001111101111110_0101101101101010"; -- 0.12302180600999917
	pesos_i(11412) := b"0000000000000000_0000000000000000_0001010110101010_0010111100000011"; -- 0.08462804614669851
	pesos_i(11413) := b"0000000000000000_0000000000000000_0010010010100100_0110011000100111"; -- 0.14313353011733654
	pesos_i(11414) := b"0000000000000000_0000000000000000_0000101011110100_0010111000011100"; -- 0.04278839280128982
	pesos_i(11415) := b"0000000000000000_0000000000000000_0000001111111001_0110101011111000"; -- 0.015524564259283946
	pesos_i(11416) := b"0000000000000000_0000000000000000_0001000011001010_1101110010001110"; -- 0.06559542137868946
	pesos_i(11417) := b"1111111111111111_1111111111111111_1110010100111001_0011101010111110"; -- -0.10459549764737718
	pesos_i(11418) := b"0000000000000000_0000000000000000_0000101111101111_1101011001011111"; -- 0.04662837820641831
	pesos_i(11419) := b"0000000000000000_0000000000000000_0000100010110000_0111000111111001"; -- 0.033942340138206246
	pesos_i(11420) := b"1111111111111111_1111111111111111_1110110100110011_1100001101100001"; -- -0.07342890625044672
	pesos_i(11421) := b"0000000000000000_0000000000000000_0001110010011111_1100101001000001"; -- 0.1118132026949599
	pesos_i(11422) := b"0000000000000000_0000000000000000_0001110000010101_1110001101010001"; -- 0.10970898357728863
	pesos_i(11423) := b"0000000000000000_0000000000000000_0010010101011011_0101101011101111"; -- 0.14592521996901092
	pesos_i(11424) := b"1111111111111111_1111111111111111_1110111101100100_0001010110111000"; -- -0.06487907648485906
	pesos_i(11425) := b"0000000000000000_0000000000000000_0001001101101010_1101001000010100"; -- 0.07584870318730554
	pesos_i(11426) := b"1111111111111111_1111111111111111_1110111011101000_1110011010101101"; -- -0.06675871156437087
	pesos_i(11427) := b"0000000000000000_0000000000000000_0001000010101010_1000101101111000"; -- 0.06510230707449823
	pesos_i(11428) := b"0000000000000000_0000000000000000_0000011110100010_0010101100101001"; -- 0.02981824626465508
	pesos_i(11429) := b"0000000000000000_0000000000000000_0001011100101010_1011011001001010"; -- 0.0904954843188839
	pesos_i(11430) := b"1111111111111111_1111111111111111_1111001100111010_0011101110000101"; -- -0.04989269265567713
	pesos_i(11431) := b"1111111111111111_1111111111111111_1111100111011011_1101010110110111"; -- -0.023989336695740972
	pesos_i(11432) := b"0000000000000000_0000000000000000_0001100011000000_1110111101111001"; -- 0.09669396129302626
	pesos_i(11433) := b"1111111111111111_1111111111111111_1110001011110010_0000111110010111"; -- -0.11349394383240964
	pesos_i(11434) := b"0000000000000000_0000000000000000_0001100101011010_1011010111010010"; -- 0.0990403782474627
	pesos_i(11435) := b"0000000000000000_0000000000000000_0001101011001110_0110110101100100"; -- 0.10471233084325847
	pesos_i(11436) := b"1111111111111111_1111111111111111_1110100101111000_1111001001101011"; -- -0.08799824613303109
	pesos_i(11437) := b"0000000000000000_0000000000000000_0001100001100111_0001111011011101"; -- 0.095323494921783
	pesos_i(11438) := b"1111111111111111_1111111111111111_1110010111100001_0010100011011000"; -- -0.1020330879228893
	pesos_i(11439) := b"1111111111111111_1111111111111111_1111110101011111_1000011110100110"; -- -0.010261079754520553
	pesos_i(11440) := b"0000000000000000_0000000000000000_0001001101010100_1010111101001110"; -- 0.0755109373412471
	pesos_i(11441) := b"1111111111111111_1111111111111111_1110111100110110_1001111101100011"; -- -0.0655727752276549
	pesos_i(11442) := b"0000000000000000_0000000000000000_0001111010010101_1011101101111010"; -- 0.11947223409936465
	pesos_i(11443) := b"1111111111111111_1111111111111111_1111001100100101_1001010110000011"; -- -0.0502077632423724
	pesos_i(11444) := b"0000000000000000_0000000000000000_0010001111100100_0010111110001110"; -- 0.14020058846854497
	pesos_i(11445) := b"1111111111111111_1111111111111111_1101101000111111_0101000110001000"; -- -0.14747133670072113
	pesos_i(11446) := b"0000000000000000_0000000000000000_0001011010110010_1011010101011010"; -- 0.08866437390033759
	pesos_i(11447) := b"0000000000000000_0000000000000000_0001111100111001_0110011000000110"; -- 0.12196958215042794
	pesos_i(11448) := b"0000000000000000_0000000000000000_0000001010010110_0100110001101001"; -- 0.010105872862639297
	pesos_i(11449) := b"1111111111111111_1111111111111111_1111111010000110_0101111010100100"; -- -0.005762181186279142
	pesos_i(11450) := b"0000000000000000_0000000000000000_0001110110100001_0001010010001111"; -- 0.11573914049486202
	pesos_i(11451) := b"1111111111111111_1111111111111111_1101111111011011_0000100010001000"; -- -0.12556406661581648
	pesos_i(11452) := b"0000000000000000_0000000000000000_0010001011111000_0111111010011011"; -- 0.13660422600495228
	pesos_i(11453) := b"0000000000000000_0000000000000000_0000101100101101_1000000010100111"; -- 0.04366306390008404
	pesos_i(11454) := b"0000000000000000_0000000000000000_0000010000010000_0001011011111011"; -- 0.015870510300158288
	pesos_i(11455) := b"1111111111111111_1111111111111111_1111001011111101_1001010101011111"; -- -0.05081812304782561
	pesos_i(11456) := b"0000000000000000_0000000000000000_0000000011101100_1111101010110100"; -- 0.0036160172334809637
	pesos_i(11457) := b"1111111111111111_1111111111111111_1101101111110100_0101011110110110"; -- -0.14080287750932952
	pesos_i(11458) := b"1111111111111111_1111111111111111_1111101111000111_0100100010110101"; -- -0.016490417323550374
	pesos_i(11459) := b"0000000000000000_0000000000000000_0000001111011101_1001011111111011"; -- 0.01510000106371631
	pesos_i(11460) := b"1111111111111111_1111111111111111_1110110010010011_0000100100101111"; -- -0.07588141056934766
	pesos_i(11461) := b"1111111111111111_1111111111111111_1110000011011101_1110001001011111"; -- -0.1216143148277987
	pesos_i(11462) := b"0000000000000000_0000000000000000_0001000011001001_1111101101010010"; -- 0.06558199637421427
	pesos_i(11463) := b"0000000000000000_0000000000000000_0001011011100111_0100001001110111"; -- 0.08946624198805257
	pesos_i(11464) := b"1111111111111111_1111111111111111_1111100110111010_0011000011101010"; -- -0.024502699733499535
	pesos_i(11465) := b"0000000000000000_0000000000000000_0001100010010111_0101110000001100"; -- 0.09605956347462201
	pesos_i(11466) := b"1111111111111111_1111111111111111_1110011001100110_0100111111100010"; -- -0.10000134204988265
	pesos_i(11467) := b"1111111111111111_1111111111111111_1111000001010111_1111111101010010"; -- -0.06115726710198189
	pesos_i(11468) := b"1111111111111111_1111111111111111_1111011000000000_1001011101111101"; -- -0.039053470629110895
	pesos_i(11469) := b"1111111111111111_1111111111111111_1111111010010101_1111000100110000"; -- -0.005524564552888688
	pesos_i(11470) := b"1111111111111111_1111111111111111_1101111111000010_1000101110000011"; -- -0.12593772947058582
	pesos_i(11471) := b"0000000000000000_0000000000000000_0000110100001011_0101000001001010"; -- 0.05095388236304456
	pesos_i(11472) := b"0000000000000000_0000000000000000_0010100101001100_1001001010001100"; -- 0.1613246529195874
	pesos_i(11473) := b"1111111111111111_1111111111111111_1111100000010100_1111111100001000"; -- -0.03092962307042159
	pesos_i(11474) := b"0000000000000000_0000000000000000_0000110100001100_1110100000100110"; -- 0.050978192487689644
	pesos_i(11475) := b"1111111111111111_1111111111111111_1110110010110000_0001010010010101"; -- -0.0754382262822358
	pesos_i(11476) := b"1111111111111111_1111111111111111_1101011111110011_0011100000100011"; -- -0.15644501813444592
	pesos_i(11477) := b"0000000000000000_0000000000000000_0010000001010110_1011101100000000"; -- 0.12632340181805574
	pesos_i(11478) := b"0000000000000000_0000000000000000_0001110001110001_1000010000011100"; -- 0.11110711745307156
	pesos_i(11479) := b"1111111111111111_1111111111111111_1101101001110101_1001011101010111"; -- -0.14664320118349167
	pesos_i(11480) := b"0000000000000000_0000000000000000_0000010011010101_1110001110101001"; -- 0.018888691761555387
	pesos_i(11481) := b"0000000000000000_0000000000000000_0001000110111011_1111010010100110"; -- 0.06927422563261817
	pesos_i(11482) := b"0000000000000000_0000000000000000_0000110101000011_0110000010100010"; -- 0.0518093485515035
	pesos_i(11483) := b"1111111111111111_1111111111111111_1101101100000110_1110010011111001"; -- -0.14442604943697826
	pesos_i(11484) := b"0000000000000000_0000000000000000_0010000011000101_1011010001011100"; -- 0.12801673159972685
	pesos_i(11485) := b"1111111111111111_1111111111111111_1111011101111101_0000110011001010"; -- -0.03324813910025214
	pesos_i(11486) := b"1111111111111111_1111111111111111_1110000000000011_1111100110011100"; -- -0.12493934581947756
	pesos_i(11487) := b"1111111111111111_1111111111111111_1101110010001011_0011101111011110"; -- -0.13850045989619333
	pesos_i(11488) := b"1111111111111111_1111111111111111_1110010101010110_0011101011010101"; -- -0.10415298739599989
	pesos_i(11489) := b"0000000000000000_0000000000000000_0001110110011111_0101111011100101"; -- 0.11571305356739402
	pesos_i(11490) := b"1111111111111111_1111111111111111_1101100111000000_0011000001111000"; -- -0.14941117352101052
	pesos_i(11491) := b"1111111111111111_1111111111111111_1110011001110001_0000100011011000"; -- -0.09983772973807373
	pesos_i(11492) := b"1111111111111111_1111111111111111_1111111110000110_1011110110001101"; -- -0.0018502742371878068
	pesos_i(11493) := b"1111111111111111_1111111111111111_1110101100110011_1000100001001111"; -- -0.08124492702822846
	pesos_i(11494) := b"0000000000000000_0000000000000000_0000111000101111_1100100100011000"; -- 0.05541664922827133
	pesos_i(11495) := b"0000000000000000_0000000000000000_0000001100110101_0011101101010010"; -- 0.0125310014883208
	pesos_i(11496) := b"0000000000000000_0000000000000000_0000000110111011_0110000011110001"; -- 0.006765421630126379
	pesos_i(11497) := b"0000000000000000_0000000000000000_0000111010101111_1011001000111111"; -- 0.057368412362171814
	pesos_i(11498) := b"0000000000000000_0000000000000000_0001001111011101_1010110110010000"; -- 0.07760128743491787
	pesos_i(11499) := b"1111111111111111_1111111111111111_1101101111101011_0101011001010100"; -- -0.14094028905206507
	pesos_i(11500) := b"1111111111111111_1111111111111111_1111011000100110_0110001001001010"; -- -0.03847680749525893
	pesos_i(11501) := b"0000000000000000_0000000000000000_0001100010110001_0101001001000001"; -- 0.09645570846416919
	pesos_i(11502) := b"0000000000000000_0000000000000000_0001001111011001_1011111011101000"; -- 0.07754128616143204
	pesos_i(11503) := b"0000000000000000_0000000000000000_0001010100001001_0000000010111010"; -- 0.08216862234557663
	pesos_i(11504) := b"1111111111111111_1111111111111111_1111111010010111_1111101000010011"; -- -0.005493517258766958
	pesos_i(11505) := b"1111111111111111_1111111111111111_1111010001010100_1001100110111101"; -- -0.0455840982184593
	pesos_i(11506) := b"0000000000000000_0000000000000000_0001111100010001_1101100100110011"; -- 0.12136609558730137
	pesos_i(11507) := b"0000000000000000_0000000000000000_0001010000100011_1001011100100001"; -- 0.07866806554895889
	pesos_i(11508) := b"0000000000000000_0000000000000000_0001010000101100_1001111110110110"; -- 0.07880590625469612
	pesos_i(11509) := b"1111111111111111_1111111111111111_1110101000100111_1101101000100000"; -- -0.08532940585568465
	pesos_i(11510) := b"1111111111111111_1111111111111111_1110000110000000_1111110000101010"; -- -0.11912559474593824
	pesos_i(11511) := b"1111111111111111_1111111111111111_1111110000101011_1100110011001000"; -- -0.014956666142846343
	pesos_i(11512) := b"1111111111111111_1111111111111111_1110110110010010_0010001001101101"; -- -0.07198891485650043
	pesos_i(11513) := b"0000000000000000_0000000000000000_0000101000001100_1110110101011101"; -- 0.03925975342502816
	pesos_i(11514) := b"1111111111111111_1111111111111111_1101110000011111_1110111111010010"; -- -0.14013768303730575
	pesos_i(11515) := b"0000000000000000_0000000000000000_0000110001000111_1111010000010010"; -- 0.04797292174321041
	pesos_i(11516) := b"0000000000000000_0000000000000000_0001000101000100_1010110110101101"; -- 0.06745419954041973
	pesos_i(11517) := b"1111111111111111_1111111111111111_1110011001101001_1111010011010100"; -- -0.09994573420695278
	pesos_i(11518) := b"1111111111111111_1111111111111111_1111111001110000_1001110110000110"; -- -0.006094126451803963
	pesos_i(11519) := b"0000000000000000_0000000000000000_0000100100001001_0001101110111111"; -- 0.035295232935774204
	pesos_i(11520) := b"0000000000000000_0000000000000000_0001011011100110_0110011010001010"; -- 0.08945313326553073
	pesos_i(11521) := b"0000000000000000_0000000000000000_0001011101010001_1010010001011011"; -- 0.09108950834673082
	pesos_i(11522) := b"0000000000000000_0000000000000000_0010011001011001_0001110000111011"; -- 0.1497972149285466
	pesos_i(11523) := b"0000000000000000_0000000000000000_0001011101110001_0101001101101011"; -- 0.09157296531293245
	pesos_i(11524) := b"1111111111111111_1111111111111111_1101100000011101_1111110111110011"; -- -0.15579235852440057
	pesos_i(11525) := b"0000000000000000_0000000000000000_0010100001110110_1110101011111001"; -- 0.15806454250892274
	pesos_i(11526) := b"0000000000000000_0000000000000000_0001101010100100_1011101100010100"; -- 0.1040760920532412
	pesos_i(11527) := b"0000000000000000_0000000000000000_0001001110000000_0110000100000111"; -- 0.07617765834882241
	pesos_i(11528) := b"0000000000000000_0000000000000000_0000000001011100_0001110100101001"; -- 0.0014055467866217154
	pesos_i(11529) := b"1111111111111111_1111111111111111_1111110011111010_0111000010100100"; -- -0.011803588946043778
	pesos_i(11530) := b"0000000000000000_0000000000000000_0000101001110111_1101000100110100"; -- 0.040890765277516915
	pesos_i(11531) := b"0000000000000000_0000000000000000_0001101100000011_1101011000011111"; -- 0.10552728906672035
	pesos_i(11532) := b"0000000000000000_0000000000000000_0000101011011011_0000101110001110"; -- 0.042404863538003976
	pesos_i(11533) := b"1111111111111111_1111111111111111_1111010100111000_0011111000010100"; -- -0.04211055762228263
	pesos_i(11534) := b"0000000000000000_0000000000000000_0010010000110010_0001001001100100"; -- 0.14138903561479718
	pesos_i(11535) := b"1111111111111111_1111111111111111_1110001111100100_1010110100111110"; -- -0.10979191994694841
	pesos_i(11536) := b"1111111111111111_1111111111111111_1110011011001000_0001110101010010"; -- -0.09850899445055783
	pesos_i(11537) := b"0000000000000000_0000000000000000_0001110111110100_1100001001111010"; -- 0.11701598628378528
	pesos_i(11538) := b"1111111111111111_1111111111111111_1111110010001100_1101101110100110"; -- -0.013475677379624068
	pesos_i(11539) := b"0000000000000000_0000000000000000_0001101101011001_1110010001010000"; -- 0.10684039074541062
	pesos_i(11540) := b"0000000000000000_0000000000000000_0001000101001100_1001011111000010"; -- 0.06757496337981034
	pesos_i(11541) := b"1111111111111111_1111111111111111_1110100001100001_0010000011101010"; -- -0.09226793565083953
	pesos_i(11542) := b"1111111111111111_1111111111111111_1110000011111001_0110001100010001"; -- -0.12119465670007583
	pesos_i(11543) := b"0000000000000000_0000000000000000_0001010000001101_1110110010101101"; -- 0.0783374712791226
	pesos_i(11544) := b"1111111111111111_1111111111111111_1111000000110000_1010100001010001"; -- -0.06175754570635369
	pesos_i(11545) := b"1111111111111111_1111111111111111_1101001111011001_1011100011101100"; -- -0.17245907059858084
	pesos_i(11546) := b"1111111111111111_1111111111111111_1101101100011000_1010101111110110"; -- -0.1441547893386517
	pesos_i(11547) := b"0000000000000000_0000000000000000_0001101000011111_0010010111000110"; -- 0.10203777397467133
	pesos_i(11548) := b"1111111111111111_1111111111111111_1111011001111100_0101000110111101"; -- -0.03716553818638188
	pesos_i(11549) := b"0000000000000000_0000000000000000_0001011110011000_0010001101101100"; -- 0.09216519735062004
	pesos_i(11550) := b"1111111111111111_1111111111111111_1111101100111101_0100111101100111"; -- -0.018595731229362693
	pesos_i(11551) := b"1111111111111111_1111111111111111_1101100111001010_0000111000000011"; -- -0.14926063947221996
	pesos_i(11552) := b"1111111111111111_1111111111111111_1111000001001100_0010100011011011"; -- -0.061337896796213216
	pesos_i(11553) := b"1111111111111111_1111111111111111_1111110110011001_1011001100101000"; -- -0.009373476841305947
	pesos_i(11554) := b"1111111111111111_1111111111111111_1110110011100110_0011111101000011"; -- -0.07461170783248824
	pesos_i(11555) := b"0000000000000000_0000000000000000_0010001011100100_1000111101110010"; -- 0.13630005392776282
	pesos_i(11556) := b"0000000000000000_0000000000000000_0010011001100100_1011111111111001"; -- 0.14997482147242763
	pesos_i(11557) := b"1111111111111111_1111111111111111_1110101000011101_1101100111100011"; -- -0.08548200809115081
	pesos_i(11558) := b"0000000000000000_0000000000000000_0000111101010110_1011100011111001"; -- 0.059917031042290465
	pesos_i(11559) := b"1111111111111111_1111111111111111_1111100001100000_1000111110100100"; -- -0.029776594712898546
	pesos_i(11560) := b"1111111111111111_1111111111111111_1110100110000000_1100010000111001"; -- -0.08787892926411653
	pesos_i(11561) := b"1111111111111111_1111111111111111_1111010010001011_1010011011110000"; -- -0.044744078147357376
	pesos_i(11562) := b"1111111111111111_1111111111111111_1110101011110011_0100101110110010"; -- -0.0822251023828962
	pesos_i(11563) := b"0000000000000000_0000000000000000_0001100100000111_0101111111011011"; -- 0.09776877497657335
	pesos_i(11564) := b"1111111111111111_1111111111111111_1101100110001110_1011010001000110"; -- -0.15016625671342396
	pesos_i(11565) := b"0000000000000000_0000000000000000_0000011101001010_0000011101111001"; -- 0.028473345857909328
	pesos_i(11566) := b"0000000000000000_0000000000000000_0000100110110001_1101110010101001"; -- 0.037870207963439484
	pesos_i(11567) := b"0000000000000000_0000000000000000_0000110101101010_1110101010110100"; -- 0.05241267094569466
	pesos_i(11568) := b"1111111111111111_1111111111111111_1111110101101010_1111000111010000"; -- -0.010086905261618146
	pesos_i(11569) := b"0000000000000000_0000000000000000_0001111010011011_0000000001000010"; -- 0.11955262766241365
	pesos_i(11570) := b"1111111111111111_1111111111111111_1101110111111110_1000000000111010"; -- -0.13283537456659872
	pesos_i(11571) := b"0000000000000000_0000000000000000_0001000001110111_0000100010101001"; -- 0.06431631217302242
	pesos_i(11572) := b"1111111111111111_1111111111111111_1111101011100101_0101011010111101"; -- -0.019938067284154717
	pesos_i(11573) := b"0000000000000000_0000000000000000_0010001100101011_0101101011101101"; -- 0.13738029741736318
	pesos_i(11574) := b"0000000000000000_0000000000000000_0001100101000011_1100001011101010"; -- 0.09869020660822322
	pesos_i(11575) := b"0000000000000000_0000000000000000_0000100011101110_0100111010111000"; -- 0.03488628371399906
	pesos_i(11576) := b"0000000000000000_0000000000000000_0000100010111101_0010001010101111"; -- 0.03413597850649165
	pesos_i(11577) := b"1111111111111111_1111111111111111_1110101011011010_0110000101111110"; -- -0.08260527308741275
	pesos_i(11578) := b"1111111111111111_1111111111111111_1101100101010100_1100111011010101"; -- -0.1510496834837467
	pesos_i(11579) := b"0000000000000000_0000000000000000_0000001000111011_0111110111111000"; -- 0.008720276874958846
	pesos_i(11580) := b"1111111111111111_1111111111111111_1110111100110010_0110011100011000"; -- -0.06563716569306137
	pesos_i(11581) := b"0000000000000000_0000000000000000_0000111110001100_0110011100001101"; -- 0.0607361228250911
	pesos_i(11582) := b"1111111111111111_1111111111111111_1110100010010000_1011000000011010"; -- -0.091542237864204
	pesos_i(11583) := b"0000000000000000_0000000000000000_0001110111101011_0011011111110111"; -- 0.1168704011056504
	pesos_i(11584) := b"0000000000000000_0000000000000000_0010011001001001_0010101010001111"; -- 0.14955392829010872
	pesos_i(11585) := b"1111111111111111_1111111111111111_1110001100011101_1000000111101011"; -- -0.11283100134230566
	pesos_i(11586) := b"0000000000000000_0000000000000000_0000110011101011_1001011110110111"; -- 0.050469858340345286
	pesos_i(11587) := b"1111111111111111_1111111111111111_1110000011111101_1010010100100100"; -- -0.12112968328414019
	pesos_i(11588) := b"1111111111111111_1111111111111111_1110011110111011_0110101101001001"; -- -0.09479646184551341
	pesos_i(11589) := b"0000000000000000_0000000000000000_0000111110111110_1010100101010010"; -- 0.06150301228097602
	pesos_i(11590) := b"0000000000000000_0000000000000000_0010000001110010_0000010101010111"; -- 0.12673982032860906
	pesos_i(11591) := b"1111111111111111_1111111111111111_1110110011000110_0011001011100101"; -- -0.0751007261077681
	pesos_i(11592) := b"0000000000000000_0000000000000000_0000001001111010_1110111010110110"; -- 0.00968830062690811
	pesos_i(11593) := b"1111111111111111_1111111111111111_1111000001011111_0101001000100101"; -- -0.06104551892003983
	pesos_i(11594) := b"1111111111111111_1111111111111111_1110111000100110_1001001111100101"; -- -0.0697238508613086
	pesos_i(11595) := b"0000000000000000_0000000000000000_0000110010111110_1100110001001001"; -- 0.04978634622162534
	pesos_i(11596) := b"0000000000000000_0000000000000000_0010000100000100_1111000110100111"; -- 0.1289816886793333
	pesos_i(11597) := b"1111111111111111_1111111111111111_1111001111111011_0001011100111001"; -- -0.04694990972676859
	pesos_i(11598) := b"0000000000000000_0000000000000000_0000010000111101_1011010101100111"; -- 0.016566598536635186
	pesos_i(11599) := b"0000000000000000_0000000000000000_0000010110100001_0101001111010101"; -- 0.021992911843995978
	pesos_i(11600) := b"0000000000000000_0000000000000000_0000000101010011_1111110100111111"; -- 0.005187824251534486
	pesos_i(11601) := b"1111111111111111_1111111111111111_1111011001001111_0010101110101111"; -- -0.03785445180514202
	pesos_i(11602) := b"0000000000000000_0000000000000000_0000110100010101_1011111101010110"; -- 0.05111308899703405
	pesos_i(11603) := b"0000000000000000_0000000000000000_0010000100001111_0101001110101110"; -- 0.12914011954754545
	pesos_i(11604) := b"0000000000000000_0000000000000000_0000010100100001_1111100001111000"; -- 0.02004959987183605
	pesos_i(11605) := b"1111111111111111_1111111111111111_1110111010011000_1110000111101100"; -- -0.06797969815453136
	pesos_i(11606) := b"0000000000000000_0000000000000000_0001110110111100_1101101101111110"; -- 0.11616298502258676
	pesos_i(11607) := b"1111111111111111_1111111111111111_1111000110000000_1000101011010011"; -- -0.0566323504951531
	pesos_i(11608) := b"1111111111111111_1111111111111111_1111001110111010_1101110011010101"; -- -0.04792995267930031
	pesos_i(11609) := b"1111111111111111_1111111111111111_1111111100100111_1001000001101101"; -- -0.003302548742876844
	pesos_i(11610) := b"0000000000000000_0000000000000000_0001110101001000_0001001111010100"; -- 0.11438106474141053
	pesos_i(11611) := b"0000000000000000_0000000000000000_0001110011100100_1010001011000111"; -- 0.11286370630213276
	pesos_i(11612) := b"0000000000000000_0000000000000000_0001101100011001_0101111001100011"; -- 0.10585584562684952
	pesos_i(11613) := b"1111111111111111_1111111111111111_1101110010010100_0001000111100010"; -- -0.13836563336841534
	pesos_i(11614) := b"0000000000000000_0000000000000000_0010001010100111_0111011101001010"; -- 0.13536782794441507
	pesos_i(11615) := b"0000000000000000_0000000000000000_0000100110111101_0110001011000110"; -- 0.03804604847923616
	pesos_i(11616) := b"0000000000000000_0000000000000000_0000101110111010_0100001101100100"; -- 0.04581090145644387
	pesos_i(11617) := b"1111111111111111_1111111111111111_1110101001010111_1011100010110010"; -- -0.0845989766143949
	pesos_i(11618) := b"0000000000000000_0000000000000000_0001110100100101_1001111100100101"; -- 0.11385531103676387
	pesos_i(11619) := b"0000000000000000_0000000000000000_0000100010001001_0111010110001110"; -- 0.03334746096839456
	pesos_i(11620) := b"0000000000000000_0000000000000000_0001011101100001_1011111111000011"; -- 0.09133528245947053
	pesos_i(11621) := b"1111111111111111_1111111111111111_1111111001111111_0100010011000001"; -- -0.005870535719013465
	pesos_i(11622) := b"1111111111111111_1111111111111111_1110111010111110_1111100001011111"; -- -0.06739852593481432
	pesos_i(11623) := b"1111111111111111_1111111111111111_1110000001011000_0011101111010100"; -- -0.12365366051030406
	pesos_i(11624) := b"1111111111111111_1111111111111111_1110001100011000_1100110011011011"; -- -0.11290282878193005
	pesos_i(11625) := b"0000000000000000_0000000000000000_0000111010101100_1100100001010101"; -- 0.05732395250675504
	pesos_i(11626) := b"0000000000000000_0000000000000000_0001010100010111_1001110011011101"; -- 0.08239155186490983
	pesos_i(11627) := b"1111111111111111_1111111111111111_1111100100111000_1110100100111001"; -- -0.026475356606751876
	pesos_i(11628) := b"1111111111111111_1111111111111111_1101111100111010_0100101101010001"; -- -0.12801675113369845
	pesos_i(11629) := b"0000000000000000_0000000000000000_0000011111000010_0110111010111010"; -- 0.030310554941124092
	pesos_i(11630) := b"0000000000000000_0000000000000000_0001010110110010_0001111101001010"; -- 0.08474917934428401
	pesos_i(11631) := b"0000000000000000_0000000000000000_0000100110101011_1100000101011010"; -- 0.03777702747527681
	pesos_i(11632) := b"0000000000000000_0000000000000000_0000101101010111_0111100010001111"; -- 0.04430345054607673
	pesos_i(11633) := b"1111111111111111_1111111111111111_1111000101001111_0111100100100000"; -- -0.057381086152717795
	pesos_i(11634) := b"0000000000000000_0000000000000000_0001110100001000_0011010010010000"; -- 0.11340645322329622
	pesos_i(11635) := b"0000000000000000_0000000000000000_0000100100010110_0110010111100000"; -- 0.035498015622616994
	pesos_i(11636) := b"0000000000000000_0000000000000000_0001010001001110_1011001111100011"; -- 0.07932590757651342
	pesos_i(11637) := b"0000000000000000_0000000000000000_0000011010100011_1000110010011100"; -- 0.02593306354402677
	pesos_i(11638) := b"0000000000000000_0000000000000000_0010100110000111_0111010001111111"; -- 0.16222313018768292
	pesos_i(11639) := b"0000000000000000_0000000000000000_0000100100110110_1101001100100000"; -- 0.03599280864810676
	pesos_i(11640) := b"1111111111111111_1111111111111111_1110000011010001_1000110001111111"; -- -0.12180253880143592
	pesos_i(11641) := b"1111111111111111_1111111111111111_1110111110010110_0100000111100101"; -- -0.06411350400171179
	pesos_i(11642) := b"1111111111111111_1111111111111111_1110011000110011_0100001100000001"; -- -0.10078030803767885
	pesos_i(11643) := b"0000000000000000_0000000000000000_0000001111111110_1010110000101010"; -- 0.015604744313210477
	pesos_i(11644) := b"1111111111111111_1111111111111111_1111101000100010_0010110111001000"; -- -0.022915972373626012
	pesos_i(11645) := b"1111111111111111_1111111111111111_1110010011001100_0001011111010001"; -- -0.10626078738526337
	pesos_i(11646) := b"0000000000000000_0000000000000000_0000010100010110_0111100101011100"; -- 0.019874176960175655
	pesos_i(11647) := b"0000000000000000_0000000000000000_0001110100001011_0111111101110111"; -- 0.1134566942264744
	pesos_i(11648) := b"1111111111111111_1111111111111111_1110011110000110_1000001000000101"; -- -0.09560382252421527
	pesos_i(11649) := b"0000000000000000_0000000000000000_0000100110110000_1111100011101100"; -- 0.03785663384665233
	pesos_i(11650) := b"0000000000000000_0000000000000000_0000010110101000_1110100111110011"; -- 0.022108670909467967
	pesos_i(11651) := b"0000000000000000_0000000000000000_0000111001111011_0101011110010000"; -- 0.05656955012557648
	pesos_i(11652) := b"0000000000000000_0000000000000000_0000001011001101_1010011010110111"; -- 0.010950488668790174
	pesos_i(11653) := b"1111111111111111_1111111111111111_1111100100001010_1101000011011011"; -- -0.027178713383417964
	pesos_i(11654) := b"0000000000000000_0000000000000000_0010000010011000_0111000000100010"; -- 0.12732601966664722
	pesos_i(11655) := b"0000000000000000_0000000000000000_0000001101011111_0010101100011110"; -- 0.013170904838353785
	pesos_i(11656) := b"1111111111111111_1111111111111111_1111011000001110_0000110011111011"; -- -0.038848103216849846
	pesos_i(11657) := b"1111111111111111_1111111111111111_1101111010000001_1111011110011101"; -- -0.13082935729877262
	pesos_i(11658) := b"0000000000000000_0000000000000000_0000001000110001_0101111110100010"; -- 0.008565880834945085
	pesos_i(11659) := b"1111111111111111_1111111111111111_1111010011100101_0101110111010100"; -- -0.04337514473102305
	pesos_i(11660) := b"1111111111111111_1111111111111111_1110010010011110_0010111010100000"; -- -0.10696133233496638
	pesos_i(11661) := b"1111111111111111_1111111111111111_1101100100011110_0000101011010011"; -- -0.1518853411141135
	pesos_i(11662) := b"0000000000000000_0000000000000000_0001110000010110_1010101010110001"; -- 0.10972086727005903
	pesos_i(11663) := b"0000000000000000_0000000000000000_0000111100011001_1001101101101011"; -- 0.058984483373163
	pesos_i(11664) := b"1111111111111111_1111111111111111_1111110111110101_1010101111100001"; -- -0.007970101908171028
	pesos_i(11665) := b"1111111111111111_1111111111111111_1110000000110111_0000001101011111"; -- -0.12416056560685644
	pesos_i(11666) := b"1111111111111111_1111111111111111_1111111000010000_1111011011100111"; -- -0.007553642941349239
	pesos_i(11667) := b"1111111111111111_1111111111111111_1110001001000000_1101001010011111"; -- -0.11619838344457137
	pesos_i(11668) := b"0000000000000000_0000000000000000_0001110100111000_0000001100010010"; -- 0.1141359251793466
	pesos_i(11669) := b"0000000000000000_0000000000000000_0001010100111100_1011001100111110"; -- 0.08295746089544967
	pesos_i(11670) := b"0000000000000000_0000000000000000_0001101011001000_1110101010100111"; -- 0.1046282442897819
	pesos_i(11671) := b"0000000000000000_0000000000000000_0010010101001110_0100011101011100"; -- 0.1457256889932434
	pesos_i(11672) := b"1111111111111111_1111111111111111_1111110100100010_0000000000110000"; -- -0.011199939959341485
	pesos_i(11673) := b"0000000000000000_0000000000000000_0001110001110101_1000010011010101"; -- 0.11116819573141212
	pesos_i(11674) := b"0000000000000000_0000000000000000_0001111100100111_0001111000001000"; -- 0.12169063266926788
	pesos_i(11675) := b"0000000000000000_0000000000000000_0001011011101100_0001011001101111"; -- 0.08953991146953547
	pesos_i(11676) := b"0000000000000000_0000000000000000_0001111101001111_1110001000100110"; -- 0.12231267376126653
	pesos_i(11677) := b"0000000000000000_0000000000000000_0000010100001010_0000100101011001"; -- 0.019684395055161646
	pesos_i(11678) := b"1111111111111111_1111111111111111_1111010101111010_1110100101010010"; -- -0.04109327075367255
	pesos_i(11679) := b"0000000000000000_0000000000000000_0001010101111001_0100011100111000"; -- 0.08388180848899843
	pesos_i(11680) := b"1111111111111111_1111111111111111_1110101110110001_1011000000101001"; -- -0.07931994430114957
	pesos_i(11681) := b"0000000000000000_0000000000000000_0001100000110010_1110111010011001"; -- 0.09452716105015756
	pesos_i(11682) := b"1111111111111111_1111111111111111_1111110111110010_1111111001001111"; -- -0.008010965009115663
	pesos_i(11683) := b"0000000000000000_0000000000000000_0001011110000110_0110111111111100"; -- 0.09189510242205733
	pesos_i(11684) := b"1111111111111111_1111111111111111_1111101110000100_1001100110111001"; -- -0.017507927273160546
	pesos_i(11685) := b"0000000000000000_0000000000000000_0000000000000011_1110000101110000"; -- 5.921345213002915e-05
	pesos_i(11686) := b"1111111111111111_1111111111111111_1110111101111010_1100001011101110"; -- -0.06453305895380787
	pesos_i(11687) := b"0000000000000000_0000000000000000_0000011110010001_1110100101110100"; -- 0.02957018932516779
	pesos_i(11688) := b"0000000000000000_0000000000000000_0000011100000110_1011100000000110"; -- 0.027446271467827566
	pesos_i(11689) := b"0000000000000000_0000000000000000_0010000001111000_0101001010010011"; -- 0.126835976518402
	pesos_i(11690) := b"0000000000000000_0000000000000000_0000011011001111_1101011010111100"; -- 0.026608868461701414
	pesos_i(11691) := b"1111111111111111_1111111111111111_1110100001101011_0011100111011011"; -- -0.09211386106746816
	pesos_i(11692) := b"0000000000000000_0000000000000000_0001101101101001_1100111000001000"; -- 0.1070832033183709
	pesos_i(11693) := b"0000000000000000_0000000000000000_0001111100011001_1011101000010111"; -- 0.121486311582177
	pesos_i(11694) := b"0000000000000000_0000000000000000_0000111110101111_0011101001011110"; -- 0.061267516926832515
	pesos_i(11695) := b"1111111111111111_1111111111111111_1111111000010010_0100100011011111"; -- -0.007533498328702823
	pesos_i(11696) := b"0000000000000000_0000000000000000_0010000011101011_0111010011010010"; -- 0.1285927784795824
	pesos_i(11697) := b"1111111111111111_1111111111111111_1111101000100000_0010001100010010"; -- -0.022947128376396224
	pesos_i(11698) := b"0000000000000000_0000000000000000_0000111010010110_1101110111011001"; -- 0.05698954154530939
	pesos_i(11699) := b"1111111111111111_1111111111111111_1101111001001011_0010101011101111"; -- -0.13166553188013377
	pesos_i(11700) := b"1111111111111111_1111111111111111_1110100000111100_0001010110001111"; -- -0.09283318757564366
	pesos_i(11701) := b"1111111111111111_1111111111111111_1101100011010001_0101100010100101"; -- -0.1530556294135332
	pesos_i(11702) := b"1111111111111111_1111111111111111_1110110000111011_1110101100100000"; -- -0.07721071701369155
	pesos_i(11703) := b"1111111111111111_1111111111111111_1111011110000100_1100101111101000"; -- -0.03312993619828674
	pesos_i(11704) := b"1111111111111111_1111111111111111_1101110011111110_1110010011011100"; -- -0.1367356266011507
	pesos_i(11705) := b"0000000000000000_0000000000000000_0001111001101111_1011101011100110"; -- 0.11889236561904072
	pesos_i(11706) := b"0000000000000000_0000000000000000_0000111101011100_0101011111010000"; -- 0.060002792546381946
	pesos_i(11707) := b"0000000000000000_0000000000000000_0000011010000110_1011001011000010"; -- 0.02549283243968448
	pesos_i(11708) := b"1111111111111111_1111111111111111_1110100101100011_0100000011110000"; -- -0.08832925930125209
	pesos_i(11709) := b"0000000000000000_0000000000000000_0000111000110000_0111000001001000"; -- 0.0554266143982142
	pesos_i(11710) := b"0000000000000000_0000000000000000_0010010101000000_0001011110000001"; -- 0.14550921334720843
	pesos_i(11711) := b"1111111111111111_1111111111111111_1110011110000100_1100101111001100"; -- -0.09562994257721885
	pesos_i(11712) := b"0000000000000000_0000000000000000_0000001000001011_1011000011010111"; -- 0.007990887096794267
	pesos_i(11713) := b"0000000000000000_0000000000000000_0010010111001001_0011000101111011"; -- 0.14760121593972236
	pesos_i(11714) := b"1111111111111111_1111111111111111_1110110011111100_0000000100001010"; -- -0.07427972319259063
	pesos_i(11715) := b"1111111111111111_1111111111111111_1110110111110010_0011100111010100"; -- -0.0705226762672351
	pesos_i(11716) := b"0000000000000000_0000000000000000_0001001011100001_0000000110110001"; -- 0.07374582834433499
	pesos_i(11717) := b"1111111111111111_1111111111111111_1111010011000000_0010100110011011"; -- -0.04394283269197921
	pesos_i(11718) := b"1111111111111111_1111111111111111_1101110111010101_0000100011101000"; -- -0.13346809696354311
	pesos_i(11719) := b"1111111111111111_1111111111111111_1110111110101101_0010011000110110"; -- -0.06376420189243125
	pesos_i(11720) := b"1111111111111111_1111111111111111_1111110111010000_0000100000010100"; -- -0.008544440423096909
	pesos_i(11721) := b"1111111111111111_1111111111111111_1111100110011100_1011111100111001"; -- -0.024951981050236056
	pesos_i(11722) := b"1111111111111111_1111111111111111_1101111000100010_1000001011001001"; -- -0.13228590586820274
	pesos_i(11723) := b"1111111111111111_1111111111111111_1110001011001010_0110001010010010"; -- -0.11409934926919948
	pesos_i(11724) := b"0000000000000000_0000000000000000_0010001101111011_1101111110101101"; -- 0.13860891310313572
	pesos_i(11725) := b"1111111111111111_1111111111111111_1110010110010000_1111110010011000"; -- -0.10325642870319886
	pesos_i(11726) := b"0000000000000000_0000000000000000_0010000110011101_0110000111000000"; -- 0.1313077061750099
	pesos_i(11727) := b"1111111111111111_1111111111111111_1111000000011110_0101110000100101"; -- -0.06203674408988069
	pesos_i(11728) := b"0000000000000000_0000000000000000_0001101110001001_1110100101101011"; -- 0.1075731168550013
	pesos_i(11729) := b"0000000000000000_0000000000000000_0001001110011011_0010110110110001"; -- 0.07658658583421098
	pesos_i(11730) := b"0000000000000000_0000000000000000_0010001001100011_1110010101001001"; -- 0.13433678656255105
	pesos_i(11731) := b"1111111111111111_1111111111111111_1111100111110111_1100101100001001"; -- -0.023562727347983977
	pesos_i(11732) := b"1111111111111111_1111111111111111_1110001101011100_0000111010010011"; -- -0.11187657266165257
	pesos_i(11733) := b"1111111111111111_1111111111111111_1110011100010101_1001100100011001"; -- -0.0973266901521679
	pesos_i(11734) := b"0000000000000000_0000000000000000_0010010100111000_0000100010001000"; -- 0.14538625065706937
	pesos_i(11735) := b"1111111111111111_1111111111111111_1101111011001000_1001111100001010"; -- -0.12975126278857158
	pesos_i(11736) := b"0000000000000000_0000000000000000_0000100011011110_0000011001000010"; -- 0.034637824175274556
	pesos_i(11737) := b"1111111111111111_1111111111111111_1111000001110000_1101100100110001"; -- -0.06077807001580607
	pesos_i(11738) := b"0000000000000000_0000000000000000_0000000101101100_1111111111101100"; -- 0.0055694533908005025
	pesos_i(11739) := b"0000000000000000_0000000000000000_0001111011000100_1111111011110001"; -- 0.12019341840955969
	pesos_i(11740) := b"1111111111111111_1111111111111111_1110100100101101_1100001111111111"; -- -0.08914542232618519
	pesos_i(11741) := b"1111111111111111_1111111111111111_1111100011100110_1110110110110101"; -- -0.02772631016176747
	pesos_i(11742) := b"1111111111111111_1111111111111111_1110011011001111_1010011110100110"; -- -0.09839393799798264
	pesos_i(11743) := b"1111111111111111_1111111111111111_1101110101011101_1000111101011000"; -- -0.13529113855471042
	pesos_i(11744) := b"0000000000000000_0000000000000000_0001000110001010_1010010000000110"; -- 0.06852173948364708
	pesos_i(11745) := b"1111111111111111_1111111111111111_1110100100000001_0001110010011001"; -- -0.08982678659488279
	pesos_i(11746) := b"0000000000000000_0000000000000000_0000011010010011_0101110101000100"; -- 0.02568610106268169
	pesos_i(11747) := b"1111111111111111_1111111111111111_1111101011010111_1001101010100010"; -- -0.02014764346061736
	pesos_i(11748) := b"1111111111111111_1111111111111111_1111111110001110_0111000100000000"; -- -0.0017327666469241557
	pesos_i(11749) := b"0000000000000000_0000000000000000_0000100011010100_0011110001010110"; -- 0.03448845947368277
	pesos_i(11750) := b"0000000000000000_0000000000000000_0001100110000100_1100110110001001"; -- 0.0996826609105239
	pesos_i(11751) := b"0000000000000000_0000000000000000_0000101110100110_0010010011011011"; -- 0.04550390576401469
	pesos_i(11752) := b"1111111111111111_1111111111111111_1111010101011011_1011001101110001"; -- -0.041569504554522234
	pesos_i(11753) := b"0000000000000000_0000000000000000_0010010100001010_1110000001101100"; -- 0.14469721457400242
	pesos_i(11754) := b"0000000000000000_0000000000000000_0001001110011011_0011101001010110"; -- 0.0765873394896764
	pesos_i(11755) := b"1111111111111111_1111111111111111_1110111100011100_1000100110100110"; -- -0.06597079946247704
	pesos_i(11756) := b"0000000000000000_0000000000000000_0000011100011100_0000000110110100"; -- 0.02777109764322281
	pesos_i(11757) := b"0000000000000000_0000000000000000_0001100110100100_0010101110000110"; -- 0.1001612855311135
	pesos_i(11758) := b"1111111111111111_1111111111111111_1110010110110001_1001111111010011"; -- -0.10275841805157702
	pesos_i(11759) := b"1111111111111111_1111111111111111_1110011011110110_0101001111011100"; -- -0.09780383939435737
	pesos_i(11760) := b"0000000000000000_0000000000000000_0010010100011111_0010100011000110"; -- 0.1450067026791301
	pesos_i(11761) := b"0000000000000000_0000000000000000_0001010001010110_1001111101000000"; -- 0.07944674778467438
	pesos_i(11762) := b"0000000000000000_0000000000000000_0001100111110101_0110111011010110"; -- 0.10140125968627449
	pesos_i(11763) := b"0000000000000000_0000000000000000_0010011110000111_0110000001001000"; -- 0.15440942542483266
	pesos_i(11764) := b"0000000000000000_0000000000000000_0001001000110111_1001000110000010"; -- 0.0711604062910898
	pesos_i(11765) := b"1111111111111111_1111111111111111_1110111011011100_0001011101101010"; -- -0.06695417074616855
	pesos_i(11766) := b"1111111111111111_1111111111111111_1111011101000000_1101101110010001"; -- -0.034166600407471236
	pesos_i(11767) := b"0000000000000000_0000000000000000_0010000111101111_1100100111011110"; -- 0.13256513281395507
	pesos_i(11768) := b"1111111111111111_1111111111111111_1110101100011101_0100111101010110"; -- -0.08158401639957143
	pesos_i(11769) := b"0000000000000000_0000000000000000_0000011110100111_1111111101111100"; -- 0.029907195762154015
	pesos_i(11770) := b"0000000000000000_0000000000000000_0000100001001001_0010101001010101"; -- 0.03236641483150139
	pesos_i(11771) := b"0000000000000000_0000000000000000_0001011011000110_0110110001001110"; -- 0.0889651957456747
	pesos_i(11772) := b"1111111111111111_1111111111111111_1110101110011111_1100000000011001"; -- -0.07959365267269637
	pesos_i(11773) := b"0000000000000000_0000000000000000_0010010000011011_1100101000101110"; -- 0.14104903824824416
	pesos_i(11774) := b"1111111111111111_1111111111111111_1110110001100011_0011110110011100"; -- -0.07661070758947236
	pesos_i(11775) := b"1111111111111111_1111111111111111_1111000000110010_1001000000010010"; -- -0.0617284733655389
	pesos_i(11776) := b"1111111111111111_1111111111111111_1111111100000101_1010110001111101"; -- -0.003819674990183015
	pesos_i(11777) := b"1111111111111111_1111111111111111_1111010100001011_0111110100011000"; -- -0.0427934471831212
	pesos_i(11778) := b"1111111111111111_1111111111111111_1111100010010101_0100110010110101"; -- -0.028971868351057056
	pesos_i(11779) := b"1111111111111111_1111111111111111_1111111110001100_1011011011010101"; -- -0.001759121859529665
	pesos_i(11780) := b"1111111111111111_1111111111111111_1110001011000011_0101001010001100"; -- -0.11420711596886172
	pesos_i(11781) := b"0000000000000000_0000000000000000_0000001110110100_0001111110001001"; -- 0.014467211610312407
	pesos_i(11782) := b"0000000000000000_0000000000000000_0010001000110100_0110000011000111"; -- 0.1336117253035036
	pesos_i(11783) := b"1111111111111111_1111111111111111_1111100101010010_1000100001010110"; -- -0.02608440295938095
	pesos_i(11784) := b"1111111111111111_1111111111111111_1110110001111001_0011010110111001"; -- -0.07627548434930721
	pesos_i(11785) := b"0000000000000000_0000000000000000_0001110110010011_0101101101001011"; -- 0.11552973359002004
	pesos_i(11786) := b"1111111111111111_1111111111111111_1111001101111111_0110010110100100"; -- -0.04883732549757585
	pesos_i(11787) := b"1111111111111111_1111111111111111_1110110001111111_1000100001111110"; -- -0.07617899815782658
	pesos_i(11788) := b"1111111111111111_1111111111111111_1101110000010001_1011111000101001"; -- -0.1403542662441046
	pesos_i(11789) := b"1111111111111111_1111111111111111_1111111111001001_1100011010111001"; -- -0.0008273886253494552
	pesos_i(11790) := b"0000000000000000_0000000000000000_0001000110100010_1110100111001110"; -- 0.06889210971129554
	pesos_i(11791) := b"0000000000000000_0000000000000000_0000001110010111_0101101100010000"; -- 0.014028254994019256
	pesos_i(11792) := b"0000000000000000_0000000000000000_0001101010010000_0111110111010001"; -- 0.10376726491766379
	pesos_i(11793) := b"1111111111111111_1111111111111111_1111010011101010_1111011100100000"; -- -0.04328971359524903
	pesos_i(11794) := b"1111111111111111_1111111111111111_1111010001001101_1010100100111011"; -- -0.045689986435954816
	pesos_i(11795) := b"0000000000000000_0000000000000000_0001101001010011_1011010110110010"; -- 0.1028398094157264
	pesos_i(11796) := b"1111111111111111_1111111111111111_1111000100100100_1101010000010010"; -- -0.05803179316079299
	pesos_i(11797) := b"0000000000000000_0000000000000000_0001010001010000_1011001011011101"; -- 0.07935636424538456
	pesos_i(11798) := b"1111111111111111_1111111111111111_1111100101100110_1100111010100101"; -- -0.025775036442365312
	pesos_i(11799) := b"0000000000000000_0000000000000000_0010001011100001_1111001010100110"; -- 0.13626019050982552
	pesos_i(11800) := b"0000000000000000_0000000000000000_0000011000111111_0010100111011010"; -- 0.024401298244387443
	pesos_i(11801) := b"1111111111111111_1111111111111111_1111101101100011_1000100101110111"; -- -0.018012436355026883
	pesos_i(11802) := b"0000000000000000_0000000000000000_0000000100000101_1101010000110100"; -- 0.003995192336261268
	pesos_i(11803) := b"0000000000000000_0000000000000000_0000100110010101_1111011110110110"; -- 0.0374445742780697
	pesos_i(11804) := b"1111111111111111_1111111111111111_1111101110001011_1001001010111000"; -- -0.017401533278292983
	pesos_i(11805) := b"1111111111111111_1111111111111111_1110010011000010_0011000000110110"; -- -0.10641192132594653
	pesos_i(11806) := b"1111111111111111_1111111111111111_1101110010001010_0011000100011011"; -- -0.13851636019420682
	pesos_i(11807) := b"0000000000000000_0000000000000000_0001101000000001_0001111100111101"; -- 0.10157962074584369
	pesos_i(11808) := b"0000000000000000_0000000000000000_0001100001111111_0100010000000111"; -- 0.09569192096932616
	pesos_i(11809) := b"1111111111111111_1111111111111111_1101110111100110_1110111100001001"; -- -0.13319498093470364
	pesos_i(11810) := b"1111111111111111_1111111111111111_1111000010000100_0000111010110110"; -- -0.06048496305299449
	pesos_i(11811) := b"0000000000000000_0000000000000000_0001001011101111_1000000010010110"; -- 0.07396701493020115
	pesos_i(11812) := b"0000000000000000_0000000000000000_0001000000110010_1010101111011010"; -- 0.06327318258989072
	pesos_i(11813) := b"0000000000000000_0000000000000000_0000010101101001_0101000010101010"; -- 0.021138230883435003
	pesos_i(11814) := b"0000000000000000_0000000000000000_0001100011000000_1100011100000001"; -- 0.09669154900853037
	pesos_i(11815) := b"0000000000000000_0000000000000000_0000100111110001_0111010001010010"; -- 0.03884055129991718
	pesos_i(11816) := b"0000000000000000_0000000000000000_0001110000001000_1110000111101001"; -- 0.10951053549846873
	pesos_i(11817) := b"1111111111111111_1111111111111111_1110111011111110_0101101010001010"; -- -0.06643137103245167
	pesos_i(11818) := b"0000000000000000_0000000000000000_0001011101101011_0000011110000000"; -- 0.0914768875234937
	pesos_i(11819) := b"1111111111111111_1111111111111111_1101101001011011_0011101100101001"; -- -0.14704542396695616
	pesos_i(11820) := b"0000000000000000_0000000000000000_0000100111111011_0100101111010100"; -- 0.038990725752145516
	pesos_i(11821) := b"0000000000000000_0000000000000000_0000111111000110_1001001100001001"; -- 0.061623754305467175
	pesos_i(11822) := b"0000000000000000_0000000000000000_0010000111001101_1011011000011011"; -- 0.1320451561179406
	pesos_i(11823) := b"1111111111111111_1111111111111111_1110100000010011_1110011110100100"; -- -0.09344627610192527
	pesos_i(11824) := b"0000000000000000_0000000000000000_0000001110010011_0010100010111110"; -- 0.01396422035980896
	pesos_i(11825) := b"1111111111111111_1111111111111111_1110110101001000_0100000110100011"; -- -0.07311620495252023
	pesos_i(11826) := b"0000000000000000_0000000000000000_0000111011001001_1001000001011001"; -- 0.05776312032722277
	pesos_i(11827) := b"0000000000000000_0000000000000000_0000001010010001_0011010010010000"; -- 0.010028157294488672
	pesos_i(11828) := b"1111111111111111_1111111111111111_1111010010110001_1011000011010111"; -- -0.04416365390010147
	pesos_i(11829) := b"1111111111111111_1111111111111111_1111110111111001_1000101100010110"; -- -0.00791102144164362
	pesos_i(11830) := b"1111111111111111_1111111111111111_1110000101011110_1110110000000110"; -- -0.11964535573773853
	pesos_i(11831) := b"0000000000000000_0000000000000000_0001001101110100_1010000110011001"; -- 0.07599840146490601
	pesos_i(11832) := b"0000000000000000_0000000000000000_0010000100101000_0110000011101101"; -- 0.1295223787418245
	pesos_i(11833) := b"0000000000000000_0000000000000000_0001011111011001_1011011100010110"; -- 0.0931658199580464
	pesos_i(11834) := b"1111111111111111_1111111111111111_1111101010000000_1111001001001000"; -- -0.021469933993068877
	pesos_i(11835) := b"0000000000000000_0000000000000000_0000110100110010_1100001110011101"; -- 0.051555848959287165
	pesos_i(11836) := b"1111111111111111_1111111111111111_1111000100000110_0010101101101011"; -- -0.05849960933963789
	pesos_i(11837) := b"1111111111111111_1111111111111111_1110010010001001_0001110101010100"; -- -0.10728279776315512
	pesos_i(11838) := b"1111111111111111_1111111111111111_1111100110000111_1001110101111101"; -- -0.025274426442902266
	pesos_i(11839) := b"1111111111111111_1111111111111111_1110000111010010_1011100001111111"; -- -0.11787840741870899
	pesos_i(11840) := b"1111111111111111_1111111111111111_1111110001110011_1010000000001010"; -- -0.013860700078109056
	pesos_i(11841) := b"0000000000000000_0000000000000000_0001001110111011_1100010101001100"; -- 0.07708390341468822
	pesos_i(11842) := b"0000000000000000_0000000000000000_0001011100100100_1101111011011011"; -- 0.09040634970732091
	pesos_i(11843) := b"1111111111111111_1111111111111111_1110010011000100_0110000111101000"; -- -0.10637844167067348
	pesos_i(11844) := b"0000000000000000_0000000000000000_0001000001111010_0000000011011010"; -- 0.06436162304912274
	pesos_i(11845) := b"0000000000000000_0000000000000000_0010010011100000_0001011001110010"; -- 0.14404430659949666
	pesos_i(11846) := b"0000000000000000_0000000000000000_0001110101000111_1111001101100011"; -- 0.11437913089575658
	pesos_i(11847) := b"1111111111111111_1111111111111111_1101111000011011_1100011111000101"; -- -0.1323886055476697
	pesos_i(11848) := b"1111111111111111_1111111111111111_1110010111001100_0101101101011101"; -- -0.10235051142305315
	pesos_i(11849) := b"0000000000000000_0000000000000000_0000100111110011_1000001001010110"; -- 0.03887190436352176
	pesos_i(11850) := b"1111111111111111_1111111111111111_1111101110111100_0110011101000000"; -- -0.01665644338166931
	pesos_i(11851) := b"0000000000000000_0000000000000000_0010001110100110_0011010111001001"; -- 0.13925491487056854
	pesos_i(11852) := b"1111111111111111_1111111111111111_1101111010101001_0110000001001100"; -- -0.130228024954932
	pesos_i(11853) := b"0000000000000000_0000000000000000_0001011000011000_1001101110011111"; -- 0.08631298665830832
	pesos_i(11854) := b"0000000000000000_0000000000000000_0000110101110101_1001101010100000"; -- 0.052575744784014306
	pesos_i(11855) := b"0000000000000000_0000000000000000_0001100011000010_1100100110001000"; -- 0.09672221728550752
	pesos_i(11856) := b"0000000000000000_0000000000000000_0010011100001101_1000001101101111"; -- 0.15254994838583127
	pesos_i(11857) := b"0000000000000000_0000000000000000_0001100001111110_1101010101000101"; -- 0.09568531939279044
	pesos_i(11858) := b"0000000000000000_0000000000000000_0000000100010101_0001011100011100"; -- 0.004228061905117985
	pesos_i(11859) := b"1111111111111111_1111111111111111_1101111010001011_0001101110010110"; -- -0.13068988396505674
	pesos_i(11860) := b"0000000000000000_0000000000000000_0001101001011000_0101110001100000"; -- 0.10291077942026888
	pesos_i(11861) := b"1111111111111111_1111111111111111_1110010001101111_1111000001111000"; -- -0.10766694139138464
	pesos_i(11862) := b"1111111111111111_1111111111111111_1110011110111110_1011001001101111"; -- -0.0947464445391849
	pesos_i(11863) := b"0000000000000000_0000000000000000_0010001011010011_0100011001111001"; -- 0.13603630492819815
	pesos_i(11864) := b"0000000000000000_0000000000000000_0001110000101110_0010100000101110"; -- 0.11007929913528784
	pesos_i(11865) := b"1111111111111111_1111111111111111_1111000001000100_0111110011100101"; -- -0.061454958059705314
	pesos_i(11866) := b"0000000000000000_0000000000000000_0010011001000111_0111110100001101"; -- 0.14952832772454971
	pesos_i(11867) := b"1111111111111111_1111111111111111_1111111101011110_0110010010101110"; -- -0.0024659228691422787
	pesos_i(11868) := b"1111111111111111_1111111111111111_1110011011001000_0111100010101111"; -- -0.09850354886725221
	pesos_i(11869) := b"0000000000000000_0000000000000000_0001111010011000_1010000100110100"; -- 0.11951644440505034
	pesos_i(11870) := b"0000000000000000_0000000000000000_0000100000000000_1101000101101101"; -- 0.03126248276410228
	pesos_i(11871) := b"1111111111111111_1111111111111111_1101110001011010_1011011101011100"; -- -0.13924077983683564
	pesos_i(11872) := b"0000000000000000_0000000000000000_0001010010010100_1100010011011011"; -- 0.08039503424909017
	pesos_i(11873) := b"0000000000000000_0000000000000000_0000010010011011_0001100100000101"; -- 0.017991603657133814
	pesos_i(11874) := b"0000000000000000_0000000000000000_0001010001100110_0101101010101110"; -- 0.07968680143888279
	pesos_i(11875) := b"1111111111111111_1111111111111111_1101001111100101_0100101001101111"; -- -0.17228255079344082
	pesos_i(11876) := b"1111111111111111_1111111111111111_1111011010111111_0101110101110011"; -- -0.03614250125028033
	pesos_i(11877) := b"0000000000000000_0000000000000000_0000010110100100_1111100111101100"; -- 0.02204858798962489
	pesos_i(11878) := b"1111111111111111_1111111111111111_1101011011000110_0111011010001000"; -- -0.16103419469218713
	pesos_i(11879) := b"1111111111111111_1111111111111111_1111010100110101_0110110000011100"; -- -0.04215359043997021
	pesos_i(11880) := b"1111111111111111_1111111111111111_1111010000101010_1100110100101001"; -- -0.04622190239013499
	pesos_i(11881) := b"1111111111111111_1111111111111111_1101101110011010_1100000110101101"; -- -0.14216985253658404
	pesos_i(11882) := b"1111111111111111_1111111111111111_1110010110001110_0011011011101111"; -- -0.10329872754521366
	pesos_i(11883) := b"1111111111111111_1111111111111111_1111100001010000_1010001110000101"; -- -0.03001955031204337
	pesos_i(11884) := b"1111111111111111_1111111111111111_1111100001011010_0101010010010100"; -- -0.02987166776290008
	pesos_i(11885) := b"0000000000000000_0000000000000000_0010010101110001_0010011001100001"; -- 0.14625778072151766
	pesos_i(11886) := b"1111111111111111_1111111111111111_1101010110111100_1111010100001100"; -- -0.16508549180064586
	pesos_i(11887) := b"0000000000000000_0000000000000000_0001100100000101_0110000111110011"; -- 0.09773838227469658
	pesos_i(11888) := b"1111111111111111_1111111111111111_1111101100111010_1011111111010100"; -- -0.018634806377726253
	pesos_i(11889) := b"1111111111111111_1111111111111111_1110110111010101_0110010100110011"; -- -0.07096259597260592
	pesos_i(11890) := b"1111111111111111_1111111111111111_1110011110100001_1100111111110111"; -- -0.0951871892831147
	pesos_i(11891) := b"0000000000000000_0000000000000000_0001001011111011_0100000011011000"; -- 0.07414632112278624
	pesos_i(11892) := b"0000000000000000_0000000000000000_0000010111111001_0001111000000101"; -- 0.023332477678407463
	pesos_i(11893) := b"1111111111111111_1111111111111111_1101111001100101_0101110110101011"; -- -0.13126577921555938
	pesos_i(11894) := b"0000000000000000_0000000000000000_0010001010000011_0101000110010000"; -- 0.1348162627829117
	pesos_i(11895) := b"0000000000000000_0000000000000000_0010111001010001_0100000000000101"; -- 0.1809272778819544
	pesos_i(11896) := b"0000000000000000_0000000000000000_0000100100100110_0011100111000111"; -- 0.03573952770406333
	pesos_i(11897) := b"0000000000000000_0000000000000000_0000100011001111_0101011011101011"; -- 0.034413750003489736
	pesos_i(11898) := b"1111111111111111_1111111111111111_1111000010000110_0000011101110011"; -- -0.060454878156587205
	pesos_i(11899) := b"1111111111111111_1111111111111111_1111011110011001_1000100010010111"; -- -0.032813513904072604
	pesos_i(11900) := b"1111111111111111_1111111111111111_1110100001010100_0001001001000101"; -- -0.09246717288145831
	pesos_i(11901) := b"1111111111111111_1111111111111111_1111000001101110_0110001011111010"; -- -0.06081563374623079
	pesos_i(11902) := b"0000000000000000_0000000000000000_0010000111101011_1001001101110101"; -- 0.13250085459316246
	pesos_i(11903) := b"0000000000000000_0000000000000000_0001001011010000_1110001101001010"; -- 0.07349987561983423
	pesos_i(11904) := b"1111111111111111_1111111111111111_1101101111011110_1101111100110110"; -- -0.1411304945033962
	pesos_i(11905) := b"1111111111111111_1111111111111111_1110101001010110_1100010000010010"; -- -0.08461355746646164
	pesos_i(11906) := b"1111111111111111_1111111111111111_1110100100101000_0011100001001001"; -- -0.08923004364231238
	pesos_i(11907) := b"1111111111111111_1111111111111111_1111100011101101_0100001011101100"; -- -0.02762967810253031
	pesos_i(11908) := b"0000000000000000_0000000000000000_0000010100100110_1010001010111010"; -- 0.02012078327343388
	pesos_i(11909) := b"1111111111111111_1111111111111111_1111111001011011_0010101111010001"; -- -0.006421338435348219
	pesos_i(11910) := b"0000000000000000_0000000000000000_0001110100101011_1011100100111011"; -- 0.11394841844942169
	pesos_i(11911) := b"1111111111111111_1111111111111111_1101111011011100_1100101110110010"; -- -0.12944342530072114
	pesos_i(11912) := b"1111111111111111_1111111111111111_1111101001101010_1010101111101000"; -- -0.02180982193211673
	pesos_i(11913) := b"0000000000000000_0000000000000000_0000110010000110_1100000010100100"; -- 0.048931159894639954
	pesos_i(11914) := b"1111111111111111_1111111111111111_1101110111001101_0101101111110011"; -- -0.13358521773499632
	pesos_i(11915) := b"1111111111111111_1111111111111111_1110010011101111_1000011001101111"; -- -0.10572013657840668
	pesos_i(11916) := b"0000000000000000_0000000000000000_0010001101000011_1111000111010000"; -- 0.13775550190043473
	pesos_i(11917) := b"0000000000000000_0000000000000000_0000000000101000_0111000100000010"; -- 0.0006170873948403938
	pesos_i(11918) := b"0000000000000000_0000000000000000_0001101110110101_1011111000011101"; -- 0.10824192247023248
	pesos_i(11919) := b"1111111111111111_1111111111111111_1110100001010000_0001100010110101"; -- -0.092527824196278
	pesos_i(11920) := b"0000000000000000_0000000000000000_0010011111101010_1011000000110000"; -- 0.1559248083349565
	pesos_i(11921) := b"0000000000000000_0000000000000000_0000111101111101_0111101001111000"; -- 0.06050839844797193
	pesos_i(11922) := b"0000000000000000_0000000000000000_0001100101101011_1011010100010101"; -- 0.09929973365369432
	pesos_i(11923) := b"0000000000000000_0000000000000000_0010000111111011_1011111111100010"; -- 0.13274764310383128
	pesos_i(11924) := b"0000000000000000_0000000000000000_0000010111001010_1101101101011111"; -- 0.022626600841316076
	pesos_i(11925) := b"0000000000000000_0000000000000000_0000110111101001_0010001100111111"; -- 0.054338648708728315
	pesos_i(11926) := b"0000000000000000_0000000000000000_0000010101000000_0100001011010100"; -- 0.020511795785685166
	pesos_i(11927) := b"1111111111111111_1111111111111111_1111110000001100_0010010110101101"; -- -0.015439648852324683
	pesos_i(11928) := b"1111111111111111_1111111111111111_1111011100101111_1001110001100010"; -- -0.03442976584235017
	pesos_i(11929) := b"1111111111111111_1111111111111111_1111011001001111_0101100111000101"; -- -0.03785170495252122
	pesos_i(11930) := b"1111111111111111_1111111111111111_1111000000010111_1000000100111001"; -- -0.062141345493894294
	pesos_i(11931) := b"1111111111111111_1111111111111111_1101101001100110_0010010011100111"; -- -0.14687890394652975
	pesos_i(11932) := b"0000000000000000_0000000000000000_0001101110011000_1000010001001011"; -- 0.10779597129316872
	pesos_i(11933) := b"0000000000000000_0000000000000000_0001010111000000_0010111100011100"; -- 0.08496374545936985
	pesos_i(11934) := b"1111111111111111_1111111111111111_1110110000110001_0110010010000110"; -- -0.07737132774591804
	pesos_i(11935) := b"1111111111111111_1111111111111111_1111101110000000_0111001011001010"; -- -0.01757128305025233
	pesos_i(11936) := b"1111111111111111_1111111111111111_1110110010100011_1101010100111001"; -- -0.07562510838716317
	pesos_i(11937) := b"0000000000000000_0000000000000000_0000001101001110_1010111111110101"; -- 0.012919423468530785
	pesos_i(11938) := b"1111111111111111_1111111111111111_1111111110100001_1110101111011100"; -- -0.0014355266109588112
	pesos_i(11939) := b"0000000000000000_0000000000000000_0010011100010010_0011111101011110"; -- 0.15262218527094476
	pesos_i(11940) := b"1111111111111111_1111111111111111_1111011100101111_0100110110100011"; -- -0.03443445944594495
	pesos_i(11941) := b"1111111111111111_1111111111111111_1101100101000100_0000000110110110"; -- -0.15130605038152856
	pesos_i(11942) := b"1111111111111111_1111111111111111_1101110110000011_0101100011011100"; -- -0.1347145521744167
	pesos_i(11943) := b"0000000000000000_0000000000000000_0000010010110100_0101001101111101"; -- 0.018376558432902337
	pesos_i(11944) := b"0000000000000000_0000000000000000_0000100000000111_0001010111010111"; -- 0.03135811329860355
	pesos_i(11945) := b"0000000000000000_0000000000000000_0001110010011111_1011010110101111"; -- 0.11181197658121159
	pesos_i(11946) := b"1111111111111111_1111111111111111_1101101111011111_1010100100110010"; -- -0.1411184551840828
	pesos_i(11947) := b"0000000000000000_0000000000000000_0000000111110101_0011011100000101"; -- 0.007647932759723306
	pesos_i(11948) := b"0000000000000000_0000000000000000_0001101001101110_0110000101100000"; -- 0.10324677077898693
	pesos_i(11949) := b"0000000000000000_0000000000000000_0000110111100011_1110000110001100"; -- 0.05425843869731283
	pesos_i(11950) := b"1111111111111111_1111111111111111_1110100011110010_1000111001101010"; -- -0.0900488846028641
	pesos_i(11951) := b"0000000000000000_0000000000000000_0001100010111111_0111011100010001"; -- 0.09667152567915044
	pesos_i(11952) := b"0000000000000000_0000000000000000_0001111011001010_0100001101001111"; -- 0.1202737874032639
	pesos_i(11953) := b"0000000000000000_0000000000000000_0001010000001001_0010111011000100"; -- 0.0782651164711226
	pesos_i(11954) := b"1111111111111111_1111111111111111_1110000011110101_1011001001110011"; -- -0.12125096021503588
	pesos_i(11955) := b"0000000000000000_0000000000000000_0000111001110000_0111000110111001"; -- 0.056403262736228976
	pesos_i(11956) := b"1111111111111111_1111111111111111_1111111111100100_1110010010100010"; -- -0.0004136186152156999
	pesos_i(11957) := b"1111111111111111_1111111111111111_1111010110001100_0110111110010111"; -- -0.040825868206846104
	pesos_i(11958) := b"0000000000000000_0000000000000000_0000111010110001_0000011000010010"; -- 0.05738866743976928
	pesos_i(11959) := b"0000000000000000_0000000000000000_0001110101010100_0110111110011000"; -- 0.11456963968819231
	pesos_i(11960) := b"1111111111111111_1111111111111111_1110001101001100_0011001001011000"; -- -0.1121185812454701
	pesos_i(11961) := b"0000000000000000_0000000000000000_0001111101110101_1100010100100100"; -- 0.12289077881003521
	pesos_i(11962) := b"1111111111111111_1111111111111111_1110111011110100_0101010000011000"; -- -0.06658434311336378
	pesos_i(11963) := b"0000000000000000_0000000000000000_0001100001001110_1001011111100110"; -- 0.09494923930367204
	pesos_i(11964) := b"0000000000000000_0000000000000000_0010000111010101_1010010001111010"; -- 0.1321661757427848
	pesos_i(11965) := b"1111111111111111_1111111111111111_1110100111100101_1101101100110111"; -- -0.08633642098718004
	pesos_i(11966) := b"1111111111111111_1111111111111111_1101101111101010_1010110111110111"; -- -0.14095032424162585
	pesos_i(11967) := b"0000000000000000_0000000000000000_0000101100001001_1010001000100011"; -- 0.043115743299989254
	pesos_i(11968) := b"0000000000000000_0000000000000000_0000111000110001_1010000110001101"; -- 0.05544480973714384
	pesos_i(11969) := b"1111111111111111_1111111111111111_1101111010001010_1010011000010001"; -- -0.13069688878574348
	pesos_i(11970) := b"0000000000000000_0000000000000000_0000101010000100_1011010101011010"; -- 0.04108746955175348
	pesos_i(11971) := b"0000000000000000_0000000000000000_0000111000100101_0001010101100001"; -- 0.05525334958732623
	pesos_i(11972) := b"0000000000000000_0000000000000000_0010010110010110_1111110101110000"; -- 0.14683517432603582
	pesos_i(11973) := b"0000000000000000_0000000000000000_0001101100100110_0010011101000001"; -- 0.10605092381340525
	pesos_i(11974) := b"1111111111111111_1111111111111111_1111111111000000_0111001000111111"; -- -0.0009697529657116038
	pesos_i(11975) := b"1111111111111111_1111111111111111_1111101111110010_1100011110111010"; -- -0.015826718306573655
	pesos_i(11976) := b"1111111111111111_1111111111111111_1101111101101101_1101011011101110"; -- -0.12723023113889548
	pesos_i(11977) := b"1111111111111111_1111111111111111_1111101100010100_0010011101111011"; -- -0.01922372111043633
	pesos_i(11978) := b"0000000000000000_0000000000000000_0001100000101100_0000011110000010"; -- 0.09442183432857476
	pesos_i(11979) := b"0000000000000000_0000000000000000_0000010111001011_1101011011000000"; -- 0.022641584315404046
	pesos_i(11980) := b"1111111111111111_1111111111111111_1101110000011101_1011101111111111"; -- -0.14017128960342604
	pesos_i(11981) := b"0000000000000000_0000000000000000_0000100011110010_1000101110101011"; -- 0.03495095184193696
	pesos_i(11982) := b"1111111111111111_1111111111111111_1110110100111000_0111111101011100"; -- -0.07335666654248457
	pesos_i(11983) := b"0000000000000000_0000000000000000_0001111101011110_0101011101100110"; -- 0.12253328550333986
	pesos_i(11984) := b"0000000000000000_0000000000000000_0000001000110011_0111101100000100"; -- 0.008598030463727476
	pesos_i(11985) := b"0000000000000000_0000000000000000_0000100111101000_1101101111011110"; -- 0.03870939410845901
	pesos_i(11986) := b"0000000000000000_0000000000000000_0001101100000011_1010011010110011"; -- 0.10552446238672737
	pesos_i(11987) := b"1111111111111111_1111111111111111_1110111110101010_0001111110110000"; -- -0.06381036712691424
	pesos_i(11988) := b"1111111111111111_1111111111111111_1111100001000011_1000111100100011"; -- -0.030219129598242654
	pesos_i(11989) := b"1111111111111111_1111111111111111_1111101000100100_1001101001111101"; -- -0.022878975403596024
	pesos_i(11990) := b"0000000000000000_0000000000000000_0001010110100001_1111101000101010"; -- 0.08450282603808895
	pesos_i(11991) := b"1111111111111111_1111111111111111_1111101111100110_1111100111100011"; -- -0.016006834163949536
	pesos_i(11992) := b"0000000000000000_0000000000000000_0001100110101010_0000111111110100"; -- 0.10025119504850039
	pesos_i(11993) := b"0000000000000000_0000000000000000_0010110101110101_1001001011010101"; -- 0.17757528023004457
	pesos_i(11994) := b"1111111111111111_1111111111111111_1110001010001111_0000011001011111"; -- -0.11500511347370115
	pesos_i(11995) := b"1111111111111111_1111111111111111_1111011000001100_0111001100000100"; -- -0.03887253913307758
	pesos_i(11996) := b"0000000000000000_0000000000000000_0000010111100100_1110110101100110"; -- 0.023024403893436293
	pesos_i(11997) := b"0000000000000000_0000000000000000_0000111100100110_0010101100011111"; -- 0.05917615420561375
	pesos_i(11998) := b"0000000000000000_0000000000000000_0000111111011101_1011100011111001"; -- 0.061976967628266634
	pesos_i(11999) := b"1111111111111111_1111111111111111_1101011100101001_0111001010000111"; -- -0.15952381325504011
	pesos_i(12000) := b"0000000000000000_0000000000000000_0001110010110110_0111010011101010"; -- 0.11215906833941894
	pesos_i(12001) := b"1111111111111111_1111111111111111_1101110110011001_0101100011010011"; -- -0.13437886083130396
	pesos_i(12002) := b"1111111111111111_1111111111111111_1101110010011110_1111000011101010"; -- -0.1381997518026701
	pesos_i(12003) := b"0000000000000000_0000000000000000_0000111111011010_0110001110011010"; -- 0.06192610269039859
	pesos_i(12004) := b"0000000000000000_0000000000000000_0000010100110000_0101001100000101"; -- 0.020268620115594688
	pesos_i(12005) := b"0000000000000000_0000000000000000_0000010101110101_0101101011110010"; -- 0.021321949139813032
	pesos_i(12006) := b"0000000000000000_0000000000000000_0000000000111011_0100011111011011"; -- 0.0009045515760702753
	pesos_i(12007) := b"1111111111111111_1111111111111111_1101101000011001_0110000101100101"; -- -0.14805022519765101
	pesos_i(12008) := b"0000000000000000_0000000000000000_0000010010110110_0100011100101000"; -- 0.01840634082172484
	pesos_i(12009) := b"1111111111111111_1111111111111111_1101111110010110_0000110001110101"; -- -0.12661668914859286
	pesos_i(12010) := b"1111111111111111_1111111111111111_1101110001101100_1110001100110101"; -- -0.13896350809403674
	pesos_i(12011) := b"1111111111111111_1111111111111111_1111111101001001_0010010000100100"; -- -0.002790204267794976
	pesos_i(12012) := b"1111111111111111_1111111111111111_1110001111110000_0001011111000101"; -- -0.10961772392926529
	pesos_i(12013) := b"0000000000000000_0000000000000000_0001000011101001_1110101111011011"; -- 0.06606935603004097
	pesos_i(12014) := b"1111111111111111_1111111111111111_1111100000101101_0001100101111001"; -- -0.03056183611425747
	pesos_i(12015) := b"1111111111111111_1111111111111111_1110011111001000_0111000000000100"; -- -0.09459781564686846
	pesos_i(12016) := b"0000000000000000_0000000000000000_0001100110000111_1100011000100000"; -- 0.09972799563889242
	pesos_i(12017) := b"0000000000000000_0000000000000000_0001001010100101_1011011011000000"; -- 0.07284109284720669
	pesos_i(12018) := b"0000000000000000_0000000000000000_0000000010000000_0000110000011011"; -- 0.001953846570656523
	pesos_i(12019) := b"0000000000000000_0000000000000000_0000000111010001_0010011010100111"; -- 0.007097640727932226
	pesos_i(12020) := b"0000000000000000_0000000000000000_0000001101010100_1000001001011101"; -- 0.013008258598037423
	pesos_i(12021) := b"1111111111111111_1111111111111111_1110010101100111_0000010011100000"; -- -0.10389680419692401
	pesos_i(12022) := b"0000000000000000_0000000000000000_0010001011000001_1001001100010111"; -- 0.1357662135538415
	pesos_i(12023) := b"0000000000000000_0000000000000000_0000101001110110_0111100110010101"; -- 0.04087028393851524
	pesos_i(12024) := b"1111111111111111_1111111111111111_1111111010111001_0100011001111011"; -- -0.004985423071938966
	pesos_i(12025) := b"1111111111111111_1111111111111111_1110110101110101_1000101111010111"; -- -0.07242513665840353
	pesos_i(12026) := b"0000000000000000_0000000000000000_0001000101111101_1101100101110000"; -- 0.0683265589462962
	pesos_i(12027) := b"1111111111111111_1111111111111111_1110010011110000_0101100001110100"; -- -0.10570761838546279
	pesos_i(12028) := b"1111111111111111_1111111111111111_1111001100111001_0000011011100000"; -- -0.04991108919484738
	pesos_i(12029) := b"0000000000000000_0000000000000000_0000010000110110_0110100110001111"; -- 0.016455266325539595
	pesos_i(12030) := b"1111111111111111_1111111111111111_1111000001111000_0010111100111111"; -- -0.06066612916359832
	pesos_i(12031) := b"0000000000000000_0000000000000000_0001101100010000_0000111001001111"; -- 0.10571374348716203
	pesos_i(12032) := b"0000000000000000_0000000000000000_0001110010111110_1001010100110100"; -- 0.11228306311997625
	pesos_i(12033) := b"1111111111111111_1111111111111111_1110101111011100_0000100011111100"; -- -0.07867378087209474
	pesos_i(12034) := b"0000000000000000_0000000000000000_0000100001111010_1011010001100011"; -- 0.03312232406743086
	pesos_i(12035) := b"1111111111111111_1111111111111111_1110000110111110_0101001010101000"; -- -0.11818965328629051
	pesos_i(12036) := b"0000000000000000_0000000000000000_0000110011100110_0011010011010010"; -- 0.05038766981761442
	pesos_i(12037) := b"0000000000000000_0000000000000000_0001101001010000_1111110010101111"; -- 0.1027982643354638
	pesos_i(12038) := b"0000000000000000_0000000000000000_0010100010101010_1001111010101001"; -- 0.15885345110931606
	pesos_i(12039) := b"1111111111111111_1111111111111111_1111011100010110_0001110011110111"; -- -0.03481883010113666
	pesos_i(12040) := b"0000000000000000_0000000000000000_0001110000111100_1111010001000000"; -- 0.11030508573247677
	pesos_i(12041) := b"1111111111111111_1111111111111111_1110010010101010_0100001101101111"; -- -0.10677698639665038
	pesos_i(12042) := b"1111111111111111_1111111111111111_1111000000101110_1111110001101100"; -- -0.061783050089458245
	pesos_i(12043) := b"1111111111111111_1111111111111111_1110101111110001_1001001001101111"; -- -0.07834515364075713
	pesos_i(12044) := b"1111111111111111_1111111111111111_1111000001010111_0011100011001011"; -- -0.061169100237948006
	pesos_i(12045) := b"1111111111111111_1111111111111111_1111111000100001_1100000011101111"; -- -0.007297460283900836
	pesos_i(12046) := b"0000000000000000_0000000000000000_0000001000100100_1010100010010100"; -- 0.008371864367905279
	pesos_i(12047) := b"1111111111111111_1111111111111111_1110000010111011_0010100110100010"; -- -0.12214412499454402
	pesos_i(12048) := b"0000000000000000_0000000000000000_0000000111000110_0010100100010011"; -- 0.006929938374764569
	pesos_i(12049) := b"0000000000000000_0000000000000000_0000111101010110_1010010111000001"; -- 0.059915885531293435
	pesos_i(12050) := b"0000000000000000_0000000000000000_0001001001001010_0000000011101101"; -- 0.0714417054910333
	pesos_i(12051) := b"1111111111111111_1111111111111111_1111011011000101_1101100111011101"; -- -0.036043532876975475
	pesos_i(12052) := b"1111111111111111_1111111111111111_1110110111101101_1100010101010011"; -- -0.07059065549275531
	pesos_i(12053) := b"1111111111111111_1111111111111111_1110100111010110_0111011100011111"; -- -0.0865712690492626
	pesos_i(12054) := b"1111111111111111_1111111111111111_1111101010110101_0100100101100010"; -- -0.02067128533251314
	pesos_i(12055) := b"1111111111111111_1111111111111111_1110010001101101_1011001010110101"; -- -0.10770114013986665
	pesos_i(12056) := b"1111111111111111_1111111111111111_1111010111000011_0000110110010011"; -- -0.03999247709805852
	pesos_i(12057) := b"1111111111111111_1111111111111111_1101111010100011_0111010100001100"; -- -0.1303183408003294
	pesos_i(12058) := b"1111111111111111_1111111111111111_1110100111010110_1110011011010101"; -- -0.08656461036513452
	pesos_i(12059) := b"0000000000000000_0000000000000000_0000010111001001_1011011000010010"; -- 0.022609118785682832
	pesos_i(12060) := b"1111111111111111_1111111111111111_1111011101110111_1101000010010010"; -- -0.03332802229587576
	pesos_i(12061) := b"1111111111111111_1111111111111111_1101101011010110_1001001101000110"; -- -0.14516334086805754
	pesos_i(12062) := b"1111111111111111_1111111111111111_1110010000101001_0010100001100111"; -- -0.10874698142844158
	pesos_i(12063) := b"0000000000000000_0000000000000000_0001000010111000_0001011111000111"; -- 0.06530903449995239
	pesos_i(12064) := b"0000000000000000_0000000000000000_0001101000001100_0110001101111011"; -- 0.10175153492686571
	pesos_i(12065) := b"1111111111111111_1111111111111111_1101111011110011_1111110000110011"; -- -0.12908958196780582
	pesos_i(12066) := b"0000000000000000_0000000000000000_0000000000011000_0101001010010100"; -- 0.00037113306690558285
	pesos_i(12067) := b"0000000000000000_0000000000000000_0000110011101001_1010111000101101"; -- 0.05044067954511411
	pesos_i(12068) := b"1111111111111111_1111111111111111_1111011100001101_0001101000001000"; -- -0.03495633410262192
	pesos_i(12069) := b"0000000000000000_0000000000000000_0001101111100000_0100111011100010"; -- 0.10889142055124088
	pesos_i(12070) := b"0000000000000000_0000000000000000_0010110110000000_1011011100011101"; -- 0.17774528940567125
	pesos_i(12071) := b"0000000000000000_0000000000000000_0001111001111001_0011101111110100"; -- 0.11903738694653479
	pesos_i(12072) := b"0000000000000000_0000000000000000_0001011110010100_1011000011010111"; -- 0.09211259114359868
	pesos_i(12073) := b"0000000000000000_0000000000000000_0000010000011111_1011001110000001"; -- 0.01610872180399297
	pesos_i(12074) := b"0000000000000000_0000000000000000_0000110100000011_1010110110010000"; -- 0.05083737146482018
	pesos_i(12075) := b"0000000000000000_0000000000000000_0010001011100111_1101000101011011"; -- 0.13634975890813364
	pesos_i(12076) := b"1111111111111111_1111111111111111_1101100111000110_1010010011101101"; -- -0.14931267950436589
	pesos_i(12077) := b"1111111111111111_1111111111111111_1110011110101011_0111001101011001"; -- -0.09504012180250139
	pesos_i(12078) := b"1111111111111111_1111111111111111_1110101101100101_1000101111110001"; -- -0.0804817711433655
	pesos_i(12079) := b"0000000000000000_0000000000000000_0000110010000010_1111110100100010"; -- 0.04887373040684226
	pesos_i(12080) := b"1111111111111111_1111111111111111_1110110011110010_0101011100010111"; -- -0.07442718204804702
	pesos_i(12081) := b"0000000000000000_0000000000000000_0010011001010001_0100101100010011"; -- 0.14967793661557002
	pesos_i(12082) := b"1111111111111111_1111111111111111_1110000010101010_1111000101011110"; -- -0.12239161916949634
	pesos_i(12083) := b"1111111111111111_1111111111111111_1111001010101010_1000101100100110"; -- -0.0520852119307511
	pesos_i(12084) := b"0000000000000000_0000000000000000_0000100110001001_1001010110100101"; -- 0.037255623511548715
	pesos_i(12085) := b"0000000000000000_0000000000000000_0001101111111010_1010001011110101"; -- 0.10929316015197435
	pesos_i(12086) := b"0000000000000000_0000000000000000_0010011101000101_1111101100001011"; -- 0.1534115697715161
	pesos_i(12087) := b"0000000000000000_0000000000000000_0001001011011011_1001011001001001"; -- 0.07366313244728966
	pesos_i(12088) := b"1111111111111111_1111111111111111_1111101010110011_1111001100110110"; -- -0.020691680141457006
	pesos_i(12089) := b"1111111111111111_1111111111111111_1110100110101010_0101001001011101"; -- -0.08724484665970653
	pesos_i(12090) := b"0000000000000000_0000000000000000_0000101110011101_1000100101110111"; -- 0.045372573505590916
	pesos_i(12091) := b"1111111111111111_1111111111111111_1111010001011001_0100010111100001"; -- -0.045512802636437893
	pesos_i(12092) := b"0000000000000000_0000000000000000_0000011100111100_1010011111100011"; -- 0.028269284274867787
	pesos_i(12093) := b"0000000000000000_0000000000000000_0001011101110100_1001000000011100"; -- 0.09162235900907623
	pesos_i(12094) := b"1111111111111111_1111111111111111_1111101011101011_0000010101100100"; -- -0.01985136336855247
	pesos_i(12095) := b"0000000000000000_0000000000000000_0001100101111100_1010110100111001"; -- 0.09955866460794006
	pesos_i(12096) := b"1111111111111111_1111111111111111_1110011011011111_1010111010010000"; -- -0.09814938519759174
	pesos_i(12097) := b"0000000000000000_0000000000000000_0001100100000100_1010110110110001"; -- 0.09772763794195574
	pesos_i(12098) := b"1111111111111111_1111111111111111_1101101011111000_0000111011111100"; -- -0.14465242711449822
	pesos_i(12099) := b"1111111111111111_1111111111111111_1111111110000101_1101001110011101"; -- -0.001864217913899417
	pesos_i(12100) := b"0000000000000000_0000000000000000_0001001100010001_1100100100100101"; -- 0.07449013860158751
	pesos_i(12101) := b"0000000000000000_0000000000000000_0001000101100000_1100110101101011"; -- 0.06788333767499737
	pesos_i(12102) := b"1111111111111111_1111111111111111_1110000000010100_0111010101010010"; -- -0.12468783138384555
	pesos_i(12103) := b"0000000000000000_0000000000000000_0000101100000110_0000000011110001"; -- 0.04306035887836453
	pesos_i(12104) := b"1111111111111111_1111111111111111_1101011110100010_0011010111000000"; -- -0.15768112246220065
	pesos_i(12105) := b"1111111111111111_1111111111111111_1110100010000110_1110010001000011"; -- -0.09169171674881499
	pesos_i(12106) := b"1111111111111111_1111111111111111_1110010100010010_0011111101010111"; -- -0.10519031639392629
	pesos_i(12107) := b"1111111111111111_1111111111111111_1111000101010011_0010011100100110"; -- -0.057324936976506355
	pesos_i(12108) := b"1111111111111111_1111111111111111_1111010000101111_0110001000110010"; -- -0.04615198396920333
	pesos_i(12109) := b"0000000000000000_0000000000000000_0000001101000101_0100100111010101"; -- 0.012776007280406313
	pesos_i(12110) := b"1111111111111111_1111111111111111_1110011111010010_1000111001101101"; -- -0.09444341517031597
	pesos_i(12111) := b"1111111111111111_1111111111111111_1111101100100110_0001010001011001"; -- -0.018950203140680327
	pesos_i(12112) := b"0000000000000000_0000000000000000_0001011100011010_0110010110010100"; -- 0.09024653299047405
	pesos_i(12113) := b"0000000000000000_0000000000000000_0001111011010011_1001111011110001"; -- 0.12041657822027917
	pesos_i(12114) := b"0000000000000000_0000000000000000_0000101010100111_0010010110111011"; -- 0.041612966652458463
	pesos_i(12115) := b"0000000000000000_0000000000000000_0001100100101001_1110011011011100"; -- 0.09829562064961914
	pesos_i(12116) := b"1111111111111111_1111111111111111_1111110001100000_1111001000000101"; -- -0.01414573077828051
	pesos_i(12117) := b"0000000000000000_0000000000000000_0001000100011100_1111111100110010"; -- 0.06684870700062016
	pesos_i(12118) := b"0000000000000000_0000000000000000_0010000100111110_0100001011010100"; -- 0.1298562782004319
	pesos_i(12119) := b"0000000000000000_0000000000000000_0000000110110111_0100011100001010"; -- 0.006702842703978691
	pesos_i(12120) := b"0000000000000000_0000000000000000_0000010011100010_0101001011100001"; -- 0.019078426216966475
	pesos_i(12121) := b"1111111111111111_1111111111111111_1101110100111101_1100101001101101"; -- -0.1357758982680071
	pesos_i(12122) := b"0000000000000000_0000000000000000_0000100111101000_0110101110001010"; -- 0.03870269895341889
	pesos_i(12123) := b"0000000000000000_0000000000000000_0010011000000110_0111010001001011"; -- 0.14853598431105716
	pesos_i(12124) := b"1111111111111111_1111111111111111_1101111101100010_1111111010111100"; -- -0.12739570523118282
	pesos_i(12125) := b"0000000000000000_0000000000000000_0001010010101111_1100010110001111"; -- 0.0808070634469265
	pesos_i(12126) := b"0000000000000000_0000000000000000_0001010000001110_0011101111101101"; -- 0.07834219500878027
	pesos_i(12127) := b"1111111111111111_1111111111111111_1110000101010010_0000001000001110"; -- -0.11984240690674497
	pesos_i(12128) := b"0000000000000000_0000000000000000_0001011000000000_1101010000010011"; -- 0.08595014061504175
	pesos_i(12129) := b"0000000000000000_0000000000000000_0000000101000101_0001110001100000"; -- 0.004960797775788746
	pesos_i(12130) := b"1111111111111111_1111111111111111_1101110010010111_0100110101001010"; -- -0.13831631605260994
	pesos_i(12131) := b"0000000000000000_0000000000000000_0000001110011101_1010100110111010"; -- 0.014124496400400663
	pesos_i(12132) := b"0000000000000000_0000000000000000_0001010100010100_1011010010101101"; -- 0.08234719499036806
	pesos_i(12133) := b"1111111111111111_1111111111111111_1110101011010111_1110111000100110"; -- -0.08264266553719048
	pesos_i(12134) := b"0000000000000000_0000000000000000_0000011110101001_1001000100001101"; -- 0.029931131027055958
	pesos_i(12135) := b"1111111111111111_1111111111111111_1101111000101011_0000111001011101"; -- -0.13215551591318903
	pesos_i(12136) := b"0000000000000000_0000000000000000_0001001100101001_1010101100010001"; -- 0.07485455676550122
	pesos_i(12137) := b"0000000000000000_0000000000000000_0010010000011100_0000111001001111"; -- 0.14105309884613226
	pesos_i(12138) := b"1111111111111111_1111111111111111_1111100110110111_0101101000110110"; -- -0.024546014552138992
	pesos_i(12139) := b"1111111111111111_1111111111111111_1110100110000101_0100001001111110"; -- -0.08781036782226602
	pesos_i(12140) := b"1111111111111111_1111111111111111_1111001111110100_0011010010000010"; -- -0.047054975683200995
	pesos_i(12141) := b"1111111111111111_1111111111111111_1110001001101101_0111000010111111"; -- -0.11551757170161536
	pesos_i(12142) := b"0000000000000000_0000000000000000_0000000100111010_0101100000011010"; -- 0.004796511085920344
	pesos_i(12143) := b"1111111111111111_1111111111111111_1111111100110001_0011111111011100"; -- -0.0031547630269739392
	pesos_i(12144) := b"1111111111111111_1111111111111111_1111011100001010_1101001011010000"; -- -0.034991096657014276
	pesos_i(12145) := b"0000000000000000_0000000000000000_0000010011010000_1001001001110110"; -- 0.01880755785593074
	pesos_i(12146) := b"0000000000000000_0000000000000000_0000111110000110_1000101100011110"; -- 0.06064671965100886
	pesos_i(12147) := b"1111111111111111_1111111111111111_1110111000000101_1010110000010101"; -- -0.07022594912143369
	pesos_i(12148) := b"0000000000000000_0000000000000000_0000001111100100_0001110101111001"; -- 0.015199510691772682
	pesos_i(12149) := b"1111111111111111_1111111111111111_1111000100101111_1101010111000101"; -- -0.057863845224725596
	pesos_i(12150) := b"1111111111111111_1111111111111111_1111011001111111_1001011100011110"; -- -0.037115626485853474
	pesos_i(12151) := b"1111111111111111_1111111111111111_1111011110111011_1010001010010111"; -- -0.0322931653368699
	pesos_i(12152) := b"0000000000000000_0000000000000000_0001001001000001_1110111111000001"; -- 0.07131861163957527
	pesos_i(12153) := b"0000000000000000_0000000000000000_0000111100100010_1100011101010111"; -- 0.059124430324291995
	pesos_i(12154) := b"1111111111111111_1111111111111111_1111000101000110_1010001010001011"; -- -0.05751594635661405
	pesos_i(12155) := b"0000000000000000_0000000000000000_0001111101100011_0001010001111011"; -- 0.12260559085989975
	pesos_i(12156) := b"1111111111111111_1111111111111111_1111100010110111_1010001111001011"; -- -0.028447878806225735
	pesos_i(12157) := b"0000000000000000_0000000000000000_0000011111010001_0100010100100101"; -- 0.030536958321691707
	pesos_i(12158) := b"0000000000000000_0000000000000000_0000011000100011_1101101011110011"; -- 0.02398460802328941
	pesos_i(12159) := b"1111111111111111_1111111111111111_1110010010010110_0000001110011100"; -- -0.1070859665518683
	pesos_i(12160) := b"1111111111111111_1111111111111111_1110000100111100_1000001010101111"; -- -0.12017043332782293
	pesos_i(12161) := b"0000000000000000_0000000000000000_0000000101001101_0010111110001101"; -- 0.005084011071764602
	pesos_i(12162) := b"1111111111111111_1111111111111111_1110101001110110_1010100101001000"; -- -0.08412687291611397
	pesos_i(12163) := b"0000000000000000_0000000000000000_0001011000111100_1001110111000101"; -- 0.08686243120889918
	pesos_i(12164) := b"0000000000000000_0000000000000000_0001011010101000_0011110000111111"; -- 0.08850456744867968
	pesos_i(12165) := b"0000000000000000_0000000000000000_0000011001010011_0000111011000110"; -- 0.0247048600265272
	pesos_i(12166) := b"0000000000000000_0000000000000000_0010010000111110_0001100000111011"; -- 0.1415724890825055
	pesos_i(12167) := b"0000000000000000_0000000000000000_0000000011000001_1101000101010100"; -- 0.0029574232217761663
	pesos_i(12168) := b"1111111111111111_1111111111111111_1110101111111011_0110110011111100"; -- -0.07819479792718893
	pesos_i(12169) := b"0000000000000000_0000000000000000_0001111001001001_1001111100101010"; -- 0.11831087842600742
	pesos_i(12170) := b"0000000000000000_0000000000000000_0001001100000100_0100101011011001"; -- 0.07428424630893055
	pesos_i(12171) := b"1111111111111111_1111111111111111_1110100101000010_0000010101011111"; -- -0.08883634981915758
	pesos_i(12172) := b"0000000000000000_0000000000000000_0001011110000101_0111010001100001"; -- 0.09188010570872844
	pesos_i(12173) := b"0000000000000000_0000000000000000_0000110001101011_0011101101011001"; -- 0.048511227908772006
	pesos_i(12174) := b"1111111111111111_1111111111111111_1110110001001110_1101010010111100"; -- -0.07692213451567237
	pesos_i(12175) := b"1111111111111111_1111111111111111_1110100100010100_0110000111100100"; -- -0.0895327395537297
	pesos_i(12176) := b"1111111111111111_1111111111111111_1111100100001100_1100100101101011"; -- -0.027148639042790485
	pesos_i(12177) := b"1111111111111111_1111111111111111_1101110001000001_1101111001010010"; -- -0.13961992739395424
	pesos_i(12178) := b"0000000000000000_0000000000000000_0010001110111011_1100100010011101"; -- 0.1395841010736134
	pesos_i(12179) := b"1111111111111111_1111111111111111_1110011101100101_0001101110110011"; -- -0.09611346131908931
	pesos_i(12180) := b"1111111111111111_1111111111111111_1111101011001011_0010100110010000"; -- -0.020337488536143103
	pesos_i(12181) := b"1111111111111111_1111111111111111_1110111000001101_0110110101010101"; -- -0.07010761912900325
	pesos_i(12182) := b"1111111111111111_1111111111111111_1110101011110001_1100101110010110"; -- -0.08224799714039734
	pesos_i(12183) := b"1111111111111111_1111111111111111_1111011100101101_1101011111001111"; -- -0.03445674120664164
	pesos_i(12184) := b"1111111111111111_1111111111111111_1110110111101111_1111001111110011"; -- -0.07055735899168708
	pesos_i(12185) := b"1111111111111111_1111111111111111_1110010001010010_0011000110000100"; -- -0.10812082782284334
	pesos_i(12186) := b"0000000000000000_0000000000000000_0001000110001100_1101010001101011"; -- 0.06855514150606688
	pesos_i(12187) := b"0000000000000000_0000000000000000_0000010001000000_1101101100010101"; -- 0.016614620906008248
	pesos_i(12188) := b"0000000000000000_0000000000000000_0010100010001110_0000110010001110"; -- 0.15841749642698205
	pesos_i(12189) := b"0000000000000000_0000000000000000_0001010100101100_1101000010010110"; -- 0.08271506936659238
	pesos_i(12190) := b"0000000000000000_0000000000000000_0001111100011111_1000110101101110"; -- 0.12157520232119619
	pesos_i(12191) := b"1111111111111111_1111111111111111_1101111010100011_0011000000010111"; -- -0.1303224509617378
	pesos_i(12192) := b"0000000000000000_0000000000000000_0000111110011100_0111001111001011"; -- 0.06098102280517946
	pesos_i(12193) := b"0000000000000000_0000000000000000_0000001101011011_1101000100010000"; -- 0.013119760928274616
	pesos_i(12194) := b"0000000000000000_0000000000000000_0000001010001001_0110011001100000"; -- 0.00990905605152313
	pesos_i(12195) := b"0000000000000000_0000000000000000_0001011000111001_0011001010011000"; -- 0.08681026660972657
	pesos_i(12196) := b"1111111111111111_1111111111111111_1110110101000111_1101011111111000"; -- -0.07312250327039861
	pesos_i(12197) := b"1111111111111111_1111111111111111_1110100000011010_0011000101100101"; -- -0.09335032724170203
	pesos_i(12198) := b"0000000000000000_0000000000000000_0000011111001110_1001111000111110"; -- 0.03049649250148432
	pesos_i(12199) := b"0000000000000000_0000000000000000_0000001110010100_0101010111000000"; -- 0.013982161887306931
	pesos_i(12200) := b"1111111111111111_1111111111111111_1111101111000001_1011110111000101"; -- -0.016574992610769904
	pesos_i(12201) := b"1111111111111111_1111111111111111_1110011100101101_1101100000010010"; -- -0.09695672568043952
	pesos_i(12202) := b"1111111111111111_1111111111111111_1101111000100000_0010000011000011"; -- -0.1323222660126613
	pesos_i(12203) := b"0000000000000000_0000000000000000_0001011110100110_0111101000000000"; -- 0.09238398085915202
	pesos_i(12204) := b"1111111111111111_1111111111111111_1111010110010010_0101101000000111"; -- -0.04073560075762536
	pesos_i(12205) := b"0000000000000000_0000000000000000_0000001000101000_1010110110000100"; -- 0.008433193816472265
	pesos_i(12206) := b"1111111111111111_1111111111111111_1101110111110100_0001111001000100"; -- -0.13299380152142062
	pesos_i(12207) := b"0000000000000000_0000000000000000_0000110110010001_1101110010101111"; -- 0.053006928235653145
	pesos_i(12208) := b"1111111111111111_1111111111111111_1111111101100001_1110011110111010"; -- -0.002412335467785139
	pesos_i(12209) := b"1111111111111111_1111111111111111_1110001100001101_0000011111010011"; -- -0.11308241941603182
	pesos_i(12210) := b"1111111111111111_1111111111111111_1111100000010111_1111000010000001"; -- -0.03088471272083238
	pesos_i(12211) := b"1111111111111111_1111111111111111_1101100110110100_0011001011001110"; -- -0.14959413980049552
	pesos_i(12212) := b"0000000000000000_0000000000000000_0000011010111010_0111101111110010"; -- 0.02628302240968885
	pesos_i(12213) := b"1111111111111111_1111111111111111_1110000101011100_0110000001101110"; -- -0.11968419371496558
	pesos_i(12214) := b"1111111111111111_1111111111111111_1110111000000011_1001110010001111"; -- -0.07025739210065299
	pesos_i(12215) := b"0000000000000000_0000000000000000_0001101000010111_0110110111001100"; -- 0.10191999647313647
	pesos_i(12216) := b"0000000000000000_0000000000000000_0010001001000111_0110110011101111"; -- 0.133902367022776
	pesos_i(12217) := b"1111111111111111_1111111111111111_1110010001000100_0000011001101101"; -- -0.10833701939012252
	pesos_i(12218) := b"1111111111111111_1111111111111111_1101100100110010_0010011100010010"; -- -0.1515784817359846
	pesos_i(12219) := b"0000000000000000_0000000000000000_0000110000100100_0011011110101011"; -- 0.04742763454634612
	pesos_i(12220) := b"0000000000000000_0000000000000000_0000111010011000_1110011111100010"; -- 0.05702065733178873
	pesos_i(12221) := b"1111111111111111_1111111111111111_1111111100001101_0101101111011100"; -- -0.0037024105779541864
	pesos_i(12222) := b"0000000000000000_0000000000000000_0010001100000000_0101011111001010"; -- 0.1367239826030549
	pesos_i(12223) := b"0000000000000000_0000000000000000_0000110101111001_0100011000101111"; -- 0.052631746850725615
	pesos_i(12224) := b"1111111111111111_1111111111111111_1111000001100000_1011010110010110"; -- -0.06102433288062013
	pesos_i(12225) := b"0000000000000000_0000000000000000_0000000110000001_0010100110001110"; -- 0.005877110679414437
	pesos_i(12226) := b"0000000000000000_0000000000000000_0001011001110100_1011101100011101"; -- 0.08771867224471477
	pesos_i(12227) := b"0000000000000000_0000000000000000_0001010111111110_0011101100010101"; -- 0.08591050390491324
	pesos_i(12228) := b"1111111111111111_1111111111111111_1110001001110101_1110011101101111"; -- -0.11538842721004454
	pesos_i(12229) := b"1111111111111111_1111111111111111_1110110010110110_0111001100110000"; -- -0.07534103466274607
	pesos_i(12230) := b"0000000000000000_0000000000000000_0001111000001000_1111000111101010"; -- 0.11732398940875793
	pesos_i(12231) := b"0000000000000000_0000000000000000_0010001001111100_0110000101001001"; -- 0.13471038839915825
	pesos_i(12232) := b"0000000000000000_0000000000000000_0001111101101110_0010011100111101"; -- 0.12277455555753014
	pesos_i(12233) := b"1111111111111111_1111111111111111_1101101101000101_0100100000000001"; -- -0.1434741016911302
	pesos_i(12234) := b"1111111111111111_1111111111111111_1111110110011111_0010100111101111"; -- -0.00929010308681773
	pesos_i(12235) := b"1111111111111111_1111111111111111_1111000111011101_0100101100010010"; -- -0.05521708309923191
	pesos_i(12236) := b"0000000000000000_0000000000000000_0000011010001101_1010110010101110"; -- 0.025599281878222413
	pesos_i(12237) := b"1111111111111111_1111111111111111_1110010001001111_0101001011111011"; -- -0.10816460960455829
	pesos_i(12238) := b"1111111111111111_1111111111111111_1110100111111111_1110010011111101"; -- -0.08593910991925051
	pesos_i(12239) := b"1111111111111111_1111111111111111_1111001011110001_1101100001110110"; -- -0.05099722971666511
	pesos_i(12240) := b"1111111111111111_1111111111111111_1111011001000010_0000000011001000"; -- -0.03805537328934442
	pesos_i(12241) := b"0000000000000000_0000000000000000_0000110100011001_0110101111110110"; -- 0.051169154662442255
	pesos_i(12242) := b"0000000000000000_0000000000000000_0001000100111101_0000000101100011"; -- 0.0673371188374157
	pesos_i(12243) := b"1111111111111111_1111111111111111_1110111100100000_1000101100110001"; -- -0.06590967228103863
	pesos_i(12244) := b"1111111111111111_1111111111111111_1101011111101010_1100101101011011"; -- -0.15657357235538058
	pesos_i(12245) := b"1111111111111111_1111111111111111_1111111000101000_1101111010011010"; -- -0.007188880267029294
	pesos_i(12246) := b"0000000000000000_0000000000000000_0010000010001101_1110010100011011"; -- 0.12716514494066072
	pesos_i(12247) := b"0000000000000000_0000000000000000_0000100000010011_0000101000110011"; -- 0.031540525021912576
	pesos_i(12248) := b"1111111111111111_1111111111111111_1101110100011011_0100101000101111"; -- -0.13630234100216337
	pesos_i(12249) := b"0000000000000000_0000000000000000_0000100100110011_1011110001100110"; -- 0.03594567777998205
	pesos_i(12250) := b"1111111111111111_1111111111111111_1110001001110111_0011010001111111"; -- -0.11536857508388175
	pesos_i(12251) := b"0000000000000000_0000000000000000_0001100011101001_1100011111001010"; -- 0.09731720620289681
	pesos_i(12252) := b"1111111111111111_1111111111111111_1101110111010100_1110000100001011"; -- -0.13347047307786175
	pesos_i(12253) := b"1111111111111111_1111111111111111_1110011110111000_1011001110101000"; -- -0.0948379245171228
	pesos_i(12254) := b"1111111111111111_1111111111111111_1111001001101110_1011101001110010"; -- -0.05299792019396904
	pesos_i(12255) := b"1111111111111111_1111111111111111_1101100101100000_1000011011011001"; -- -0.1508708686236615
	pesos_i(12256) := b"1111111111111111_1111111111111111_1110110111110101_0111011011110001"; -- -0.07047325730092957
	pesos_i(12257) := b"0000000000000000_0000000000000000_0010000011111010_0101100101000010"; -- 0.12882001755487724
	pesos_i(12258) := b"1111111111111111_1111111111111111_1110100000100001_0100010000010110"; -- -0.093242401681139
	pesos_i(12259) := b"1111111111111111_1111111111111111_1110011010001010_1001100011001010"; -- -0.0994476802558275
	pesos_i(12260) := b"0000000000000000_0000000000000000_0001011100011011_1100110011111110"; -- 0.09026795573180148
	pesos_i(12261) := b"1111111111111111_1111111111111111_1110001001100110_1011001010011010"; -- -0.11562045795491808
	pesos_i(12262) := b"0000000000000000_0000000000000000_0000000100010111_1000011111000011"; -- 0.004265294203350103
	pesos_i(12263) := b"1111111111111111_1111111111111111_1110000111101011_0100101110001110"; -- -0.11750343119014338
	pesos_i(12264) := b"0000000000000000_0000000000000000_0000100000111100_0001100001010000"; -- 0.03216697637790336
	pesos_i(12265) := b"0000000000000000_0000000000000000_0001101001010110_0011000111001110"; -- 0.10287772439516235
	pesos_i(12266) := b"1111111111111111_1111111111111111_1110110010101001_0100011000000001"; -- -0.07554209210038443
	pesos_i(12267) := b"0000000000000000_0000000000000000_0001101100001010_0001100011001000"; -- 0.10562281501033455
	pesos_i(12268) := b"1111111111111111_1111111111111111_1111101111000111_1111111011001101"; -- -0.016479563762263758
	pesos_i(12269) := b"0000000000000000_0000000000000000_0001000101100111_1010000110100011"; -- 0.0679875395681787
	pesos_i(12270) := b"1111111111111111_1111111111111111_1111110000110001_1000000100110111"; -- -0.014869617632809135
	pesos_i(12271) := b"0000000000000000_0000000000000000_0001110110010100_0110100000100010"; -- 0.11554575765328172
	pesos_i(12272) := b"1111111111111111_1111111111111111_1101101110001011_0011110010010010"; -- -0.14240666797833357
	pesos_i(12273) := b"1111111111111111_1111111111111111_1111101100111110_1111011000010110"; -- -0.018570537324749486
	pesos_i(12274) := b"0000000000000000_0000000000000000_0000010111010001_0111001110101011"; -- 0.022727231254517533
	pesos_i(12275) := b"0000000000000000_0000000000000000_0000010101001000_1100110100000001"; -- 0.020642102035562233
	pesos_i(12276) := b"1111111111111111_1111111111111111_1111011000110100_0110100100111110"; -- -0.03826277015292656
	pesos_i(12277) := b"1111111111111111_1111111111111111_1111000001100111_0000001001001100"; -- -0.06092820785063461
	pesos_i(12278) := b"0000000000000000_0000000000000000_0001111000001110_0000000000100010"; -- 0.11740113103721632
	pesos_i(12279) := b"1111111111111111_1111111111111111_1110011110011000_0011101101010110"; -- -0.0953333773969376
	pesos_i(12280) := b"0000000000000000_0000000000000000_0001110111110110_1101101000111010"; -- 0.11704791939832923
	pesos_i(12281) := b"0000000000000000_0000000000000000_0010000111101010_0010110011000100"; -- 0.13247947483385883
	pesos_i(12282) := b"1111111111111111_1111111111111111_1101111001000100_1000111111011000"; -- -0.13176632851354125
	pesos_i(12283) := b"0000000000000000_0000000000000000_0001000101111000_0100110111111111"; -- 0.06824195351203086
	pesos_i(12284) := b"0000000000000000_0000000000000000_0000111010101100_1011111011001011"; -- 0.05732338389424794
	pesos_i(12285) := b"1111111111111111_1111111111111111_1111001100100101_1110111100110100"; -- -0.050202417163620845
	pesos_i(12286) := b"1111111111111111_1111111111111111_1110111110101001_0010000010010101"; -- -0.06382557269996296
	pesos_i(12287) := b"1111111111111111_1111111111111111_1101111110000101_1111100001011011"; -- -0.12686202792109427
	pesos_i(12288) := b"1111111111111111_1111111111111111_1111111000001111_0001111001100110"; -- -0.007581806253492949
	pesos_i(12289) := b"1111111111111111_1111111111111111_1101101111011101_1011101000000001"; -- -0.14114797094608064
	pesos_i(12290) := b"0000000000000000_0000000000000000_0001111000000101_0101100010011111"; -- 0.11726907618276686
	pesos_i(12291) := b"0000000000000000_0000000000000000_0000010001100111_1001001001110100"; -- 0.017205384587937102
	pesos_i(12292) := b"0000000000000000_0000000000000000_0001111110010110_0110010000110001"; -- 0.12338854032687382
	pesos_i(12293) := b"1111111111111111_1111111111111111_1110011010010011_0010000000011110"; -- -0.09931754366301317
	pesos_i(12294) := b"0000000000000000_0000000000000000_0001111011011111_0010111101010111"; -- 0.12059303171236822
	pesos_i(12295) := b"0000000000000000_0000000000000000_0001100000110110_1101010110010010"; -- 0.09458670439090315
	pesos_i(12296) := b"0000000000000000_0000000000000000_0001010000111000_1101001100000110"; -- 0.07899207005297258
	pesos_i(12297) := b"1111111111111111_1111111111111111_1111111111010110_0011111001100010"; -- -0.000637150769997358
	pesos_i(12298) := b"1111111111111111_1111111111111111_1101101110000110_1010111011111111"; -- -0.14247614179578838
	pesos_i(12299) := b"0000000000000000_0000000000000000_0001010110111000_0101011001100101"; -- 0.0848440167226867
	pesos_i(12300) := b"1111111111111111_1111111111111111_1101110100011110_1000001011000101"; -- -0.13625319193342963
	pesos_i(12301) := b"1111111111111111_1111111111111111_1101110101011001_0111110001111111"; -- -0.13535329725140213
	pesos_i(12302) := b"0000000000000000_0000000000000000_0000001001100011_0011100111101101"; -- 0.009326572648123945
	pesos_i(12303) := b"1111111111111111_1111111111111111_1110011000100110_0110010011000110"; -- -0.10097665937860327
	pesos_i(12304) := b"1111111111111111_1111111111111111_1111100100110010_0000011011110001"; -- -0.026580396812511425
	pesos_i(12305) := b"0000000000000000_0000000000000000_0001100001000110_0000101100000001"; -- 0.09481877108960207
	pesos_i(12306) := b"1111111111111111_1111111111111111_1110100110000000_0110000001000001"; -- -0.0878848877840795
	pesos_i(12307) := b"1111111111111111_1111111111111111_1111111101101101_0111100000111010"; -- -0.002235875943353188
	pesos_i(12308) := b"1111111111111111_1111111111111111_1111111100111110_0111000111000101"; -- -0.0029534239483162005
	pesos_i(12309) := b"1111111111111111_1111111111111111_1110100000110011_0000110100010000"; -- -0.09297102308669468
	pesos_i(12310) := b"0000000000000000_0000000000000000_0001110100000001_1100101111010010"; -- 0.11330865751933361
	pesos_i(12311) := b"0000000000000000_0000000000000000_0010010011001110_1100001011101010"; -- 0.1437799283350829
	pesos_i(12312) := b"0000000000000000_0000000000000000_0010000010100000_0001101111000001"; -- 0.12744306041122805
	pesos_i(12313) := b"1111111111111111_1111111111111111_1101110000101011_1000100110101000"; -- -0.1399606671813439
	pesos_i(12314) := b"1111111111111111_1111111111111111_1101111110010110_1110100010001101"; -- -0.126603570630449
	pesos_i(12315) := b"1111111111111111_1111111111111111_1111011100110010_0001000100000001"; -- -0.03439229699868075
	pesos_i(12316) := b"1111111111111111_1111111111111111_1110001100101101_0100110110011001"; -- -0.11258997933962632
	pesos_i(12317) := b"1111111111111111_1111111111111111_1111101010110101_0001000101011011"; -- -0.020674624714576737
	pesos_i(12318) := b"1111111111111111_1111111111111111_1110010010101111_0110101100010010"; -- -0.10669833008840439
	pesos_i(12319) := b"1111111111111111_1111111111111111_1110110010110100_0100000011000011"; -- -0.07537455795710661
	pesos_i(12320) := b"0000000000000000_0000000000000000_0001110110110010_1011100011011110"; -- 0.11600833330447104
	pesos_i(12321) := b"0000000000000000_0000000000000000_0001101100101100_1111100000111001"; -- 0.10615493187357976
	pesos_i(12322) := b"1111111111111111_1111111111111111_1111101101001101_1000001000111011"; -- -0.018348560807709198
	pesos_i(12323) := b"1111111111111111_1111111111111111_1110011110000010_1101011010111011"; -- -0.09565980839211483
	pesos_i(12324) := b"0000000000000000_0000000000000000_0000011110110010_0010101000110001"; -- 0.030062329251957884
	pesos_i(12325) := b"0000000000000000_0000000000000000_0010011001000000_0010010100011110"; -- 0.14941627487109915
	pesos_i(12326) := b"0000000000000000_0000000000000000_0000111100111000_1010011000000111"; -- 0.05945813814456492
	pesos_i(12327) := b"0000000000000000_0000000000000000_0001000111111011_0000100010100010"; -- 0.07023672053438283
	pesos_i(12328) := b"0000000000000000_0000000000000000_0000100101111000_1111110101100010"; -- 0.037002407396782545
	pesos_i(12329) := b"1111111111111111_1111111111111111_1110110010000111_0100101000101001"; -- -0.0760606432790236
	pesos_i(12330) := b"0000000000000000_0000000000000000_0000001011000010_1001001011111011"; -- 0.010781465840402946
	pesos_i(12331) := b"0000000000000000_0000000000000000_0000111010101111_0001011010001001"; -- 0.05735913122415708
	pesos_i(12332) := b"0000000000000000_0000000000000000_0001110111001001_1111110111110110"; -- 0.11636340377444898
	pesos_i(12333) := b"1111111111111111_1111111111111111_1110000010010011_1110111110101101"; -- -0.12274267219492853
	pesos_i(12334) := b"0000000000000000_0000000000000000_0000100011110011_0001000101100111"; -- 0.034958923036485144
	pesos_i(12335) := b"0000000000000000_0000000000000000_0001000110000010_0101010100000101"; -- 0.06839496005396142
	pesos_i(12336) := b"0000000000000000_0000000000000000_0001001110000100_0011100000010001"; -- 0.07623625203542052
	pesos_i(12337) := b"1111111111111111_1111111111111111_1110001110100011_1011011100000001"; -- -0.11078315947422297
	pesos_i(12338) := b"1111111111111111_1111111111111111_1110101010010100_1100111110000100"; -- -0.08366683043427335
	pesos_i(12339) := b"1111111111111111_1111111111111111_1101111111111011_1111110000011010"; -- -0.12506126749549912
	pesos_i(12340) := b"1111111111111111_1111111111111111_1101100000011010_1011100110100011"; -- -0.15584220675557348
	pesos_i(12341) := b"1111111111111111_1111111111111111_1110001100110010_1000001110110011"; -- -0.11251046054995345
	pesos_i(12342) := b"0000000000000000_0000000000000000_0010000111010000_0011001110000011"; -- 0.13208314846242208
	pesos_i(12343) := b"1111111111111111_1111111111111111_1111010101100011_0111101110000100"; -- -0.041450767877210866
	pesos_i(12344) := b"0000000000000000_0000000000000000_0000001111010110_1110111100110001"; -- 0.014998387775927912
	pesos_i(12345) := b"0000000000000000_0000000000000000_0001011111010111_1001101011001001"; -- 0.09313361555621423
	pesos_i(12346) := b"1111111111111111_1111111111111111_1111010011001001_0101011000110100"; -- -0.04380284536421285
	pesos_i(12347) := b"1111111111111111_1111111111111111_1111110101111110_0010101011001110"; -- -0.009793591243829364
	pesos_i(12348) := b"1111111111111111_1111111111111111_1110011001111011_0011100111100011"; -- -0.09968221860233153
	pesos_i(12349) := b"1111111111111111_1111111111111111_1111101111101110_1110001100110010"; -- -0.015886116295769484
	pesos_i(12350) := b"1111111111111111_1111111111111111_1111110100010101_1101000110001100"; -- -0.011385825368316808
	pesos_i(12351) := b"1111111111111111_1111111111111111_1111000110101000_1101011111110000"; -- -0.056017402635563006
	pesos_i(12352) := b"0000000000000000_0000000000000000_0010000101011001_0011000011011100"; -- 0.13026719438663326
	pesos_i(12353) := b"0000000000000000_0000000000000000_0001100100011010_0001011001001000"; -- 0.09805430657395996
	pesos_i(12354) := b"1111111111111111_1111111111111111_1110010110101010_1111111101111011"; -- -0.10285952812215497
	pesos_i(12355) := b"1111111111111111_1111111111111111_1101101000011101_1100000001111010"; -- -0.14798352257777972
	pesos_i(12356) := b"1111111111111111_1111111111111111_1111111000010011_1011001011111000"; -- -0.00751191552270244
	pesos_i(12357) := b"0000000000000000_0000000000000000_0000100001010010_1100000010100101"; -- 0.0325127031311815
	pesos_i(12358) := b"1111111111111111_1111111111111111_1110100010000101_1101000101100010"; -- -0.09170810075138004
	pesos_i(12359) := b"0000000000000000_0000000000000000_0000001101110010_0111100010110001"; -- 0.013465445626159837
	pesos_i(12360) := b"0000000000000000_0000000000000000_0001111000011010_0000100100111111"; -- 0.11758477971997353
	pesos_i(12361) := b"0000000000000000_0000000000000000_0010001001110001_0110110011111010"; -- 0.13454323865383797
	pesos_i(12362) := b"0000000000000000_0000000000000000_0001010100110100_1110111100010001"; -- 0.08283895646687134
	pesos_i(12363) := b"0000000000000000_0000000000000000_0000101111011001_0000100111101111"; -- 0.04628049931935365
	pesos_i(12364) := b"1111111111111111_1111111111111111_1101101111011011_0111000001100111"; -- -0.1411828753961096
	pesos_i(12365) := b"1111111111111111_1111111111111111_1101101110011110_0101100101110101"; -- -0.14211502917059587
	pesos_i(12366) := b"1111111111111111_1111111111111111_1111011110010001_0000001100100000"; -- -0.03294353925247379
	pesos_i(12367) := b"1111111111111111_1111111111111111_1110011000011000_1101000011000001"; -- -0.10118384635806522
	pesos_i(12368) := b"1111111111111111_1111111111111111_1111100100100000_1111100100010001"; -- -0.026840623217378772
	pesos_i(12369) := b"1111111111111111_1111111111111111_1111100110101001_1100000010011001"; -- -0.024753535003610085
	pesos_i(12370) := b"1111111111111111_1111111111111111_1101111010011010_0001110100010001"; -- -0.13046091410513838
	pesos_i(12371) := b"1111111111111111_1111111111111111_1111000010110001_1011101000101110"; -- -0.05978809710210118
	pesos_i(12372) := b"1111111111111111_1111111111111111_1111100100110011_1111100010111001"; -- -0.026550726684823382
	pesos_i(12373) := b"0000000000000000_0000000000000000_0001101100010111_0010011100011101"; -- 0.10582203356815138
	pesos_i(12374) := b"1111111111111111_1111111111111111_1111001000100111_1110101011011110"; -- -0.05407840815697748
	pesos_i(12375) := b"1111111111111111_1111111111111111_1101111000100111_1000110010111010"; -- -0.13220901937246704
	pesos_i(12376) := b"0000000000000000_0000000000000000_0000111111110100_1110100100011010"; -- 0.062330788459479494
	pesos_i(12377) := b"1111111111111111_1111111111111111_1110000110010100_0101011101110011"; -- -0.1188302367565297
	pesos_i(12378) := b"1111111111111111_1111111111111111_1101110100010100_1001111100000011"; -- -0.1364040962712076
	pesos_i(12379) := b"1111111111111111_1111111111111111_1111011101000110_0011111111001011"; -- -0.034084332494155996
	pesos_i(12380) := b"0000000000000000_0000000000000000_0000100110010011_1000110110111101"; -- 0.03740774033971224
	pesos_i(12381) := b"0000000000000000_0000000000000000_0000110100000011_0010110101010110"; -- 0.0508297285979787
	pesos_i(12382) := b"0000000000000000_0000000000000000_0010001101011000_0000000001000110"; -- 0.13806153962493506
	pesos_i(12383) := b"1111111111111111_1111111111111111_1111100010101100_1101011011111011"; -- -0.028612674448541358
	pesos_i(12384) := b"0000000000000000_0000000000000000_0001100110011100_1111010001001101"; -- 0.10005118262478832
	pesos_i(12385) := b"0000000000000000_0000000000000000_0001010100101001_1010001100001001"; -- 0.08266657795544421
	pesos_i(12386) := b"1111111111111111_1111111111111111_1110001010011011_1011101110101010"; -- -0.11481120205881444
	pesos_i(12387) := b"1111111111111111_1111111111111111_1110000111001000_1100100001001111"; -- -0.11803005294586226
	pesos_i(12388) := b"0000000000000000_0000000000000000_0010000000111011_0101111101011010"; -- 0.12590595206285127
	pesos_i(12389) := b"1111111111111111_1111111111111111_1101011111110110_0110110111011000"; -- -0.15639604066773247
	pesos_i(12390) := b"0000000000000000_0000000000000000_0000101111111001_1111111010011010"; -- 0.04678336389097091
	pesos_i(12391) := b"1111111111111111_1111111111111111_1111011110110111_1101000100111100"; -- -0.03235142017589184
	pesos_i(12392) := b"0000000000000000_0000000000000000_0000100010010000_0100010010011101"; -- 0.03345135519604346
	pesos_i(12393) := b"1111111111111111_1111111111111111_1110000110111111_0011010111111010"; -- -0.11817610402439074
	pesos_i(12394) := b"1111111111111111_1111111111111111_1101111000100000_0100010101011100"; -- -0.13232008450716862
	pesos_i(12395) := b"1111111111111111_1111111111111111_1110011000100000_0110000101010001"; -- -0.101068418202141
	pesos_i(12396) := b"0000000000000000_0000000000000000_0000111001001001_0110011110010000"; -- 0.05580756450960852
	pesos_i(12397) := b"1111111111111111_1111111111111111_1101111001101101_0111011000110110"; -- -0.1311422459915711
	pesos_i(12398) := b"0000000000000000_0000000000000000_0000100011001100_1011011001011110"; -- 0.034373662840085424
	pesos_i(12399) := b"0000000000000000_0000000000000000_0010001101110001_1110100100111010"; -- 0.13845689463277377
	pesos_i(12400) := b"1111111111111111_1111111111111111_1111010110001000_0110110111101010"; -- -0.04088700336675945
	pesos_i(12401) := b"1111111111111111_1111111111111111_1110110010100100_0001111101000110"; -- -0.0756206946460708
	pesos_i(12402) := b"0000000000000000_0000000000000000_0000111100101010_0010001101000000"; -- 0.05923672024734029
	pesos_i(12403) := b"1111111111111111_1111111111111111_1111101100011110_0100111100101001"; -- -0.01906876803149228
	pesos_i(12404) := b"1111111111111111_1111111111111111_1111000101110101_0101011110000101"; -- -0.05680325514446225
	pesos_i(12405) := b"1111111111111111_1111111111111111_1111010111000110_1111111001001100"; -- -0.039932352470175236
	pesos_i(12406) := b"0000000000000000_0000000000000000_0001001111100110_1011111110110111"; -- 0.07773969850107156
	pesos_i(12407) := b"1111111111111111_1111111111111111_1110000100110000_0100100011101000"; -- -0.12035698262012831
	pesos_i(12408) := b"0000000000000000_0000000000000000_0000010000110101_0101101001011101"; -- 0.016439101919361
	pesos_i(12409) := b"1111111111111111_1111111111111111_1111110111010101_1001111000111000"; -- -0.008459197376261876
	pesos_i(12410) := b"0000000000000000_0000000000000000_0000000011011100_1011111011111010"; -- 0.003368316601156665
	pesos_i(12411) := b"1111111111111111_1111111111111111_1101101111111001_1101011001001101"; -- -0.1407190381328282
	pesos_i(12412) := b"0000000000000000_0000000000000000_0001000000110001_1000011010001111"; -- 0.06325570106113153
	pesos_i(12413) := b"1111111111111111_1111111111111111_1101111010110011_1001101100110001"; -- -0.13007192651719857
	pesos_i(12414) := b"1111111111111111_1111111111111111_1110000011010111_1010110101010010"; -- -0.1217090296537096
	pesos_i(12415) := b"0000000000000000_0000000000000000_0010010000110101_0110101011110001"; -- 0.14144009001317667
	pesos_i(12416) := b"1111111111111111_1111111111111111_1111110010101111_1100111101101111"; -- -0.012942348009828127
	pesos_i(12417) := b"0000000000000000_0000000000000000_0000101010110111_1001101001011111"; -- 0.041864059556045156
	pesos_i(12418) := b"0000000000000000_0000000000000000_0001100001000101_1101100010111000"; -- 0.0948157739096753
	pesos_i(12419) := b"1111111111111111_1111111111111111_1111011011001101_0110100000010011"; -- -0.03592824492450159
	pesos_i(12420) := b"1111111111111111_1111111111111111_1111101010011100_0101110110010010"; -- -0.02105155165643128
	pesos_i(12421) := b"0000000000000000_0000000000000000_0001001101101001_0000001111001100"; -- 0.0758211491684478
	pesos_i(12422) := b"1111111111111111_1111111111111111_1110101100011000_1010111001110000"; -- -0.08165464173110311
	pesos_i(12423) := b"1111111111111111_1111111111111111_1110111001101000_0011010110100110"; -- -0.06872238824897747
	pesos_i(12424) := b"1111111111111111_1111111111111111_1110110000111000_1001011000110110"; -- -0.07726155452128719
	pesos_i(12425) := b"1111111111111111_1111111111111111_1110010011010000_1011001000011110"; -- -0.10619055527359685
	pesos_i(12426) := b"0000000000000000_0000000000000000_0010000101000100_0011001100100000"; -- 0.1299468948786741
	pesos_i(12427) := b"0000000000000000_0000000000000000_0001111101111101_0011111000001001"; -- 0.12300479627891894
	pesos_i(12428) := b"0000000000000000_0000000000000000_0001001010100000_0110011101001001"; -- 0.0727600624788384
	pesos_i(12429) := b"0000000000000000_0000000000000000_0001110001000101_1010011100000001"; -- 0.11043781069245114
	pesos_i(12430) := b"1111111111111111_1111111111111111_1101110010010101_0000001100101001"; -- -0.13835125205994997
	pesos_i(12431) := b"0000000000000000_0000000000000000_0000100010111011_1011010101111010"; -- 0.034114210434209924
	pesos_i(12432) := b"1111111111111111_1111111111111111_1101110001001010_1101011101000001"; -- -0.13948301941635902
	pesos_i(12433) := b"0000000000000000_0000000000000000_0001101000110100_0001100110000011"; -- 0.10235747755814166
	pesos_i(12434) := b"0000000000000000_0000000000000000_0000000110101000_0001000010001110"; -- 0.006470713228330118
	pesos_i(12435) := b"1111111111111111_1111111111111111_1110000110010000_0100001010101101"; -- -0.11889251010588718
	pesos_i(12436) := b"0000000000000000_0000000000000000_0000010000100111_0111001011110010"; -- 0.016226944115737253
	pesos_i(12437) := b"0000000000000000_0000000000000000_0000010100011010_1001000101001000"; -- 0.01993663791931539
	pesos_i(12438) := b"0000000000000000_0000000000000000_0010100100010001_1010101011110010"; -- 0.16042583853847225
	pesos_i(12439) := b"0000000000000000_0000000000000000_0000010111110010_1110100110101110"; -- 0.023237805340791725
	pesos_i(12440) := b"1111111111111111_1111111111111111_1111000001001011_1111101011110011"; -- -0.06134063312348629
	pesos_i(12441) := b"1111111111111111_1111111111111111_1110011011101100_1110100001100010"; -- -0.09794757478297535
	pesos_i(12442) := b"1111111111111111_1111111111111111_1110010011111010_1001011010001101"; -- -0.10555132913308046
	pesos_i(12443) := b"1111111111111111_1111111111111111_1101101100110011_0111000001011000"; -- -0.1437463556491095
	pesos_i(12444) := b"0000000000000000_0000000000000000_0001110000000111_1101011001110101"; -- 0.10949459424904924
	pesos_i(12445) := b"0000000000000000_0000000000000000_0001011001011110_0010010100100001"; -- 0.08737403918459374
	pesos_i(12446) := b"0000000000000000_0000000000000000_0010001001100100_0111010010010011"; -- 0.13434532735691665
	pesos_i(12447) := b"0000000000000000_0000000000000000_0010100000001000_0110011010011110"; -- 0.15637818669263276
	pesos_i(12448) := b"1111111111111111_1111111111111111_1111101000100110_1110110110110001"; -- -0.022843498440031362
	pesos_i(12449) := b"0000000000000000_0000000000000000_0001110011011000_1010110101101101"; -- 0.1126812355034081
	pesos_i(12450) := b"1111111111111111_1111111111111111_1111100100110010_1100110111000101"; -- -0.02656854569417288
	pesos_i(12451) := b"0000000000000000_0000000000000000_0000010011011011_0001101010001110"; -- 0.018968257537566792
	pesos_i(12452) := b"0000000000000000_0000000000000000_0000110011011101_1010100110110000"; -- 0.05025730651437003
	pesos_i(12453) := b"0000000000000000_0000000000000000_0000111010000101_1101001010100010"; -- 0.05672947360075288
	pesos_i(12454) := b"1111111111111111_1111111111111111_1111101111011111_1010100100101111"; -- -0.016118455868902093
	pesos_i(12455) := b"0000000000000000_0000000000000000_0000101101101100_0000100101111111"; -- 0.044617265166880214
	pesos_i(12456) := b"0000000000000000_0000000000000000_0001100000111110_0011010100110000"; -- 0.09469921521147677
	pesos_i(12457) := b"0000000000000000_0000000000000000_0001100011101001_1001000000111010"; -- 0.09731389436959685
	pesos_i(12458) := b"0000000000000000_0000000000000000_0000011010110101_0011110110110011"; -- 0.026203018349746504
	pesos_i(12459) := b"1111111111111111_1111111111111111_1111110011100101_1101010000101010"; -- -0.012118091266388674
	pesos_i(12460) := b"0000000000000000_0000000000000000_0000011001000101_1101001101111001"; -- 0.02450296115550275
	pesos_i(12461) := b"1111111111111111_1111111111111111_1110100011110101_0010111110101011"; -- -0.09000875544121419
	pesos_i(12462) := b"0000000000000000_0000000000000000_0001111001100001_1001011001100001"; -- 0.11867656591137801
	pesos_i(12463) := b"0000000000000000_0000000000000000_0010010111000010_0101110001100000"; -- 0.14749696098783796
	pesos_i(12464) := b"0000000000000000_0000000000000000_0000110101011000_1011011010000110"; -- 0.052134902674221884
	pesos_i(12465) := b"1111111111111111_1111111111111111_1101111000011100_1101001101100101"; -- -0.1323726536975901
	pesos_i(12466) := b"0000000000000000_0000000000000000_0001100110010000_0111111111100101"; -- 0.09986113871396876
	pesos_i(12467) := b"1111111111111111_1111111111111111_1110100111010000_0011110110010100"; -- -0.08666625160071043
	pesos_i(12468) := b"1111111111111111_1111111111111111_1111111111001110_1001010000100010"; -- -0.0007541099777478891
	pesos_i(12469) := b"0000000000000000_0000000000000000_0001000001000101_0010101110010001"; -- 0.06355545316821713
	pesos_i(12470) := b"0000000000000000_0000000000000000_0000111110111110_0111101011010100"; -- 0.06150024107213145
	pesos_i(12471) := b"1111111111111111_1111111111111111_1111010110100001_0110101110110101"; -- -0.040505665130106824
	pesos_i(12472) := b"1111111111111111_1111111111111111_1110000011100101_1101000111011000"; -- -0.12149322962071482
	pesos_i(12473) := b"0000000000000000_0000000000000000_0000011010100010_0111000101101010"; -- 0.025916183809126928
	pesos_i(12474) := b"0000000000000000_0000000000000000_0001000110010101_1010101011110001"; -- 0.06868999838693299
	pesos_i(12475) := b"1111111111111111_1111111111111111_1111111101111111_1111011100000010"; -- -0.0019536609662388097
	pesos_i(12476) := b"0000000000000000_0000000000000000_0000010101111100_1110100100010111"; -- 0.021437233092336284
	pesos_i(12477) := b"0000000000000000_0000000000000000_0000111101001010_0100010111111100"; -- 0.05972707183094766
	pesos_i(12478) := b"1111111111111111_1111111111111111_1111001111001000_1110111011010100"; -- -0.0477152569516644
	pesos_i(12479) := b"1111111111111111_1111111111111111_1110111111001101_1111000011001011"; -- -0.0632638457523866
	pesos_i(12480) := b"0000000000000000_0000000000000000_0000100000011100_0101110011110011"; -- 0.03168278622731897
	pesos_i(12481) := b"0000000000000000_0000000000000000_0001011011011011_0110000101100111"; -- 0.08928498054242653
	pesos_i(12482) := b"0000000000000000_0000000000000000_0010000110011010_1000100010000101"; -- 0.1312642407770611
	pesos_i(12483) := b"0000000000000000_0000000000000000_0000101101010011_1010101101111000"; -- 0.04424544991138849
	pesos_i(12484) := b"0000000000000000_0000000000000000_0001100110000101_0011111101011110"; -- 0.09968944602949673
	pesos_i(12485) := b"0000000000000000_0000000000000000_0010001011000111_1000011111001100"; -- 0.13585709306393176
	pesos_i(12486) := b"1111111111111111_1111111111111111_1101111000110010_1011011010100000"; -- -0.13203867533059635
	pesos_i(12487) := b"1111111111111111_1111111111111111_1101110111100001_0001000011111100"; -- -0.13328451009891748
	pesos_i(12488) := b"0000000000000000_0000000000000000_0001011001100101_0101100101101110"; -- 0.08748396819510022
	pesos_i(12489) := b"1111111111111111_1111111111111111_1111100011000010_0111110010000111"; -- -0.028282372422591046
	pesos_i(12490) := b"0000000000000000_0000000000000000_0000101001100111_0100001010111000"; -- 0.04063813203329125
	pesos_i(12491) := b"1111111111111111_1111111111111111_1110010101010110_1110111000000000"; -- -0.10414230825563052
	pesos_i(12492) := b"1111111111111111_1111111111111111_1101100001100100_1011010010111010"; -- -0.15471334889321203
	pesos_i(12493) := b"0000000000000000_0000000000000000_0001100000011111_1110110101001100"; -- 0.09423716648887186
	pesos_i(12494) := b"0000000000000000_0000000000000000_0000010000111011_1111111011001110"; -- 0.016540455982633494
	pesos_i(12495) := b"0000000000000000_0000000000000000_0001010001001100_0101010100101010"; -- 0.07928974410976698
	pesos_i(12496) := b"0000000000000000_0000000000000000_0000000101010111_1010100000110100"; -- 0.0052437904093943204
	pesos_i(12497) := b"0000000000000000_0000000000000000_0001100101001010_0111011010000011"; -- 0.09879246430022551
	pesos_i(12498) := b"1111111111111111_1111111111111111_1110110101100100_1111111111101010"; -- -0.07267761750447099
	pesos_i(12499) := b"0000000000000000_0000000000000000_0010001000011000_0001000111011100"; -- 0.13317977548283252
	pesos_i(12500) := b"1111111111111111_1111111111111111_1110001101101101_1110011101100111"; -- -0.1116042492512241
	pesos_i(12501) := b"0000000000000000_0000000000000000_0000011101000011_1000000110101001"; -- 0.02837381716823244
	pesos_i(12502) := b"0000000000000000_0000000000000000_0001111010111011_0001011000011110"; -- 0.12004221184708208
	pesos_i(12503) := b"1111111111111111_1111111111111111_1110110011111001_1100000010011100"; -- -0.07431408109071294
	pesos_i(12504) := b"1111111111111111_1111111111111111_1111001110100000_0011011000001001"; -- -0.04833662293365181
	pesos_i(12505) := b"0000000000000000_0000000000000000_0001011111001010_1100110001101111"; -- 0.09293821058620973
	pesos_i(12506) := b"0000000000000000_0000000000000000_0010101001011100_0000011101001101"; -- 0.16546674371795586
	pesos_i(12507) := b"1111111111111111_1111111111111111_1111100011111011_0111000000100110"; -- -0.027413359361291127
	pesos_i(12508) := b"1111111111111111_1111111111111111_1110010000111101_1100110001010111"; -- -0.10843203421252226
	pesos_i(12509) := b"1111111111111111_1111111111111111_1110000100010000_1001001111110011"; -- -0.12084079098811515
	pesos_i(12510) := b"1111111111111111_1111111111111111_1111110110010100_1001100111010111"; -- -0.009451279606098584
	pesos_i(12511) := b"1111111111111111_1111111111111111_1110000000100110_0110000000110100"; -- -0.1244144318745196
	pesos_i(12512) := b"1111111111111111_1111111111111111_1111011110001000_1111011101001110"; -- -0.03306631410565761
	pesos_i(12513) := b"1111111111111111_1111111111111111_1110101000011111_0010100100001111"; -- -0.08546203015721048
	pesos_i(12514) := b"1111111111111111_1111111111111111_1101100110011100_1000110011011010"; -- -0.14995498356804138
	pesos_i(12515) := b"0000000000000000_0000000000000000_0001010100111110_0001101111000010"; -- 0.08297894950063359
	pesos_i(12516) := b"1111111111111111_1111111111111111_1111110000010111_1101010001110100"; -- -0.01526138477052349
	pesos_i(12517) := b"0000000000000000_0000000000000000_0010001100110011_0011111111010110"; -- 0.1375007530690125
	pesos_i(12518) := b"0000000000000000_0000000000000000_0001011110011000_0111011000000011"; -- 0.09217012007115721
	pesos_i(12519) := b"1111111111111111_1111111111111111_1111101001001101_0111100010101111"; -- -0.022255379920609376
	pesos_i(12520) := b"1111111111111111_1111111111111111_1111100001100111_1010101111111101"; -- -0.029668093386226706
	pesos_i(12521) := b"0000000000000000_0000000000000000_0000111000101101_1010000011010101"; -- 0.0553837317618668
	pesos_i(12522) := b"1111111111111111_1111111111111111_1110100101101111_0100111001101010"; -- -0.08814535065451855
	pesos_i(12523) := b"1111111111111111_1111111111111111_1101110010101010_1101110010010000"; -- -0.13801785920450316
	pesos_i(12524) := b"0000000000000000_0000000000000000_0000010010100001_0101110001110001"; -- 0.018087175025694773
	pesos_i(12525) := b"1111111111111111_1111111111111111_1111100101101000_1010011101000111"; -- -0.02574686546241374
	pesos_i(12526) := b"1111111111111111_1111111111111111_1111111101100001_1000000110111000"; -- -0.002418415644978003
	pesos_i(12527) := b"0000000000000000_0000000000000000_0001001111101000_1111000111001111"; -- 0.07777320203145892
	pesos_i(12528) := b"1111111111111111_1111111111111111_1110100000100100_0111001010100101"; -- -0.09319385019864855
	pesos_i(12529) := b"0000000000000000_0000000000000000_0010011001010100_1001001110111100"; -- 0.14972804387728142
	pesos_i(12530) := b"0000000000000000_0000000000000000_0000111110001000_0000111001001000"; -- 0.0606697964504957
	pesos_i(12531) := b"1111111111111111_1111111111111111_1101111010100101_1100011010011100"; -- -0.13028296179997448
	pesos_i(12532) := b"0000000000000000_0000000000000000_0001111100011100_1100101100001011"; -- 0.12153309843948705
	pesos_i(12533) := b"1111111111111111_1111111111111111_1110000011101111_0001110011111100"; -- -0.12135142182538101
	pesos_i(12534) := b"0000000000000000_0000000000000000_0010000110011111_1000001101000000"; -- 0.131340220468213
	pesos_i(12535) := b"1111111111111111_1111111111111111_1110110010001100_0010000111010010"; -- -0.07598675370823739
	pesos_i(12536) := b"0000000000000000_0000000000000000_0001100101000010_1011110100110101"; -- 0.09867460763258654
	pesos_i(12537) := b"0000000000000000_0000000000000000_0001111010001100_0101111111010111"; -- 0.11932944303288935
	pesos_i(12538) := b"0000000000000000_0000000000000000_0001110110101110_0000100111100110"; -- 0.11593686921355145
	pesos_i(12539) := b"1111111111111111_1111111111111111_1110011000111110_0111110011110001"; -- -0.10060900809399585
	pesos_i(12540) := b"1111111111111111_1111111111111111_1111111010110111_0011011011110001"; -- -0.005016866913966831
	pesos_i(12541) := b"0000000000000000_0000000000000000_0001101100111101_0111100011001101"; -- 0.10640673645085408
	pesos_i(12542) := b"0000000000000000_0000000000000000_0001100110111010_1111011010011011"; -- 0.1005090835886639
	pesos_i(12543) := b"1111111111111111_1111111111111111_1110011011111110_0001111111010010"; -- -0.09768487085875834
	pesos_i(12544) := b"1111111111111111_1111111111111111_1111101000001111_0011010111101011"; -- -0.02320540431829377
	pesos_i(12545) := b"1111111111111111_1111111111111111_1101101101001101_1010000111100101"; -- -0.14334667359356465
	pesos_i(12546) := b"1111111111111111_1111111111111111_1110111110110011_1011100111110000"; -- -0.06366384392596115
	pesos_i(12547) := b"0000000000000000_0000000000000000_0000001110110110_0000100010000101"; -- 0.014496357505202557
	pesos_i(12548) := b"1111111111111111_1111111111111111_1110010000101101_1001110001110001"; -- -0.1086790298026676
	pesos_i(12549) := b"1111111111111111_1111111111111111_1111010100001011_1000110100000101"; -- -0.04279249790757689
	pesos_i(12550) := b"0000000000000000_0000000000000000_0010001011100010_0111000000000011"; -- 0.13626766276552588
	pesos_i(12551) := b"1111111111111111_1111111111111111_1101011010000111_1110100110010001"; -- -0.1619886417508685
	pesos_i(12552) := b"1111111111111111_1111111111111111_1111111110010110_0011000001111010"; -- -0.0016145421566520842
	pesos_i(12553) := b"1111111111111111_1111111111111111_1111000110010011_1100111100011100"; -- -0.05633836335646465
	pesos_i(12554) := b"0000000000000000_0000000000000000_0000000110110101_0000010011011101"; -- 0.006668380618680299
	pesos_i(12555) := b"0000000000000000_0000000000000000_0001100001010101_0101011100000111"; -- 0.09505218432055644
	pesos_i(12556) := b"0000000000000000_0000000000000000_0000111010101001_0000101111100001"; -- 0.05726694344293257
	pesos_i(12557) := b"1111111111111111_1111111111111111_1111000101110001_1010101111101100"; -- -0.056859259525149836
	pesos_i(12558) := b"0000000000000000_0000000000000000_0000011001110100_0001001011001100"; -- 0.025208639890725727
	pesos_i(12559) := b"0000000000000000_0000000000000000_0010001001011010_0111011001100001"; -- 0.13419284684881333
	pesos_i(12560) := b"0000000000000000_0000000000000000_0000110101111101_0101110000111101"; -- 0.05269409657829148
	pesos_i(12561) := b"0000000000000000_0000000000000000_0010010000011011_0010011000110111"; -- 0.14103926503989783
	pesos_i(12562) := b"0000000000000000_0000000000000000_0000000111101010_0110110000011001"; -- 0.007483249808951569
	pesos_i(12563) := b"1111111111111111_1111111111111111_1110001101000001_1011101000111110"; -- -0.11227832783770647
	pesos_i(12564) := b"1111111111111111_1111111111111111_1111010111110110_0110001001101010"; -- -0.039209221963590654
	pesos_i(12565) := b"1111111111111111_1111111111111111_1110100101000000_1011110111010001"; -- -0.08885587355295291
	pesos_i(12566) := b"1111111111111111_1111111111111111_1110011011001101_0101000110110011"; -- -0.09842957858766423
	pesos_i(12567) := b"0000000000000000_0000000000000000_0000101001110000_1101000111100011"; -- 0.04078399467012734
	pesos_i(12568) := b"0000000000000000_0000000000000000_0001001011110000_1001001110011010"; -- 0.07398340715824123
	pesos_i(12569) := b"0000000000000000_0000000000000000_0001000111111111_1000101000101000"; -- 0.0703054759906954
	pesos_i(12570) := b"1111111111111111_1111111111111111_1111011010100001_1101111011100000"; -- -0.036592550669343894
	pesos_i(12571) := b"0000000000000000_0000000000000000_0001010111100011_0010000010111101"; -- 0.08549694656109709
	pesos_i(12572) := b"0000000000000000_0000000000000000_0010000110000110_1110110001110101"; -- 0.1309650216738665
	pesos_i(12573) := b"0000000000000000_0000000000000000_0000101001001101_0001100000111111"; -- 0.040238871842769336
	pesos_i(12574) := b"0000000000000000_0000000000000000_0000101000000001_0000100100100000"; -- 0.039078302724256254
	pesos_i(12575) := b"0000000000000000_0000000000000000_0010000101110000_0110010100010111"; -- 0.130621259718358
	pesos_i(12576) := b"1111111111111111_1111111111111111_1110010110110100_0000010000011111"; -- -0.10272192236069959
	pesos_i(12577) := b"0000000000000000_0000000000000000_0001110110000100_1101111000101010"; -- 0.11530865210787627
	pesos_i(12578) := b"0000000000000000_0000000000000000_0000101001011001_1101111010011001"; -- 0.04043380003266253
	pesos_i(12579) := b"0000000000000000_0000000000000000_0001100111011111_0000000110000101"; -- 0.10105905058694198
	pesos_i(12580) := b"0000000000000000_0000000000000000_0001100100011001_1111011100101110"; -- 0.09805245289476848
	pesos_i(12581) := b"0000000000000000_0000000000000000_0001101100100001_1000010000101101"; -- 0.10598016843842396
	pesos_i(12582) := b"0000000000000000_0000000000000000_0001010011000011_0011010001101101"; -- 0.08110358868600759
	pesos_i(12583) := b"0000000000000000_0000000000000000_0001111101011111_0010010100011111"; -- 0.12254554755929209
	pesos_i(12584) := b"1111111111111111_1111111111111111_1111100111011110_0101001010010110"; -- -0.023951376350274965
	pesos_i(12585) := b"0000000000000000_0000000000000000_0001110111001011_0110101100001011"; -- 0.11638516446697553
	pesos_i(12586) := b"1111111111111111_1111111111111111_1110000000000001_0110110100010101"; -- -0.12497823933168747
	pesos_i(12587) := b"0000000000000000_0000000000000000_0000101001101111_1111010001001000"; -- 0.040770785998901715
	pesos_i(12588) := b"1111111111111111_1111111111111111_1111000010011110_0011001100001001"; -- -0.06008606936473504
	pesos_i(12589) := b"1111111111111111_1111111111111111_1111110100000000_0100000010100000"; -- -0.011714897985427953
	pesos_i(12590) := b"1111111111111111_1111111111111111_1110010111010111_0001110100011010"; -- -0.10218637575104617
	pesos_i(12591) := b"0000000000000000_0000000000000000_0000101010111110_1111101111110001"; -- 0.041976686877636414
	pesos_i(12592) := b"0000000000000000_0000000000000000_0010001110010001_0110110011000101"; -- 0.13893775748275905
	pesos_i(12593) := b"1111111111111111_1111111111111111_1110110110011011_0000010101000101"; -- -0.07185332367977713
	pesos_i(12594) := b"1111111111111111_1111111111111111_1111111111110100_0110000000100001"; -- -0.00017737578330123747
	pesos_i(12595) := b"1111111111111111_1111111111111111_1111010010001100_1010100000100101"; -- -0.044728747437566475
	pesos_i(12596) := b"0000000000000000_0000000000000000_0001011110001010_0011011111010000"; -- 0.09195278961340857
	pesos_i(12597) := b"1111111111111111_1111111111111111_1110010010000110_0010100010001000"; -- -0.10732790647587492
	pesos_i(12598) := b"0000000000000000_0000000000000000_0000110010100101_0000000011101110"; -- 0.04939275558934903
	pesos_i(12599) := b"1111111111111111_1111111111111111_1110110110001110_1000011111101001"; -- -0.072043901070341
	pesos_i(12600) := b"1111111111111111_1111111111111111_1111101110111111_0000001011010100"; -- -0.016616652833583247
	pesos_i(12601) := b"1111111111111111_1111111111111111_1111000101100011_1111110011111001"; -- -0.057068051553394616
	pesos_i(12602) := b"1111111111111111_1111111111111111_1111101101011001_0110100000111010"; -- -0.018167005496233235
	pesos_i(12603) := b"0000000000000000_0000000000000000_0010001000011010_0110100010110011"; -- 0.1332154690053867
	pesos_i(12604) := b"0000000000000000_0000000000000000_0001001001100010_1101100100101111"; -- 0.07182080643815841
	pesos_i(12605) := b"0000000000000000_0000000000000000_0010010001011001_0011011110001001"; -- 0.14198634234724142
	pesos_i(12606) := b"0000000000000000_0000000000000000_0001101000111101_1011111101010010"; -- 0.1025046896386655
	pesos_i(12607) := b"1111111111111111_1111111111111111_1101110001010010_1001010011010001"; -- -0.1393649092215843
	pesos_i(12608) := b"0000000000000000_0000000000000000_0010000011111100_0010100011001110"; -- 0.12884764707128007
	pesos_i(12609) := b"0000000000000000_0000000000000000_0000100011010100_0101001100111010"; -- 0.03448982408534045
	pesos_i(12610) := b"1111111111111111_1111111111111111_1110111110110111_0101011101101011"; -- -0.06360868112989697
	pesos_i(12611) := b"1111111111111111_1111111111111111_1101101101010000_1100001111001011"; -- -0.1432988766813199
	pesos_i(12612) := b"0000000000000000_0000000000000000_0010001111010110_0001001011100011"; -- 0.13998525668093878
	pesos_i(12613) := b"1111111111111111_1111111111111111_1101110100001111_1110101011000110"; -- -0.1364758746742203
	pesos_i(12614) := b"0000000000000000_0000000000000000_0001101111101000_1000000001000001"; -- 0.10901643366501677
	pesos_i(12615) := b"0000000000000000_0000000000000000_0010001001100010_1011110101001011"; -- 0.13431914403404296
	pesos_i(12616) := b"0000000000000000_0000000000000000_0001101110001101_1010011000100010"; -- 0.10763014153654325
	pesos_i(12617) := b"1111111111111111_1111111111111111_1110001111111011_1101110101111111"; -- -0.10943809165888058
	pesos_i(12618) := b"1111111111111111_1111111111111111_1110000111001001_1000110010100101"; -- -0.11801835022164264
	pesos_i(12619) := b"0000000000000000_0000000000000000_0001010010110000_0010110010101000"; -- 0.08081320857171947
	pesos_i(12620) := b"0000000000000000_0000000000000000_0010001001010101_1110111011011000"; -- 0.13412373328797128
	pesos_i(12621) := b"0000000000000000_0000000000000000_0001000011010011_1000001011111111"; -- 0.0657274124968351
	pesos_i(12622) := b"1111111111111111_1111111111111111_1110101000110110_0001101010011011"; -- -0.08511193961994913
	pesos_i(12623) := b"1111111111111111_1111111111111111_1101101100010111_0111000000011101"; -- -0.14417361547464055
	pesos_i(12624) := b"0000000000000000_0000000000000000_0000000001110010_1111011010011110"; -- 0.0017542014569440442
	pesos_i(12625) := b"1111111111111111_1111111111111111_1111110011100000_0000010111101001"; -- -0.012206678921055914
	pesos_i(12626) := b"1111111111111111_1111111111111111_1110110000001100_1010100101100011"; -- -0.07793179833423064
	pesos_i(12627) := b"1111111111111111_1111111111111111_1101011000010011_0001011101011110"; -- -0.16377119016191483
	pesos_i(12628) := b"0000000000000000_0000000000000000_0001011111010010_0101111111111110"; -- 0.09305381734137738
	pesos_i(12629) := b"1111111111111111_1111111111111111_1110100110001110_0111001111011100"; -- -0.08767009618098763
	pesos_i(12630) := b"1111111111111111_1111111111111111_1111100101100011_1101000010001101"; -- -0.02582069922174418
	pesos_i(12631) := b"0000000000000000_0000000000000000_0001111010101110_0101011110011001"; -- 0.11984775044931935
	pesos_i(12632) := b"1111111111111111_1111111111111111_1110010011001011_0111000100000111"; -- -0.1062707288611069
	pesos_i(12633) := b"1111111111111111_1111111111111111_1101111110001100_0101100001100111"; -- -0.12676475041523722
	pesos_i(12634) := b"1111111111111111_1111111111111111_1110110001101111_0001000110100100"; -- -0.07643022304832521
	pesos_i(12635) := b"0000000000000000_0000000000000000_0010000001100001_0101100111101110"; -- 0.12648546277892733
	pesos_i(12636) := b"0000000000000000_0000000000000000_0000111010011010_1001111000010011"; -- 0.057046775427732205
	pesos_i(12637) := b"0000000000000000_0000000000000000_0001110110011011_1000001111110111"; -- 0.11565422791633884
	pesos_i(12638) := b"1111111111111111_1111111111111111_1101101110011011_0000110011010000"; -- -0.14216537394732504
	pesos_i(12639) := b"1111111111111111_1111111111111111_1101101110100001_1000111010011011"; -- -0.14206608499281628
	pesos_i(12640) := b"0000000000000000_0000000000000000_0001001111101001_0111100101101001"; -- 0.07778128455224735
	pesos_i(12641) := b"1111111111111111_1111111111111111_1110010110111001_1010110001000101"; -- -0.10263560595842547
	pesos_i(12642) := b"1111111111111111_1111111111111111_1111010111000111_1000011110000000"; -- -0.039924174636588254
	pesos_i(12643) := b"0000000000000000_0000000000000000_0001011010110011_1010010001010000"; -- 0.08867861704688162
	pesos_i(12644) := b"0000000000000000_0000000000000000_0000001001100110_0111011111101000"; -- 0.00937604352974242
	pesos_i(12645) := b"1111111111111111_1111111111111111_1110010100111101_0111111010101001"; -- -0.10453041436557639
	pesos_i(12646) := b"1111111111111111_1111111111111111_1101110011100000_0111001000011000"; -- -0.13720023065223477
	pesos_i(12647) := b"0000000000000000_0000000000000000_0001000000110100_0010010110010101"; -- 0.06329569714283341
	pesos_i(12648) := b"0000000000000000_0000000000000000_0001011100010110_0100011010111000"; -- 0.09018365847896556
	pesos_i(12649) := b"1111111111111111_1111111111111111_1110010100000011_0010110000000100"; -- -0.10542035019646054
	pesos_i(12650) := b"1111111111111111_1111111111111111_1111001010010001_1010110010100010"; -- -0.05246468594941612
	pesos_i(12651) := b"1111111111111111_1111111111111111_1110011101100010_0010111100000101"; -- -0.09615808598928728
	pesos_i(12652) := b"0000000000000000_0000000000000000_0000110100110001_1110000001101010"; -- 0.051542306681155066
	pesos_i(12653) := b"1111111111111111_1111111111111111_1110100010110111_1110010100110101"; -- -0.09094397979458832
	pesos_i(12654) := b"0000000000000000_0000000000000000_0001110010011101_1111101011110110"; -- 0.11178558829788422
	pesos_i(12655) := b"0000000000000000_0000000000000000_0010010011101011_1100100101001011"; -- 0.14422281332362755
	pesos_i(12656) := b"0000000000000000_0000000000000000_0000001010110101_0000110101000110"; -- 0.010575131944635519
	pesos_i(12657) := b"1111111111111111_1111111111111111_1111111110111000_1011100110010011"; -- -0.0010875716773944735
	pesos_i(12658) := b"0000000000000000_0000000000000000_0001011110001101_1101011101010011"; -- 0.09200807347514221
	pesos_i(12659) := b"0000000000000000_0000000000000000_0000110011110111_1110110000101110"; -- 0.05065799839585174
	pesos_i(12660) := b"1111111111111111_1111111111111111_1111101010001001_1010011010001111"; -- -0.021337118237166858
	pesos_i(12661) := b"0000000000000000_0000000000000000_0000001110011101_1010000010000100"; -- 0.01412394729688834
	pesos_i(12662) := b"0000000000000000_0000000000000000_0000000000111101_0111111110101100"; -- 0.0009383958627992965
	pesos_i(12663) := b"1111111111111111_1111111111111111_1111100110101111_1100000011011101"; -- -0.024661966312748414
	pesos_i(12664) := b"0000000000000000_0000000000000000_0000011011110011_1000011011001100"; -- 0.027153420373497418
	pesos_i(12665) := b"0000000000000000_0000000000000000_0000110010110101_0111110101000001"; -- 0.0496443065704559
	pesos_i(12666) := b"0000000000000000_0000000000000000_0001100001000011_1001001001100000"; -- 0.09478106342612291
	pesos_i(12667) := b"0000000000000000_0000000000000000_0000100001000001_0011010110100000"; -- 0.032245017585233425
	pesos_i(12668) := b"1111111111111111_1111111111111111_1101110000000001_0010010001111001"; -- -0.1406075672356876
	pesos_i(12669) := b"1111111111111111_1111111111111111_1111010010011000_1010010111010100"; -- -0.04454578001984279
	pesos_i(12670) := b"0000000000000000_0000000000000000_0001011100000101_0000100100010110"; -- 0.08992058549785155
	pesos_i(12671) := b"0000000000000000_0000000000000000_0000101111101101_0111111010111110"; -- 0.0465926374738946
	pesos_i(12672) := b"0000000000000000_0000000000000000_0000001101011111_1100010011110111"; -- 0.013180074919168724
	pesos_i(12673) := b"1111111111111111_1111111111111111_1111100010101011_1110111110001110"; -- -0.02862646847682629
	pesos_i(12674) := b"0000000000000000_0000000000000000_0001111101101011_1010010010000111"; -- 0.12273624709816147
	pesos_i(12675) := b"0000000000000000_0000000000000000_0010011010011111_1000111111000011"; -- 0.15087221631460015
	pesos_i(12676) := b"1111111111111111_1111111111111111_1110000000001111_1011111111101011"; -- -0.12475967889001302
	pesos_i(12677) := b"0000000000000000_0000000000000000_0001111111111100_0001110010000011"; -- 0.1249406642338725
	pesos_i(12678) := b"0000000000000000_0000000000000000_0001101010111010_0101011101110000"; -- 0.10440584648853006
	pesos_i(12679) := b"0000000000000000_0000000000000000_0001001010011001_0111001101010010"; -- 0.07265396841309693
	pesos_i(12680) := b"1111111111111111_1111111111111111_1111011001100111_0110110010011011"; -- -0.03748437133826553
	pesos_i(12681) := b"1111111111111111_1111111111111111_1110100011011101_1100100010101111"; -- -0.090365845830324
	pesos_i(12682) := b"1111111111111111_1111111111111111_1110100000101110_0010000110100101"; -- -0.09304609044171243
	pesos_i(12683) := b"1111111111111111_1111111111111111_1111001000100010_1111010010110001"; -- -0.05415411631895374
	pesos_i(12684) := b"1111111111111111_1111111111111111_1101110111000001_1100101110010011"; -- -0.13376166979314205
	pesos_i(12685) := b"0000000000000000_0000000000000000_0010010000110000_1010001001111101"; -- 0.14136710687849274
	pesos_i(12686) := b"1111111111111111_1111111111111111_1111100110011001_0010110101011110"; -- -0.025006451191232956
	pesos_i(12687) := b"1111111111111111_1111111111111111_1110110001100110_1111010110100010"; -- -0.07655396273422477
	pesos_i(12688) := b"0000000000000000_0000000000000000_0001100011010101_1001010101001101"; -- 0.09700902109960652
	pesos_i(12689) := b"1111111111111111_1111111111111111_1101111100101100_0110011010110001"; -- -0.12822874235073223
	pesos_i(12690) := b"0000000000000000_0000000000000000_0000010010110001_1110011110101011"; -- 0.018339614074317286
	pesos_i(12691) := b"1111111111111111_1111111111111111_1110110011111100_1011110110111010"; -- -0.07426847652276151
	pesos_i(12692) := b"0000000000000000_0000000000000000_0010011011011001_0100011111000001"; -- 0.1517529340754581
	pesos_i(12693) := b"0000000000000000_0000000000000000_0000110111011010_0110011011111100"; -- 0.054113804460906585
	pesos_i(12694) := b"1111111111111111_1111111111111111_1110011011001111_1000101100001110"; -- -0.0983956423644355
	pesos_i(12695) := b"1111111111111111_1111111111111111_1110010100101000_0100100010100100"; -- -0.10485406873896873
	pesos_i(12696) := b"1111111111111111_1111111111111111_1111010110101000_0100101001111101"; -- -0.04040083362129181
	pesos_i(12697) := b"1111111111111111_1111111111111111_1110000111011101_1111010001011100"; -- -0.11770699256438666
	pesos_i(12698) := b"0000000000000000_0000000000000000_0001001111101000_0011011000101011"; -- 0.07776201779369371
	pesos_i(12699) := b"0000000000000000_0000000000000000_0000010000001011_0010010110000100"; -- 0.01579508279531018
	pesos_i(12700) := b"1111111111111111_1111111111111111_1111111110101010_1100010011000010"; -- -0.0013005281995129955
	pesos_i(12701) := b"1111111111111111_1111111111111111_1110011010111100_1100111110111101"; -- -0.09868146543924622
	pesos_i(12702) := b"0000000000000000_0000000000000000_0001101111000101_1011010100011000"; -- 0.1084855254669966
	pesos_i(12703) := b"0000000000000000_0000000000000000_0010001011001000_1111110001011010"; -- 0.13587929902275478
	pesos_i(12704) := b"1111111111111111_1111111111111111_1110101110100001_0001101100111111"; -- -0.07957296105844075
	pesos_i(12705) := b"0000000000000000_0000000000000000_0000111011011101_1100101000111100"; -- 0.05807174652470992
	pesos_i(12706) := b"1111111111111111_1111111111111111_1111111100011111_1010011011001110"; -- -0.0034232850966604907
	pesos_i(12707) := b"0000000000000000_0000000000000000_0000110001111000_1111100101011110"; -- 0.04872091821865734
	pesos_i(12708) := b"0000000000000000_0000000000000000_0001100100011101_0000100100010010"; -- 0.09809929554710721
	pesos_i(12709) := b"0000000000000000_0000000000000000_0010011000001011_0110110000110110"; -- 0.14861179650917788
	pesos_i(12710) := b"0000000000000000_0000000000000000_0000110100011100_0110101001011100"; -- 0.05121483555154138
	pesos_i(12711) := b"0000000000000000_0000000000000000_0001011011000000_0010000011101111"; -- 0.08886915043317886
	pesos_i(12712) := b"0000000000000000_0000000000000000_0001000010010010_0110101100100000"; -- 0.06473416840853106
	pesos_i(12713) := b"0000000000000000_0000000000000000_0001001110110111_1001100101100110"; -- 0.07702025167020916
	pesos_i(12714) := b"1111111111111111_1111111111111111_1101111100110010_0100001011101111"; -- -0.1281393209958112
	pesos_i(12715) := b"1111111111111111_1111111111111111_1111010010010011_1000010111101100"; -- -0.044623975618308664
	pesos_i(12716) := b"1111111111111111_1111111111111111_1111010100010111_1001001001110000"; -- -0.04260906960624017
	pesos_i(12717) := b"1111111111111111_1111111111111111_1111101101011101_1001010111010011"; -- -0.018103252479056045
	pesos_i(12718) := b"1111111111111111_1111111111111111_1110100001011001_1100101100001010"; -- -0.09237986574450169
	pesos_i(12719) := b"0000000000000000_0000000000000000_0001001000100110_1111011011010100"; -- 0.07090704608140809
	pesos_i(12720) := b"1111111111111111_1111111111111111_1111001101111101_1011000101000001"; -- -0.04886333624228844
	pesos_i(12721) := b"1111111111111111_1111111111111111_1111001011110110_0001000111001010"; -- -0.0509327776908257
	pesos_i(12722) := b"1111111111111111_1111111111111111_1111010001110101_0000000011110010"; -- -0.04508966525332235
	pesos_i(12723) := b"0000000000000000_0000000000000000_0000100000110100_1001000001010000"; -- 0.032052058771447685
	pesos_i(12724) := b"0000000000000000_0000000000000000_0000000110100100_0010001110000110"; -- 0.006410808819216164
	pesos_i(12725) := b"0000000000000000_0000000000000000_0000100000000011_0101110110000001"; -- 0.0313013496246988
	pesos_i(12726) := b"0000000000000000_0000000000000000_0001111011100101_1011111001100101"; -- 0.1206931111062862
	pesos_i(12727) := b"0000000000000000_0000000000000000_0000001010010110_0001001010001111"; -- 0.010102424453348276
	pesos_i(12728) := b"0000000000000000_0000000000000000_0001001100000001_0101011000100001"; -- 0.07423914251006243
	pesos_i(12729) := b"1111111111111111_1111111111111111_1110110010001110_0111101011000011"; -- -0.07595093469208423
	pesos_i(12730) := b"1111111111111111_1111111111111111_1111110100110111_1100110101101000"; -- -0.010867273324807782
	pesos_i(12731) := b"1111111111111111_1111111111111111_1110110010110110_1110110111101111"; -- -0.07533371853152304
	pesos_i(12732) := b"1111111111111111_1111111111111111_1110010100101111_1111010001101000"; -- -0.10473701914902663
	pesos_i(12733) := b"1111111111111111_1111111111111111_1110001101100100_1100010000000101"; -- -0.11174368741647352
	pesos_i(12734) := b"1111111111111111_1111111111111111_1111110110111001_1111110111101010"; -- -0.008880739471175696
	pesos_i(12735) := b"1111111111111111_1111111111111111_1110100100011001_1110100100101001"; -- -0.08944838282355909
	pesos_i(12736) := b"1111111111111111_1111111111111111_1110010010100000_0101000000000000"; -- -0.10692882536229592
	pesos_i(12737) := b"1111111111111111_1111111111111111_1111100000110000_1101110111101100"; -- -0.030504350469514392
	pesos_i(12738) := b"1111111111111111_1111111111111111_1111110010010101_0101000111001001"; -- -0.013346565760163142
	pesos_i(12739) := b"0000000000000000_0000000000000000_0001110011011111_0100010111100011"; -- 0.11278187554209892
	pesos_i(12740) := b"1111111111111111_1111111111111111_1110110000100011_0001001001000110"; -- -0.07758985316504337
	pesos_i(12741) := b"0000000000000000_0000000000000000_0010001001011101_0000101000111101"; -- 0.13423217752549937
	pesos_i(12742) := b"1111111111111111_1111111111111111_1101101110101100_0110110101011011"; -- -0.14190022021108384
	pesos_i(12743) := b"1111111111111111_1111111111111111_1101100011000010_0011000010110100"; -- -0.15328689209753796
	pesos_i(12744) := b"1111111111111111_1111111111111111_1111001001011110_0111101100100111"; -- -0.05324583329698225
	pesos_i(12745) := b"1111111111111111_1111111111111111_1110110011011010_1000001000000001"; -- -0.07479083518305217
	pesos_i(12746) := b"0000000000000000_0000000000000000_0000011000110110_1101001111000111"; -- 0.024274097488947377
	pesos_i(12747) := b"0000000000000000_0000000000000000_0000001000100111_0011001100000010"; -- 0.008410632972477976
	pesos_i(12748) := b"0000000000000000_0000000000000000_0000110110110000_0111011111111000"; -- 0.05347394749655958
	pesos_i(12749) := b"1111111111111111_1111111111111111_1110011101001101_1100101010100111"; -- -0.09646924430724203
	pesos_i(12750) := b"1111111111111111_1111111111111111_1101110100010101_0011101000100101"; -- -0.13639484976547694
	pesos_i(12751) := b"1111111111111111_1111111111111111_1111111000111110_1000111110011010"; -- -0.0068578957004530585
	pesos_i(12752) := b"0000000000000000_0000000000000000_0000100011111011_0111000111101000"; -- 0.03508674543332101
	pesos_i(12753) := b"1111111111111111_1111111111111111_1110111011001110_0101111100111000"; -- -0.06716351389778033
	pesos_i(12754) := b"1111111111111111_1111111111111111_1111111010000111_0110000000001011"; -- -0.005746838775878647
	pesos_i(12755) := b"0000000000000000_0000000000000000_0001001110101010_0000001011101111"; -- 0.07681291890411648
	pesos_i(12756) := b"1111111111111111_1111111111111111_1111101100111111_1001100000001111"; -- -0.018560882840482323
	pesos_i(12757) := b"1111111111111111_1111111111111111_1110001111100010_1111000111011111"; -- -0.10981834706600495
	pesos_i(12758) := b"1111111111111111_1111111111111111_1110010111111111_1101000100000000"; -- -0.10156530139001434
	pesos_i(12759) := b"0000000000000000_0000000000000000_0010001111110011_1111001111010000"; -- 0.14044116808955343
	pesos_i(12760) := b"0000000000000000_0000000000000000_0010001010001100_0101001000001111"; -- 0.1349536215606849
	pesos_i(12761) := b"0000000000000000_0000000000000000_0001111100110010_1001101111001101"; -- 0.12186597588315447
	pesos_i(12762) := b"1111111111111111_1111111111111111_1110101011011011_0110001000001010"; -- -0.08258998150248953
	pesos_i(12763) := b"1111111111111111_1111111111111111_1111011000010110_1011000101010011"; -- -0.038716237200484845
	pesos_i(12764) := b"1111111111111111_1111111111111111_1110000011111010_0100010100111111"; -- -0.12118117537160387
	pesos_i(12765) := b"1111111111111111_1111111111111111_1111111010101010_0101111101011110"; -- -0.005212821477015302
	pesos_i(12766) := b"1111111111111111_1111111111111111_1101111001111001_0110100010000101"; -- -0.13095995674643557
	pesos_i(12767) := b"1111111111111111_1111111111111111_1101110100111011_0101001010110011"; -- -0.13581355213088686
	pesos_i(12768) := b"1111111111111111_1111111111111111_1111001101001010_1101010100100111"; -- -0.049639394717631735
	pesos_i(12769) := b"0000000000000000_0000000000000000_0001100100011011_1111100100010110"; -- 0.09808308396441323
	pesos_i(12770) := b"1111111111111111_1111111111111111_1110010010101100_0001101111011111"; -- -0.10674882712840181
	pesos_i(12771) := b"1111111111111111_1111111111111111_1111111011000100_1001110010101000"; -- -0.004812439814800779
	pesos_i(12772) := b"1111111111111111_1111111111111111_1110111001010010_1101000101110000"; -- -0.06904879577586172
	pesos_i(12773) := b"1111111111111111_1111111111111111_1110101100010000_1111001011101000"; -- -0.08177263097532068
	pesos_i(12774) := b"0000000000000000_0000000000000000_0000100100001000_0101000000110110"; -- 0.03528310122656584
	pesos_i(12775) := b"0000000000000000_0000000000000000_0000110101011100_0001010110010010"; -- 0.05218634427024342
	pesos_i(12776) := b"0000000000000000_0000000000000000_0001000010101111_1010110100000100"; -- 0.0651806006540955
	pesos_i(12777) := b"1111111111111111_1111111111111111_1110010011101110_1001010100110110"; -- -0.10573451462873606
	pesos_i(12778) := b"1111111111111111_1111111111111111_1111100111011110_1111100011001110"; -- -0.02394146885028124
	pesos_i(12779) := b"0000000000000000_0000000000000000_0001101001101101_1011000111110010"; -- 0.10323631431041923
	pesos_i(12780) := b"0000000000000000_0000000000000000_0001010001101110_1010110101010110"; -- 0.07981379838154302
	pesos_i(12781) := b"1111111111111111_1111111111111111_1110010110111011_0011000101011011"; -- -0.10261241466987119
	pesos_i(12782) := b"1111111111111111_1111111111111111_1110010000010000_0101101000011110"; -- -0.10912548806834667
	pesos_i(12783) := b"1111111111111111_1111111111111111_1110100101110001_0000111011010011"; -- -0.0881186231671379
	pesos_i(12784) := b"1111111111111111_1111111111111111_1101111010000100_0110110011001111"; -- -0.1307918543424327
	pesos_i(12785) := b"0000000000000000_0000000000000000_0000001010000011_0010010111101100"; -- 0.009813661756918916
	pesos_i(12786) := b"1111111111111111_1111111111111111_1110001101011111_1010000001101000"; -- -0.11182210419602248
	pesos_i(12787) := b"0000000000000000_0000000000000000_0010010010110100_0100011000100110"; -- 0.14337576312989306
	pesos_i(12788) := b"1111111111111111_1111111111111111_1101101001110110_1100011111000101"; -- -0.14662505581013924
	pesos_i(12789) := b"1111111111111111_1111111111111111_1101010101111111_0011110010111110"; -- -0.1660272631677872
	pesos_i(12790) := b"0000000000000000_0000000000000000_0000111111001100_1111011100000111"; -- 0.06172126685583016
	pesos_i(12791) := b"0000000000000000_0000000000000000_0000111101000001_0101101011001001"; -- 0.05959098248543421
	pesos_i(12792) := b"1111111111111111_1111111111111111_1111010001011010_0111111000110110"; -- -0.04549418630929236
	pesos_i(12793) := b"1111111111111111_1111111111111111_1110000110001101_1000100110110000"; -- -0.11893405388008632
	pesos_i(12794) := b"1111111111111111_1111111111111111_1110011101011110_1101011101100010"; -- -0.09620908595390634
	pesos_i(12795) := b"1111111111111111_1111111111111111_1110011001101101_0001001100011100"; -- -0.09989815302638431
	pesos_i(12796) := b"0000000000000000_0000000000000000_0000101100011001_0110101000010111"; -- 0.04335654309108668
	pesos_i(12797) := b"1111111111111111_1111111111111111_1110100101001101_0011000011111100"; -- -0.08866590357458103
	pesos_i(12798) := b"0000000000000000_0000000000000000_0000000100100000_0100000001111000"; -- 0.004398373824080084
	pesos_i(12799) := b"0000000000000000_0000000000000000_0000010100010110_1101001001101100"; -- 0.01987948555300375
	pesos_i(12800) := b"1111111111111111_1111111111111111_1110110100110100_1100111001111110"; -- -0.07341298506211846
	pesos_i(12801) := b"0000000000000000_0000000000000000_0000100111110101_0111101111010001"; -- 0.03890203346026669
	pesos_i(12802) := b"0000000000000000_0000000000000000_0001010101100000_0000110000111001"; -- 0.08349682234639698
	pesos_i(12803) := b"1111111111111111_1111111111111111_1111100110110000_1100100011111011"; -- -0.024646223802733184
	pesos_i(12804) := b"1111111111111111_1111111111111111_1110100010001110_1001110011100110"; -- -0.09157389996194042
	pesos_i(12805) := b"1111111111111111_1111111111111111_1110110101001000_0111100110100111"; -- -0.0731128661741037
	pesos_i(12806) := b"0000000000000000_0000000000000000_0000000110100111_0011010111001100"; -- 0.006457674250624576
	pesos_i(12807) := b"0000000000000000_0000000000000000_0001010000001111_1010100000001101"; -- 0.07836389845738281
	pesos_i(12808) := b"0000000000000000_0000000000000000_0000110010100101_1101101001001001"; -- 0.049405711071102594
	pesos_i(12809) := b"0000000000000000_0000000000000000_0010011000010010_0100010111100111"; -- 0.14871632460774098
	pesos_i(12810) := b"1111111111111111_1111111111111111_1110101000001001_0000001000001111"; -- -0.08580004808399831
	pesos_i(12811) := b"0000000000000000_0000000000000000_0001110101011000_0011110111101011"; -- 0.11462771411911751
	pesos_i(12812) := b"1111111111111111_1111111111111111_1111000011010111_1011110110010110"; -- -0.0592080600800859
	pesos_i(12813) := b"1111111111111111_1111111111111111_1110111110010111_0101111001001100"; -- -0.06409655241831885
	pesos_i(12814) := b"0000000000000000_0000000000000000_0010011011101101_0011100100101010"; -- 0.1520572402850078
	pesos_i(12815) := b"1111111111111111_1111111111111111_1110111100000110_0010100110101100"; -- -0.06631221340972997
	pesos_i(12816) := b"0000000000000000_0000000000000000_0001110001010111_0010011011010101"; -- 0.11070482922643445
	pesos_i(12817) := b"0000000000000000_0000000000000000_0001100111100100_0010000111011101"; -- 0.10113727224498313
	pesos_i(12818) := b"0000000000000000_0000000000000000_0000101110100010_0001111110001101"; -- 0.0454425543840027
	pesos_i(12819) := b"1111111111111111_1111111111111111_1110101100110000_0110001000010010"; -- -0.08129298260143031
	pesos_i(12820) := b"1111111111111111_1111111111111111_1101111110100100_1001110110001010"; -- -0.12639441842439592
	pesos_i(12821) := b"0000000000000000_0000000000000000_0001111001011010_1011001001110000"; -- 0.11857142677882107
	pesos_i(12822) := b"0000000000000000_0000000000000000_0000111000111101_0001011100110001"; -- 0.055619668380591916
	pesos_i(12823) := b"0000000000000000_0000000000000000_0001110110011101_1011110100100100"; -- 0.1156881535379023
	pesos_i(12824) := b"0000000000000000_0000000000000000_0001001111010000_0110110001101101"; -- 0.07739904082893956
	pesos_i(12825) := b"1111111111111111_1111111111111111_1110110011001110_1111001001111100"; -- -0.07496723629609031
	pesos_i(12826) := b"1111111111111111_1111111111111111_1111100110000110_0010111001011100"; -- -0.02529630912875113
	pesos_i(12827) := b"1111111111111111_1111111111111111_1110110011001100_0110100101011100"; -- -0.07500592717600632
	pesos_i(12828) := b"0000000000000000_0000000000000000_0000110110101011_1110011000110110"; -- 0.05340422467022527
	pesos_i(12829) := b"0000000000000000_0000000000000000_0001011010111001_0111010111001110"; -- 0.08876739776493305
	pesos_i(12830) := b"1111111111111111_1111111111111111_1111000101101010_0000111110100101"; -- -0.0569753857973209
	pesos_i(12831) := b"0000000000000000_0000000000000000_0001001000100000_0001000000100100"; -- 0.070801743276573
	pesos_i(12832) := b"1111111111111111_1111111111111111_1111010101001011_0000101111110001"; -- -0.04182362900830156
	pesos_i(12833) := b"0000000000000000_0000000000000000_0010000001100010_0110011000000100"; -- 0.12650144199141417
	pesos_i(12834) := b"0000000000000000_0000000000000000_0001010010110001_0001101111001100"; -- 0.08082746252774052
	pesos_i(12835) := b"1111111111111111_1111111111111111_1111111110001000_1110111100011111"; -- -0.0018168018850706251
	pesos_i(12836) := b"1111111111111111_1111111111111111_1111110001001101_0011011011110101"; -- -0.014446797469947953
	pesos_i(12837) := b"0000000000000000_0000000000000000_0001100001110000_1000000001011011"; -- 0.09546663497826988
	pesos_i(12838) := b"1111111111111111_1111111111111111_1111110010100101_0000100011100011"; -- -0.013106770174173174
	pesos_i(12839) := b"1111111111111111_1111111111111111_1110010110110100_1110000100001001"; -- -0.10270875491423512
	pesos_i(12840) := b"1111111111111111_1111111111111111_1111110101110111_1100000011101010"; -- -0.00989145564017884
	pesos_i(12841) := b"1111111111111111_1111111111111111_1110011101001011_0000111111000001"; -- -0.09651090190453342
	pesos_i(12842) := b"0000000000000000_0000000000000000_0001010100100010_0110010100000101"; -- 0.08255607013869423
	pesos_i(12843) := b"1111111111111111_1111111111111111_1111110010110010_1010001011011001"; -- -0.012899229133288354
	pesos_i(12844) := b"1111111111111111_1111111111111111_1111110100100111_1100011100001111"; -- -0.011111792455184311
	pesos_i(12845) := b"0000000000000000_0000000000000000_0001110001101100_0001011100001110"; -- 0.11102432343129853
	pesos_i(12846) := b"0000000000000000_0000000000000000_0000100011011010_1110000100110001"; -- 0.03458983837381917
	pesos_i(12847) := b"0000000000000000_0000000000000000_0001111100101100_1111110001001001"; -- 0.12178017418305173
	pesos_i(12848) := b"0000000000000000_0000000000000000_0000010110111101_0110111011000011"; -- 0.02242176299819117
	pesos_i(12849) := b"0000000000000000_0000000000000000_0000001101101000_0101100101000110"; -- 0.01331098514240069
	pesos_i(12850) := b"1111111111111111_1111111111111111_1110001111011101_1101010101101010"; -- -0.1098963371217739
	pesos_i(12851) := b"0000000000000000_0000000000000000_0001011011111010_1001000111100110"; -- 0.08976089351603311
	pesos_i(12852) := b"0000000000000000_0000000000000000_0000110100111011_1100111000100111"; -- 0.0516938062291544
	pesos_i(12853) := b"1111111111111111_1111111111111111_1111001011010111_0001110100111111"; -- -0.051405117104753546
	pesos_i(12854) := b"0000000000000000_0000000000000000_0000000010001000_0100001001011101"; -- 0.0020791508590500673
	pesos_i(12855) := b"0000000000000000_0000000000000000_0001000111110110_1011111001010010"; -- 0.07017125618026675
	pesos_i(12856) := b"1111111111111111_1111111111111111_1110111001101000_0101111010011001"; -- -0.0687199474328215
	pesos_i(12857) := b"0000000000000000_0000000000000000_0010000001000001_0001001001000010"; -- 0.12599290953953693
	pesos_i(12858) := b"1111111111111111_1111111111111111_1111111001110001_0111111111100110"; -- -0.0060806335913042775
	pesos_i(12859) := b"0000000000000000_0000000000000000_0001101101011000_0101010000011000"; -- 0.1068165359242181
	pesos_i(12860) := b"1111111111111111_1111111111111111_1100110011001011_0110010111100011"; -- -0.2000213928585825
	pesos_i(12861) := b"1111111111111111_1111111111111111_1110101101100110_1100011101111111"; -- -0.08046296271683713
	pesos_i(12862) := b"0000000000000000_0000000000000000_0000001001010001_1010011011010010"; -- 0.009058405086750506
	pesos_i(12863) := b"0000000000000000_0000000000000000_0001111010011000_0011000101110010"; -- 0.11950978307317109
	pesos_i(12864) := b"1111111111111111_1111111111111111_1110111001101011_0010110101010001"; -- -0.06867710846886174
	pesos_i(12865) := b"0000000000000000_0000000000000000_0000100011001100_1111000110101000"; -- 0.03437719680349708
	pesos_i(12866) := b"0000000000000000_0000000000000000_0010010000111100_0110111111101110"; -- 0.14154719894194548
	pesos_i(12867) := b"0000000000000000_0000000000000000_0010110010000011_1000101011111101"; -- 0.17388218563322402
	pesos_i(12868) := b"0000000000000000_0000000000000000_0000111011100010_1100101110000001"; -- 0.058148116208119674
	pesos_i(12869) := b"1111111111111111_1111111111111111_1111011001001010_0011001010001001"; -- -0.03793033759012689
	pesos_i(12870) := b"1111111111111111_1111111111111111_1111000110101000_0011101111011101"; -- -0.05602670520410149
	pesos_i(12871) := b"1111111111111111_1111111111111111_1111000111000111_1000010011001100"; -- -0.05554933559961615
	pesos_i(12872) := b"0000000000000000_0000000000000000_0001111011110001_0010111101101010"; -- 0.12086769424386679
	pesos_i(12873) := b"0000000000000000_0000000000000000_0001000101010011_0010101011010010"; -- 0.06767528184619356
	pesos_i(12874) := b"1111111111111111_1111111111111111_1111100000000011_0110101100101101"; -- -0.031197835499826684
	pesos_i(12875) := b"0000000000000000_0000000000000000_0000000101000010_0111001001110111"; -- 0.004920152661508026
	pesos_i(12876) := b"0000000000000000_0000000000000000_0000011011010101_1000110110111001"; -- 0.026696069506792836
	pesos_i(12877) := b"0000000000000000_0000000000000000_0001001101010111_1110100001110001"; -- 0.07556011927459128
	pesos_i(12878) := b"1111111111111111_1111111111111111_1110000010110101_1101110010101100"; -- -0.1222250062063164
	pesos_i(12879) := b"0000000000000000_0000000000000000_0000001100111001_0011000000000011"; -- 0.01259136269421005
	pesos_i(12880) := b"1111111111111111_1111111111111111_1101110010111101_0010111111101100"; -- -0.13773823254192433
	pesos_i(12881) := b"1111111111111111_1111111111111111_1110000011101011_1011100000111010"; -- -0.1214032037031073
	pesos_i(12882) := b"0000000000000000_0000000000000000_0010001110001111_0110011011011011"; -- 0.1389068875891627
	pesos_i(12883) := b"1111111111111111_1111111111111111_1110100011110010_1011101100100001"; -- -0.09004621938928828
	pesos_i(12884) := b"0000000000000000_0000000000000000_0010000001001111_1111111111100100"; -- 0.12622069658313603
	pesos_i(12885) := b"0000000000000000_0000000000000000_0001110011001110_1001111110110000"; -- 0.1125278287224022
	pesos_i(12886) := b"0000000000000000_0000000000000000_0001000111100110_1000100110000100"; -- 0.06992396813114395
	pesos_i(12887) := b"0000000000000000_0000000000000000_0010000000101101_1011101111000001"; -- 0.12569783656996408
	pesos_i(12888) := b"1111111111111111_1111111111111111_1110111000000001_1101110111110001"; -- -0.07028401258530556
	pesos_i(12889) := b"0000000000000000_0000000000000000_0001101010000010_1010011100100110"; -- 0.1035561054184796
	pesos_i(12890) := b"0000000000000000_0000000000000000_0000100000010011_1110111000101111"; -- 0.03155411383326804
	pesos_i(12891) := b"0000000000000000_0000000000000000_0000001010010010_0010111001000100"; -- 0.010043040740564233
	pesos_i(12892) := b"0000000000000000_0000000000000000_0000111100110010_1111111011101101"; -- 0.05937188412443612
	pesos_i(12893) := b"1111111111111111_1111111111111111_1110111100010001_1001110001010110"; -- -0.06613753232022278
	pesos_i(12894) := b"1111111111111111_1111111111111111_1110011100010100_1011010101101000"; -- -0.09734026165179373
	pesos_i(12895) := b"0000000000000000_0000000000000000_0000100011110001_1111000010110011"; -- 0.03494171496020148
	pesos_i(12896) := b"0000000000000000_0000000000000000_0001010100100100_1100110001100000"; -- 0.08259274803193087
	pesos_i(12897) := b"0000000000000000_0000000000000000_0000110011011100_1000111010011010"; -- 0.05024043330791839
	pesos_i(12898) := b"1111111111111111_1111111111111111_1101101000100011_1110011000010100"; -- -0.14788972862941782
	pesos_i(12899) := b"0000000000000000_0000000000000000_0001010000001000_0111001001100110"; -- 0.0782538890918036
	pesos_i(12900) := b"0000000000000000_0000000000000000_0000101001010010_0101011011001100"; -- 0.040318894087154805
	pesos_i(12901) := b"1111111111111111_1111111111111111_1110010000011110_1000110001110011"; -- -0.10890886485061319
	pesos_i(12902) := b"0000000000000000_0000000000000000_0000110000011000_1010000101101011"; -- 0.04725083217028277
	pesos_i(12903) := b"1111111111111111_1111111111111111_1101001111100111_1101101111001101"; -- -0.17224336853519456
	pesos_i(12904) := b"1111111111111111_1111111111111111_1110101000000100_0000111000110011"; -- -0.08587561859501854
	pesos_i(12905) := b"0000000000000000_0000000000000000_0001011101100101_0100000111010001"; -- 0.0913888106280253
	pesos_i(12906) := b"1111111111111111_1111111111111111_1111000000001110_0101100001010101"; -- -0.06228111196876836
	pesos_i(12907) := b"0000000000000000_0000000000000000_0000000101000001_1111011110110001"; -- 0.004912834914245755
	pesos_i(12908) := b"0000000000000000_0000000000000000_0001111001100111_1010000010010001"; -- 0.11876872571996983
	pesos_i(12909) := b"1111111111111111_1111111111111111_1110001010100011_0101011011000111"; -- -0.11469514501800215
	pesos_i(12910) := b"1111111111111111_1111111111111111_1110110000111101_1000010100101100"; -- -0.07718627621121357
	pesos_i(12911) := b"1111111111111111_1111111111111111_1111110110011111_1110000011000010"; -- -0.009279206023586103
	pesos_i(12912) := b"0000000000000000_0000000000000000_0000011100001010_0001100101000011"; -- 0.027497843621967628
	pesos_i(12913) := b"0000000000000000_0000000000000000_0000110101101110_1110010011101001"; -- 0.0524733610106778
	pesos_i(12914) := b"1111111111111111_1111111111111111_1111001110101010_1101010011101001"; -- -0.04817456546829892
	pesos_i(12915) := b"0000000000000000_0000000000000000_0000101110101110_0101011000011010"; -- 0.04562891144509149
	pesos_i(12916) := b"0000000000000000_0000000000000000_0001001111101101_1100101011110101"; -- 0.07784718029332935
	pesos_i(12917) := b"0000000000000000_0000000000000000_0000100000001100_0101001101101010"; -- 0.031438077241043506
	pesos_i(12918) := b"1111111111111111_1111111111111111_1101111101010101_0001100011011000"; -- -0.127607772145673
	pesos_i(12919) := b"0000000000000000_0000000000000000_0010001011011110_1110111101110011"; -- 0.13621422350191503
	pesos_i(12920) := b"1111111111111111_1111111111111111_1111101000100000_0111111000011101"; -- -0.022941701838051876
	pesos_i(12921) := b"0000000000000000_0000000000000000_0001100001101110_0100110110000001"; -- 0.09543308633247966
	pesos_i(12922) := b"1111111111111111_1111111111111111_1111001101001000_1011111110001101"; -- -0.04967119988242067
	pesos_i(12923) := b"1111111111111111_1111111111111111_1110000100000001_1000001001101100"; -- -0.12107071742745645
	pesos_i(12924) := b"0000000000000000_0000000000000000_0001110110101110_0100010000101100"; -- 0.11594034275769506
	pesos_i(12925) := b"0000000000000000_0000000000000000_0000011001100101_1111111000100101"; -- 0.024993785811104154
	pesos_i(12926) := b"0000000000000000_0000000000000000_0000110100110011_0011101100001010"; -- 0.051562967322467526
	pesos_i(12927) := b"1111111111111111_1111111111111111_1110110110100010_0011111101101001"; -- -0.07174304659717994
	pesos_i(12928) := b"1111111111111111_1111111111111111_1101110001111110_1111000100100110"; -- -0.1386880189849296
	pesos_i(12929) := b"0000000000000000_0000000000000000_0010100101110011_0100100010100111"; -- 0.16191534121622
	pesos_i(12930) := b"0000000000000000_0000000000000000_0000110000001111_0001101110101010"; -- 0.04710553065191846
	pesos_i(12931) := b"0000000000000000_0000000000000000_0001000001101100_0110010110110110"; -- 0.06415401168858659
	pesos_i(12932) := b"1111111111111111_1111111111111111_1110000001111111_1110000001011000"; -- -0.12304876192156036
	pesos_i(12933) := b"1111111111111111_1111111111111111_1110000001010111_0111011100011101"; -- -0.12366538561460112
	pesos_i(12934) := b"0000000000000000_0000000000000000_0000110010001101_0101010010000100"; -- 0.04903152683709301
	pesos_i(12935) := b"1111111111111111_1111111111111111_1111111101011000_0111100111010010"; -- -0.002556215496847076
	pesos_i(12936) := b"0000000000000000_0000000000000000_0000111100000111_1011100001101110"; -- 0.058711554470043434
	pesos_i(12937) := b"1111111111111111_1111111111111111_1110101001100001_0010011011011000"; -- -0.08445508208745926
	pesos_i(12938) := b"1111111111111111_1111111111111111_1110011101110101_0000000001000101"; -- -0.0958709556388534
	pesos_i(12939) := b"1111111111111111_1111111111111111_1101110110101111_1011011100011111"; -- -0.13403754714295404
	pesos_i(12940) := b"1111111111111111_1111111111111111_1110100101001100_1000101101110101"; -- -0.0886757696889608
	pesos_i(12941) := b"0000000000000000_0000000000000000_0001101110111010_0100110001011101"; -- 0.1083114363240414
	pesos_i(12942) := b"1111111111111111_1111111111111111_1110001100010100_0111011111101110"; -- -0.11296892590512851
	pesos_i(12943) := b"1111111111111111_1111111111111111_1101111011001111_1101011010001110"; -- -0.12964114231155324
	pesos_i(12944) := b"1111111111111111_1111111111111111_1111001001110011_1101011000110010"; -- -0.052919972215131526
	pesos_i(12945) := b"1111111111111111_1111111111111111_1111100111001010_0111001111001011"; -- -0.024254572833125262
	pesos_i(12946) := b"1111111111111111_1111111111111111_1110001010001000_1100000011011011"; -- -0.11510080964497964
	pesos_i(12947) := b"1111111111111111_1111111111111111_1101111110000001_0100110101010101"; -- -0.12693325687876497
	pesos_i(12948) := b"1111111111111111_1111111111111111_1111100011111000_0111101001011100"; -- -0.027458527059407774
	pesos_i(12949) := b"0000000000000000_0000000000000000_0001001010101011_0001011101100101"; -- 0.07292314730091298
	pesos_i(12950) := b"0000000000000000_0000000000000000_0010000100101000_1010100010100000"; -- 0.1295266524842883
	pesos_i(12951) := b"0000000000000000_0000000000000000_0001010000111101_0001111100100011"; -- 0.07905764205738858
	pesos_i(12952) := b"1111111111111111_1111111111111111_1111001100101011_0011110000010010"; -- -0.050121541680662594
	pesos_i(12953) := b"0000000000000000_0000000000000000_0001011101000010_1111000110100001"; -- 0.09086523228507173
	pesos_i(12954) := b"1111111111111111_1111111111111111_1111101110001000_1010100101111101"; -- -0.017445952451415017
	pesos_i(12955) := b"1111111111111111_1111111111111111_1111101001100111_0000101001010011"; -- -0.021865229433070756
	pesos_i(12956) := b"0000000000000000_0000000000000000_0000100001100100_0000100001011110"; -- 0.032776377630070866
	pesos_i(12957) := b"0000000000000000_0000000000000000_0001011000111000_0101000111000100"; -- 0.08679686584144398
	pesos_i(12958) := b"1111111111111111_1111111111111111_1101110010010110_0101010000101010"; -- -0.13833116504881462
	pesos_i(12959) := b"0000000000000000_0000000000000000_0000111101100110_1011011011111111"; -- 0.0601610537882015
	pesos_i(12960) := b"0000000000000000_0000000000000000_0001001001011100_1011100111000110"; -- 0.07172738144881229
	pesos_i(12961) := b"1111111111111111_1111111111111111_1101110101011010_0001101101000001"; -- -0.13534383441397035
	pesos_i(12962) := b"1111111111111111_1111111111111111_1101101111100000_0111010000101000"; -- -0.1411063579116912
	pesos_i(12963) := b"0000000000000000_0000000000000000_0010000011111111_0001011010000000"; -- 0.12889233232944966
	pesos_i(12964) := b"1111111111111111_1111111111111111_1101100001100010_1011010001000100"; -- -0.15474389409422945
	pesos_i(12965) := b"1111111111111111_1111111111111111_1101101011011100_1011000110101101"; -- -0.14506997600640295
	pesos_i(12966) := b"0000000000000000_0000000000000000_0000110011010111_0010101111111000"; -- 0.050158260434279185
	pesos_i(12967) := b"1111111111111111_1111111111111111_1110100011000100_1110001101011000"; -- -0.09074572667033676
	pesos_i(12968) := b"1111111111111111_1111111111111111_1111101110011010_1011110011111001"; -- -0.01717013292727411
	pesos_i(12969) := b"0000000000000000_0000000000000000_0010001011010010_0000101010111101"; -- 0.1360174857102167
	pesos_i(12970) := b"1111111111111111_1111111111111111_1110000111111000_0111010011011100"; -- -0.11730260493572327
	pesos_i(12971) := b"0000000000000000_0000000000000000_0000111010110100_0011010101100010"; -- 0.05743726389469098
	pesos_i(12972) := b"1111111111111111_1111111111111111_1111111100110101_0111011001000000"; -- -0.003090485961134312
	pesos_i(12973) := b"0000000000000000_0000000000000000_0000001001101000_0001110000101001"; -- 0.009401092510937447
	pesos_i(12974) := b"0000000000000000_0000000000000000_0010000000010000_0000000000001000"; -- 0.12524414247500998
	pesos_i(12975) := b"0000000000000000_0000000000000000_0010010000010100_0110011111110001"; -- 0.1409363711356146
	pesos_i(12976) := b"1111111111111111_1111111111111111_1110010011100101_1101100011100110"; -- -0.10586780923565016
	pesos_i(12977) := b"1111111111111111_1111111111111111_1110000001111001_0100110111100111"; -- -0.12314904315050079
	pesos_i(12978) := b"1111111111111111_1111111111111111_1110000100010110_0110000011101011"; -- -0.12075227984648736
	pesos_i(12979) := b"0000000000000000_0000000000000000_0001101101000110_1111100111010110"; -- 0.10655175658925103
	pesos_i(12980) := b"1111111111111111_1111111111111111_1111111100101101_0110110000111001"; -- -0.0032131538840547095
	pesos_i(12981) := b"0000000000000000_0000000000000000_0000011111000100_0101010110111011"; -- 0.03033958267741672
	pesos_i(12982) := b"1111111111111111_1111111111111111_1110101001110100_0010010000111011"; -- -0.08416532094014123
	pesos_i(12983) := b"1111111111111111_1111111111111111_1111011110010011_0000111010110100"; -- -0.03291233164799844
	pesos_i(12984) := b"0000000000000000_0000000000000000_0001111101110001_1111011101001001"; -- 0.12283273255450383
	pesos_i(12985) := b"1111111111111111_1111111111111111_1110111110100001_1001110001010110"; -- -0.06394026653645099
	pesos_i(12986) := b"1111111111111111_1111111111111111_1111100100101100_1010100110001010"; -- -0.02666225792496816
	pesos_i(12987) := b"1111111111111111_1111111111111111_1111001011011000_0010111000101100"; -- -0.05138884945180229
	pesos_i(12988) := b"0000000000000000_0000000000000000_0001101001000010_0110100111101110"; -- 0.10257589387717188
	pesos_i(12989) := b"0000000000000000_0000000000000000_0000111011111010_1010011011110111"; -- 0.05851214923760307
	pesos_i(12990) := b"0000000000000000_0000000000000000_0000110100000101_1101000101100111"; -- 0.050870025290636535
	pesos_i(12991) := b"0000000000000000_0000000000000000_0000011101010010_0000011001001000"; -- 0.028595345210814645
	pesos_i(12992) := b"0000000000000000_0000000000000000_0000000010000101_1100001011001101"; -- 0.0020410298661154565
	pesos_i(12993) := b"0000000000000000_0000000000000000_0001110011000110_0000111100001110"; -- 0.11239713757538879
	pesos_i(12994) := b"0000000000000000_0000000000000000_0000110010001101_1100001010100110"; -- 0.049038091279595346
	pesos_i(12995) := b"0000000000000000_0000000000000000_0000101100111010_0100011111100001"; -- 0.043858044054367606
	pesos_i(12996) := b"0000000000000000_0000000000000000_0000101010011100_1110001010010000"; -- 0.04145637518725221
	pesos_i(12997) := b"1111111111111111_1111111111111111_1110000001111111_1101001000101001"; -- -0.12304960738174042
	pesos_i(12998) := b"1111111111111111_1111111111111111_1111110101001110_0110010010100100"; -- -0.010522565866110365
	pesos_i(12999) := b"0000000000000000_0000000000000000_0001011100001011_0010101010011101"; -- 0.09001413669063923
	pesos_i(13000) := b"1111111111111111_1111111111111111_1110000110001101_0110011110001111"; -- -0.11893608814949079
	pesos_i(13001) := b"0000000000000000_0000000000000000_0000111001101001_1010010110000110"; -- 0.05629953877006069
	pesos_i(13002) := b"0000000000000000_0000000000000000_0000111000101100_0000111101111101"; -- 0.055359809803125166
	pesos_i(13003) := b"0000000000000000_0000000000000000_0000001111001110_0011111001010110"; -- 0.014865775997156659
	pesos_i(13004) := b"0000000000000000_0000000000000000_0010010011011000_1101111001111010"; -- 0.14393415903425083
	pesos_i(13005) := b"1111111111111111_1111111111111111_1111000001101111_1100000011000000"; -- -0.06079478551997015
	pesos_i(13006) := b"1111111111111111_1111111111111111_1111011110100101_1000001001010110"; -- -0.03263078120537977
	pesos_i(13007) := b"1111111111111111_1111111111111111_1101101110101001_1101001001110111"; -- -0.1419399698520111
	pesos_i(13008) := b"1111111111111111_1111111111111111_1101100000010110_1010010010101001"; -- -0.15590449206406032
	pesos_i(13009) := b"0000000000000000_0000000000000000_0001100100010100_0001111001000111"; -- 0.09796323035065006
	pesos_i(13010) := b"1111111111111111_1111111111111111_1111111101101000_0011000101110000"; -- -0.002316389150973332
	pesos_i(13011) := b"1111111111111111_1111111111111111_1111100111101111_1010010011100001"; -- -0.02368707194440241
	pesos_i(13012) := b"1111111111111111_1111111111111111_1110010001110100_0110010001001101"; -- -0.107599002019954
	pesos_i(13013) := b"1111111111111111_1111111111111111_1101100101001110_0111110100000000"; -- -0.15114611390200966
	pesos_i(13014) := b"1111111111111111_1111111111111111_1111001000011101_0100111111111010"; -- -0.05424022813671091
	pesos_i(13015) := b"0000000000000000_0000000000000000_0010000001111101_0011111000001100"; -- 0.12691104685643936
	pesos_i(13016) := b"1111111111111111_1111111111111111_1111100111101100_1010100000100111"; -- -0.023732653169722836
	pesos_i(13017) := b"1111111111111111_1111111111111111_1110001010110010_0011100110111001"; -- -0.11446799495234192
	pesos_i(13018) := b"1111111111111111_1111111111111111_1101110110110101_1000110001000101"; -- -0.13394854841040627
	pesos_i(13019) := b"0000000000000000_0000000000000000_0000110001111111_1010101101111011"; -- 0.048823087154206066
	pesos_i(13020) := b"1111111111111111_1111111111111111_1111101011000010_1110110000111010"; -- -0.020463214802843962
	pesos_i(13021) := b"1111111111111111_1111111111111111_1111100101000110_1111100011110000"; -- -0.026260796837838135
	pesos_i(13022) := b"1111111111111111_1111111111111111_1111010011110111_0100010100110001"; -- -0.04310195499010929
	pesos_i(13023) := b"1111111111111111_1111111111111111_1110110111111100_0110101110000101"; -- -0.0703671264698059
	pesos_i(13024) := b"1111111111111111_1111111111111111_1101011000111110_1100101101000100"; -- -0.1631043394371438
	pesos_i(13025) := b"1111111111111111_1111111111111111_1110100101110011_1111001101100010"; -- -0.08807448256515399
	pesos_i(13026) := b"1111111111111111_1111111111111111_1110011010001010_1100010010010101"; -- -0.09944506986509359
	pesos_i(13027) := b"0000000000000000_0000000000000000_0000111111010100_1101100110101010"; -- 0.061841587114299434
	pesos_i(13028) := b"1111111111111111_1111111111111111_1110000101011010_0110010100101111"; -- -0.11971442795088992
	pesos_i(13029) := b"0000000000000000_0000000000000000_0001110000000111_0011101110100010"; -- 0.10948536592450439
	pesos_i(13030) := b"0000000000000000_0000000000000000_0001001010001101_0100110010100011"; -- 0.07246855723530157
	pesos_i(13031) := b"0000000000000000_0000000000000000_0001010111010010_1100101111101010"; -- 0.08524774984135113
	pesos_i(13032) := b"0000000000000000_0000000000000000_0010000100100011_0011111011100000"; -- 0.12944405526935557
	pesos_i(13033) := b"1111111111111111_1111111111111111_1111101010110011_0111000111011111"; -- -0.0206993895542305
	pesos_i(13034) := b"1111111111111111_1111111111111111_1101111001100001_1110111001000101"; -- -0.13131819558795818
	pesos_i(13035) := b"0000000000000000_0000000000000000_0000101000011000_1010000000111110"; -- 0.03943826217463313
	pesos_i(13036) := b"1111111111111111_1111111111111111_1110000101001000_0000010001110010"; -- -0.11999485217207272
	pesos_i(13037) := b"1111111111111111_1111111111111111_1111010011010011_1101010101101110"; -- -0.04364267406785756
	pesos_i(13038) := b"0000000000000000_0000000000000000_0001110011001101_1100110111100001"; -- 0.11251532304026322
	pesos_i(13039) := b"0000000000000000_0000000000000000_0001111100000101_0001000001000110"; -- 0.12117101386024996
	pesos_i(13040) := b"1111111111111111_1111111111111111_1111000111111011_0110100001110011"; -- -0.05475756829323128
	pesos_i(13041) := b"1111111111111111_1111111111111111_1110111100100001_1000111100100011"; -- -0.06589417832123146
	pesos_i(13042) := b"1111111111111111_1111111111111111_1110110110010000_1110000100000101"; -- -0.07200807215790145
	pesos_i(13043) := b"1111111111111111_1111111111111111_1111001011000001_0110110001100010"; -- -0.05173609349432174
	pesos_i(13044) := b"0000000000000000_0000000000000000_0001100010001110_0011001011011000"; -- 0.0959197785254381
	pesos_i(13045) := b"0000000000000000_0000000000000000_0001001111110100_1110011110100100"; -- 0.07795570140578767
	pesos_i(13046) := b"1111111111111111_1111111111111111_1110010001100100_1101000111011111"; -- -0.10783661180547013
	pesos_i(13047) := b"0000000000000000_0000000000000000_0000010011100000_0101110111101010"; -- 0.01904856638302764
	pesos_i(13048) := b"0000000000000000_0000000000000000_0001001011011110_1011110011011111"; -- 0.07371120873813651
	pesos_i(13049) := b"0000000000000000_0000000000000000_0000011000110101_0100000101101011"; -- 0.02425011504016458
	pesos_i(13050) := b"0000000000000000_0000000000000000_0001100001100000_0110011111110011"; -- 0.09522103965916125
	pesos_i(13051) := b"1111111111111111_1111111111111111_1110001000111101_1110100000101011"; -- -0.11624287562260584
	pesos_i(13052) := b"0000000000000000_0000000000000000_0010000000010110_1111110101110101"; -- 0.1253508005755964
	pesos_i(13053) := b"0000000000000000_0000000000000000_0001011010111011_0110110011011111"; -- 0.08879738284298395
	pesos_i(13054) := b"0000000000000000_0000000000000000_0000010110000001_0110101100000010"; -- 0.021506012047549476
	pesos_i(13055) := b"0000000000000000_0000000000000000_0001001101110111_1001100010000000"; -- 0.076043635713395
	pesos_i(13056) := b"0000000000000000_0000000000000000_0000101100010001_0101101010101101"; -- 0.043233554197056816
	pesos_i(13057) := b"0000000000000000_0000000000000000_0000101010010101_0110100010110100"; -- 0.04134230045572328
	pesos_i(13058) := b"0000000000000000_0000000000000000_0001000110000011_0000111111101010"; -- 0.06840609986411786
	pesos_i(13059) := b"1111111111111111_1111111111111111_1111011100111111_0111001101110110"; -- -0.034188064375595115
	pesos_i(13060) := b"0000000000000000_0000000000000000_0000000110010110_0001111011110000"; -- 0.006196912470422888
	pesos_i(13061) := b"0000000000000000_0000000000000000_0001000001010001_0001100101111010"; -- 0.0637374805290119
	pesos_i(13062) := b"1111111111111111_1111111111111111_1110011001001001_1101000100001110"; -- -0.10043614769076156
	pesos_i(13063) := b"1111111111111111_1111111111111111_1111001100110111_0101100010111000"; -- -0.049936728471702094
	pesos_i(13064) := b"0000000000000000_0000000000000000_0010011101111101_0100111100001010"; -- 0.15425580975223535
	pesos_i(13065) := b"1111111111111111_1111111111111111_1110001101100000_1011101100001011"; -- -0.1118052577109324
	pesos_i(13066) := b"0000000000000000_0000000000000000_0001010011101011_0100111110010111"; -- 0.08171555943779017
	pesos_i(13067) := b"0000000000000000_0000000000000000_0001010011010111_1100111110110100"; -- 0.08141801963847745
	pesos_i(13068) := b"1111111111111111_1111111111111111_1101100110010110_0000001001010100"; -- -0.1500547928916839
	pesos_i(13069) := b"0000000000000000_0000000000000000_0000111010010101_0011111011110101"; -- 0.05696481217744295
	pesos_i(13070) := b"1111111111111111_1111111111111111_1110000101100010_0100010011100001"; -- -0.11959428312274138
	pesos_i(13071) := b"1111111111111111_1111111111111111_1110100100111000_1101001001000111"; -- -0.08897672441866589
	pesos_i(13072) := b"0000000000000000_0000000000000000_0001111011001110_1010000011001110"; -- 0.12034039524666128
	pesos_i(13073) := b"1111111111111111_1111111111111111_1110011010100110_1000011101100110"; -- -0.09902147067037417
	pesos_i(13074) := b"1111111111111111_1111111111111111_1110111000011001_0010011101110000"; -- -0.06992867968762655
	pesos_i(13075) := b"1111111111111111_1111111111111111_1110101110101011_1001101110011010"; -- -0.0794127224205933
	pesos_i(13076) := b"1111111111111111_1111111111111111_1110011001000000_0011011010000110"; -- -0.10058268775099174
	pesos_i(13077) := b"1111111111111111_1111111111111111_1111101010011110_1111011101110110"; -- -0.021011861533329766
	pesos_i(13078) := b"1111111111111111_1111111111111111_1110101000111001_0101011110001111"; -- -0.08506253007137256
	pesos_i(13079) := b"0000000000000000_0000000000000000_0001111110001111_1100111111010100"; -- 0.1232881443054646
	pesos_i(13080) := b"1111111111111111_1111111111111111_1110110011101100_1110101101010011"; -- -0.0745098994354403
	pesos_i(13081) := b"1111111111111111_1111111111111111_1111010011000011_0001000100101010"; -- -0.043898513104297175
	pesos_i(13082) := b"0000000000000000_0000000000000000_0010000001011010_0011001110010110"; -- 0.12637636570545802
	pesos_i(13083) := b"0000000000000000_0000000000000000_0000110001110110_1010001001001011"; -- 0.04868521041295268
	pesos_i(13084) := b"1111111111111111_1111111111111111_1111001010101101_1100111011010011"; -- -0.052035401867240066
	pesos_i(13085) := b"0000000000000000_0000000000000000_0000111110101001_1001010101001101"; -- 0.06118138447431376
	pesos_i(13086) := b"1111111111111111_1111111111111111_1111000110100100_1101110000110001"; -- -0.056078184247816965
	pesos_i(13087) := b"0000000000000000_0000000000000000_0001001011100100_0111000001110111"; -- 0.07379820739189613
	pesos_i(13088) := b"1111111111111111_1111111111111111_1110011101100101_0010100000110001"; -- -0.09611271665083233
	pesos_i(13089) := b"0000000000000000_0000000000000000_0000010110001000_0011000000100010"; -- 0.021609314190744473
	pesos_i(13090) := b"0000000000000000_0000000000000000_0001101010110010_0101100100010111"; -- 0.10428387465283474
	pesos_i(13091) := b"1111111111111111_1111111111111111_1110001000100001_0011111111011000"; -- -0.11668015455850786
	pesos_i(13092) := b"0000000000000000_0000000000000000_0001001011011100_0010100000100010"; -- 0.07367182568029558
	pesos_i(13093) := b"0000000000000000_0000000000000000_0000001110010100_0100011000111000"; -- 0.013981236243850103
	pesos_i(13094) := b"1111111111111111_1111111111111111_1111111010111100_0011001000101001"; -- -0.004940857894060613
	pesos_i(13095) := b"0000000000000000_0000000000000000_0001001100101111_1110100100101110"; -- 0.074949811659513
	pesos_i(13096) := b"1111111111111111_1111111111111111_1110110011011111_0011001111011000"; -- -0.0747191999754981
	pesos_i(13097) := b"0000000000000000_0000000000000000_0000000111100110_0000000111010011"; -- 0.00741588022774195
	pesos_i(13098) := b"1111111111111111_1111111111111111_1110011111110100_0011110100110010"; -- -0.09392945792463757
	pesos_i(13099) := b"0000000000000000_0000000000000000_0000100011010100_1011010111011100"; -- 0.03449570283068331
	pesos_i(13100) := b"1111111111111111_1111111111111111_1111011101111100_0000001110110100"; -- -0.03326393935416839
	pesos_i(13101) := b"1111111111111111_1111111111111111_1111011010001011_1001011000001111"; -- -0.036932584085679954
	pesos_i(13102) := b"0000000000000000_0000000000000000_0000101001101000_0001101010000000"; -- 0.04065099363428966
	pesos_i(13103) := b"0000000000000000_0000000000000000_0000000011010010_1011101001110001"; -- 0.0032154585857925503
	pesos_i(13104) := b"1111111111111111_1111111111111111_1111011111111101_0101011001000111"; -- -0.03129063390625142
	pesos_i(13105) := b"1111111111111111_1111111111111111_1110011000111000_0000100111000011"; -- -0.10070742588234384
	pesos_i(13106) := b"0000000000000000_0000000000000000_0010000110100000_0111101101010101"; -- 0.13135500751894524
	pesos_i(13107) := b"0000000000000000_0000000000000000_0001001001100100_0101111101010001"; -- 0.07184406030195775
	pesos_i(13108) := b"1111111111111111_1111111111111111_1110001100001111_0000110101011110"; -- -0.11305157135281066
	pesos_i(13109) := b"0000000000000000_0000000000000000_0001101101100111_1100110101101000"; -- 0.10705264851984592
	pesos_i(13110) := b"1111111111111111_1111111111111111_1110001010010111_1000010111000101"; -- -0.11487544945685953
	pesos_i(13111) := b"0000000000000000_0000000000000000_0001000111101110_1010101110010100"; -- 0.07004806873343351
	pesos_i(13112) := b"1111111111111111_1111111111111111_1110110111011101_1011101101111100"; -- -0.07083538267722612
	pesos_i(13113) := b"0000000000000000_0000000000000000_0001111011010011_0001011010101001"; -- 0.12040845519163994
	pesos_i(13114) := b"0000000000000000_0000000000000000_0001101011111000_0111111110110111"; -- 0.10535429203657698
	pesos_i(13115) := b"1111111111111111_1111111111111111_1111000001000101_0100001000110001"; -- -0.06144319817722389
	pesos_i(13116) := b"0000000000000000_0000000000000000_0001001100101100_0101100010101101"; -- 0.07489542226932602
	pesos_i(13117) := b"0000000000000000_0000000000000000_0001100101100011_1101000101111000"; -- 0.09917935532840381
	pesos_i(13118) := b"1111111111111111_1111111111111111_1110110101010000_1011011010001101"; -- -0.07298716601384163
	pesos_i(13119) := b"1111111111111111_1111111111111111_1110010110000001_0100010011101011"; -- -0.1034962584831375
	pesos_i(13120) := b"0000000000000000_0000000000000000_0000111011110000_0010100110010011"; -- 0.05835208735773415
	pesos_i(13121) := b"1111111111111111_1111111111111111_1111000100010011_1001000111011101"; -- -0.058295138876380735
	pesos_i(13122) := b"1111111111111111_1111111111111111_1111001010001100_0100111101111001"; -- -0.05254653259658215
	pesos_i(13123) := b"0000000000000000_0000000000000000_0001111001000000_0111001010110000"; -- 0.11817089834939365
	pesos_i(13124) := b"0000000000000000_0000000000000000_0001110111110100_1101111111111101"; -- 0.11701774534666447
	pesos_i(13125) := b"1111111111111111_1111111111111111_1110100101001010_1111000110000101"; -- -0.08870020396157145
	pesos_i(13126) := b"0000000000000000_0000000000000000_0001000101010001_1110000101100111"; -- 0.06765564686666783
	pesos_i(13127) := b"0000000000000000_0000000000000000_0001101111011010_1111000100010110"; -- 0.10880953592125532
	pesos_i(13128) := b"1111111111111111_1111111111111111_1110011001000010_1010010101010000"; -- -0.10054556647024102
	pesos_i(13129) := b"1111111111111111_1111111111111111_1111100000101101_1110110100101001"; -- -0.030549218605579468
	pesos_i(13130) := b"0000000000000000_0000000000000000_0010100000110100_1110000101000110"; -- 0.1570568843957601
	pesos_i(13131) := b"0000000000000000_0000000000000000_0000010111000000_1001001110101000"; -- 0.02246973859353326
	pesos_i(13132) := b"0000000000000000_0000000000000000_0000001100110000_0000100000110001"; -- 0.012451660192629747
	pesos_i(13133) := b"1111111111111111_1111111111111111_1101110110111101_0111111100101100"; -- -0.1338272588409882
	pesos_i(13134) := b"1111111111111111_1111111111111111_1110000101011101_1001001111110110"; -- -0.11966586355867552
	pesos_i(13135) := b"1111111111111111_1111111111111111_1110001000101011_1100000111010011"; -- -0.11651981921640281
	pesos_i(13136) := b"0000000000000000_0000000000000000_0001111110110101_0001100010101101"; -- 0.12385706162213314
	pesos_i(13137) := b"0000000000000000_0000000000000000_0000000100011101_1001000100110111"; -- 0.00435741047426015
	pesos_i(13138) := b"0000000000000000_0000000000000000_0001011010110011_1001101011010101"; -- 0.08867805202491517
	pesos_i(13139) := b"1111111111111111_1111111111111111_1101011100011011_0010010000101011"; -- -0.15974210682358814
	pesos_i(13140) := b"1111111111111111_1111111111111111_1110110011110001_1011101101101001"; -- -0.07443646138899297
	pesos_i(13141) := b"1111111111111111_1111111111111111_1110000000101101_1100101101011100"; -- -0.12430123340574133
	pesos_i(13142) := b"0000000000000000_0000000000000000_0001001100010011_0110100000111000"; -- 0.07451487895591055
	pesos_i(13143) := b"1111111111111111_1111111111111111_1111011010011110_1000100000000101"; -- -0.036643503918116674
	pesos_i(13144) := b"0000000000000000_0000000000000000_0000010011111110_1110110110101111"; -- 0.019514899572000415
	pesos_i(13145) := b"1111111111111111_1111111111111111_1111010000100111_0001010000110001"; -- -0.04627870367405489
	pesos_i(13146) := b"1111111111111111_1111111111111111_1101110101101011_0000000010011101"; -- -0.13508602301538983
	pesos_i(13147) := b"0000000000000000_0000000000000000_0000100111001011_1101001110010111"; -- 0.03826639596330596
	pesos_i(13148) := b"1111111111111111_1111111111111111_1111011000011001_1111110010100010"; -- -0.03866597217953084
	pesos_i(13149) := b"1111111111111111_1111111111111111_1111011011101010_1110110111001000"; -- -0.03547777038245357
	pesos_i(13150) := b"0000000000000000_0000000000000000_0010010010101111_1000011111101010"; -- 0.1433033892412765
	pesos_i(13151) := b"0000000000000000_0000000000000000_0010001011001100_0110011000110000"; -- 0.13593138372987792
	pesos_i(13152) := b"0000000000000000_0000000000000000_0010001100000010_1010110011111111"; -- 0.13675957894676435
	pesos_i(13153) := b"1111111111111111_1111111111111111_1111110100000111_1110010010110101"; -- -0.011598306572300406
	pesos_i(13154) := b"1111111111111111_1111111111111111_1110001100100001_0101101111010100"; -- -0.11277223656688633
	pesos_i(13155) := b"1111111111111111_1111111111111111_1110111100010000_0101001011111111"; -- -0.06615716245943494
	pesos_i(13156) := b"0000000000000000_0000000000000000_0001010011011100_0100001111110101"; -- 0.08148598405532119
	pesos_i(13157) := b"1111111111111111_1111111111111111_1110001001110010_0111111111011111"; -- -0.11544037639056347
	pesos_i(13158) := b"1111111111111111_1111111111111111_1110101011110100_1110111110101000"; -- -0.08220007082421472
	pesos_i(13159) := b"1111111111111111_1111111111111111_1111001001111110_1000000111100001"; -- -0.05275715126535808
	pesos_i(13160) := b"1111111111111111_1111111111111111_1110010111000000_1001011101000110"; -- -0.10253004585198197
	pesos_i(13161) := b"1111111111111111_1111111111111111_1110110001100110_0101101010101000"; -- -0.07656320006964688
	pesos_i(13162) := b"0000000000000000_0000000000000000_0000101101010100_1100110110111010"; -- 0.04426275046330167
	pesos_i(13163) := b"1111111111111111_1111111111111111_1110011000100011_0100111111010100"; -- -0.1010236841563139
	pesos_i(13164) := b"0000000000000000_0000000000000000_0010000011001110_0100011000011001"; -- 0.12814748880717355
	pesos_i(13165) := b"1111111111111111_1111111111111111_1110010111001100_1110010010000001"; -- -0.10234233702437917
	pesos_i(13166) := b"0000000000000000_0000000000000000_0010101010011111_1011011100111000"; -- 0.16649956804686145
	pesos_i(13167) := b"0000000000000000_0000000000000000_0010001110101000_1011101100010011"; -- 0.13929337710132142
	pesos_i(13168) := b"1111111111111111_1111111111111111_1101011111110001_0110011011100101"; -- -0.15647274874823436
	pesos_i(13169) := b"0000000000000000_0000000000000000_0000101011111010_1111011000111000"; -- 0.04289187310887525
	pesos_i(13170) := b"0000000000000000_0000000000000000_0000010010000100_0100100011000100"; -- 0.01764349733084686
	pesos_i(13171) := b"1111111111111111_1111111111111111_1111011100101011_0100000000110100"; -- -0.03449629518019725
	pesos_i(13172) := b"0000000000000000_0000000000000000_0000011101000110_0110001011011111"; -- 0.028417758373733143
	pesos_i(13173) := b"0000000000000000_0000000000000000_0000100110111111_0001000010011010"; -- 0.03807166818546997
	pesos_i(13174) := b"1111111111111111_1111111111111111_1110101111110101_0100101010000111"; -- -0.07828840448589391
	pesos_i(13175) := b"0000000000000000_0000000000000000_0010000010110000_1001001000110001"; -- 0.12769426045886761
	pesos_i(13176) := b"0000000000000000_0000000000000000_0000011011000011_0011111011110001"; -- 0.02641671547067931
	pesos_i(13177) := b"1111111111111111_1111111111111111_1111011100000111_0111001000011111"; -- -0.03504263639532141
	pesos_i(13178) := b"0000000000000000_0000000000000000_0001100010100000_0010001110101100"; -- 0.09619353251768752
	pesos_i(13179) := b"0000000000000000_0000000000000000_0000010111110111_1000100011100110"; -- 0.023308330628807158
	pesos_i(13180) := b"1111111111111111_1111111111111111_1111000000010011_0101100100011011"; -- -0.06220477200583712
	pesos_i(13181) := b"1111111111111111_1111111111111111_1111100101000010_0000110110011110"; -- -0.02633585838475247
	pesos_i(13182) := b"1111111111111111_1111111111111111_1110111000100000_1110001101111110"; -- -0.06981065913761812
	pesos_i(13183) := b"0000000000000000_0000000000000000_0001110010110101_1010111000110101"; -- 0.1121472244707769
	pesos_i(13184) := b"1111111111111111_1111111111111111_1111100101101110_0101011100011110"; -- -0.02566009052317405
	pesos_i(13185) := b"0000000000000000_0000000000000000_0001011100010000_0111010010000010"; -- 0.09009483499126945
	pesos_i(13186) := b"1111111111111111_1111111111111111_1110101001100111_0111110110111111"; -- -0.08435834963143402
	pesos_i(13187) := b"0000000000000000_0000000000000000_0010000000000010_0011111000110101"; -- 0.12503422534734057
	pesos_i(13188) := b"1111111111111111_1111111111111111_1101111111000100_0010110001000111"; -- -0.12591288826377303
	pesos_i(13189) := b"1111111111111111_1111111111111111_1111100011110011_1000111100100011"; -- -0.02753358264607086
	pesos_i(13190) := b"1111111111111111_1111111111111111_1111001011000111_1101011001111001"; -- -0.0516382175056086
	pesos_i(13191) := b"1111111111111111_1111111111111111_1110000101011100_1010010000110100"; -- -0.11968015413786098
	pesos_i(13192) := b"1111111111111111_1111111111111111_1110001110000001_0000010110000000"; -- -0.11131253831482203
	pesos_i(13193) := b"1111111111111111_1111111111111111_1111010110100110_1001101011111111"; -- -0.04042655259585527
	pesos_i(13194) := b"0000000000000000_0000000000000000_0000000001111011_1101011010101000"; -- 0.0018896254612928071
	pesos_i(13195) := b"0000000000000000_0000000000000000_0001100100010110_1110000010100111"; -- 0.09800533374671774
	pesos_i(13196) := b"1111111111111111_1111111111111111_1101110100001111_1110110010000011"; -- -0.13647577087943316
	pesos_i(13197) := b"0000000000000000_0000000000000000_0010001101110110_0010010011010110"; -- 0.13852148261328034
	pesos_i(13198) := b"1111111111111111_1111111111111111_1111010100100111_1100100010001010"; -- -0.0423617040944343
	pesos_i(13199) := b"1111111111111111_1111111111111111_1101111110011000_0111011010101110"; -- -0.12657984016186752
	pesos_i(13200) := b"1111111111111111_1111111111111111_1110101010011001_0000011000000011"; -- -0.08360254689327289
	pesos_i(13201) := b"1111111111111111_1111111111111111_1110101011010000_1001000100110001"; -- -0.08275501790313346
	pesos_i(13202) := b"1111111111111111_1111111111111111_1110000111110101_0001111000101111"; -- -0.11735354749468238
	pesos_i(13203) := b"0000000000000000_0000000000000000_0000101010101011_1100001111001011"; -- 0.041683423029073255
	pesos_i(13204) := b"1111111111111111_1111111111111111_1110010010001011_0011010110001111"; -- -0.10725083593942562
	pesos_i(13205) := b"1111111111111111_1111111111111111_1110011001100100_0001000111111111"; -- -0.10003554838181425
	pesos_i(13206) := b"1111111111111111_1111111111111111_1111000011101110_0100000000001101"; -- -0.05886459054445797
	pesos_i(13207) := b"1111111111111111_1111111111111111_1111110000110111_1011011000110100"; -- -0.014774906384431923
	pesos_i(13208) := b"1111111111111111_1111111111111111_1111010001100000_1010101110011001"; -- -0.0453999283380931
	pesos_i(13209) := b"1111111111111111_1111111111111111_1110100000001010_1100000000000011"; -- -0.0935859672498483
	pesos_i(13210) := b"1111111111111111_1111111111111111_1111010011001101_0111101110001011"; -- -0.04373958441957653
	pesos_i(13211) := b"0000000000000000_0000000000000000_0010001011110111_1001101000010011"; -- 0.13659060433453596
	pesos_i(13212) := b"0000000000000000_0000000000000000_0001011000101010_1100000010010011"; -- 0.08658984753178967
	pesos_i(13213) := b"1111111111111111_1111111111111111_1101100100001110_0000001100011101"; -- -0.15212994145789116
	pesos_i(13214) := b"0000000000000000_0000000000000000_0010010100110111_0001100010000001"; -- 0.14537194404265172
	pesos_i(13215) := b"0000000000000000_0000000000000000_0000001110111111_1001010011011101"; -- 0.014642051721713574
	pesos_i(13216) := b"1111111111111111_1111111111111111_1110011010101111_1110010010100110"; -- -0.09887858330951282
	pesos_i(13217) := b"1111111111111111_1111111111111111_1110111101111100_0100001000111000"; -- -0.06451021312697834
	pesos_i(13218) := b"0000000000000000_0000000000000000_0000001001110010_0111100010110100"; -- 0.009559196435320608
	pesos_i(13219) := b"1111111111111111_1111111111111111_1101111111010110_0010010001011000"; -- -0.12563870287182025
	pesos_i(13220) := b"0000000000000000_0000000000000000_0000011100001010_1010000100101111"; -- 0.027505945099956512
	pesos_i(13221) := b"1111111111111111_1111111111111111_1110001000000001_0101000011011010"; -- -0.11716742202039611
	pesos_i(13222) := b"1111111111111111_1111111111111111_1110001110100000_0001011000100110"; -- -0.11083852369249758
	pesos_i(13223) := b"1111111111111111_1111111111111111_1110011011101011_1111110101100001"; -- -0.0979615820838639
	pesos_i(13224) := b"1111111111111111_1111111111111111_1111100100000110_1110011011010011"; -- -0.02723843902194417
	pesos_i(13225) := b"0000000000000000_0000000000000000_0001010010110011_0101011101111101"; -- 0.08086153794233111
	pesos_i(13226) := b"1111111111111111_1111111111111111_1110110101100101_0010001010111010"; -- -0.07267554234463953
	pesos_i(13227) := b"0000000000000000_0000000000000000_0001110000000100_0101010011101101"; -- 0.10944109715403352
	pesos_i(13228) := b"1111111111111111_1111111111111111_1110010111100010_0011100100010000"; -- -0.1020168625684894
	pesos_i(13229) := b"0000000000000000_0000000000000000_0000000101101100_1011010000110100"; -- 0.005564940088273399
	pesos_i(13230) := b"0000000000000000_0000000000000000_0001111011110100_0101000101011000"; -- 0.12091549289833402
	pesos_i(13231) := b"1111111111111111_1111111111111111_1101100000010111_0001111111001011"; -- -0.15589715292092698
	pesos_i(13232) := b"1111111111111111_1111111111111111_1111011101110011_1100111110000001"; -- -0.03338912100679376
	pesos_i(13233) := b"1111111111111111_1111111111111111_1111001111100101_0110111100101110"; -- -0.047280360573375146
	pesos_i(13234) := b"0000000000000000_0000000000000000_0010000101100010_0011110011011111"; -- 0.1304052396286619
	pesos_i(13235) := b"1111111111111111_1111111111111111_1111101001101010_1101010111001001"; -- -0.02180732587687993
	pesos_i(13236) := b"0000000000000000_0000000000000000_0001011001100100_0110101001000101"; -- 0.0874697131121057
	pesos_i(13237) := b"0000000000000000_0000000000000000_0010010001000011_1110110101110111"; -- 0.14166149298096978
	pesos_i(13238) := b"0000000000000000_0000000000000000_0010100101011010_0010101110000110"; -- 0.16153213527602375
	pesos_i(13239) := b"1111111111111111_1111111111111111_1101110001111100_1110011011111001"; -- -0.13871914320910875
	pesos_i(13240) := b"1111111111111111_1111111111111111_1111101010000110_1011000111110001"; -- -0.021382216211052452
	pesos_i(13241) := b"1111111111111111_1111111111111111_1110001011111011_0101101001111101"; -- -0.11335215041087311
	pesos_i(13242) := b"0000000000000000_0000000000000000_0001000111010100_1110011010111101"; -- 0.06965486634606559
	pesos_i(13243) := b"1111111111111111_1111111111111111_1101111110111110_0101001001011011"; -- -0.12600217142027892
	pesos_i(13244) := b"1111111111111111_1111111111111111_1110101111111110_0101000101101101"; -- -0.07815066431672747
	pesos_i(13245) := b"1111111111111111_1111111111111111_1110000001110000_0110000110000001"; -- -0.1232852040414269
	pesos_i(13246) := b"1111111111111111_1111111111111111_1110100011100001_0011101001001001"; -- -0.09031329835430053
	pesos_i(13247) := b"1111111111111111_1111111111111111_1110101010000110_1010110000000100"; -- -0.08388256934503066
	pesos_i(13248) := b"1111111111111111_1111111111111111_1101111010010010_0000110111100110"; -- -0.13058388839297333
	pesos_i(13249) := b"0000000000000000_0000000000000000_0001111010011101_0000011011011010"; -- 0.11958353826416879
	pesos_i(13250) := b"1111111111111111_1111111111111111_1110111111000100_0001101110011001"; -- -0.06341388238650182
	pesos_i(13251) := b"1111111111111111_1111111111111111_1111101011111010_0000011100100111"; -- -0.019622376495533025
	pesos_i(13252) := b"0000000000000000_0000000000000000_0001010011110110_0110000010111001"; -- 0.08188442723577846
	pesos_i(13253) := b"0000000000000000_0000000000000000_0000110010001110_1101010001010010"; -- 0.04905440329043747
	pesos_i(13254) := b"0000000000000000_0000000000000000_0001100010000001_0011011100100101"; -- 0.09572167058111518
	pesos_i(13255) := b"0000000000000000_0000000000000000_0001100111100101_1000100110000101"; -- 0.10115870940224476
	pesos_i(13256) := b"1111111111111111_1111111111111111_1111011011001110_1101111110111000"; -- -0.035905854811722066
	pesos_i(13257) := b"1111111111111111_1111111111111111_1101101000000110_1010101101011100"; -- -0.148335733361973
	pesos_i(13258) := b"1111111111111111_1111111111111111_1111001101101111_0011111101100011"; -- -0.049083746214068094
	pesos_i(13259) := b"0000000000000000_0000000000000000_0001111011000010_1001001101011111"; -- 0.12015648904449154
	pesos_i(13260) := b"0000000000000000_0000000000000000_0001111110001100_1101011101100010"; -- 0.12324281821019323
	pesos_i(13261) := b"0000000000000000_0000000000000000_0010010001101000_1000001100111110"; -- 0.14221973680074665
	pesos_i(13262) := b"0000000000000000_0000000000000000_0001000111110011_1111101000100110"; -- 0.07012904570180974
	pesos_i(13263) := b"1111111111111111_1111111111111111_1101110100011001_1010011000100100"; -- -0.13632737760773847
	pesos_i(13264) := b"1111111111111111_1111111111111111_1101111111101001_1101100100110010"; -- -0.12533800635300754
	pesos_i(13265) := b"1111111111111111_1111111111111111_1111001110001010_1011011111111000"; -- -0.04866457169246839
	pesos_i(13266) := b"1111111111111111_1111111111111111_1111101011010001_1111001101001011"; -- -0.020233911613708785
	pesos_i(13267) := b"0000000000000000_0000000000000000_0010000000110111_1100001001100011"; -- 0.1258508196550381
	pesos_i(13268) := b"0000000000000000_0000000000000000_0001100101111011_0001011011001011"; -- 0.09953443966672594
	pesos_i(13269) := b"1111111111111111_1111111111111111_1110001000000011_0000001111011101"; -- -0.11714149331518624
	pesos_i(13270) := b"0000000000000000_0000000000000000_0000011010011100_1010101111100010"; -- 0.0258281161910485
	pesos_i(13271) := b"0000000000000000_0000000000000000_0001101110101101_0101010110101000"; -- 0.10811362598261942
	pesos_i(13272) := b"1111111111111111_1111111111111111_1110011100100010_0011001101000010"; -- -0.09713439587876131
	pesos_i(13273) := b"1111111111111111_1111111111111111_1101011110000110_1111110110111110"; -- -0.1580964480735825
	pesos_i(13274) := b"0000000000000000_0000000000000000_0000001001111101_1011111001011011"; -- 0.009731194793664157
	pesos_i(13275) := b"0000000000000000_0000000000000000_0010011011111000_1111110011011000"; -- 0.15223675024084216
	pesos_i(13276) := b"0000000000000000_0000000000000000_0000110001001110_1001101111101110"; -- 0.04807447959893115
	pesos_i(13277) := b"1111111111111111_1111111111111111_1111101100111010_0100001000100110"; -- -0.018642297475311934
	pesos_i(13278) := b"0000000000000000_0000000000000000_0000010110100001_1001011111101111"; -- 0.021996970968593592
	pesos_i(13279) := b"0000000000000000_0000000000000000_0000010110010110_1010010011000100"; -- 0.02182988908345234
	pesos_i(13280) := b"1111111111111111_1111111111111111_1110001111010101_1111101001101111"; -- -0.11001620086749402
	pesos_i(13281) := b"0000000000000000_0000000000000000_0000001111101001_1101001110111000"; -- 0.01528666728533008
	pesos_i(13282) := b"1111111111111111_1111111111111111_1110110001010110_1001000100011011"; -- -0.07680409527074941
	pesos_i(13283) := b"0000000000000000_0000000000000000_0001100001000101_1111100100110010"; -- 0.09481770959410658
	pesos_i(13284) := b"1111111111111111_1111111111111111_1101111000001001_0011000000101001"; -- -0.13267230028550606
	pesos_i(13285) := b"0000000000000000_0000000000000000_0000000111011111_1111000101111010"; -- 0.007323353076958361
	pesos_i(13286) := b"0000000000000000_0000000000000000_0000010100001000_1010110110100001"; -- 0.019663669364640493
	pesos_i(13287) := b"0000000000000000_0000000000000000_0001011100110100_1010000101111110"; -- 0.09064683282101482
	pesos_i(13288) := b"0000000000000000_0000000000000000_0000110000000110_0110111010100111"; -- 0.04697314815154211
	pesos_i(13289) := b"0000000000000000_0000000000000000_0001001011110111_0010111011011001"; -- 0.0740842132841951
	pesos_i(13290) := b"1111111111111111_1111111111111111_1110001101110011_0001001001110111"; -- -0.11152538860490488
	pesos_i(13291) := b"1111111111111111_1111111111111111_1111101100100001_1010110101100110"; -- -0.01901737463329222
	pesos_i(13292) := b"1111111111111111_1111111111111111_1110001111101001_0000110100110111"; -- -0.10972516438960643
	pesos_i(13293) := b"1111111111111111_1111111111111111_1101110110010100_1111001011111110"; -- -0.13444596580454016
	pesos_i(13294) := b"0000000000000000_0000000000000000_0000110110101110_0100101010111101"; -- 0.05344073402549289
	pesos_i(13295) := b"0000000000000000_0000000000000000_0001011010101011_1000100000101001"; -- 0.08855486879439449
	pesos_i(13296) := b"0000000000000000_0000000000000000_0000101000101011_1001111101110100"; -- 0.03972813201069545
	pesos_i(13297) := b"0000000000000000_0000000000000000_0001101100111101_1010101000011111"; -- 0.10640967623694968
	pesos_i(13298) := b"1111111111111111_1111111111111111_1101110100010100_0111101010101011"; -- -0.136406262578916
	pesos_i(13299) := b"0000000000000000_0000000000000000_0001111001011001_1101111010010011"; -- 0.11855879877957179
	pesos_i(13300) := b"0000000000000000_0000000000000000_0001101011110010_0101000011010101"; -- 0.10525994482752724
	pesos_i(13301) := b"1111111111111111_1111111111111111_1110111000110110_0011101110011101"; -- -0.06948497218853521
	pesos_i(13302) := b"1111111111111111_1111111111111111_1110101001110110_1011011100110000"; -- -0.08412604406334352
	pesos_i(13303) := b"0000000000000000_0000000000000000_0000000011011110_0110100101001100"; -- 0.003393727309457086
	pesos_i(13304) := b"0000000000000000_0000000000000000_0010000101001011_1101110100111110"; -- 0.13006384615361608
	pesos_i(13305) := b"0000000000000000_0000000000000000_0000001110001010_0101110011011101"; -- 0.013829997882106638
	pesos_i(13306) := b"1111111111111111_1111111111111111_1111010111110101_1001011000110010"; -- -0.03922139434249548
	pesos_i(13307) := b"1111111111111111_1111111111111111_1111010110100011_1111000010101011"; -- -0.04046722247294726
	pesos_i(13308) := b"0000000000000000_0000000000000000_0001101000010011_0101111011010110"; -- 0.10185806962943657
	pesos_i(13309) := b"1111111111111111_1111111111111111_1111100110100010_0011101011010101"; -- -0.024868319595055203
	pesos_i(13310) := b"1111111111111111_1111111111111111_1110011101010100_0100011111001001"; -- -0.09637023300053542
	pesos_i(13311) := b"0000000000000000_0000000000000000_0001010111100110_0111000110110010"; -- 0.08554754826194776
	pesos_i(13312) := b"1111111111111111_1111111111111111_1110000100011010_0001111001011100"; -- -0.1206952119180925
	pesos_i(13313) := b"0000000000000000_0000000000000000_0000100110111101_1001001101110001"; -- 0.038048949363579776
	pesos_i(13314) := b"1111111111111111_1111111111111111_1101111110110101_1000100101011111"; -- -0.12613622115848117
	pesos_i(13315) := b"1111111111111111_1111111111111111_1110011001100000_0010101010001011"; -- -0.1000951204711049
	pesos_i(13316) := b"0000000000000000_0000000000000000_0001100001010000_1000111001111100"; -- 0.09497919587305577
	pesos_i(13317) := b"1111111111111111_1111111111111111_1110011011111010_1011010110101100"; -- -0.09773697419005284
	pesos_i(13318) := b"0000000000000000_0000000000000000_0001110011011110_1110100000100111"; -- 0.11277628849922734
	pesos_i(13319) := b"0000000000000000_0000000000000000_0001010111010100_1100001011101111"; -- 0.08527773222056932
	pesos_i(13320) := b"1111111111111111_1111111111111111_1111000100001011_0011110001101001"; -- -0.058422302643589774
	pesos_i(13321) := b"0000000000000000_0000000000000000_0001111011110000_0001111000111110"; -- 0.12085141185455468
	pesos_i(13322) := b"1111111111111111_1111111111111111_1110100001101000_0000101001110111"; -- -0.0921624621771236
	pesos_i(13323) := b"1111111111111111_1111111111111111_1111000111001001_0101100101100100"; -- -0.0555214052562215
	pesos_i(13324) := b"1111111111111111_1111111111111111_1110010111111101_1100010001111010"; -- -0.10159656556247999
	pesos_i(13325) := b"1111111111111111_1111111111111111_1111100010100111_1101111011010110"; -- -0.02868850025731335
	pesos_i(13326) := b"1111111111111111_1111111111111111_1101111111100001_0110100110011100"; -- -0.12546672770774756
	pesos_i(13327) := b"0000000000000000_0000000000000000_0001110011001100_0110111111101111"; -- 0.11249446471283876
	pesos_i(13328) := b"0000000000000000_0000000000000000_0001101100101010_0101000111111101"; -- 0.10611450597310418
	pesos_i(13329) := b"0000000000000000_0000000000000000_0000110110111100_1001110001111110"; -- 0.05365922994398691
	pesos_i(13330) := b"1111111111111111_1111111111111111_1101100101111110_1110010010111000"; -- -0.15040750991374954
	pesos_i(13331) := b"0000000000000000_0000000000000000_0010001000100100_1011000000011110"; -- 0.13337231385255274
	pesos_i(13332) := b"1111111111111111_1111111111111111_1111001101010000_1100110000100101"; -- -0.04954837880573538
	pesos_i(13333) := b"0000000000000000_0000000000000000_0000010111110101_1101000100110100"; -- 0.023282122706090855
	pesos_i(13334) := b"1111111111111111_1111111111111111_1111110001000010_1110100010001100"; -- -0.014604058995364677
	pesos_i(13335) := b"1111111111111111_1111111111111111_1111010001010000_0010001101010011"; -- -0.04565219143762304
	pesos_i(13336) := b"0000000000000000_0000000000000000_0000101001101110_0001111110101000"; -- 0.04074285363787703
	pesos_i(13337) := b"0000000000000000_0000000000000000_0001110100111110_0010011110011011"; -- 0.11422965570503081
	pesos_i(13338) := b"1111111111111111_1111111111111111_1111010101010111_1000111011100010"; -- -0.041632718941918286
	pesos_i(13339) := b"1111111111111111_1111111111111111_1101111000011101_0011010101011000"; -- -0.13236681551644255
	pesos_i(13340) := b"0000000000000000_0000000000000000_0000110010110100_0000010111010010"; -- 0.049621928927550234
	pesos_i(13341) := b"0000000000000000_0000000000000000_0000100001000101_0100000001001010"; -- 0.03230668839766703
	pesos_i(13342) := b"0000000000000000_0000000000000000_0000101101110011_0000111011111111"; -- 0.044724404621746316
	pesos_i(13343) := b"1111111111111111_1111111111111111_1110010001000011_1110010000100010"; -- -0.10833906343034967
	pesos_i(13344) := b"0000000000000000_0000000000000000_0010000000101011_1010000110000011"; -- 0.12566575487469023
	pesos_i(13345) := b"0000000000000000_0000000000000000_0001000100011001_1111101111001100"; -- 0.06680272798265481
	pesos_i(13346) := b"0000000000000000_0000000000000000_0010001100110110_1100001111101110"; -- 0.13755440295976468
	pesos_i(13347) := b"0000000000000000_0000000000000000_0001100001101000_0110011111110100"; -- 0.09534311010846577
	pesos_i(13348) := b"0000000000000000_0000000000000000_0001010101001011_1101000001001010"; -- 0.08318807416750189
	pesos_i(13349) := b"1111111111111111_1111111111111111_1110011110110010_0000000101011000"; -- -0.0949401054212499
	pesos_i(13350) := b"1111111111111111_1111111111111111_1110100010011111_1000101111011100"; -- -0.09131551620583134
	pesos_i(13351) := b"1111111111111111_1111111111111111_1110111000110011_1011111110111110"; -- -0.06952287301247263
	pesos_i(13352) := b"0000000000000000_0000000000000000_0001011111111000_0000111110111100"; -- 0.09362886751240296
	pesos_i(13353) := b"1111111111111111_1111111111111111_1111100100000110_1010100110001011"; -- -0.02724209171836372
	pesos_i(13354) := b"0000000000000000_0000000000000000_0000001000011100_1011101111111110"; -- 0.008250951240009814
	pesos_i(13355) := b"0000000000000000_0000000000000000_0000100111100100_1111100010101101"; -- 0.03865007610767062
	pesos_i(13356) := b"0000000000000000_0000000000000000_0001011001101110_1011001101110001"; -- 0.08762666229946804
	pesos_i(13357) := b"0000000000000000_0000000000000000_0001111001101001_1101000011011101"; -- 0.11880212202382673
	pesos_i(13358) := b"1111111111111111_1111111111111111_1111000110011110_0111111110011011"; -- -0.056175255481499924
	pesos_i(13359) := b"0000000000000000_0000000000000000_0000010101001011_0110110001011001"; -- 0.020682117310444587
	pesos_i(13360) := b"1111111111111111_1111111111111111_1110010000101100_1111101011111101"; -- -0.10868865315317093
	pesos_i(13361) := b"1111111111111111_1111111111111111_1111100101000011_0110011111001010"; -- -0.026315224852724094
	pesos_i(13362) := b"1111111111111111_1111111111111111_1110100000011010_0111100111100110"; -- -0.09334600580324896
	pesos_i(13363) := b"1111111111111111_1111111111111111_1101111100111000_0010001100101111"; -- -0.12804966082074776
	pesos_i(13364) := b"0000000000000000_0000000000000000_0001110100010001_0110011000111101"; -- 0.11354674322496305
	pesos_i(13365) := b"0000000000000000_0000000000000000_0001010110111001_0110000101100111"; -- 0.08485993149256128
	pesos_i(13366) := b"0000000000000000_0000000000000000_0001010011101001_0111011001111101"; -- 0.08168736035289681
	pesos_i(13367) := b"0000000000000000_0000000000000000_0001111110100110_1011110110110001"; -- 0.1236380154146335
	pesos_i(13368) := b"1111111111111111_1111111111111111_1110010011011101_1010000011000100"; -- -0.10599322523542146
	pesos_i(13369) := b"1111111111111111_1111111111111111_1101101001001010_0000110010100111"; -- -0.14730759549092057
	pesos_i(13370) := b"0000000000000000_0000000000000000_0000100001001010_1101101101001001"; -- 0.03239222073091016
	pesos_i(13371) := b"0000000000000000_0000000000000000_0001110001011001_1100000111001110"; -- 0.1107445838720997
	pesos_i(13372) := b"0000000000000000_0000000000000000_0000111011011111_0000100111110000"; -- 0.058090802301189515
	pesos_i(13373) := b"0000000000000000_0000000000000000_0000110101010100_0101101101001000"; -- 0.05206842917144267
	pesos_i(13374) := b"0000000000000000_0000000000000000_0000001111101001_0111100000000110"; -- 0.015281201694198355
	pesos_i(13375) := b"0000000000000000_0000000000000000_0000110000000010_1100011000001110"; -- 0.04691732248052116
	pesos_i(13376) := b"1111111111111111_1111111111111111_1111001111001100_0011011000110100"; -- -0.04766522624360177
	pesos_i(13377) := b"1111111111111111_1111111111111111_1110111010101111_1001110001001110"; -- -0.0676328953495919
	pesos_i(13378) := b"0000000000000000_0000000000000000_0001001101111100_0101110000100001"; -- 0.07611633107768284
	pesos_i(13379) := b"1111111111111111_1111111111111111_1111101111111001_1111100101011010"; -- -0.01571694890230132
	pesos_i(13380) := b"0000000000000000_0000000000000000_0001000101001011_1000111111011001"; -- 0.06755923315837341
	pesos_i(13381) := b"0000000000000000_0000000000000000_0000110110110100_0110101101001010"; -- 0.05353422688343793
	pesos_i(13382) := b"1111111111111111_1111111111111111_1110011101110100_0000000001101101"; -- -0.09588620518898491
	pesos_i(13383) := b"0000000000000000_0000000000000000_0001100111110001_0101000110000101"; -- 0.10133847703067747
	pesos_i(13384) := b"0000000000000000_0000000000000000_0001111001110011_1111100011010101"; -- 0.11895709218918422
	pesos_i(13385) := b"1111111111111111_1111111111111111_1110111000000100_1110110111001110"; -- -0.07023729048745192
	pesos_i(13386) := b"1111111111111111_1111111111111111_1101110000000100_1110001110010101"; -- -0.140550399831326
	pesos_i(13387) := b"0000000000000000_0000000000000000_0000100100101111_0100101000101010"; -- 0.0358778335983819
	pesos_i(13388) := b"0000000000000000_0000000000000000_0001110010001001_0000001011101001"; -- 0.11146562753980677
	pesos_i(13389) := b"1111111111111111_1111111111111111_1101100100111001_1001100011000101"; -- -0.15146489330417193
	pesos_i(13390) := b"0000000000000000_0000000000000000_0001001011011000_1000110011001000"; -- 0.07361678972575635
	pesos_i(13391) := b"0000000000000000_0000000000000000_0001001101011101_1001011110010110"; -- 0.07564685252479257
	pesos_i(13392) := b"1111111111111111_1111111111111111_1110110101110011_0110111000100111"; -- -0.07245742359685003
	pesos_i(13393) := b"1111111111111111_1111111111111111_1110101011001101_1110101100111101"; -- -0.08279542698574453
	pesos_i(13394) := b"0000000000000000_0000000000000000_0000011000110001_1010001111000111"; -- 0.024194942530816457
	pesos_i(13395) := b"0000000000000000_0000000000000000_0001110110111011_1011001010100111"; -- 0.11614529194941425
	pesos_i(13396) := b"1111111111111111_1111111111111111_1111000000111101_1101110111101101"; -- -0.06155598596547955
	pesos_i(13397) := b"0000000000000000_0000000000000000_0001010110001100_1001010011101111"; -- 0.0841763577124809
	pesos_i(13398) := b"0000000000000000_0000000000000000_0001001101111011_1100111110001110"; -- 0.07610795229705973
	pesos_i(13399) := b"1111111111111111_1111111111111111_1111100001001011_0010000011010010"; -- -0.030103634546111886
	pesos_i(13400) := b"1111111111111111_1111111111111111_1110011101111000_1000101111010101"; -- -0.09581686076543765
	pesos_i(13401) := b"0000000000000000_0000000000000000_0000011010100010_1011011101101111"; -- 0.025920357378398273
	pesos_i(13402) := b"0000000000000000_0000000000000000_0001000100000000_1000101111100010"; -- 0.06641458768782392
	pesos_i(13403) := b"1111111111111111_1111111111111111_1110001100100001_0110110101100010"; -- -0.11277119020665516
	pesos_i(13404) := b"0000000000000000_0000000000000000_0000000100000000_1100010001101100"; -- 0.003917957625943224
	pesos_i(13405) := b"1111111111111111_1111111111111111_1110011110010101_0000010000000111"; -- -0.0953824503036837
	pesos_i(13406) := b"1111111111111111_1111111111111111_1111011100011000_0111001010011000"; -- -0.034783208767384055
	pesos_i(13407) := b"1111111111111111_1111111111111111_1110110011111110_0010001011001111"; -- -0.0742471927727091
	pesos_i(13408) := b"1111111111111111_1111111111111111_1111110001000101_0101011100001010"; -- -0.01456695557952826
	pesos_i(13409) := b"0000000000000000_0000000000000000_0000011111001110_1010111000011100"; -- 0.030497438210062774
	pesos_i(13410) := b"1111111111111111_1111111111111111_1111100011111010_1011101100110011"; -- -0.027424144865287457
	pesos_i(13411) := b"1111111111111111_1111111111111111_1110111010000111_0111100110111001"; -- -0.06824530817141364
	pesos_i(13412) := b"1111111111111111_1111111111111111_1111000000110111_1101000000010011"; -- -0.061648364443327164
	pesos_i(13413) := b"1111111111111111_1111111111111111_1110010000011001_0011101111001111"; -- -0.10898996548443757
	pesos_i(13414) := b"0000000000000000_0000000000000000_0000110011001100_0110111111110101"; -- 0.04999446621631721
	pesos_i(13415) := b"0000000000000000_0000000000000000_0001000011110110_0010110101001111"; -- 0.06625636261844117
	pesos_i(13416) := b"1111111111111111_1111111111111111_1111001001000011_0111101100010010"; -- -0.05365782551932106
	pesos_i(13417) := b"0000000000000000_0000000000000000_0001101100010001_1100000111101111"; -- 0.10573970864826368
	pesos_i(13418) := b"0000000000000000_0000000000000000_0001110000001100_1110011000100010"; -- 0.10957182238446057
	pesos_i(13419) := b"1111111111111111_1111111111111111_1110001100111111_1100010101000011"; -- -0.11230818858971163
	pesos_i(13420) := b"1111111111111111_1111111111111111_1110100111101001_0001011000010011"; -- -0.08628713645925366
	pesos_i(13421) := b"1111111111111111_1111111111111111_1101110101110110_0001101110111000"; -- -0.13491656070171348
	pesos_i(13422) := b"1111111111111111_1111111111111111_1110001000110000_1101011110110010"; -- -0.1164422216546361
	pesos_i(13423) := b"1111111111111111_1111111111111111_1111110001000000_0100111001111100"; -- -0.01464375942882413
	pesos_i(13424) := b"1111111111111111_1111111111111111_1110110001111000_1101001110101011"; -- -0.07628132891552118
	pesos_i(13425) := b"0000000000000000_0000000000000000_0001110111101110_0011001111001010"; -- 0.11691592861174144
	pesos_i(13426) := b"0000000000000000_0000000000000000_0000101000001110_0100010100101011"; -- 0.039280245689220464
	pesos_i(13427) := b"0000000000000000_0000000000000000_0001101110011011_1100100110011100"; -- 0.10784587924079413
	pesos_i(13428) := b"0000000000000000_0000000000000000_0010000110000000_1010001011011101"; -- 0.1308690823657009
	pesos_i(13429) := b"0000000000000000_0000000000000000_0000101010100101_1000101011111110"; -- 0.041588484685801966
	pesos_i(13430) := b"1111111111111111_1111111111111111_1110001110111011_1110000100110101"; -- -0.11041443306476141
	pesos_i(13431) := b"1111111111111111_1111111111111111_1110001001000011_1010010000000110"; -- -0.11615538448148253
	pesos_i(13432) := b"0000000000000000_0000000000000000_0010001000011010_1000011110001011"; -- 0.133217307565836
	pesos_i(13433) := b"1111111111111111_1111111111111111_1110011000100111_1100000011110001"; -- -0.10095590700189735
	pesos_i(13434) := b"0000000000000000_0000000000000000_0001101110011010_1110011011000100"; -- 0.1078323581160313
	pesos_i(13435) := b"1111111111111111_1111111111111111_1110000100010100_0100101100010101"; -- -0.12078409893954252
	pesos_i(13436) := b"1111111111111111_1111111111111111_1110100011000011_1011001000011001"; -- -0.09076392076367462
	pesos_i(13437) := b"1111111111111111_1111111111111111_1111011110010110_0010000101111110"; -- -0.03286543530785228
	pesos_i(13438) := b"0000000000000000_0000000000000000_0001000010011010_1110101100101101"; -- 0.06486387106952594
	pesos_i(13439) := b"1111111111111111_1111111111111111_1101110001010110_0100111101100111"; -- -0.13930801129567266
	pesos_i(13440) := b"0000000000000000_0000000000000000_0000010010011011_0110100100001010"; -- 0.017996373168782415
	pesos_i(13441) := b"0000000000000000_0000000000000000_0010000110000111_1110101101011111"; -- 0.13098021574183993
	pesos_i(13442) := b"0000000000000000_0000000000000000_0000101001100011_0011011011100000"; -- 0.04057639094286441
	pesos_i(13443) := b"0000000000000000_0000000000000000_0000101100000101_0100111001010001"; -- 0.04304971190111272
	pesos_i(13444) := b"1111111111111111_1111111111111111_1110110110111001_0000001000110010"; -- -0.0713957430731959
	pesos_i(13445) := b"1111111111111111_1111111111111111_1111101000110011_0111011010001100"; -- -0.02265223572161076
	pesos_i(13446) := b"0000000000000000_0000000000000000_0001010010110000_1001101001000100"; -- 0.08081974175717865
	pesos_i(13447) := b"0000000000000000_0000000000000000_0010011100101001_0011011001000111"; -- 0.1529725956176205
	pesos_i(13448) := b"0000000000000000_0000000000000000_0001001110110000_1111111001100111"; -- 0.07691946041134369
	pesos_i(13449) := b"0000000000000000_0000000000000000_0001011100110011_0111110110010001"; -- 0.09062943265976331
	pesos_i(13450) := b"0000000000000000_0000000000000000_0001111111110011_1110110001000101"; -- 0.12481571847280483
	pesos_i(13451) := b"0000000000000000_0000000000000000_0000100111001001_0011010101100001"; -- 0.03822644818151814
	pesos_i(13452) := b"0000000000000000_0000000000000000_0001001100111001_1110010011000000"; -- 0.07510213561209653
	pesos_i(13453) := b"1111111111111111_1111111111111111_1110000110001101_1010110000011111"; -- -0.1189320015861722
	pesos_i(13454) := b"0000000000000000_0000000000000000_0001101011001110_0111010000010000"; -- 0.10471272833924536
	pesos_i(13455) := b"0000000000000000_0000000000000000_0010011100010101_0110100011001101"; -- 0.15267043123258678
	pesos_i(13456) := b"0000000000000000_0000000000000000_0000101001110100_1000011011001100"; -- 0.04084055393518339
	pesos_i(13457) := b"0000000000000000_0000000000000000_0000011110101001_1100000010000010"; -- 0.029933959773391174
	pesos_i(13458) := b"1111111111111111_1111111111111111_1111010000101110_1101010000100101"; -- -0.04616045090750341
	pesos_i(13459) := b"1111111111111111_1111111111111111_1110110100000001_1000001010010101"; -- -0.0741957080284669
	pesos_i(13460) := b"0000000000000000_0000000000000000_0000110100001100_0000100110110000"; -- 0.05096493286135634
	pesos_i(13461) := b"0000000000000000_0000000000000000_0001000100000110_1000001111000010"; -- 0.06650565608610164
	pesos_i(13462) := b"0000000000000000_0000000000000000_0000010011011000_0110011001011100"; -- 0.018926999426956834
	pesos_i(13463) := b"0000000000000000_0000000000000000_0000110010110100_1110001101110001"; -- 0.049635138534907766
	pesos_i(13464) := b"0000000000000000_0000000000000000_0001111000001110_1100101111101110"; -- 0.11741327821699842
	pesos_i(13465) := b"1111111111111111_1111111111111111_1111100111000101_1011100100001101"; -- -0.024326738646090133
	pesos_i(13466) := b"0000000000000000_0000000000000000_0000010111101001_1000010101001111"; -- 0.023094493724039405
	pesos_i(13467) := b"1111111111111111_1111111111111111_1101111101011001_0101010100001001"; -- -0.12754314933773125
	pesos_i(13468) := b"1111111111111111_1111111111111111_1110101000101010_1010111101011000"; -- -0.08528617966876603
	pesos_i(13469) := b"1111111111111111_1111111111111111_1101110011100101_1000000011001101"; -- -0.13712306028496887
	pesos_i(13470) := b"0000000000000000_0000000000000000_0010001101001111_1100011011101100"; -- 0.13793605095708059
	pesos_i(13471) := b"0000000000000000_0000000000000000_0000110001101001_1011101110110110"; -- 0.04848836123353992
	pesos_i(13472) := b"0000000000000000_0000000000000000_0010011000111001_1100111010111101"; -- 0.14931957343868152
	pesos_i(13473) := b"1111111111111111_1111111111111111_1111001011111001_1000110111001000"; -- -0.05087961079278955
	pesos_i(13474) := b"1111111111111111_1111111111111111_1101101111010110_0110111000101101"; -- -0.14125930210707655
	pesos_i(13475) := b"1111111111111111_1111111111111111_1111011100100101_0001010100011111"; -- -0.03459041590331664
	pesos_i(13476) := b"0000000000000000_0000000000000000_0001000001111111_1011001101101100"; -- 0.06444856060994324
	pesos_i(13477) := b"0000000000000000_0000000000000000_0001101101011010_0110110100000100"; -- 0.10684853874753647
	pesos_i(13478) := b"0000000000000000_0000000000000000_0001100001101111_0110001010000011"; -- 0.0954495973173347
	pesos_i(13479) := b"0000000000000000_0000000000000000_0010000000111001_1011011111001010"; -- 0.12588070569847162
	pesos_i(13480) := b"1111111111111111_1111111111111111_1110110110110011_1000101110010101"; -- -0.07147910706968945
	pesos_i(13481) := b"1111111111111111_1111111111111111_1110001101000100_1101110000000001"; -- -0.11223053912727621
	pesos_i(13482) := b"0000000000000000_0000000000000000_0001011111010010_0000100000110001"; -- 0.09304858394548968
	pesos_i(13483) := b"1111111111111111_1111111111111111_1111011110000101_0010100111111101"; -- -0.03312432836992178
	pesos_i(13484) := b"1111111111111111_1111111111111111_1111000010001101_1110000000011111"; -- -0.06033515209269169
	pesos_i(13485) := b"0000000000000000_0000000000000000_0001010000110101_0000010111001101"; -- 0.07893406146796458
	pesos_i(13486) := b"1111111111111111_1111111111111111_1111110100000001_0000111101000111"; -- -0.011702580718926008
	pesos_i(13487) := b"0000000000000000_0000000000000000_0001011001001101_1010011111001011"; -- 0.08712242794994447
	pesos_i(13488) := b"0000000000000000_0000000000000000_0000101010110011_0010010001111010"; -- 0.04179599743848463
	pesos_i(13489) := b"1111111111111111_1111111111111111_1110001000101100_1001111001001101"; -- -0.11650667774601665
	pesos_i(13490) := b"1111111111111111_1111111111111111_1110001011110000_0001101000100000"; -- -0.113523833507422
	pesos_i(13491) := b"0000000000000000_0000000000000000_0001001011011001_1111100011011110"; -- 0.07363849090656445
	pesos_i(13492) := b"1111111111111111_1111111111111111_1111100010011010_0100000110000001"; -- -0.028896242182895937
	pesos_i(13493) := b"1111111111111111_1111111111111111_1101111111100011_1001011100111010"; -- -0.12543349116623204
	pesos_i(13494) := b"0000000000000000_0000000000000000_0000101110001001_1001111011000011"; -- 0.04506866703677369
	pesos_i(13495) := b"0000000000000000_0000000000000000_0001011110011111_1000111101010110"; -- 0.09227844084206743
	pesos_i(13496) := b"1111111111111111_1111111111111111_1101101101011010_0110101001000010"; -- -0.14315162563949616
	pesos_i(13497) := b"1111111111111111_1111111111111111_1111111010001001_1111111011101100"; -- -0.005706851333559652
	pesos_i(13498) := b"1111111111111111_1111111111111111_1110100101100000_1111011100010010"; -- -0.08836417967774593
	pesos_i(13499) := b"0000000000000000_0000000000000000_0001010101110100_1010010110110111"; -- 0.08381114701958503
	pesos_i(13500) := b"1111111111111111_1111111111111111_1101100001111101_1111010101110000"; -- -0.15432802204556037
	pesos_i(13501) := b"0000000000000000_0000000000000000_0001100110010100_0100010100101101"; -- 0.09991867396850242
	pesos_i(13502) := b"1111111111111111_1111111111111111_1111110111100111_1001011010001111"; -- -0.00818499583744061
	pesos_i(13503) := b"1111111111111111_1111111111111111_1111011100000110_0111001010100101"; -- -0.035057863895384796
	pesos_i(13504) := b"0000000000000000_0000000000000000_0001110011100100_0011100110000000"; -- 0.11285743126206271
	pesos_i(13505) := b"0000000000000000_0000000000000000_0000001110000000_0011010011101011"; -- 0.013675029238856105
	pesos_i(13506) := b"1111111111111111_1111111111111111_1110110011010010_0111100011100111"; -- -0.07491344790322486
	pesos_i(13507) := b"0000000000000000_0000000000000000_0001010001000000_1011011010001111"; -- 0.07911244384004217
	pesos_i(13508) := b"1111111111111111_1111111111111111_1111101001000100_1000011011101100"; -- -0.022391860325042166
	pesos_i(13509) := b"0000000000000000_0000000000000000_0000111000110101_0000010110001110"; -- 0.05549654680621071
	pesos_i(13510) := b"1111111111111111_1111111111111111_1111110101001101_0100101001010000"; -- -0.010539393817357428
	pesos_i(13511) := b"1111111111111111_1111111111111111_1110000001001001_1001000100111010"; -- -0.12387745215446298
	pesos_i(13512) := b"0000000000000000_0000000000000000_0000111100010100_1110101101110011"; -- 0.05891295962091613
	pesos_i(13513) := b"1111111111111111_1111111111111111_1110001101101011_0001110000111001"; -- -0.11164687726304118
	pesos_i(13514) := b"0000000000000000_0000000000000000_0010000001111100_0101101001011110"; -- 0.12689747619142114
	pesos_i(13515) := b"1111111111111111_1111111111111111_1110010100111111_0001110000100110"; -- -0.10450576858592166
	pesos_i(13516) := b"1111111111111111_1111111111111111_1111111011000101_0100010101010111"; -- -0.00480238559929982
	pesos_i(13517) := b"0000000000000000_0000000000000000_0000100110101001_1011101000001111"; -- 0.037746075249574115
	pesos_i(13518) := b"0000000000000000_0000000000000000_0010000010100110_0000100001010011"; -- 0.12753345525193882
	pesos_i(13519) := b"1111111111111111_1111111111111111_1110110010110100_0000111001111010"; -- -0.07537755512841476
	pesos_i(13520) := b"1111111111111111_1111111111111111_1111111000010110_1110110010101010"; -- -0.007462700346907336
	pesos_i(13521) := b"0000000000000000_0000000000000000_0001001100010111_1010110100011011"; -- 0.07458002008144697
	pesos_i(13522) := b"1111111111111111_1111111111111111_1110000010100111_1100100100101011"; -- -0.12243979163539555
	pesos_i(13523) := b"1111111111111111_1111111111111111_1101111000000111_0101001110011000"; -- -0.13270070591069874
	pesos_i(13524) := b"1111111111111111_1111111111111111_1110000100011110_1101100111101110"; -- -0.12062299674898685
	pesos_i(13525) := b"1111111111111111_1111111111111111_1111110101101111_1000000110100010"; -- -0.010017297671146137
	pesos_i(13526) := b"0000000000000000_0000000000000000_0010011001111011_0000001110111000"; -- 0.15031455273301111
	pesos_i(13527) := b"0000000000000000_0000000000000000_0000101111111011_1111000000010011"; -- 0.04681301566143051
	pesos_i(13528) := b"0000000000000000_0000000000000000_0010011000111001_1101111010000001"; -- 0.1493205133577137
	pesos_i(13529) := b"1111111111111111_1111111111111111_1101111001010110_0110100111110011"; -- -0.1314939291386304
	pesos_i(13530) := b"0000000000000000_0000000000000000_0000100101110100_1110111010010000"; -- 0.0369404890094846
	pesos_i(13531) := b"0000000000000000_0000000000000000_0010010110010000_0101000011000001"; -- 0.14673332893770455
	pesos_i(13532) := b"1111111111111111_1111111111111111_1111000110111010_1000111011001111"; -- -0.05574710315308132
	pesos_i(13533) := b"0000000000000000_0000000000000000_0001011000101111_1010001100100101"; -- 0.0866643873489466
	pesos_i(13534) := b"1111111111111111_1111111111111111_1101111111101110_1000111010010000"; -- -0.12526616072974892
	pesos_i(13535) := b"0000000000000000_0000000000000000_0000011101011111_1101110010100101"; -- 0.028806486330118376
	pesos_i(13536) := b"1111111111111111_1111111111111111_1111001101100110_0011110100100010"; -- -0.049221209812435614
	pesos_i(13537) := b"1111111111111111_1111111111111111_1111110011001010_1110100001100100"; -- -0.012528872934042612
	pesos_i(13538) := b"0000000000000000_0000000000000000_0001110100100110_0100101100001100"; -- 0.11386555713778673
	pesos_i(13539) := b"0000000000000000_0000000000000000_0000011000111011_0000010110000110"; -- 0.02433809788137677
	pesos_i(13540) := b"1111111111111111_1111111111111111_1101100110010101_1111011101011100"; -- -0.15005544665719903
	pesos_i(13541) := b"1111111111111111_1111111111111111_1111101010111010_1000100111011111"; -- -0.020591147527946108
	pesos_i(13542) := b"0000000000000000_0000000000000000_0010001001111000_1011001001100000"; -- 0.13465418656565947
	pesos_i(13543) := b"1111111111111111_1111111111111111_1110101101001001_0000000100000000"; -- -0.08091729869907735
	pesos_i(13544) := b"1111111111111111_1111111111111111_1111110101011000_0011000100110100"; -- -0.010373043794467856
	pesos_i(13545) := b"1111111111111111_1111111111111111_1110110000011011_1111000001010100"; -- -0.07769868803010693
	pesos_i(13546) := b"1111111111111111_1111111111111111_1111100101111111_0100101111110011"; -- -0.025401356951478753
	pesos_i(13547) := b"0000000000000000_0000000000000000_0010001110111010_0000111010011100"; -- 0.1395577555579154
	pesos_i(13548) := b"0000000000000000_0000000000000000_0001100000110010_1000101010010101"; -- 0.0945211996555037
	pesos_i(13549) := b"1111111111111111_1111111111111111_1110001111011010_1100000011100010"; -- -0.10994333734782821
	pesos_i(13550) := b"1111111111111111_1111111111111111_1111001001100110_0101001111011010"; -- -0.053126105537711264
	pesos_i(13551) := b"1111111111111111_1111111111111111_1110101101000110_1111000100001101"; -- -0.0809487670140255
	pesos_i(13552) := b"1111111111111111_1111111111111111_1101111111001000_1010000111111101"; -- -0.12584483694613124
	pesos_i(13553) := b"1111111111111111_1111111111111111_1110010010101100_0101011100111001"; -- -0.10674528943398498
	pesos_i(13554) := b"1111111111111111_1111111111111111_1110101101001001_1001000100010110"; -- -0.0809087104905828
	pesos_i(13555) := b"0000000000000000_0000000000000000_0000000010110000_0011101011110010"; -- 0.00268906024330331
	pesos_i(13556) := b"0000000000000000_0000000000000000_0000011111001010_1100001100110010"; -- 0.030437660032402655
	pesos_i(13557) := b"0000000000000000_0000000000000000_0001110101000010_1011100110110100"; -- 0.11429939882714393
	pesos_i(13558) := b"0000000000000000_0000000000000000_0000100010011100_1000101100000001"; -- 0.0336386562898602
	pesos_i(13559) := b"1111111111111111_1111111111111111_1110100111001010_0010001110011101"; -- -0.08675935194640422
	pesos_i(13560) := b"0000000000000000_0000000000000000_0001000010001010_0111100111111101"; -- 0.06461298396077693
	pesos_i(13561) := b"1111111111111111_1111111111111111_1111110100111111_0111100011111010"; -- -0.010750235617463579
	pesos_i(13562) := b"1111111111111111_1111111111111111_1111110101101110_0101000111111000"; -- -0.010035397395075347
	pesos_i(13563) := b"1111111111111111_1111111111111111_1110101111110100_0001111101111001"; -- -0.07830622943990956
	pesos_i(13564) := b"1111111111111111_1111111111111111_1110010001111110_1000000100110001"; -- -0.10744469205918547
	pesos_i(13565) := b"0000000000000000_0000000000000000_0000010100111000_0111000100001111"; -- 0.020392480994685373
	pesos_i(13566) := b"0000000000000000_0000000000000000_0001001001000001_0000100010001110"; -- 0.0713048311743229
	pesos_i(13567) := b"1111111111111111_1111111111111111_1110110101011010_0011111100011011"; -- -0.07284169766896247
	pesos_i(13568) := b"1111111111111111_1111111111111111_1110101100110110_1101011100001101"; -- -0.08119445739108551
	pesos_i(13569) := b"1111111111111111_1111111111111111_1110101000010011_0110100111000110"; -- -0.0856412783310198
	pesos_i(13570) := b"0000000000000000_0000000000000000_0000101010110010_0101010001100110"; -- 0.041783594887366604
	pesos_i(13571) := b"0000000000000000_0000000000000000_0001110000100111_0011111101101110"; -- 0.10997387350498448
	pesos_i(13572) := b"0000000000000000_0000000000000000_0000100001011010_0010011110100011"; -- 0.03262565354878482
	pesos_i(13573) := b"1111111111111111_1111111111111111_1101010110010010_0101010010100101"; -- -0.165735921481137
	pesos_i(13574) := b"1111111111111111_1111111111111111_1101111000110101_0001110010001110"; -- -0.13200208227112195
	pesos_i(13575) := b"0000000000000000_0000000000000000_0000011100110111_1000010111010101"; -- 0.028190960424963784
	pesos_i(13576) := b"1111111111111111_1111111111111111_1110010001000001_1011110010011001"; -- -0.1083719373090461
	pesos_i(13577) := b"0000000000000000_0000000000000000_0000010110101001_0010110101101101"; -- 0.022112693035815457
	pesos_i(13578) := b"1111111111111111_1111111111111111_1110100000110100_1110101011000101"; -- -0.09294254964590676
	pesos_i(13579) := b"0000000000000000_0000000000000000_0010000001111001_1101001010011011"; -- 0.1268588664708083
	pesos_i(13580) := b"1111111111111111_1111111111111111_1110110101101000_1111000001001110"; -- -0.07261751263323345
	pesos_i(13581) := b"0000000000000000_0000000000000000_0001000000000000_1000000111010000"; -- 0.06250773743958453
	pesos_i(13582) := b"1111111111111111_1111111111111111_1101111011101001_0010010110011111"; -- -0.12925495973037734
	pesos_i(13583) := b"0000000000000000_0000000000000000_0010000100111111_1000010111010111"; -- 0.12987553127312992
	pesos_i(13584) := b"1111111111111111_1111111111111111_1111110010101111_0000101010100100"; -- -0.012954077728962262
	pesos_i(13585) := b"0000000000000000_0000000000000000_0000011100001100_1110101110001101"; -- 0.027540895320833765
	pesos_i(13586) := b"0000000000000000_0000000000000000_0000100101111111_0101101110011100"; -- 0.03709957647531154
	pesos_i(13587) := b"1111111111111111_1111111111111111_1110101111111101_1111100011000110"; -- -0.07815594822895275
	pesos_i(13588) := b"1111111111111111_1111111111111111_1111000110000111_1001010111010010"; -- -0.05652488348516818
	pesos_i(13589) := b"1111111111111111_1111111111111111_1101101110101110_0100011110010100"; -- -0.14187195442894443
	pesos_i(13590) := b"0000000000000000_0000000000000000_0000001001100010_0000110001010111"; -- 0.009308596945373457
	pesos_i(13591) := b"0000000000000000_0000000000000000_0000111000011000_0010101100010011"; -- 0.05505627836414692
	pesos_i(13592) := b"0000000000000000_0000000000000000_0000010011011110_1010101100110011"; -- 0.019022655469127896
	pesos_i(13593) := b"1111111111111111_1111111111111111_1110000001111000_1100100010011110"; -- -0.12315698756070526
	pesos_i(13594) := b"0000000000000000_0000000000000000_0001111101011101_1101000111011001"; -- 0.12252532526050526
	pesos_i(13595) := b"0000000000000000_0000000000000000_0001010100001010_1101001110011001"; -- 0.08219645009566093
	pesos_i(13596) := b"0000000000000000_0000000000000000_0010001001000000_0100100010001111"; -- 0.13379338734495608
	pesos_i(13597) := b"1111111111111111_1111111111111111_1101101011100101_1100101110111000"; -- -0.14493109468317844
	pesos_i(13598) := b"1111111111111111_1111111111111111_1110010001000110_1010010000000010"; -- -0.10829710903170224
	pesos_i(13599) := b"0000000000000000_0000000000000000_0000110010100110_0001011100100110"; -- 0.049409338848543954
	pesos_i(13600) := b"0000000000000000_0000000000000000_0001111010100001_0111011111101010"; -- 0.11965131250055401
	pesos_i(13601) := b"0000000000000000_0000000000000000_0000111110011101_1101000001111111"; -- 0.06100180713443802
	pesos_i(13602) := b"0000000000000000_0000000000000000_0000100110011000_1001011001101001"; -- 0.03748455099621498
	pesos_i(13603) := b"0000000000000000_0000000000000000_0010000101101100_1001001000111110"; -- 0.1305629159841527
	pesos_i(13604) := b"0000000000000000_0000000000000000_0001011111011111_0010000100110001"; -- 0.09324843829740583
	pesos_i(13605) := b"0000000000000000_0000000000000000_0000000001100110_1111101100010101"; -- 0.0015713620656772423
	pesos_i(13606) := b"0000000000000000_0000000000000000_0000011001101000_0011111010111101"; -- 0.02502815362743286
	pesos_i(13607) := b"1111111111111111_1111111111111111_1110111100000010_1110001010011000"; -- -0.06636222638776038
	pesos_i(13608) := b"1111111111111111_1111111111111111_1111010001010001_0001011111101110"; -- -0.04563761172890514
	pesos_i(13609) := b"1111111111111111_1111111111111111_1101101111110100_0110101011100101"; -- -0.1408017339791118
	pesos_i(13610) := b"1111111111111111_1111111111111111_1101110011111000_0000101101011110"; -- -0.13684014276470102
	pesos_i(13611) := b"1111111111111111_1111111111111111_1111100100101110_1000111011111101"; -- -0.02663332298116758
	pesos_i(13612) := b"1111111111111111_1111111111111111_1111010110010110_1111011001111011"; -- -0.04066524030432619
	pesos_i(13613) := b"0000000000000000_0000000000000000_0010001000111011_1111010101111100"; -- 0.13372740061336777
	pesos_i(13614) := b"0000000000000000_0000000000000000_0000111011100010_1100011101111111"; -- 0.05814787720842273
	pesos_i(13615) := b"0000000000000000_0000000000000000_0000100011110111_0001101001100110"; -- 0.03502049442255051
	pesos_i(13616) := b"1111111111111111_1111111111111111_1111011001111010_1010000101100110"; -- -0.03719130760130589
	pesos_i(13617) := b"0000000000000000_0000000000000000_0001001110010100_0101011110000011"; -- 0.07648226697854173
	pesos_i(13618) := b"0000000000000000_0000000000000000_0000011111001111_1100101010101011"; -- 0.030514399331200818
	pesos_i(13619) := b"0000000000000000_0000000000000000_0000101111111101_1101010001110001"; -- 0.04684188613362216
	pesos_i(13620) := b"1111111111111111_1111111111111111_1101101100110100_0001010101111010"; -- -0.14373651275951724
	pesos_i(13621) := b"1111111111111111_1111111111111111_1111101110110100_1011011010110100"; -- -0.01677377808520586
	pesos_i(13622) := b"0000000000000000_0000000000000000_0000010100000100_1101010100000011"; -- 0.01960498153034521
	pesos_i(13623) := b"0000000000000000_0000000000000000_0001010100110110_0000100111110010"; -- 0.08285581736017943
	pesos_i(13624) := b"1111111111111111_1111111111111111_1111110011010010_1110000000000000"; -- -0.012407302753936141
	pesos_i(13625) := b"1111111111111111_1111111111111111_1101110110100101_0000000011011000"; -- -0.1342009995718311
	pesos_i(13626) := b"1111111111111111_1111111111111111_1110101001000000_1010000110010100"; -- -0.08495130668118757
	pesos_i(13627) := b"0000000000000000_0000000000000000_0010010010111000_0101000100111100"; -- 0.14343745919300127
	pesos_i(13628) := b"0000000000000000_0000000000000000_0001000000001000_1101010111101011"; -- 0.0626348208377263
	pesos_i(13629) := b"1111111111111111_1111111111111111_1111001011101100_0000111101100001"; -- -0.051085509173723474
	pesos_i(13630) := b"0000000000000000_0000000000000000_0010001011101110_1111000000001111"; -- 0.13645840049654287
	pesos_i(13631) := b"1111111111111111_1111111111111111_1110110000111010_1110010111001101"; -- -0.07722629292646836
	pesos_i(13632) := b"0000000000000000_0000000000000000_0001101101110000_1011110000011000"; -- 0.10718894558215929
	pesos_i(13633) := b"0000000000000000_0000000000000000_0000010000000010_0001110011010111"; -- 0.0156572366266453
	pesos_i(13634) := b"1111111111111111_1111111111111111_1111110100001100_0100001110000100"; -- -0.011531620246694848
	pesos_i(13635) := b"1111111111111111_1111111111111111_1110111010101100_1111111011100001"; -- -0.06767279638265469
	pesos_i(13636) := b"0000000000000000_0000000000000000_0001101000011111_1100011011101010"; -- 0.1020473785987833
	pesos_i(13637) := b"0000000000000000_0000000000000000_0000100001110001_0010001110010101"; -- 0.032976363941532964
	pesos_i(13638) := b"1111111111111111_1111111111111111_1101011011101100_0011101101110001"; -- -0.16045788288028465
	pesos_i(13639) := b"0000000000000000_0000000000000000_0000111101000011_1110001001010000"; -- 0.05962957816740587
	pesos_i(13640) := b"0000000000000000_0000000000000000_0010010000110001_0111010100111011"; -- 0.14137966808203337
	pesos_i(13641) := b"1111111111111111_1111111111111111_1111101000001000_0111100010010100"; -- -0.023308242784522423
	pesos_i(13642) := b"0000000000000000_0000000000000000_0001111101001001_1101100001101001"; -- 0.12222054054113198
	pesos_i(13643) := b"0000000000000000_0000000000000000_0000100110100010_0001111010000010"; -- 0.03762999217722158
	pesos_i(13644) := b"1111111111111111_1111111111111111_1111101001100111_1110000100011001"; -- -0.021852427858936964
	pesos_i(13645) := b"0000000000000000_0000000000000000_0010011100100110_0011011000011111"; -- 0.15292680986228502
	pesos_i(13646) := b"1111111111111111_1111111111111111_1110011000001111_1111011101111001"; -- -0.10131886759670117
	pesos_i(13647) := b"1111111111111111_1111111111111111_1110010011110001_0110011001100110"; -- -0.1056915283838871
	pesos_i(13648) := b"0000000000000000_0000000000000000_0000010010010011_1110010101001101"; -- 0.017881709380774952
	pesos_i(13649) := b"1111111111111111_1111111111111111_1110101111101100_1101111011111100"; -- -0.07841688485221966
	pesos_i(13650) := b"1111111111111111_1111111111111111_1111000111011101_0100001100011010"; -- -0.05521755794805712
	pesos_i(13651) := b"1111111111111111_1111111111111111_1111000110010001_1001101000111111"; -- -0.05637203171026911
	pesos_i(13652) := b"1111111111111111_1111111111111111_1110000000011011_0000010011100111"; -- -0.12458772055349975
	pesos_i(13653) := b"1111111111111111_1111111111111111_1110111000010101_0011110101000110"; -- -0.06998841327012857
	pesos_i(13654) := b"1111111111111111_1111111111111111_1101110101011101_1101101101101000"; -- -0.13528660497657488
	pesos_i(13655) := b"1111111111111111_1111111111111111_1110110001011000_1100101100011111"; -- -0.0767701195565844
	pesos_i(13656) := b"0000000000000000_0000000000000000_0001110111010100_1011101011101000"; -- 0.11652725380634611
	pesos_i(13657) := b"0000000000000000_0000000000000000_0001111100111110_1111000110110000"; -- 0.1220542006467236
	pesos_i(13658) := b"1111111111111111_1111111111111111_1111011001011111_0110010100110010"; -- -0.03760688343045557
	pesos_i(13659) := b"1111111111111111_1111111111111111_1111100010110111_0010110011110001"; -- -0.02845496286554012
	pesos_i(13660) := b"0000000000000000_0000000000000000_0010010101001010_0010001011011000"; -- 0.14566247720075765
	pesos_i(13661) := b"1111111111111111_1111111111111111_1101111100101000_0011010110110101"; -- -0.12829269720970632
	pesos_i(13662) := b"0000000000000000_0000000000000000_0000000100001010_1010000100010010"; -- 0.00406843834621291
	pesos_i(13663) := b"1111111111111111_1111111111111111_1111011100110111_1110011011110110"; -- -0.03430325019039468
	pesos_i(13664) := b"1111111111111111_1111111111111111_1110111011011000_1110000010101100"; -- -0.06700321008395252
	pesos_i(13665) := b"0000000000000000_0000000000000000_0000100101000011_1010010101110100"; -- 0.03618845066173347
	pesos_i(13666) := b"1111111111111111_1111111111111111_1111111010000001_0101110110011011"; -- -0.005838536859528589
	pesos_i(13667) := b"1111111111111111_1111111111111111_1110000010110001_0100010001010001"; -- -0.12229512240218471
	pesos_i(13668) := b"1111111111111111_1111111111111111_1111010111101100_0100001001110010"; -- -0.039363715420565965
	pesos_i(13669) := b"0000000000000000_0000000000000000_0001101000100100_1001100101111001"; -- 0.10212096400045823
	pesos_i(13670) := b"1111111111111111_1111111111111111_1101101111011110_0001011110101101"; -- -0.14114238756062258
	pesos_i(13671) := b"1111111111111111_1111111111111111_1110011011001000_0011111001001011"; -- -0.09850702930801396
	pesos_i(13672) := b"0000000000000000_0000000000000000_0000110011001110_1101000001110010"; -- 0.0500307348663002
	pesos_i(13673) := b"0000000000000000_0000000000000000_0010000010010011_0110010001111010"; -- 0.12724903082202074
	pesos_i(13674) := b"0000000000000000_0000000000000000_0000001000101000_0011111010101010"; -- 0.0084265867101987
	pesos_i(13675) := b"0000000000000000_0000000000000000_0010011110000111_1000101000011011"; -- 0.1544119181835997
	pesos_i(13676) := b"0000000000000000_0000000000000000_0010001100111110_1000000100000100"; -- 0.1376724848800819
	pesos_i(13677) := b"1111111111111111_1111111111111111_1101100101010111_1101101111001101"; -- -0.15100313426023593
	pesos_i(13678) := b"1111111111111111_1111111111111111_1111000101111010_0100000001010001"; -- -0.05672834408660182
	pesos_i(13679) := b"1111111111111111_1111111111111111_1110000101110000_1000110011001010"; -- -0.11937637400419646
	pesos_i(13680) := b"1111111111111111_1111111111111111_1111100111000010_0011101000011111"; -- -0.024380080682369933
	pesos_i(13681) := b"0000000000000000_0000000000000000_0001000100100111_0111000011001011"; -- 0.06700806568177667
	pesos_i(13682) := b"0000000000000000_0000000000000000_0010001110011101_0010111010011011"; -- 0.13911715770084027
	pesos_i(13683) := b"1111111111111111_1111111111111111_1110010101110100_0100101000100000"; -- -0.10369431235712116
	pesos_i(13684) := b"1111111111111111_1111111111111111_1101100111100001_0000110110110000"; -- -0.14890970668031517
	pesos_i(13685) := b"0000000000000000_0000000000000000_0001101111100000_1101100001110000"; -- 0.10889961945107024
	pesos_i(13686) := b"1111111111111111_1111111111111111_1110100001111101_1111100101101100"; -- -0.0918277847377069
	pesos_i(13687) := b"1111111111111111_1111111111111111_1111011111010010_1100011111001011"; -- -0.0319399957451429
	pesos_i(13688) := b"0000000000000000_0000000000000000_0010001110111000_0101011110000101"; -- 0.1395315836621172
	pesos_i(13689) := b"0000000000000000_0000000000000000_0000010101000110_0010010110010001"; -- 0.020601604332424552
	pesos_i(13690) := b"1111111111111111_1111111111111111_1110001100100101_0111110100111111"; -- -0.11270920945674606
	pesos_i(13691) := b"1111111111111111_1111111111111111_1110110000011001_1010011000100000"; -- -0.07773362850644612
	pesos_i(13692) := b"1111111111111111_1111111111111111_1110100000001011_1001011011010011"; -- -0.09357316346234934
	pesos_i(13693) := b"0000000000000000_0000000000000000_0001010010010110_0000111100000001"; -- 0.08041471260815299
	pesos_i(13694) := b"1111111111111111_1111111111111111_1111001001111110_0000101000100000"; -- -0.05276428911158167
	pesos_i(13695) := b"1111111111111111_1111111111111111_1110010010011000_0110010101001000"; -- -0.10704962720551406
	pesos_i(13696) := b"1111111111111111_1111111111111111_1101101100001100_1100010101111011"; -- -0.14433637388926795
	pesos_i(13697) := b"1111111111111111_1111111111111111_1111111100010011_0111111111011000"; -- -0.0036087128594735484
	pesos_i(13698) := b"1111111111111111_1111111111111111_1110110010010010_1101110100010000"; -- -0.07588404051817757
	pesos_i(13699) := b"0000000000000000_0000000000000000_0010000110011000_1111011001001101"; -- 0.13124026669302366
	pesos_i(13700) := b"0000000000000000_0000000000000000_0001111000011001_0011101001000101"; -- 0.11757244296351275
	pesos_i(13701) := b"0000000000000000_0000000000000000_0000000011111100_0011000100110011"; -- 0.0038481473058438022
	pesos_i(13702) := b"0000000000000000_0000000000000000_0000111100111100_0100100100111100"; -- 0.05951364253829935
	pesos_i(13703) := b"0000000000000000_0000000000000000_0000111011111100_0011110011011001"; -- 0.0585363416112053
	pesos_i(13704) := b"0000000000000000_0000000000000000_0000000011000110_0111110101011101"; -- 0.0030287123812433674
	pesos_i(13705) := b"0000000000000000_0000000000000000_0001111110100100_1001010110011100"; -- 0.12360510878316405
	pesos_i(13706) := b"1111111111111111_1111111111111111_1111110000110011_1110110100100010"; -- -0.014832667638266154
	pesos_i(13707) := b"0000000000000000_0000000000000000_0000001101000000_1001000100100010"; -- 0.012703963093626112
	pesos_i(13708) := b"0000000000000000_0000000000000000_0000101001110001_0011011010110011"; -- 0.040790003504001505
	pesos_i(13709) := b"0000000000000000_0000000000000000_0001101101001111_0101111001011101"; -- 0.10667981878497174
	pesos_i(13710) := b"0000000000000000_0000000000000000_0010001011101000_0110010001010001"; -- 0.13635851836346197
	pesos_i(13711) := b"0000000000000000_0000000000000000_0010010111100101_0010000011010000"; -- 0.14802746841835326
	pesos_i(13712) := b"0000000000000000_0000000000000000_0001000000101110_1010111110001010"; -- 0.06321236722387778
	pesos_i(13713) := b"0000000000000000_0000000000000000_0001110101011000_0000100111001110"; -- 0.11462460784811115
	pesos_i(13714) := b"0000000000000000_0000000000000000_0001100101110000_1101010101100001"; -- 0.09937795285117482
	pesos_i(13715) := b"0000000000000000_0000000000000000_0001010000101110_1111110100010110"; -- 0.07884198941841772
	pesos_i(13716) := b"1111111111111111_1111111111111111_1111111010001011_1100001110111000"; -- -0.0056798626128406575
	pesos_i(13717) := b"1111111111111111_1111111111111111_1110010110010110_1101011010111001"; -- -0.10316713307443764
	pesos_i(13718) := b"1111111111111111_1111111111111111_1111000111000100_1001101001100100"; -- -0.05559382501606774
	pesos_i(13719) := b"1111111111111111_1111111111111111_1111011010010100_0111001101111100"; -- -0.03679731580399145
	pesos_i(13720) := b"0000000000000000_0000000000000000_0001111000011011_0000110110010110"; -- 0.11760029712252767
	pesos_i(13721) := b"1111111111111111_1111111111111111_1111110010100000_1001110010110000"; -- -0.013174254505545263
	pesos_i(13722) := b"1111111111111111_1111111111111111_1110101000010010_0000111011100011"; -- -0.08566195455006838
	pesos_i(13723) := b"1111111111111111_1111111111111111_1110001001100011_1111100101110101"; -- -0.11566201104343134
	pesos_i(13724) := b"1111111111111111_1111111111111111_1101110010001011_0100011111111011"; -- -0.13849973792952744
	pesos_i(13725) := b"1111111111111111_1111111111111111_1111011010011000_0010101110110010"; -- -0.03674055967965869
	pesos_i(13726) := b"1111111111111111_1111111111111111_1111111101110011_1111110100101110"; -- -0.0021363985213489105
	pesos_i(13727) := b"1111111111111111_1111111111111111_1111011001111110_1100110101000001"; -- -0.03712765854059031
	pesos_i(13728) := b"0000000000000000_0000000000000000_0001000110011001_0000110001110100"; -- 0.06874158698232864
	pesos_i(13729) := b"0000000000000000_0000000000000000_0000000111001011_1000001010000000"; -- 0.007011562668576986
	pesos_i(13730) := b"1111111111111111_1111111111111111_1111101011000011_1011011000010111"; -- -0.020451182706079013
	pesos_i(13731) := b"0000000000000000_0000000000000000_0001110110010110_1010011000010110"; -- 0.11557996783178869
	pesos_i(13732) := b"0000000000000000_0000000000000000_0000100110010100_1001110101110010"; -- 0.03742393526311814
	pesos_i(13733) := b"0000000000000000_0000000000000000_0001111101111100_1101111100001001"; -- 0.1229991337495613
	pesos_i(13734) := b"0000000000000000_0000000000000000_0000000000110010_1100010010010100"; -- 0.0007746563332372931
	pesos_i(13735) := b"0000000000000000_0000000000000000_0010001100010001_0100101010110110"; -- 0.13698260262455167
	pesos_i(13736) := b"0000000000000000_0000000000000000_0000110100110100_0000101011011000"; -- 0.051575353467556685
	pesos_i(13737) := b"0000000000000000_0000000000000000_0001111110111000_1101110101010001"; -- 0.12391455876595504
	pesos_i(13738) := b"1111111111111111_1111111111111111_1110011010000101_1000100111001001"; -- -0.09952486851420783
	pesos_i(13739) := b"0000000000000000_0000000000000000_0001100110001111_1100011100111110"; -- 0.09985013252537725
	pesos_i(13740) := b"1111111111111111_1111111111111111_1110100110010101_0011101100010001"; -- -0.08756666987625068
	pesos_i(13741) := b"1111111111111111_1111111111111111_1111111001011001_1111010111110110"; -- -0.00643980724895503
	pesos_i(13742) := b"0000000000000000_0000000000000000_0001101011010010_1110001010000100"; -- 0.10478034700585784
	pesos_i(13743) := b"0000000000000000_0000000000000000_0010001100010110_0111100111011011"; -- 0.13706170656236796
	pesos_i(13744) := b"0000000000000000_0000000000000000_0010010111000100_1100000110110110"; -- 0.14753351862183564
	pesos_i(13745) := b"1111111111111111_1111111111111111_1111000110101101_1011001000010011"; -- -0.05594336555200648
	pesos_i(13746) := b"1111111111111111_1111111111111111_1111000111111000_1101110101111001"; -- -0.05479636950904464
	pesos_i(13747) := b"0000000000000000_0000000000000000_0001110110100100_1111000100101011"; -- 0.11579806612016168
	pesos_i(13748) := b"1111111111111111_1111111111111111_1111101111110101_0001010110111100"; -- -0.015791551140151763
	pesos_i(13749) := b"1111111111111111_1111111111111111_1111100100010000_1011001000101001"; -- -0.027088990199954213
	pesos_i(13750) := b"1111111111111111_1111111111111111_1110011101101100_1100011101000110"; -- -0.09599642312399546
	pesos_i(13751) := b"0000000000000000_0000000000000000_0001000011101101_1110101011011011"; -- 0.06613033152429681
	pesos_i(13752) := b"1111111111111111_1111111111111111_1111100100000111_0101100001111010"; -- -0.02723166487037905
	pesos_i(13753) := b"0000000000000000_0000000000000000_0001001001110000_1011000011010111"; -- 0.07203202485544179
	pesos_i(13754) := b"1111111111111111_1111111111111111_1101110000010111_1001100100110100"; -- -0.1402649163123725
	pesos_i(13755) := b"1111111111111111_1111111111111111_1110000111000111_1011011010110000"; -- -0.11804636203414651
	pesos_i(13756) := b"0000000000000000_0000000000000000_0010011000000011_0010101011001100"; -- 0.14848582724785267
	pesos_i(13757) := b"0000000000000000_0000000000000000_0000101010001100_1111011100110001"; -- 0.041213464189748354
	pesos_i(13758) := b"0000000000000000_0000000000000000_0001000010000000_1101000100010100"; -- 0.06446558691382265
	pesos_i(13759) := b"0000000000000000_0000000000000000_0001110100011110_0111100100110101"; -- 0.11374623816651834
	pesos_i(13760) := b"1111111111111111_1111111111111111_1111110011100110_0010010100101010"; -- -0.012113263452878024
	pesos_i(13761) := b"0000000000000000_0000000000000000_0001010110001101_0001010101011010"; -- 0.08418401200585247
	pesos_i(13762) := b"1111111111111111_1111111111111111_1101111110010000_0100001111101111"; -- -0.12670493521960935
	pesos_i(13763) := b"1111111111111111_1111111111111111_1111100001100100_1000100010111000"; -- -0.02971597190802002
	pesos_i(13764) := b"1111111111111111_1111111111111111_1110011101011011_0010111110111000"; -- -0.09626485597676078
	pesos_i(13765) := b"0000000000000000_0000000000000000_0010000001100010_0101110101101111"; -- 0.12650093041288088
	pesos_i(13766) := b"1111111111111111_1111111111111111_1101100101111101_1000001110011011"; -- -0.1504285571682039
	pesos_i(13767) := b"0000000000000000_0000000000000000_0001101001101011_0100111111111101"; -- 0.10319995820814021
	pesos_i(13768) := b"0000000000000000_0000000000000000_0010001111010110_1110100001000011"; -- 0.13999797483594575
	pesos_i(13769) := b"1111111111111111_1111111111111111_1111110100111001_0010110001000101"; -- -0.010846360338223072
	pesos_i(13770) := b"1111111111111111_1111111111111111_1110101100000000_1000111111010000"; -- -0.08202267807294457
	pesos_i(13771) := b"1111111111111111_1111111111111111_1110110001000000_1110001001000111"; -- -0.07713495035087718
	pesos_i(13772) := b"0000000000000000_0000000000000000_0001101110010000_0011011100100011"; -- 0.10766930209114267
	pesos_i(13773) := b"0000000000000000_0000000000000000_0000111010101010_0011101101001000"; -- 0.057285027570289485
	pesos_i(13774) := b"1111111111111111_1111111111111111_1110110001110010_1101001011000101"; -- -0.07637293514074638
	pesos_i(13775) := b"1111111111111111_1111111111111111_1110010000011000_1010100111101011"; -- -0.10899866117119113
	pesos_i(13776) := b"0000000000000000_0000000000000000_0000011010011010_1100111011010000"; -- 0.025799680402564078
	pesos_i(13777) := b"1111111111111111_1111111111111111_1110111010000000_0011111001000001"; -- -0.0683556643330231
	pesos_i(13778) := b"1111111111111111_1111111111111111_1111000010001111_0001110000000110"; -- -0.06031632291725516
	pesos_i(13779) := b"0000000000000000_0000000000000000_0000110001111011_0111011001011010"; -- 0.04875888542890878
	pesos_i(13780) := b"0000000000000000_0000000000000000_0001101100100000_0111101000101110"; -- 0.10596431373048507
	pesos_i(13781) := b"1111111111111111_1111111111111111_1111001101011101_1101001011010001"; -- -0.0493496168923437
	pesos_i(13782) := b"0000000000000000_0000000000000000_0000001111001000_1000100110100011"; -- 0.014778711633161233
	pesos_i(13783) := b"0000000000000000_0000000000000000_0010011000100100_1011000001101011"; -- 0.14899733165249907
	pesos_i(13784) := b"1111111111111111_1111111111111111_1111100100101101_0011011011011111"; -- -0.02665383395119058
	pesos_i(13785) := b"0000000000000000_0000000000000000_0000000110010110_0001010100001010"; -- 0.00619632235642099
	pesos_i(13786) := b"1111111111111111_1111111111111111_1110111110000101_0111001010110010"; -- -0.064369994638525
	pesos_i(13787) := b"0000000000000000_0000000000000000_0000010110010001_1110011111000101"; -- 0.021757588846572164
	pesos_i(13788) := b"1111111111111111_1111111111111111_1111110110110011_0100100110110000"; -- -0.008983034628424652
	pesos_i(13789) := b"0000000000000000_0000000000000000_0000101001011000_0100011000100010"; -- 0.0404094537402936
	pesos_i(13790) := b"1111111111111111_1111111111111111_1110100100011110_1001110101101001"; -- -0.08937660401417846
	pesos_i(13791) := b"0000000000000000_0000000000000000_0010001001011010_0101100000101010"; -- 0.13419104595116593
	pesos_i(13792) := b"0000000000000000_0000000000000000_0000110101101011_1011011111000001"; -- 0.05242489297536632
	pesos_i(13793) := b"0000000000000000_0000000000000000_0001110000110010_0111110111111100"; -- 0.11014544880587038
	pesos_i(13794) := b"0000000000000000_0000000000000000_0001001100000100_1010100111000101"; -- 0.07428990427583189
	pesos_i(13795) := b"0000000000000000_0000000000000000_0000011101000010_0000011101100111"; -- 0.02835127117816823
	pesos_i(13796) := b"0000000000000000_0000000000000000_0001101010010110_0101111111011000"; -- 0.10385703118509058
	pesos_i(13797) := b"1111111111111111_1111111111111111_1110111011101000_1111011010110100"; -- -0.06675775633897418
	pesos_i(13798) := b"1111111111111111_1111111111111111_1101111011001010_0000101100110101"; -- -0.12972955656616655
	pesos_i(13799) := b"1111111111111111_1111111111111111_1111101001011101_0000100100001110"; -- -0.02201789286668959
	pesos_i(13800) := b"1111111111111111_1111111111111111_1101110010101110_1001100110000010"; -- -0.13796082084539205
	pesos_i(13801) := b"1111111111111111_1111111111111111_1110010111111110_1100100101011001"; -- -0.10158101629732139
	pesos_i(13802) := b"0000000000000000_0000000000000000_0010011000100001_0011011011000001"; -- 0.14894430363467695
	pesos_i(13803) := b"1111111111111111_1111111111111111_1110000100101100_0000110010010010"; -- -0.12042161405111526
	pesos_i(13804) := b"1111111111111111_1111111111111111_1111100100101101_0101100010110001"; -- -0.02665181799842637
	pesos_i(13805) := b"1111111111111111_1111111111111111_1111001000100000_1010111111010011"; -- -0.05418873870411932
	pesos_i(13806) := b"0000000000000000_0000000000000000_0000101100100111_0010111010101010"; -- 0.043566624243799985
	pesos_i(13807) := b"1111111111111111_1111111111111111_1111010101100110_1000000111001110"; -- -0.04140461658558104
	pesos_i(13808) := b"0000000000000000_0000000000000000_0001101101011010_0011111101000000"; -- 0.10684581102397604
	pesos_i(13809) := b"1111111111111111_1111111111111111_1110011011010100_1000010010001000"; -- -0.09831973712502677
	pesos_i(13810) := b"0000000000000000_0000000000000000_0001011110011001_0001100010001101"; -- 0.09217980809787871
	pesos_i(13811) := b"0000000000000000_0000000000000000_0001110100110010_0001101100100111"; -- 0.11404580784701944
	pesos_i(13812) := b"0000000000000000_0000000000000000_0000110110001110_0101000001010001"; -- 0.05295278522843706
	pesos_i(13813) := b"0000000000000000_0000000000000000_0000000010001010_0000100000111010"; -- 0.002106203267421319
	pesos_i(13814) := b"1111111111111111_1111111111111111_1110110001100000_1000011001000010"; -- -0.07665215381804291
	pesos_i(13815) := b"0000000000000000_0000000000000000_0001010011000110_1000110100001100"; -- 0.08115464726993742
	pesos_i(13816) := b"1111111111111111_1111111111111111_1111000000010010_0001111101100001"; -- -0.06222347140537883
	pesos_i(13817) := b"1111111111111111_1111111111111111_1111100011111011_1000000110100011"; -- -0.02741231710310819
	pesos_i(13818) := b"0000000000000000_0000000000000000_0010001101110011_0010101101010100"; -- 0.13847609337063635
	pesos_i(13819) := b"1111111111111111_1111111111111111_1110111100101001_0100010110110010"; -- -0.06577648539811211
	pesos_i(13820) := b"0000000000000000_0000000000000000_0001010011100000_1010001111100111"; -- 0.08155273818212318
	pesos_i(13821) := b"1111111111111111_1111111111111111_1110111101001101_0111101110010001"; -- -0.06522395805528831
	pesos_i(13822) := b"1111111111111111_1111111111111111_1101110010010010_1001001010011111"; -- -0.13838847750926683
	pesos_i(13823) := b"1111111111111111_1111111111111111_1111100101101110_1111010001001111"; -- -0.025650721313862444
	pesos_i(13824) := b"0000000000000000_0000000000000000_0000101111111011_1101010001111110"; -- 0.04681137158649383
	pesos_i(13825) := b"0000000000000000_0000000000000000_0000001111001000_1011100101100110"; -- 0.014781558501373405
	pesos_i(13826) := b"1111111111111111_1111111111111111_1110000001000011_0100001010011011"; -- -0.12397369124716207
	pesos_i(13827) := b"1111111111111111_1111111111111111_1110111001001001_0111001010011110"; -- -0.06919177678114978
	pesos_i(13828) := b"0000000000000000_0000000000000000_0000101100101001_0110001010111010"; -- 0.04360024484442503
	pesos_i(13829) := b"0000000000000000_0000000000000000_0000011111011111_0101100011110011"; -- 0.030751761826793043
	pesos_i(13830) := b"1111111111111111_1111111111111111_1101101100111011_0100001000001011"; -- -0.14362704505730212
	pesos_i(13831) := b"0000000000000000_0000000000000000_0000111110110001_1000101011111010"; -- 0.06130283940551357
	pesos_i(13832) := b"0000000000000000_0000000000000000_0001011101100001_1010011111011001"; -- 0.09133385704277283
	pesos_i(13833) := b"1111111111111111_1111111111111111_1111011101001000_1010110101000010"; -- -0.03404729011111077
	pesos_i(13834) := b"1111111111111111_1111111111111111_1110100101011001_1101001101010111"; -- -0.088473120970144
	pesos_i(13835) := b"0000000000000000_0000000000000000_0001000000101111_1110010001101010"; -- 0.06323077771249769
	pesos_i(13836) := b"1111111111111111_1111111111111111_1111000001100110_0101011101110111"; -- -0.060938390247148755
	pesos_i(13837) := b"1111111111111111_1111111111111111_1110001110001111_1001101111000101"; -- -0.11108995860173401
	pesos_i(13838) := b"0000000000000000_0000000000000000_0001000111110101_0111111000110101"; -- 0.07015217582260275
	pesos_i(13839) := b"0000000000000000_0000000000000000_0010010110010001_0101111011110111"; -- 0.14674943465680543
	pesos_i(13840) := b"0000000000000000_0000000000000000_0000011000000101_0001000011011101"; -- 0.023514799015081796
	pesos_i(13841) := b"1111111111111111_1111111111111111_1101110001011111_1110011000011000"; -- -0.1391617004128082
	pesos_i(13842) := b"1111111111111111_1111111111111111_1111110100101010_1111011001000001"; -- -0.011063202894193004
	pesos_i(13843) := b"1111111111111111_1111111111111111_1111101011011111_1001101100111010"; -- -0.020025537720745116
	pesos_i(13844) := b"1111111111111111_1111111111111111_1111001000101000_1001011000101111"; -- -0.05406819673438495
	pesos_i(13845) := b"1111111111111111_1111111111111111_1110000010101101_0111110111010110"; -- -0.12235272910670843
	pesos_i(13846) := b"0000000000000000_0000000000000000_0000011011010011_0001001000100100"; -- 0.026658185750997328
	pesos_i(13847) := b"0000000000000000_0000000000000000_0001100011110100_0011100101111111"; -- 0.09747657159800277
	pesos_i(13848) := b"1111111111111111_1111111111111111_1111110110001110_1101111000110100"; -- -0.009538757567811865
	pesos_i(13849) := b"1111111111111111_1111111111111111_1101101110000101_1110011011001111"; -- -0.14248807374522998
	pesos_i(13850) := b"0000000000000000_0000000000000000_0001100110000011_1010110110000101"; -- 0.0996654940305059
	pesos_i(13851) := b"1111111111111111_1111111111111111_1111000111011011_0110101100100101"; -- -0.05524568883187937
	pesos_i(13852) := b"1111111111111111_1111111111111111_1111011010110000_0011101110000011"; -- -0.03637340583716218
	pesos_i(13853) := b"1111111111111111_1111111111111111_1111010010111110_0111011110101010"; -- -0.04396869758706833
	pesos_i(13854) := b"1111111111111111_1111111111111111_1111011111101101_0000001001101011"; -- -0.03153977279348697
	pesos_i(13855) := b"0000000000000000_0000000000000000_0001001101110101_1101100100111110"; -- 0.07601697693805473
	pesos_i(13856) := b"0000000000000000_0000000000000000_0000010100010100_1110011011110011"; -- 0.01985019146284075
	pesos_i(13857) := b"1111111111111111_1111111111111111_1111100110101001_1110100011001000"; -- -0.024751139858239807
	pesos_i(13858) := b"1111111111111111_1111111111111111_1110001101101010_1101011111101011"; -- -0.11165094857643142
	pesos_i(13859) := b"1111111111111111_1111111111111111_1111011001001010_0101100010010101"; -- -0.037928069819943164
	pesos_i(13860) := b"1111111111111111_1111111111111111_1110110110010100_1001111100100100"; -- -0.07195096381045708
	pesos_i(13861) := b"0000000000000000_0000000000000000_0010000000010110_1001111111001110"; -- 0.1253452184109224
	pesos_i(13862) := b"1111111111111111_1111111111111111_1110100001111001_1110010110010100"; -- -0.09189000267234375
	pesos_i(13863) := b"1111111111111111_1111111111111111_1110010011101110_0010001001111000"; -- -0.10574135381102336
	pesos_i(13864) := b"0000000000000000_0000000000000000_0001010010111101_0011100010110100"; -- 0.08101229084893131
	pesos_i(13865) := b"1111111111111111_1111111111111111_1110001010001100_1111100000111111"; -- -0.11503647288531758
	pesos_i(13866) := b"0000000000000000_0000000000000000_0001110010100100_0101101000001011"; -- 0.11188280842543638
	pesos_i(13867) := b"0000000000000000_0000000000000000_0001110010010001_0010000001111001"; -- 0.11158946001122956
	pesos_i(13868) := b"0000000000000000_0000000000000000_0001100101110011_1010110100001111"; -- 0.09942132580694757
	pesos_i(13869) := b"0000000000000000_0000000000000000_0001110000000111_0100010101101000"; -- 0.10948594842596608
	pesos_i(13870) := b"0000000000000000_0000000000000000_0000000100101111_1011001000101010"; -- 0.004634032599516816
	pesos_i(13871) := b"1111111111111111_1111111111111111_1101111001100000_1100110001101100"; -- -0.13133547186496605
	pesos_i(13872) := b"1111111111111111_1111111111111111_1111100001010000_1000111000001101"; -- -0.030020829878227583
	pesos_i(13873) := b"0000000000000000_0000000000000000_0001010101100101_1101011110100001"; -- 0.08358524029362989
	pesos_i(13874) := b"1111111111111111_1111111111111111_1110010000101110_1101100001001010"; -- -0.1086602039177664
	pesos_i(13875) := b"0000000000000000_0000000000000000_0001111110001001_0101000011110000"; -- 0.12318902835097507
	pesos_i(13876) := b"1111111111111111_1111111111111111_1111100011001001_1111100010111111"; -- -0.028168156944118474
	pesos_i(13877) := b"1111111111111111_1111111111111111_1110010111001011_1001001110010110"; -- -0.10236241890105574
	pesos_i(13878) := b"1111111111111111_1111111111111111_1101110011000110_1000110010010000"; -- -0.1375953816002428
	pesos_i(13879) := b"0000000000000000_0000000000000000_0000100111000010_1100011111001101"; -- 0.03812836404919699
	pesos_i(13880) := b"0000000000000000_0000000000000000_0000110110011101_1000010111000001"; -- 0.053184852166710296
	pesos_i(13881) := b"0000000000000000_0000000000000000_0000000111110100_0011100000001011"; -- 0.007632734881091035
	pesos_i(13882) := b"1111111111111111_1111111111111111_1101111111010000_0110011101001000"; -- -0.1257262658632939
	pesos_i(13883) := b"1111111111111111_1111111111111111_1101101111100101_1000000101110100"; -- -0.1410292713963458
	pesos_i(13884) := b"1111111111111111_1111111111111111_1110111000010010_0100101001011010"; -- -0.07003341008451383
	pesos_i(13885) := b"0000000000000000_0000000000000000_0001100111110110_0001101100100011"; -- 0.10141152949249728
	pesos_i(13886) := b"1111111111111111_1111111111111111_1101101101110111_0101111101110110"; -- -0.14270976414003067
	pesos_i(13887) := b"0000000000000000_0000000000000000_0000011101010100_0101000001111111"; -- 0.02863028626394988
	pesos_i(13888) := b"0000000000000000_0000000000000000_0000010101001001_0000001101001100"; -- 0.02064533800427009
	pesos_i(13889) := b"1111111111111111_1111111111111111_1111111100000101_1100000001010010"; -- -0.0038184928949871466
	pesos_i(13890) := b"0000000000000000_0000000000000000_0001100111011000_1110001010111010"; -- 0.10096566229106053
	pesos_i(13891) := b"1111111111111111_1111111111111111_1110100001010011_1100110001110100"; -- -0.09247133412335151
	pesos_i(13892) := b"1111111111111111_1111111111111111_1110000010100101_0000101010101111"; -- -0.12248166307936384
	pesos_i(13893) := b"0000000000000000_0000000000000000_0000010010011111_1001011110010001"; -- 0.018060181461030576
	pesos_i(13894) := b"0000000000000000_0000000000000000_0000000100010000_0011101111111110"; -- 0.004153966438795467
	pesos_i(13895) := b"1111111111111111_1111111111111111_1101110111100101_0101000100100010"; -- -0.13321965138348185
	pesos_i(13896) := b"1111111111111111_1111111111111111_1110000011110100_1000101010101111"; -- -0.12126858925078068
	pesos_i(13897) := b"1111111111111111_1111111111111111_1111110110000100_1000110001111111"; -- -0.00969621565429778
	pesos_i(13898) := b"1111111111111111_1111111111111111_1110100100100010_0000010101001000"; -- -0.08932463636250751
	pesos_i(13899) := b"0000000000000000_0000000000000000_0000000000011100_0001011010101011"; -- 0.00042859718948421414
	pesos_i(13900) := b"1111111111111111_1111111111111111_1111010011001101_0011100110010110"; -- -0.04374351575517571
	pesos_i(13901) := b"1111111111111111_1111111111111111_1110111101011101_1110110111010011"; -- -0.06497300720743894
	pesos_i(13902) := b"1111111111111111_1111111111111111_1111110111111001_1110101001100000"; -- -0.00790534174849061
	pesos_i(13903) := b"0000000000000000_0000000000000000_0000010000001110_1011101001101010"; -- 0.015849734092577564
	pesos_i(13904) := b"1111111111111111_1111111111111111_1111110001110001_0100001110101111"; -- -0.013896722637971034
	pesos_i(13905) := b"1111111111111111_1111111111111111_1110001110111001_0111000100100100"; -- -0.11045163020454382
	pesos_i(13906) := b"0000000000000000_0000000000000000_0001101101010001_0100110100011101"; -- 0.10670930812674737
	pesos_i(13907) := b"0000000000000000_0000000000000000_0001000111111010_0100101011000011"; -- 0.0702254034265405
	pesos_i(13908) := b"1111111111111111_1111111111111111_1110011010011011_0001010011010000"; -- -0.09919614728676207
	pesos_i(13909) := b"0000000000000000_0000000000000000_0000000101000100_1000100111100011"; -- 0.004952066392094647
	pesos_i(13910) := b"1111111111111111_1111111111111111_1111111100111000_0111111000110110"; -- -0.003044235009857783
	pesos_i(13911) := b"1111111111111111_1111111111111111_1110011110001111_1100001110000111"; -- -0.09546258889928533
	pesos_i(13912) := b"1111111111111111_1111111111111111_1110011001110100_0101010001110101"; -- -0.09978744644154426
	pesos_i(13913) := b"1111111111111111_1111111111111111_1110010011011011_0110000101001101"; -- -0.10602752565504515
	pesos_i(13914) := b"0000000000000000_0000000000000000_0000101010101110_1110101101100010"; -- 0.04173155920789316
	pesos_i(13915) := b"0000000000000000_0000000000000000_0001010001101101_0110100000101101"; -- 0.07979441732438679
	pesos_i(13916) := b"0000000000000000_0000000000000000_0001011110100100_1111010100100000"; -- 0.09236080202077356
	pesos_i(13917) := b"1111111111111111_1111111111111111_1110111000011011_0011111000111101"; -- -0.06989680302462555
	pesos_i(13918) := b"0000000000000000_0000000000000000_0001010000101100_0000101010101000"; -- 0.07879702189332695
	pesos_i(13919) := b"1111111111111111_1111111111111111_1101110000010100_1010001111000011"; -- -0.14031006335926607
	pesos_i(13920) := b"0000000000000000_0000000000000000_0001111010100001_0001100010001010"; -- 0.11964562769698245
	pesos_i(13921) := b"1111111111111111_1111111111111111_1111111000101101_1010111000000001"; -- -0.007115483009384011
	pesos_i(13922) := b"1111111111111111_1111111111111111_1101101100011101_1110100111101110"; -- -0.1440748018849378
	pesos_i(13923) := b"1111111111111111_1111111111111111_1110111111110000_1100110100111101"; -- -0.06273190749817358
	pesos_i(13924) := b"0000000000000000_0000000000000000_0000010101111101_1000011001011011"; -- 0.021446606857730293
	pesos_i(13925) := b"1111111111111111_1111111111111111_1110011011001010_1110101111011100"; -- -0.09846616634947483
	pesos_i(13926) := b"1111111111111111_1111111111111111_1110101110110100_0101011000000110"; -- -0.07927954050018741
	pesos_i(13927) := b"0000000000000000_0000000000000000_0010110001110010_0001000110010111"; -- 0.17361555049545455
	pesos_i(13928) := b"1111111111111111_1111111111111111_1110011101011001_1111011101101110"; -- -0.09628346982654855
	pesos_i(13929) := b"0000000000000000_0000000000000000_0001100001111111_1100000011010000"; -- 0.09569935874468266
	pesos_i(13930) := b"0000000000000000_0000000000000000_0000111100110101_1100110110001101"; -- 0.05941471770622951
	pesos_i(13931) := b"1111111111111111_1111111111111111_1111110100100111_1101000101001111"; -- -0.011111181431898631
	pesos_i(13932) := b"0000000000000000_0000000000000000_0001011110000000_0011010100010001"; -- 0.0918000381161469
	pesos_i(13933) := b"0000000000000000_0000000000000000_0001011100001000_1110100110100110"; -- 0.08997974686402518
	pesos_i(13934) := b"1111111111111111_1111111111111111_1101111000011000_0001100001010010"; -- -0.1324448395552892
	pesos_i(13935) := b"0000000000000000_0000000000000000_0010001100010010_1101001010010010"; -- 0.1370059592741654
	pesos_i(13936) := b"0000000000000000_0000000000000000_0000111011000101_0100111110000000"; -- 0.057698220062648166
	pesos_i(13937) := b"1111111111111111_1111111111111111_1101111101111101_1011101111101111"; -- -0.12698769959367617
	pesos_i(13938) := b"0000000000000000_0000000000000000_0010011111001011_1100000100111000"; -- 0.15545280087800586
	pesos_i(13939) := b"0000000000000000_0000000000000000_0010010100110101_1101011011111101"; -- 0.14535278006894287
	pesos_i(13940) := b"1111111111111111_1111111111111111_1101111110001110_0110001110001100"; -- -0.12673356853355167
	pesos_i(13941) := b"1111111111111111_1111111111111111_1101110101101001_1000001101001100"; -- -0.13510875135473072
	pesos_i(13942) := b"1111111111111111_1111111111111111_1111111010111000_1010101100011100"; -- -0.004994683963752501
	pesos_i(13943) := b"0000000000000000_0000000000000000_0001011011100001_1000010000000100"; -- 0.08937859635207815
	pesos_i(13944) := b"0000000000000000_0000000000000000_0000110001100101_1011010000011010"; -- 0.04842687246900754
	pesos_i(13945) := b"0000000000000000_0000000000000000_0001110101111111_0111100111101010"; -- 0.11522638287130452
	pesos_i(13946) := b"1111111111111111_1111111111111111_1111000101101110_0011111011101110"; -- -0.0569115323611407
	pesos_i(13947) := b"1111111111111111_1111111111111111_1110100111111001_1101110011011011"; -- -0.08603114741628745
	pesos_i(13948) := b"0000000000000000_0000000000000000_0000110100111010_0100100100011010"; -- 0.05167061705468759
	pesos_i(13949) := b"1111111111111111_1111111111111111_1111001100100110_0011000010010010"; -- -0.05019852109675919
	pesos_i(13950) := b"1111111111111111_1111111111111111_1111010000010100_0000100100100100"; -- -0.046569279382533954
	pesos_i(13951) := b"0000000000000000_0000000000000000_0000110000111110_1011011000100111"; -- 0.047831901969897124
	pesos_i(13952) := b"0000000000000000_0000000000000000_0000101111101011_1011100110000101"; -- 0.04656562325081728
	pesos_i(13953) := b"0000000000000000_0000000000000000_0000001111111011_1001000110011100"; -- 0.015557385160596168
	pesos_i(13954) := b"0000000000000000_0000000000000000_0001101000110000_1011110111011000"; -- 0.10230623735412003
	pesos_i(13955) := b"0000000000000000_0000000000000000_0001000111010111_1001010110101100"; -- 0.06969581084409499
	pesos_i(13956) := b"0000000000000000_0000000000000000_0001010010011100_0101110100111110"; -- 0.08051092870513035
	pesos_i(13957) := b"1111111111111111_1111111111111111_1101011000100110_1011001111110110"; -- -0.16347193950724323
	pesos_i(13958) := b"1111111111111111_1111111111111111_1110110011000111_0011111010000010"; -- -0.07508477528837706
	pesos_i(13959) := b"0000000000000000_0000000000000000_0000000000011010_0011110010011100"; -- 0.0004003410435818102
	pesos_i(13960) := b"1111111111111111_1111111111111111_1111101011110101_0101001101010010"; -- -0.019694130361938397
	pesos_i(13961) := b"0000000000000000_0000000000000000_0000010110101111_0111000001100100"; -- 0.02220823706266367
	pesos_i(13962) := b"1111111111111111_1111111111111111_1101111100111001_0110000001001110"; -- -0.12803075876071277
	pesos_i(13963) := b"1111111111111111_1111111111111111_1110001010101100_0111111111010011"; -- -0.11455536946694163
	pesos_i(13964) := b"1111111111111111_1111111111111111_1110101110101011_1111010001010100"; -- -0.07940743392923248
	pesos_i(13965) := b"0000000000000000_0000000000000000_0001110011001010_1111101010000010"; -- 0.11247220690028666
	pesos_i(13966) := b"0000000000000000_0000000000000000_0000001101000101_0001011100100100"; -- 0.012772985636665717
	pesos_i(13967) := b"0000000000000000_0000000000000000_0001101001001110_1101110100011011"; -- 0.10276586440309905
	pesos_i(13968) := b"0000000000000000_0000000000000000_0010001000111101_0011110111011110"; -- 0.13374697359743307
	pesos_i(13969) := b"0000000000000000_0000000000000000_0001111001110101_0100000011001001"; -- 0.11897663977525386
	pesos_i(13970) := b"0000000000000000_0000000000000000_0010010111110110_0111001000010110"; -- 0.14829171208051342
	pesos_i(13971) := b"1111111111111111_1111111111111111_1111000001010000_1001100011000111"; -- -0.06127019057648339
	pesos_i(13972) := b"1111111111111111_1111111111111111_1111100101011011_0001000111111011"; -- -0.025954128421027574
	pesos_i(13973) := b"0000000000000000_0000000000000000_0001100001101101_0011000111110111"; -- 0.09541618615465126
	pesos_i(13974) := b"1111111111111111_1111111111111111_1110111001110110_0111100011010101"; -- -0.06850476084545984
	pesos_i(13975) := b"1111111111111111_1111111111111111_1111001111101010_0011000000110101"; -- -0.04720781999289524
	pesos_i(13976) := b"0000000000000000_0000000000000000_0000100000111011_0100110001110010"; -- 0.03215482502483768
	pesos_i(13977) := b"0000000000000000_0000000000000000_0001110011000111_0110001010111100"; -- 0.11241738403612894
	pesos_i(13978) := b"0000000000000000_0000000000000000_0010000010111100_1011011110011110"; -- 0.12787959668134494
	pesos_i(13979) := b"0000000000000000_0000000000000000_0001011011100000_0111001111111001"; -- 0.0893623812207727
	pesos_i(13980) := b"0000000000000000_0000000000000000_0001011001110110_0001111110111111"; -- 0.08773992923342926
	pesos_i(13981) := b"1111111111111111_1111111111111111_1111110011100101_1011110000010010"; -- -0.012119527549334487
	pesos_i(13982) := b"1111111111111111_1111111111111111_1110101111010110_1100111100011111"; -- -0.07875352385943031
	pesos_i(13983) := b"1111111111111111_1111111111111111_1111111000111001_0101100110101110"; -- -0.00693740378725262
	pesos_i(13984) := b"1111111111111111_1111111111111111_1111011001010111_0100110101110001"; -- -0.03773036959281536
	pesos_i(13985) := b"0000000000000000_0000000000000000_0000111000001111_0100000100100000"; -- 0.0549202636117597
	pesos_i(13986) := b"0000000000000000_0000000000000000_0010100110011101_0010010010000010"; -- 0.16255405582582214
	pesos_i(13987) := b"0000000000000000_0000000000000000_0000001110111101_0110011101011010"; -- 0.014608821284339829
	pesos_i(13988) := b"0000000000000000_0000000000000000_0010000111000100_0100001000000111"; -- 0.1319009081639369
	pesos_i(13989) := b"0000000000000000_0000000000000000_0001101100010111_0001110101000100"; -- 0.10582144645348678
	pesos_i(13990) := b"0000000000000000_0000000000000000_0001110011100111_0011000010010100"; -- 0.1129026757446633
	pesos_i(13991) := b"1111111111111111_1111111111111111_1110001001111111_0011110000101111"; -- -0.11524604665591098
	pesos_i(13992) := b"0000000000000000_0000000000000000_0010000010111111_1011100000010010"; -- 0.12792540021082155
	pesos_i(13993) := b"1111111111111111_1111111111111111_1110010001100010_1011000111011101"; -- -0.10786903723289126
	pesos_i(13994) := b"1111111111111111_1111111111111111_1101100110000001_0011011100110001"; -- -0.15037207658805582
	pesos_i(13995) := b"0000000000000000_0000000000000000_0000010001010011_0000001011111100"; -- 0.016891657450630915
	pesos_i(13996) := b"0000000000000000_0000000000000000_0000110110111010_0010111110010000"; -- 0.053622219801435174
	pesos_i(13997) := b"1111111111111111_1111111111111111_1111110001110110_0100101000001000"; -- -0.013820050331136311
	pesos_i(13998) := b"1111111111111111_1111111111111111_1111101110110100_0100101011000001"; -- -0.016780212281098307
	pesos_i(13999) := b"1111111111111111_1111111111111111_1111011001010000_0000111010111101"; -- -0.03784091842067267
	pesos_i(14000) := b"1111111111111111_1111111111111111_1101110111111001_1001111110000100"; -- -0.13290980365720279
	pesos_i(14001) := b"0000000000000000_0000000000000000_0000000100101010_1011100110100010"; -- 0.004558183714836652
	pesos_i(14002) := b"0000000000000000_0000000000000000_0010010000000100_0000010000000010"; -- 0.14068627403341355
	pesos_i(14003) := b"0000000000000000_0000000000000000_0001100000001111_0000110000000111"; -- 0.09397959861692044
	pesos_i(14004) := b"0000000000000000_0000000000000000_0000110001010100_0000101011010111"; -- 0.04815738437596294
	pesos_i(14005) := b"0000000000000000_0000000000000000_0000101101100110_1110101101010101"; -- 0.04453917347893897
	pesos_i(14006) := b"1111111111111111_1111111111111111_1101110111011111_1110011110101011"; -- -0.13330223165323793
	pesos_i(14007) := b"1111111111111111_1111111111111111_1111001111111000_0010100110110101"; -- -0.046994584487859085
	pesos_i(14008) := b"1111111111111111_1111111111111111_1110110101100100_0111110110001110"; -- -0.07268538744064229
	pesos_i(14009) := b"0000000000000000_0000000000000000_0001101100111101_1110001000010111"; -- 0.10641301207640531
	pesos_i(14010) := b"0000000000000000_0000000000000000_0000000001011111_1111111001011011"; -- 0.0014647457883580582
	pesos_i(14011) := b"0000000000000000_0000000000000000_0001100010111010_1101110001100010"; -- 0.0966012706490304
	pesos_i(14012) := b"1111111111111111_1111111111111111_1110111010011110_0001000000010111"; -- -0.06790065222370498
	pesos_i(14013) := b"0000000000000000_0000000000000000_0000011101011111_1010010000110100"; -- 0.028803122249752327
	pesos_i(14014) := b"1111111111111111_1111111111111111_1111110100000001_0011110110110100"; -- -0.01169981335841366
	pesos_i(14015) := b"0000000000000000_0000000000000000_0000110000011100_0001100111011010"; -- 0.047303786851733365
	pesos_i(14016) := b"1111111111111111_1111111111111111_1110010000001010_0100010110000111"; -- -0.10921826791683216
	pesos_i(14017) := b"0000000000000000_0000000000000000_0010001100101010_0111111001010101"; -- 0.13736714918928533
	pesos_i(14018) := b"1111111111111111_1111111111111111_1110010011101010_1000000011010010"; -- -0.10579676508685246
	pesos_i(14019) := b"0000000000000000_0000000000000000_0000100010000001_0101000011110000"; -- 0.033223207934221295
	pesos_i(14020) := b"0000000000000000_0000000000000000_0000001011010010_0001100010010100"; -- 0.011018310568657146
	pesos_i(14021) := b"0000000000000000_0000000000000000_0001001111000100_1001001010110000"; -- 0.07721821595949183
	pesos_i(14022) := b"0000000000000000_0000000000000000_0001111100000000_0000010001101010"; -- 0.12109401315414763
	pesos_i(14023) := b"1111111111111111_1111111111111111_1111011010001000_0110110001010100"; -- -0.03698084777811283
	pesos_i(14024) := b"0000000000000000_0000000000000000_0001001101010101_0111001110000001"; -- 0.07552263171477691
	pesos_i(14025) := b"1111111111111111_1111111111111111_1101111010001011_0001110010001101"; -- -0.13068982665845788
	pesos_i(14026) := b"1111111111111111_1111111111111111_1110001010110011_1000111001001100"; -- -0.11444769511436013
	pesos_i(14027) := b"0000000000000000_0000000000000000_0010010011110100_1011011010011000"; -- 0.14435902786914237
	pesos_i(14028) := b"0000000000000000_0000000000000000_0001110101111101_1010110011011101"; -- 0.11519890205619274
	pesos_i(14029) := b"1111111111111111_1111111111111111_1101111110110100_0101111100101101"; -- -0.126153995019386
	pesos_i(14030) := b"1111111111111111_1111111111111111_1110110110011110_0010010100100101"; -- -0.07180564730751934
	pesos_i(14031) := b"0000000000000000_0000000000000000_0000111001000100_0010011110001010"; -- 0.05572745438979531
	pesos_i(14032) := b"1111111111111111_1111111111111111_1101100000101000_1001000001011000"; -- -0.15563104494499255
	pesos_i(14033) := b"1111111111111111_1111111111111111_1110110011000100_1100000011101111"; -- -0.07512277768207304
	pesos_i(14034) := b"0000000000000000_0000000000000000_0000000110011100_0110011010010000"; -- 0.0062927342717865355
	pesos_i(14035) := b"0000000000000000_0000000000000000_0000100111100100_0110100010110001"; -- 0.03864149390055392
	pesos_i(14036) := b"0000000000000000_0000000000000000_0000111000111000_1100101101000000"; -- 0.0555541067415201
	pesos_i(14037) := b"1111111111111111_1111111111111111_1111111101111011_0101100011100011"; -- -0.0020241209168961314
	pesos_i(14038) := b"0000000000000000_0000000000000000_0001011110110011_1100110000111010"; -- 0.09258724613758249
	pesos_i(14039) := b"1111111111111111_1111111111111111_1101101010110101_0100100101111101"; -- -0.14567127900447274
	pesos_i(14040) := b"0000000000000000_0000000000000000_0000000101101101_0010001100001111"; -- 0.0055715475482286565
	pesos_i(14041) := b"0000000000000000_0000000000000000_0001100110110010_1100010000100000"; -- 0.10038400436049981
	pesos_i(14042) := b"1111111111111111_1111111111111111_1111101100011000_0011110010111101"; -- -0.019161418882534174
	pesos_i(14043) := b"0000000000000000_0000000000000000_0001101001000011_1001100110110111"; -- 0.10259400103048741
	pesos_i(14044) := b"1111111111111111_1111111111111111_1110101000000010_0011100001011110"; -- -0.08590362278965077
	pesos_i(14045) := b"0000000000000000_0000000000000000_0001110101111010_0000000010101110"; -- 0.11514286287484121
	pesos_i(14046) := b"1111111111111111_1111111111111111_1110010100010110_1011011100011100"; -- -0.10512214254801487
	pesos_i(14047) := b"1111111111111111_1111111111111111_1111111110001111_0000010011000001"; -- -0.0017239598310023665
	pesos_i(14048) := b"0000000000000000_0000000000000000_0000110110100110_1001001111010000"; -- 0.05332301939767735
	pesos_i(14049) := b"0000000000000000_0000000000000000_0001001101111011_0000010110010111"; -- 0.076095914263798
	pesos_i(14050) := b"0000000000000000_0000000000000000_0000010101001110_1000111101000011"; -- 0.02072997451881129
	pesos_i(14051) := b"1111111111111111_1111111111111111_1111111010101111_1101000011010011"; -- -0.0051297650119107125
	pesos_i(14052) := b"0000000000000000_0000000000000000_0000001111111110_1111011100001001"; -- 0.01560920677079142
	pesos_i(14053) := b"1111111111111111_1111111111111111_1110010010010000_0110110010011001"; -- -0.10717126147615212
	pesos_i(14054) := b"1111111111111111_1111111111111111_1110000100100111_0100110110011110"; -- -0.12049403083927668
	pesos_i(14055) := b"0000000000000000_0000000000000000_0000001110100001_0000001101111100"; -- 0.014175622765005
	pesos_i(14056) := b"1111111111111111_1111111111111111_1101111101011100_1100010011000011"; -- -0.1274907135823495
	pesos_i(14057) := b"0000000000000000_0000000000000000_0000000101000111_1110001001110101"; -- 0.005003121893423951
	pesos_i(14058) := b"1111111111111111_1111111111111111_1111000001001101_0001110010010000"; -- -0.061323370761289596
	pesos_i(14059) := b"1111111111111111_1111111111111111_1101110011001110_1000000010000001"; -- -0.13747403004608333
	pesos_i(14060) := b"0000000000000000_0000000000000000_0000110110100101_0110101010010000"; -- 0.05330530187283236
	pesos_i(14061) := b"0000000000000000_0000000000000000_0000110011000110_0111011111101000"; -- 0.04990338716924453
	pesos_i(14062) := b"1111111111111111_1111111111111111_1110111000011010_0001110000001001"; -- -0.06991410056563417
	pesos_i(14063) := b"0000000000000000_0000000000000000_0000101111101010_0111000100111010"; -- 0.046546055490242794
	pesos_i(14064) := b"1111111111111111_1111111111111111_1110000011011110_1101001111011000"; -- -0.12159992190765563
	pesos_i(14065) := b"0000000000000000_0000000000000000_0010010010110101_0101100111010001"; -- 0.14339219429501487
	pesos_i(14066) := b"1111111111111111_1111111111111111_1101110001000001_1000010110000110"; -- -0.13962522012444992
	pesos_i(14067) := b"1111111111111111_1111111111111111_1110011101101011_1010101010100111"; -- -0.09601338779756716
	pesos_i(14068) := b"1111111111111111_1111111111111111_1110011111101101_0011001011101101"; -- -0.0940368816804042
	pesos_i(14069) := b"0000000000000000_0000000000000000_0001001000101001_0101111011000010"; -- 0.0709437582523246
	pesos_i(14070) := b"0000000000000000_0000000000000000_0000100000001111_1111001110011000"; -- 0.0314934011340209
	pesos_i(14071) := b"1111111111111111_1111111111111111_1101011001000100_0010110001010010"; -- -0.1630222605413482
	pesos_i(14072) := b"0000000000000000_0000000000000000_0001101000101010_0101100110101101"; -- 0.10220871417079419
	pesos_i(14073) := b"0000000000000000_0000000000000000_0001010100111101_0010000110000000"; -- 0.08296403298012901
	pesos_i(14074) := b"1111111111111111_1111111111111111_1111101100011010_0110011101010010"; -- -0.01912836315516856
	pesos_i(14075) := b"1111111111111111_1111111111111111_1111111000100111_0101111111111010"; -- -0.0072116865501432635
	pesos_i(14076) := b"0000000000000000_0000000000000000_0001001001011111_0111001110011001"; -- 0.07176897522233754
	pesos_i(14077) := b"0000000000000000_0000000000000000_0000110111011101_0110110101011111"; -- 0.05415996144374407
	pesos_i(14078) := b"0000000000000000_0000000000000000_0001010011001111_1010101100010010"; -- 0.08129376580805764
	pesos_i(14079) := b"1111111111111111_1111111111111111_1101101110001011_0001101010001001"; -- -0.1424086967470224
	pesos_i(14080) := b"0000000000000000_0000000000000000_0010001111010000_0101100011001001"; -- 0.13989787023115458
	pesos_i(14081) := b"1111111111111111_1111111111111111_1110100001011000_0100101110011111"; -- -0.09240271912038839
	pesos_i(14082) := b"1111111111111111_1111111111111111_1111110011000000_0101001001100001"; -- -0.012690402364656947
	pesos_i(14083) := b"1111111111111111_1111111111111111_1110100110110100_1000110110111001"; -- -0.0870887206231789
	pesos_i(14084) := b"1111111111111111_1111111111111111_1110101010010011_1111011101000011"; -- -0.08367972007090442
	pesos_i(14085) := b"1111111111111111_1111111111111111_1110001100101011_1100000011011110"; -- -0.11261362619861184
	pesos_i(14086) := b"1111111111111111_1111111111111111_1101100110110000_0110010100010010"; -- -0.14965217888068091
	pesos_i(14087) := b"1111111111111111_1111111111111111_1111011111010111_0101000000111011"; -- -0.03187082835233771
	pesos_i(14088) := b"0000000000000000_0000000000000000_0001100010100010_1011000110110101"; -- 0.09623251603611761
	pesos_i(14089) := b"0000000000000000_0000000000000000_0010001111101001_1110010011011001"; -- 0.14028768821259008
	pesos_i(14090) := b"1111111111111111_1111111111111111_1110010100110001_0110111000111001"; -- -0.10471449951843517
	pesos_i(14091) := b"1111111111111111_1111111111111111_1111100110011111_0110110100100000"; -- -0.024911098254603838
	pesos_i(14092) := b"1111111111111111_1111111111111111_1110101110011001_0001010101110110"; -- -0.0796953760554045
	pesos_i(14093) := b"0000000000000000_0000000000000000_0000111011010011_0000001110001010"; -- 0.05790731538362772
	pesos_i(14094) := b"1111111111111111_1111111111111111_1101101111010101_1110000110110000"; -- -0.14126767587789144
	pesos_i(14095) := b"1111111111111111_1111111111111111_1111000010011011_0001111000110000"; -- -0.06013308835357488
	pesos_i(14096) := b"1111111111111111_1111111111111111_1111110001111100_1010111101010110"; -- -0.013722459350908132
	pesos_i(14097) := b"0000000000000000_0000000000000000_0010010101010000_0111101101100000"; -- 0.1457593069492307
	pesos_i(14098) := b"1111111111111111_1111111111111111_1110111000011101_0011001010011100"; -- -0.0698669786687997
	pesos_i(14099) := b"0000000000000000_0000000000000000_0000011000100110_1000011000100000"; -- 0.024025328479525255
	pesos_i(14100) := b"0000000000000000_0000000000000000_0001110000011111_1101011111011001"; -- 0.1098608880236208
	pesos_i(14101) := b"1111111111111111_1111111111111111_1111100011110111_1101010100111101"; -- -0.027468369168247696
	pesos_i(14102) := b"0000000000000000_0000000000000000_0001101111011010_1111000001110011"; -- 0.10880949786147733
	pesos_i(14103) := b"1111111111111111_1111111111111111_1110101011011100_1001010000001010"; -- -0.08257174262226855
	pesos_i(14104) := b"1111111111111111_1111111111111111_1101011101111101_0000010011101110"; -- -0.1582486075425881
	pesos_i(14105) := b"1111111111111111_1111111111111111_1110110101101001_0001101101011001"; -- -0.07261494716184397
	pesos_i(14106) := b"1111111111111111_1111111111111111_1110110111000100_0101110110111101"; -- -0.07122244014676277
	pesos_i(14107) := b"0000000000000000_0000000000000000_0010001110010001_1001010010111010"; -- 0.13894013930842802
	pesos_i(14108) := b"0000000000000000_0000000000000000_0010010111101101_0100010101100110"; -- 0.14815171954705222
	pesos_i(14109) := b"0000000000000000_0000000000000000_0000100010101111_0011110001100111"; -- 0.033923888428936094
	pesos_i(14110) := b"0000000000000000_0000000000000000_0010000010000000_0001001000111010"; -- 0.12695421139877008
	pesos_i(14111) := b"0000000000000000_0000000000000000_0000101101101100_1010011010001101"; -- 0.04462662648474104
	pesos_i(14112) := b"1111111111111111_1111111111111111_1110000010111100_1000100001100101"; -- -0.12212321787247062
	pesos_i(14113) := b"1111111111111111_1111111111111111_1111010110011010_1001011011001110"; -- -0.04060990772489612
	pesos_i(14114) := b"0000000000000000_0000000000000000_0000001011010100_1111001110000010"; -- 0.011061877447626848
	pesos_i(14115) := b"0000000000000000_0000000000000000_0001000100100110_0101011110011011"; -- 0.0669913056974545
	pesos_i(14116) := b"0000000000000000_0000000000000000_0001111011100101_1010010110011000"; -- 0.12069163274963704
	pesos_i(14117) := b"0000000000000000_0000000000000000_0000111010100010_0110101110011011"; -- 0.057165837504088095
	pesos_i(14118) := b"1111111111111111_1111111111111111_1110011111101101_1111010011000001"; -- -0.09402532850405014
	pesos_i(14119) := b"0000000000000000_0000000000000000_0001100001101011_1010010000001011"; -- 0.09539246806354681
	pesos_i(14120) := b"0000000000000000_0000000000000000_0000100000100101_0111110011101010"; -- 0.0318220206221544
	pesos_i(14121) := b"1111111111111111_1111111111111111_1111111010100101_0111100010100101"; -- -0.005287608854795118
	pesos_i(14122) := b"0000000000000000_0000000000000000_0000000111111111_0111011011101011"; -- 0.007804329314886246
	pesos_i(14123) := b"0000000000000000_0000000000000000_0010001110111011_0101110100110101"; -- 0.13957769915167986
	pesos_i(14124) := b"0000000000000000_0000000000000000_0001000011010001_0001001110000011"; -- 0.06569024995910534
	pesos_i(14125) := b"0000000000000000_0000000000000000_0000101010010011_1010010110010000"; -- 0.04131541027582128
	pesos_i(14126) := b"0000000000000000_0000000000000000_0001100101010011_0100001000001001"; -- 0.09892666544412806
	pesos_i(14127) := b"0000000000000000_0000000000000000_0000111001000111_1000000111011110"; -- 0.05577861460504593
	pesos_i(14128) := b"1111111111111111_1111111111111111_1110100000000010_0110011001010101"; -- -0.09371338285026971
	pesos_i(14129) := b"0000000000000000_0000000000000000_0000110000100010_1111000000000011"; -- 0.04740810463873628
	pesos_i(14130) := b"0000000000000000_0000000000000000_0000100001111001_1110111101011011"; -- 0.03311058020127977
	pesos_i(14131) := b"0000000000000000_0000000000000000_0001110101100100_1110100001101111"; -- 0.11482098313903076
	pesos_i(14132) := b"0000000000000000_0000000000000000_0001011110001110_0010110011010111"; -- 0.09201317078323101
	pesos_i(14133) := b"1111111111111111_1111111111111111_1110111001101111_1001011111100110"; -- -0.06860972052012385
	pesos_i(14134) := b"1111111111111111_1111111111111111_1101011100101111_1110000010000011"; -- -0.15942570507572473
	pesos_i(14135) := b"0000000000000000_0000000000000000_0000111111001110_1011010110100111"; -- 0.06174788788389959
	pesos_i(14136) := b"0000000000000000_0000000000000000_0001110011010101_0010110111000101"; -- 0.11262785008481574
	pesos_i(14137) := b"1111111111111111_1111111111111111_1110101011111110_0111011001000111"; -- -0.0820547178008276
	pesos_i(14138) := b"0000000000000000_0000000000000000_0000011010100101_1011111110110001"; -- 0.025966625821696034
	pesos_i(14139) := b"1111111111111111_1111111111111111_1101111111100010_1001010111010111"; -- -0.12544883246706046
	pesos_i(14140) := b"0000000000000000_0000000000000000_0001000001000111_0000010111100111"; -- 0.0635837257827775
	pesos_i(14141) := b"0000000000000000_0000000000000000_0001100110000010_0001010110010001"; -- 0.09964117813427409
	pesos_i(14142) := b"0000000000000000_0000000000000000_0000011011101101_1011010101011111"; -- 0.02706464359278413
	pesos_i(14143) := b"0000000000000000_0000000000000000_0010010110111100_1101100110010110"; -- 0.1474128715624967
	pesos_i(14144) := b"1111111111111111_1111111111111111_1111010100010101_0011110100111011"; -- -0.042644665694891705
	pesos_i(14145) := b"1111111111111111_1111111111111111_1101100110110111_0011111101110100"; -- -0.14954760944076387
	pesos_i(14146) := b"1111111111111111_1111111111111111_1110110000110101_0110111001000000"; -- -0.077309712764179
	pesos_i(14147) := b"1111111111111111_1111111111111111_1110100001110000_1000011000001110"; -- -0.09203302527188689
	pesos_i(14148) := b"0000000000000000_0000000000000000_0010001110101101_0110110101011111"; -- 0.1393650394871616
	pesos_i(14149) := b"0000000000000000_0000000000000000_0000011011001101_1100111101000001"; -- 0.026577905105523516
	pesos_i(14150) := b"0000000000000000_0000000000000000_0001011110000111_1101110101101001"; -- 0.0919168836008251
	pesos_i(14151) := b"1111111111111111_1111111111111111_1110100101101001_0100010001011111"; -- -0.08823750202692937
	pesos_i(14152) := b"1111111111111111_1111111111111111_1111011001010011_1011001110000010"; -- -0.037785321097361504
	pesos_i(14153) := b"1111111111111111_1111111111111111_1111111101000010_0100110111111100"; -- -0.00289452159539307
	pesos_i(14154) := b"1111111111111111_1111111111111111_1111011001101011_0010000101111001"; -- -0.03742781455526341
	pesos_i(14155) := b"0000000000000000_0000000000000000_0000011111000101_1011110000110011"; -- 0.030360949058011077
	pesos_i(14156) := b"1111111111111111_1111111111111111_1111001001100111_1000011010100100"; -- -0.05310781955183633
	pesos_i(14157) := b"1111111111111111_1111111111111111_1111111101000010_1010101011000010"; -- -0.002888991969077046
	pesos_i(14158) := b"0000000000000000_0000000000000000_0010010001100100_1001010011011001"; -- 0.1421597509557019
	pesos_i(14159) := b"0000000000000000_0000000000000000_0001100110100011_0100111010100110"; -- 0.10014812042753218
	pesos_i(14160) := b"0000000000000000_0000000000000000_0010010110101001_0101100000010011"; -- 0.14711523502683205
	pesos_i(14161) := b"0000000000000000_0000000000000000_0001010100101010_1000100100000111"; -- 0.08268028664992774
	pesos_i(14162) := b"0000000000000000_0000000000000000_0001100011110000_0111100001001011"; -- 0.09741927946191714
	pesos_i(14163) := b"0000000000000000_0000000000000000_0001011111011001_0111100000100111"; -- 0.09316206886686067
	pesos_i(14164) := b"1111111111111111_1111111111111111_1110100110111101_1111111000110000"; -- -0.08694468822656694
	pesos_i(14165) := b"0000000000000000_0000000000000000_0001100100101010_0011110110000001"; -- 0.09830078496350152
	pesos_i(14166) := b"1111111111111111_1111111111111111_1110100010011101_0010000010000111"; -- -0.09135243124833646
	pesos_i(14167) := b"0000000000000000_0000000000000000_0000111101000011_1011001000011111"; -- 0.05962670576767835
	pesos_i(14168) := b"0000000000000000_0000000000000000_0010001110100111_1111000011100110"; -- 0.13928132653792336
	pesos_i(14169) := b"0000000000000000_0000000000000000_0010001001010100_0101011100001000"; -- 0.13409942577916792
	pesos_i(14170) := b"0000000000000000_0000000000000000_0001111100100001_1101110000010101"; -- 0.12161040785311507
	pesos_i(14171) := b"0000000000000000_0000000000000000_0001001011101101_1011101110110100"; -- 0.07394002098675148
	pesos_i(14172) := b"0000000000000000_0000000000000000_0000101111110110_0000001111100010"; -- 0.04672264352318763
	pesos_i(14173) := b"1111111111111111_1111111111111111_1110000000001110_0001110101111011"; -- -0.12478461977143437
	pesos_i(14174) := b"1111111111111111_1111111111111111_1110001111111101_0100101111000010"; -- -0.1094162609520137
	pesos_i(14175) := b"0000000000000000_0000000000000000_0000101011010011_0010111110000100"; -- 0.04228493675121926
	pesos_i(14176) := b"1111111111111111_1111111111111111_1110100100110101_1000111001110110"; -- -0.08902654291614098
	pesos_i(14177) := b"0000000000000000_0000000000000000_0001101011101000_1100110000110111"; -- 0.10511471112435425
	pesos_i(14178) := b"1111111111111111_1111111111111111_1110111100100000_0011110101110010"; -- -0.065914306308453
	pesos_i(14179) := b"0000000000000000_0000000000000000_0010010001110011_1110111010110111"; -- 0.14239398927685137
	pesos_i(14180) := b"1111111111111111_1111111111111111_1111101010000001_0111110011001111"; -- -0.021461677055544345
	pesos_i(14181) := b"0000000000000000_0000000000000000_0000011001111001_1011000000010110"; -- 0.025294309076447856
	pesos_i(14182) := b"1111111111111111_1111111111111111_1101011101110110_1000111010010000"; -- -0.15834721539490867
	pesos_i(14183) := b"0000000000000000_0000000000000000_0000001111100110_1001110110011010"; -- 0.015237665250875157
	pesos_i(14184) := b"1111111111111111_1111111111111111_1111100000011001_1011011100101100"; -- -0.030857612482648244
	pesos_i(14185) := b"0000000000000000_0000000000000000_0000000000111111_0011100000110111"; -- 0.0009646542735071895
	pesos_i(14186) := b"1111111111111111_1111111111111111_1111010001011011_1001101110000010"; -- -0.045477181143581624
	pesos_i(14187) := b"1111111111111111_1111111111111111_1111010111010010_0100011111111100"; -- -0.03976011359936212
	pesos_i(14188) := b"0000000000000000_0000000000000000_0010010100101100_0000011000101011"; -- 0.14520300431023905
	pesos_i(14189) := b"0000000000000000_0000000000000000_0010000000010010_0101110111001110"; -- 0.12528024946606686
	pesos_i(14190) := b"1111111111111111_1111111111111111_1110100110111111_0000001110001110"; -- -0.0869291094582965
	pesos_i(14191) := b"0000000000000000_0000000000000000_0001111101111011_0111001001000011"; -- 0.12297739147698279
	pesos_i(14192) := b"1111111111111111_1111111111111111_1110010000000100_0010000100001000"; -- -0.10931199596044759
	pesos_i(14193) := b"1111111111111111_1111111111111111_1101110101010101_1000110111101111"; -- -0.13541329309090994
	pesos_i(14194) := b"1111111111111111_1111111111111111_1110110110010000_0110000111000000"; -- -0.07201565807586167
	pesos_i(14195) := b"1111111111111111_1111111111111111_1101110001001101_0111110001000011"; -- -0.13944266655642185
	pesos_i(14196) := b"0000000000000000_0000000000000000_0010001001111110_1101011001111110"; -- 0.13474789205852591
	pesos_i(14197) := b"1111111111111111_1111111111111111_1101101001100110_0011100001001001"; -- -0.14687774865705833
	pesos_i(14198) := b"0000000000000000_0000000000000000_0000100000011011_1001001100011101"; -- 0.03167075591346107
	pesos_i(14199) := b"0000000000000000_0000000000000000_0000110100011110_0010001101010100"; -- 0.051241119444786105
	pesos_i(14200) := b"1111111111111111_1111111111111111_1101101101110011_0101001010011100"; -- -0.14277156537798186
	pesos_i(14201) := b"0000000000000000_0000000000000000_0010000000011101_0000000011001011"; -- 0.12544255217263192
	pesos_i(14202) := b"1111111111111111_1111111111111111_1101101111010110_1110101000011100"; -- -0.14125191506085602
	pesos_i(14203) := b"1111111111111111_1111111111111111_1111001110111011_1111100000111100"; -- -0.047913060615839845
	pesos_i(14204) := b"0000000000000000_0000000000000000_0001000101100010_0001010111100100"; -- 0.06790291609081561
	pesos_i(14205) := b"0000000000000000_0000000000000000_0000011010110000_0100001000101000"; -- 0.026126990174188056
	pesos_i(14206) := b"1111111111111111_1111111111111111_1110100111001011_0000001011110111"; -- -0.0867460391672513
	pesos_i(14207) := b"0000000000000000_0000000000000000_0001101111111011_0010101011000110"; -- 0.10930125555241813
	pesos_i(14208) := b"0000000000000000_0000000000000000_0010001000011100_1100100011110000"; -- 0.1332517228081441
	pesos_i(14209) := b"1111111111111111_1111111111111111_1111011100111000_0100010011010110"; -- -0.034297654783011486
	pesos_i(14210) := b"0000000000000000_0000000000000000_0001001111011110_0011101101111001"; -- 0.07760974594197588
	pesos_i(14211) := b"0000000000000000_0000000000000000_0001010011100011_1010101011111010"; -- 0.08159893606653461
	pesos_i(14212) := b"1111111111111111_1111111111111111_1111101010100101_0010111001101101"; -- -0.020917032655560882
	pesos_i(14213) := b"0000000000000000_0000000000000000_0001101100101000_0110111111100100"; -- 0.10608577069370705
	pesos_i(14214) := b"1111111111111111_1111111111111111_1110000111011010_0110011100011110"; -- -0.11776118772629417
	pesos_i(14215) := b"0000000000000000_0000000000000000_0001101111101111_0001111111101101"; -- 0.10911750344278498
	pesos_i(14216) := b"0000000000000000_0000000000000000_0000010001100111_1101011111111110"; -- 0.017209529458275818
	pesos_i(14217) := b"0000000000000000_0000000000000000_0000110111110100_1100101000001110"; -- 0.05451643802516138
	pesos_i(14218) := b"0000000000000000_0000000000000000_0010000101010111_0111110110111111"; -- 0.13024125973291392
	pesos_i(14219) := b"0000000000000000_0000000000000000_0000111000101001_0101010100100011"; -- 0.05531818478495675
	pesos_i(14220) := b"1111111111111111_1111111111111111_1111110001110011_1011111001010011"; -- -0.01385889495734942
	pesos_i(14221) := b"0000000000000000_0000000000000000_0001101111011010_1111010010000101"; -- 0.10880974060502664
	pesos_i(14222) := b"0000000000000000_0000000000000000_0001011101001000_1111111010010011"; -- 0.09095755666964642
	pesos_i(14223) := b"0000000000000000_0000000000000000_0000011001011010_1000110010110101"; -- 0.024819177924052194
	pesos_i(14224) := b"1111111111111111_1111111111111111_1111110010010010_0001101101001011"; -- -0.01339559011263642
	pesos_i(14225) := b"0000000000000000_0000000000000000_0001100101000110_0100100110011011"; -- 0.09872875243852032
	pesos_i(14226) := b"1111111111111111_1111111111111111_1110111001111001_1010011111010001"; -- -0.06845618379076897
	pesos_i(14227) := b"0000000000000000_0000000000000000_0010010110101000_1011000000111110"; -- 0.14710523144026771
	pesos_i(14228) := b"0000000000000000_0000000000000000_0001001110100110_1010010100111100"; -- 0.07676155761526109
	pesos_i(14229) := b"1111111111111111_1111111111111111_1110010110101011_0100101000100100"; -- -0.102855077956891
	pesos_i(14230) := b"1111111111111111_1111111111111111_1111010000110011_1111100001010100"; -- -0.04608200033721381
	pesos_i(14231) := b"0000000000000000_0000000000000000_0000111110110111_0100101111011101"; -- 0.06139063012783451
	pesos_i(14232) := b"0000000000000000_0000000000000000_0001011001111100_1111010000000011"; -- 0.08784413414402069
	pesos_i(14233) := b"1111111111111111_1111111111111111_1110110110111001_0111010000010111"; -- -0.07138895445822428
	pesos_i(14234) := b"1111111111111111_1111111111111111_1111111000011011_0001111011100110"; -- -0.007398670995532093
	pesos_i(14235) := b"0000000000000000_0000000000000000_0000100111000001_1100110101011011"; -- 0.038113436461222304
	pesos_i(14236) := b"0000000000000000_0000000000000000_0000100111001000_1010001010110000"; -- 0.03821770476462474
	pesos_i(14237) := b"0000000000000000_0000000000000000_0000010101001101_1001110001111010"; -- 0.02071550355924535
	pesos_i(14238) := b"1111111111111111_1111111111111111_1111111010101011_1000010001010011"; -- -0.0051953598958223044
	pesos_i(14239) := b"1111111111111111_1111111111111111_1101110100000001_0110100110000011"; -- -0.13669720230284765
	pesos_i(14240) := b"1111111111111111_1111111111111111_1101101101001101_0000101111001001"; -- -0.14335562083446782
	pesos_i(14241) := b"1111111111111111_1111111111111111_1110101111000110_1000111101100010"; -- -0.07900146355957553
	pesos_i(14242) := b"1111111111111111_1111111111111111_1111110010000001_0011110001000011"; -- -0.013653024258328398
	pesos_i(14243) := b"1111111111111111_1111111111111111_1111000101011001_1110101011011011"; -- -0.057221719389986964
	pesos_i(14244) := b"0000000000000000_0000000000000000_0001011111011100_1100011010110010"; -- 0.0932125268110323
	pesos_i(14245) := b"1111111111111111_1111111111111111_1111001100110001_0000011010001010"; -- -0.0500331794768971
	pesos_i(14246) := b"1111111111111111_1111111111111111_1111010100111000_1000100010111011"; -- -0.04210610811941846
	pesos_i(14247) := b"1111111111111111_1111111111111111_1111010100100100_1110101101000001"; -- -0.04240541142137259
	pesos_i(14248) := b"1111111111111111_1111111111111111_1110111100010100_0100101111011101"; -- -0.06609655234581631
	pesos_i(14249) := b"1111111111111111_1111111111111111_1111010001011011_1111001010101110"; -- -0.04547198540693137
	pesos_i(14250) := b"0000000000000000_0000000000000000_0000010011011011_1101101001100000"; -- 0.018979691004467752
	pesos_i(14251) := b"1111111111111111_1111111111111111_1111110100110111_0101100001010000"; -- -0.010874252675163194
	pesos_i(14252) := b"1111111111111111_1111111111111111_1111111010100101_1110100101110000"; -- -0.005280885805157335
	pesos_i(14253) := b"0000000000000000_0000000000000000_0001001010101001_0011100011010100"; -- 0.07289462259067986
	pesos_i(14254) := b"1111111111111111_1111111111111111_1101101110100000_1100010001000001"; -- -0.14207814613937023
	pesos_i(14255) := b"1111111111111111_1111111111111111_1111100000111000_1001001010101010"; -- -0.030386765843046178
	pesos_i(14256) := b"1111111111111111_1111111111111111_1101111111000010_1101111011111111"; -- -0.12593275341299293
	pesos_i(14257) := b"1111111111111111_1111111111111111_1111010100100110_0111111111011111"; -- -0.042381294340244645
	pesos_i(14258) := b"1111111111111111_1111111111111111_1101101100011101_1111000010110111"; -- -0.14407439732137722
	pesos_i(14259) := b"1111111111111111_1111111111111111_1111110010010100_1001100010100111"; -- -0.013357600415213907
	pesos_i(14260) := b"1111111111111111_1111111111111111_1111111110111101_0011100100000001"; -- -0.0010189412484661149
	pesos_i(14261) := b"1111111111111111_1111111111111111_1111101011101010_0110000100101101"; -- -0.019861151310965212
	pesos_i(14262) := b"1111111111111111_1111111111111111_1101101110010100_0100111110010101"; -- -0.14226820577433544
	pesos_i(14263) := b"1111111111111111_1111111111111111_1111000101101001_1100110001000111"; -- -0.056979401196542545
	pesos_i(14264) := b"0000000000000000_0000000000000000_0001001111100011_0100111101101010"; -- 0.07768722866549706
	pesos_i(14265) := b"1111111111111111_1111111111111111_1110001111100110_1100000110101100"; -- -0.10976018482695431
	pesos_i(14266) := b"1111111111111111_1111111111111111_1110100010010100_0111011011001110"; -- -0.09148461797969175
	pesos_i(14267) := b"0000000000000000_0000000000000000_0010010111110111_0100001111010000"; -- 0.14830421280369227
	pesos_i(14268) := b"1111111111111111_1111111111111111_1111101011101011_1111010100001011"; -- -0.019837078837726896
	pesos_i(14269) := b"1111111111111111_1111111111111111_1111100010011101_0111010101111011"; -- -0.028847367775195223
	pesos_i(14270) := b"1111111111111111_1111111111111111_1111110110101110_0001101100110110"; -- -0.009062098915714628
	pesos_i(14271) := b"0000000000000000_0000000000000000_0000110100101000_0110100100110100"; -- 0.05139787215024053
	pesos_i(14272) := b"1111111111111111_1111111111111111_1111001010001110_1100010100010000"; -- -0.052509006030677714
	pesos_i(14273) := b"0000000000000000_0000000000000000_0001001011010000_1110000010001000"; -- 0.0734997112120968
	pesos_i(14274) := b"0000000000000000_0000000000000000_0000100101100110_1000001101000101"; -- 0.03672047066378679
	pesos_i(14275) := b"1111111111111111_1111111111111111_1110001111000011_1001000111010111"; -- -0.11029709336008879
	pesos_i(14276) := b"1111111111111111_1111111111111111_1110100110001100_1000111001101100"; -- -0.08769903061111273
	pesos_i(14277) := b"0000000000000000_0000000000000000_0001110001101011_0011101010100101"; -- 0.11101118595903763
	pesos_i(14278) := b"1111111111111111_1111111111111111_1111101001001001_1011110011101110"; -- -0.022312347211000793
	pesos_i(14279) := b"1111111111111111_1111111111111111_1110101011010000_0011010001111010"; -- -0.08276054412032738
	pesos_i(14280) := b"1111111111111111_1111111111111111_1111100010011001_0101110010001000"; -- -0.02890989005255864
	pesos_i(14281) := b"1111111111111111_1111111111111111_1110110001111001_1011011111010010"; -- -0.07626772996683472
	pesos_i(14282) := b"0000000000000000_0000000000000000_0010100110000100_0011111101001011"; -- 0.16217418274260154
	pesos_i(14283) := b"1111111111111111_1111111111111111_1111001110001110_1100100100101101"; -- -0.04860251099541466
	pesos_i(14284) := b"0000000000000000_0000000000000000_0001001101010010_0100011101101101"; -- 0.0754742279255829
	pesos_i(14285) := b"1111111111111111_1111111111111111_1111100011001101_0101100100010001"; -- -0.028116639388187065
	pesos_i(14286) := b"1111111111111111_1111111111111111_1110110110011010_1100110011110010"; -- -0.0718566807765062
	pesos_i(14287) := b"0000000000000000_0000000000000000_0010000000000110_0110101010001010"; -- 0.12509790299197443
	pesos_i(14288) := b"1111111111111111_1111111111111111_1110100101000100_0100011011010010"; -- -0.088801931153032
	pesos_i(14289) := b"0000000000000000_0000000000000000_0001011010111110_0011110011100010"; -- 0.08884029888155746
	pesos_i(14290) := b"1111111111111111_1111111111111111_1111111010011000_1101110011110011"; -- -0.005479994468236629
	pesos_i(14291) := b"0000000000000000_0000000000000000_0000111110100101_0100010111111001"; -- 0.061115620821650306
	pesos_i(14292) := b"0000000000000000_0000000000000000_0001010000011001_0011000111101111"; -- 0.07850944605209759
	pesos_i(14293) := b"0000000000000000_0000000000000000_0000111011001101_0111100000000000"; -- 0.057822704215436484
	pesos_i(14294) := b"1111111111111111_1111111111111111_1111001110001100_0011100111010011"; -- -0.04864157305295275
	pesos_i(14295) := b"0000000000000000_0000000000000000_0010010110000011_1110110101101100"; -- 0.14654430276729352
	pesos_i(14296) := b"1111111111111111_1111111111111111_1110101011110110_0110101000010101"; -- -0.08217751486489608
	pesos_i(14297) := b"0000000000000000_0000000000000000_0001110110010100_1110101000101000"; -- 0.11555350759004067
	pesos_i(14298) := b"0000000000000000_0000000000000000_0010001110101100_0110011001011001"; -- 0.13934936202507434
	pesos_i(14299) := b"1111111111111111_1111111111111111_1111011000000111_0001101010011011"; -- -0.03895410261018304
	pesos_i(14300) := b"1111111111111111_1111111111111111_1111000111001000_1101111000000100"; -- -0.05552875899673079
	pesos_i(14301) := b"0000000000000000_0000000000000000_0000101000001111_0101100100100000"; -- 0.039296694027012344
	pesos_i(14302) := b"0000000000000000_0000000000000000_0001001100001111_1010101001101011"; -- 0.0744577894899775
	pesos_i(14303) := b"1111111111111111_1111111111111111_1110101111101101_0011010011011101"; -- -0.07841176609662784
	pesos_i(14304) := b"1111111111111111_1111111111111111_1101101110111010_0001000100010111"; -- -0.14169209648739534
	pesos_i(14305) := b"0000000000000000_0000000000000000_0001011010110100_0111011000000000"; -- 0.08869111542899016
	pesos_i(14306) := b"0000000000000000_0000000000000000_0010011001100010_1000001101010010"; -- 0.1499406886072361
	pesos_i(14307) := b"0000000000000000_0000000000000000_0001011111101001_1001011110100011"; -- 0.09340808601527414
	pesos_i(14308) := b"0000000000000000_0000000000000000_0000000110101011_0100010111011011"; -- 0.006519666538168675
	pesos_i(14309) := b"0000000000000000_0000000000000000_0010010010011010_0010111110111011"; -- 0.14297769843245964
	pesos_i(14310) := b"1111111111111111_1111111111111111_1111010110011100_0011111110000100"; -- -0.04058459317513957
	pesos_i(14311) := b"1111111111111111_1111111111111111_1111110100110001_1100111100111000"; -- -0.010958718105904545
	pesos_i(14312) := b"1111111111111111_1111111111111111_1111001011100111_0010011110011110"; -- -0.05116035840379422
	pesos_i(14313) := b"1111111111111111_1111111111111111_1110100110011101_0001100010011011"; -- -0.08744665349718038
	pesos_i(14314) := b"1111111111111111_1111111111111111_1110110100101011_1111000010000000"; -- -0.07354828717241037
	pesos_i(14315) := b"0000000000000000_0000000000000000_0000011000011001_1110110110001011"; -- 0.02383312829417919
	pesos_i(14316) := b"0000000000000000_0000000000000000_0000000110110000_1101111001111011"; -- 0.006605057748557863
	pesos_i(14317) := b"1111111111111111_1111111111111111_1111011101110011_1111101000000000"; -- -0.03338658805477298
	pesos_i(14318) := b"0000000000000000_0000000000000000_0001100110011110_0001011111001001"; -- 0.10006855647930728
	pesos_i(14319) := b"0000000000000000_0000000000000000_0001111000001101_1101100001110001"; -- 0.11739876518250952
	pesos_i(14320) := b"0000000000000000_0000000000000000_0000001011100101_1001101111010100"; -- 0.011316050809347368
	pesos_i(14321) := b"0000000000000000_0000000000000000_0001100001110111_1110101111000110"; -- 0.09557984905419224
	pesos_i(14322) := b"1111111111111111_1111111111111111_1111010110000001_1111111110000001"; -- -0.04098513702568467
	pesos_i(14323) := b"0000000000000000_0000000000000000_0000010001111010_1010101010110001"; -- 0.017496746255933202
	pesos_i(14324) := b"0000000000000000_0000000000000000_0000010000001001_1100110101110001"; -- 0.015774574287206824
	pesos_i(14325) := b"0000000000000000_0000000000000000_0000100010101110_0110011010111101"; -- 0.03391115303567704
	pesos_i(14326) := b"1111111111111111_1111111111111111_1110101000010000_0000110110111010"; -- -0.08569254119876843
	pesos_i(14327) := b"0000000000000000_0000000000000000_0010000001000111_1001011010110101"; -- 0.12609235691989387
	pesos_i(14328) := b"0000000000000000_0000000000000000_0010000100101101_1000010100011000"; -- 0.12960082849425303
	pesos_i(14329) := b"1111111111111111_1111111111111111_1101111101000101_0011010110110111"; -- -0.1278501918126805
	pesos_i(14330) := b"1111111111111111_1111111111111111_1101100111111110_0100010000001000"; -- -0.14846396258508573
	pesos_i(14331) := b"1111111111111111_1111111111111111_1111010101100100_1111101111010010"; -- -0.04142786154337255
	pesos_i(14332) := b"0000000000000000_0000000000000000_0010001110111111_0101001101000110"; -- 0.13963814221183593
	pesos_i(14333) := b"1111111111111111_1111111111111111_1110010100101101_1111010101100000"; -- -0.10476747909861622
	pesos_i(14334) := b"1111111111111111_1111111111111111_1110010110010101_1000001010011010"; -- -0.10318740596483174
	pesos_i(14335) := b"1111111111111111_1111111111111111_1110111111111101_0011001100001001"; -- -0.06254273441176132
	pesos_i(14336) := b"0000000000000000_0000000000000000_0001010001001110_1000001100010000"; -- 0.07932299745295401
	pesos_i(14337) := b"1111111111111111_1111111111111111_1110111100101001_0111101100101111"; -- -0.06577329742611085
	pesos_i(14338) := b"0000000000000000_0000000000000000_0001001010110111_1000101100101011"; -- 0.07311315339214962
	pesos_i(14339) := b"1111111111111111_1111111111111111_1111010000101100_0010001000000000"; -- -0.04620158681514589
	pesos_i(14340) := b"1111111111111111_1111111111111111_1111111111000001_1001010111000111"; -- -0.000952376342468268
	pesos_i(14341) := b"0000000000000000_0000000000000000_0000111011110010_1000001110100110"; -- 0.05838797374265484
	pesos_i(14342) := b"0000000000000000_0000000000000000_0000110001011111_1010101100000101"; -- 0.048334778606072375
	pesos_i(14343) := b"0000000000000000_0000000000000000_0010011111110011_1000011001001011"; -- 0.1560596401684524
	pesos_i(14344) := b"1111111111111111_1111111111111111_1110000101111010_1010101011000000"; -- -0.1192220003045742
	pesos_i(14345) := b"1111111111111111_1111111111111111_1111010000110010_1100100010011110"; -- -0.04610010287121485
	pesos_i(14346) := b"0000000000000000_0000000000000000_0010000101111010_0101100011011001"; -- 0.1307731179053569
	pesos_i(14347) := b"0000000000000000_0000000000000000_0001101100011010_1111010110011010"; -- 0.10588011744972313
	pesos_i(14348) := b"1111111111111111_1111111111111111_1111111101110100_1111010100010011"; -- -0.0021216228347141377
	pesos_i(14349) := b"1111111111111111_1111111111111111_1111101101101111_0010111111100000"; -- -0.017834670755659848
	pesos_i(14350) := b"1111111111111111_1111111111111111_1101101111001011_0011111101001101"; -- -0.14142994282212482
	pesos_i(14351) := b"1111111111111111_1111111111111111_1101111111010011_0101100001110000"; -- -0.12568137416099423
	pesos_i(14352) := b"1111111111111111_1111111111111111_1110011001111111_1110110010100100"; -- -0.0996105290186201
	pesos_i(14353) := b"1111111111111111_1111111111111111_1110110101110100_0000101100111001"; -- -0.07244806161066655
	pesos_i(14354) := b"1111111111111111_1111111111111111_1101110010010000_1110010100100110"; -- -0.13841407614684828
	pesos_i(14355) := b"1111111111111111_1111111111111111_1111111111110001_0111100100000101"; -- -0.00022166862335929965
	pesos_i(14356) := b"0000000000000000_0000000000000000_0000001111001111_1001111101000010"; -- 0.014886811869617047
	pesos_i(14357) := b"1111111111111111_1111111111111111_1110101110010110_0011010010100101"; -- -0.07973929388962347
	pesos_i(14358) := b"0000000000000000_0000000000000000_0000001001001111_1010101101001101"; -- 0.009028154665418899
	pesos_i(14359) := b"1111111111111111_1111111111111111_1110001001110000_0010110010110001"; -- -0.11547585178758298
	pesos_i(14360) := b"1111111111111111_1111111111111111_1110001110110100_0001111110001111"; -- -0.11053278683735626
	pesos_i(14361) := b"0000000000000000_0000000000000000_0000011110010111_1101010100101110"; -- 0.029660533629260005
	pesos_i(14362) := b"1111111111111111_1111111111111111_1111000111000101_0111000110110111"; -- -0.05558099072814159
	pesos_i(14363) := b"0000000000000000_0000000000000000_0001011011010001_1000111011001000"; -- 0.08913509727546
	pesos_i(14364) := b"0000000000000000_0000000000000000_0001000100000000_1001000111100101"; -- 0.06641494595788491
	pesos_i(14365) := b"1111111111111111_1111111111111111_1110010100100011_1010011001000100"; -- -0.10492478218272742
	pesos_i(14366) := b"0000000000000000_0000000000000000_0010000111110010_0111000010101100"; -- 0.13260559275300796
	pesos_i(14367) := b"0000000000000000_0000000000000000_0000011100110010_0011100101111011"; -- 0.028110115468103887
	pesos_i(14368) := b"0000000000000000_0000000000000000_0001000000011000_0110100001010111"; -- 0.0628724300308787
	pesos_i(14369) := b"1111111111111111_1111111111111111_1111011010110100_0000010111000001"; -- -0.036315575041965704
	pesos_i(14370) := b"0000000000000000_0000000000000000_0001001101101101_1111010110000000"; -- 0.0758965909951861
	pesos_i(14371) := b"0000000000000000_0000000000000000_0001111010100011_0101001001011110"; -- 0.1196795920215667
	pesos_i(14372) := b"1111111111111111_1111111111111111_1101101001100110_0011100010001101"; -- -0.14687773280757258
	pesos_i(14373) := b"0000000000000000_0000000000000000_0000001010011010_0011111010010011"; -- 0.01016608319565631
	pesos_i(14374) := b"1111111111111111_1111111111111111_1110101101011100_0000010101001101"; -- -0.08062712546164469
	pesos_i(14375) := b"0000000000000000_0000000000000000_0010000101111111_0001111001111001"; -- 0.13084593258659025
	pesos_i(14376) := b"1111111111111111_1111111111111111_1111010000111100_0011010011110111"; -- -0.045956315704059246
	pesos_i(14377) := b"1111111111111111_1111111111111111_1111101110111110_0011100111000101"; -- -0.01662863680688527
	pesos_i(14378) := b"1111111111111111_1111111111111111_1111101000111000_1111000101001100"; -- -0.022568625364427906
	pesos_i(14379) := b"1111111111111111_1111111111111111_1110000101010100_1011111101010000"; -- -0.11980060862069139
	pesos_i(14380) := b"0000000000000000_0000000000000000_0010011010111110_0100111110100010"; -- 0.15134141645557153
	pesos_i(14381) := b"1111111111111111_1111111111111111_1111000000001000_0011010000011100"; -- -0.06237482379410281
	pesos_i(14382) := b"0000000000000000_0000000000000000_0010010100110111_1011110011010101"; -- 0.1453817386886717
	pesos_i(14383) := b"1111111111111111_1111111111111111_1111110010111010_0011001000000010"; -- -0.012783884560966725
	pesos_i(14384) := b"0000000000000000_0000000000000000_0001100011101001_0011001011001010"; -- 0.09730832502675514
	pesos_i(14385) := b"0000000000000000_0000000000000000_0001001101111100_1111100101001011"; -- 0.0761256989555132
	pesos_i(14386) := b"0000000000000000_0000000000000000_0010010001001100_0011010001100111"; -- 0.14178779147847206
	pesos_i(14387) := b"0000000000000000_0000000000000000_0000001001110011_0111101100110110"; -- 0.009574604744470793
	pesos_i(14388) := b"1111111111111111_1111111111111111_1111010001010010_0100010101111011"; -- -0.04561963782451667
	pesos_i(14389) := b"0000000000000000_0000000000000000_0000001010011111_0101001110110111"; -- 0.010243637176886455
	pesos_i(14390) := b"0000000000000000_0000000000000000_0001011011010011_0111111110101001"; -- 0.08916471360671856
	pesos_i(14391) := b"0000000000000000_0000000000000000_0000001010001101_0111101000110100"; -- 0.009971273053654106
	pesos_i(14392) := b"0000000000000000_0000000000000000_0010000101100010_0100011111011010"; -- 0.13040589402707975
	pesos_i(14393) := b"0000000000000000_0000000000000000_0010001001011111_0011000111100000"; -- 0.1342650576569676
	pesos_i(14394) := b"0000000000000000_0000000000000000_0001011100110001_1010100111101010"; -- 0.09060155841134843
	pesos_i(14395) := b"1111111111111111_1111111111111111_1101110011011101_1011100100111101"; -- -0.13724176654286252
	pesos_i(14396) := b"1111111111111111_1111111111111111_1111110011001011_1111010000110000"; -- -0.01251291108718754
	pesos_i(14397) := b"1111111111111111_1111111111111111_1110110010000010_0101010100000000"; -- -0.07613629102845643
	pesos_i(14398) := b"1111111111111111_1111111111111111_1110100110001101_1011111011110100"; -- -0.08768087901755657
	pesos_i(14399) := b"0000000000000000_0000000000000000_0000110111100011_1011001001011001"; -- 0.05425562541475902
	pesos_i(14400) := b"1111111111111111_1111111111111111_1101100111000101_0000001110010000"; -- -0.14933755609949223
	pesos_i(14401) := b"1111111111111111_1111111111111111_1111101000101010_1100011010011111"; -- -0.022784792003804014
	pesos_i(14402) := b"1111111111111111_1111111111111111_1111010110101011_0001000101010001"; -- -0.04035846492100174
	pesos_i(14403) := b"1111111111111111_1111111111111111_1110010100000100_1101001011111111"; -- -0.10539513851314279
	pesos_i(14404) := b"1111111111111111_1111111111111111_1111110111101100_1111011101011011"; -- -0.00810293233329396
	pesos_i(14405) := b"0000000000000000_0000000000000000_0001011100101110_0110001101101010"; -- 0.09055157990072062
	pesos_i(14406) := b"1111111111111111_1111111111111111_1110010001000001_1100001100011011"; -- -0.10837154959380754
	pesos_i(14407) := b"1111111111111111_1111111111111111_1111100110110001_0001000011111000"; -- -0.024641933004844498
	pesos_i(14408) := b"1111111111111111_1111111111111111_1110000011110110_1100110010111101"; -- -0.12123413454894771
	pesos_i(14409) := b"0000000000000000_0000000000000000_0000010011001011_1101100111111110"; -- 0.018735527557211643
	pesos_i(14410) := b"1111111111111111_1111111111111111_1110100011100000_1001110010010011"; -- -0.0903226987539845
	pesos_i(14411) := b"0000000000000000_0000000000000000_0000100110010101_1011011011011110"; -- 0.037440709402644025
	pesos_i(14412) := b"1111111111111111_1111111111111111_1111010110100110_0010110000010010"; -- -0.040433164162622215
	pesos_i(14413) := b"1111111111111111_1111111111111111_1111001001111001_0100001100101100"; -- -0.052837182877350994
	pesos_i(14414) := b"0000000000000000_0000000000000000_0000111011001111_0111000000001101"; -- 0.05785274818536026
	pesos_i(14415) := b"1111111111111111_1111111111111111_1110000000011000_1110111110011101"; -- -0.12461950709787553
	pesos_i(14416) := b"1111111111111111_1111111111111111_1110101001111101_1111111110001100"; -- -0.08401491969597905
	pesos_i(14417) := b"0000000000000000_0000000000000000_0000111010110111_1001111111001101"; -- 0.057489383231804594
	pesos_i(14418) := b"1111111111111111_1111111111111111_1110000010111101_1100011001010010"; -- -0.12210426795928395
	pesos_i(14419) := b"0000000000000000_0000000000000000_0000111101011111_1110001000001101"; -- 0.06005680856364335
	pesos_i(14420) := b"1111111111111111_1111111111111111_1101110001010010_1010010100100111"; -- -0.1393639353911866
	pesos_i(14421) := b"1111111111111111_1111111111111111_1110110011001111_1010000101110101"; -- -0.0749568071205198
	pesos_i(14422) := b"0000000000000000_0000000000000000_0000010111101101_0110000011010110"; -- 0.023153354896127458
	pesos_i(14423) := b"0000000000000000_0000000000000000_0001011001011000_0011010011100101"; -- 0.08728342629611764
	pesos_i(14424) := b"1111111111111111_1111111111111111_1110010001000001_1110011101010100"; -- -0.10836939037393753
	pesos_i(14425) := b"1111111111111111_1111111111111111_1111110110100100_1011001101000101"; -- -0.009205623358076719
	pesos_i(14426) := b"0000000000000000_0000000000000000_0010001100110000_1110100010000011"; -- 0.13746503067916432
	pesos_i(14427) := b"1111111111111111_1111111111111111_1111010111111000_0110000010111110"; -- -0.039178804020086985
	pesos_i(14428) := b"0000000000000000_0000000000000000_0001110010001010_1000111001110101"; -- 0.111489204033157
	pesos_i(14429) := b"0000000000000000_0000000000000000_0000111010011100_1001100010100111"; -- 0.057076969885735025
	pesos_i(14430) := b"0000000000000000_0000000000000000_0010000111010000_0010111111111000"; -- 0.13208293719168418
	pesos_i(14431) := b"1111111111111111_1111111111111111_1110100110011000_1011111101110100"; -- -0.08751300258799279
	pesos_i(14432) := b"1111111111111111_1111111111111111_1111111101110110_1010010011000000"; -- -0.002095893070695943
	pesos_i(14433) := b"0000000000000000_0000000000000000_0000111001010101_0010001101110010"; -- 0.05598660972873849
	pesos_i(14434) := b"1111111111111111_1111111111111111_1111000010111110_1100001100110111"; -- -0.05958919431216531
	pesos_i(14435) := b"1111111111111111_1111111111111111_1111010100111000_0001010110011011"; -- -0.04211297005004972
	pesos_i(14436) := b"0000000000000000_0000000000000000_0001001111011011_1001000010101001"; -- 0.07756904722710928
	pesos_i(14437) := b"0000000000000000_0000000000000000_0001100000110000_1000110000100010"; -- 0.09449077438236768
	pesos_i(14438) := b"1111111111111111_1111111111111111_1110010110010101_0011010001011101"; -- -0.10319206938295104
	pesos_i(14439) := b"0000000000000000_0000000000000000_0001110011111010_1000010011101000"; -- 0.11319761911116788
	pesos_i(14440) := b"1111111111111111_1111111111111111_1110001001000111_0101101110011001"; -- -0.11609866642001353
	pesos_i(14441) := b"1111111111111111_1111111111111111_1110000111100100_0110111010011110"; -- -0.11760815288387887
	pesos_i(14442) := b"1111111111111111_1111111111111111_1101101101001101_1001100000001100"; -- -0.14334726053912325
	pesos_i(14443) := b"0000000000000000_0000000000000000_0001000010101111_1011001111001010"; -- 0.06518100436222532
	pesos_i(14444) := b"0000000000000000_0000000000000000_0001110101110011_1001100111101110"; -- 0.11504518566109248
	pesos_i(14445) := b"1111111111111111_1111111111111111_1110100111011011_1010000101010010"; -- -0.08649245982346308
	pesos_i(14446) := b"1111111111111111_1111111111111111_1110001101001100_0010100100011000"; -- -0.11211913269475295
	pesos_i(14447) := b"1111111111111111_1111111111111111_1101111000100011_1010000000001011"; -- -0.13226890313228548
	pesos_i(14448) := b"1111111111111111_1111111111111111_1101110110110010_0110100011111100"; -- -0.1339964280394146
	pesos_i(14449) := b"0000000000000000_0000000000000000_0001010001000100_1111010010010000"; -- 0.07917717465253139
	pesos_i(14450) := b"1111111111111111_1111111111111111_1110101011010010_0010001111101101"; -- -0.08273101299539935
	pesos_i(14451) := b"1111111111111111_1111111111111111_1110010000101000_1010110011010001"; -- -0.10875434776779905
	pesos_i(14452) := b"0000000000000000_0000000000000000_0000001100011100_0110011111110010"; -- 0.012152191708573365
	pesos_i(14453) := b"0000000000000000_0000000000000000_0001100001110010_1011010101110111"; -- 0.09550031812008693
	pesos_i(14454) := b"0000000000000000_0000000000000000_0000100001101010_1011111110011001"; -- 0.03287885171898696
	pesos_i(14455) := b"0000000000000000_0000000000000000_0000001001110001_0110100010001101"; -- 0.009542974919507974
	pesos_i(14456) := b"1111111111111111_1111111111111111_1111100001001110_0010101110110110"; -- -0.030057209093009043
	pesos_i(14457) := b"0000000000000000_0000000000000000_0001000001100010_1101110111011110"; -- 0.06400858558609324
	pesos_i(14458) := b"1111111111111111_1111111111111111_1110011111011110_1111001110000101"; -- -0.09425428384521492
	pesos_i(14459) := b"1111111111111111_1111111111111111_1111001001010110_1010001111010011"; -- -0.05336547942933864
	pesos_i(14460) := b"0000000000000000_0000000000000000_0001011101010011_0101011010101000"; -- 0.09111539468469673
	pesos_i(14461) := b"0000000000000000_0000000000000000_0001000011111111_0000010110011011"; -- 0.0663913253038822
	pesos_i(14462) := b"1111111111111111_1111111111111111_1111011100001001_1000101011010010"; -- -0.03501064660739903
	pesos_i(14463) := b"1111111111111111_1111111111111111_1111100110000001_0111010001110100"; -- -0.025368425030969987
	pesos_i(14464) := b"1111111111111111_1111111111111111_1110001101100100_0010101101000100"; -- -0.11175279223438729
	pesos_i(14465) := b"0000000000000000_0000000000000000_0010010011100101_1001100000101100"; -- 0.14412833276772524
	pesos_i(14466) := b"1111111111111111_1111111111111111_1111010010111000_0111110111100010"; -- -0.0440598796426914
	pesos_i(14467) := b"1111111111111111_1111111111111111_1110000001100111_1000000001011101"; -- -0.12342069366899065
	pesos_i(14468) := b"0000000000000000_0000000000000000_0000100100101010_0001100000001101"; -- 0.03579855257658315
	pesos_i(14469) := b"1111111111111111_1111111111111111_1111101110100011_0110110001110100"; -- -0.017037602991987734
	pesos_i(14470) := b"0000000000000000_0000000000000000_0000001110110101_1110010000010001"; -- 0.01449418456541418
	pesos_i(14471) := b"1111111111111111_1111111111111111_1111101100000111_0001011010000000"; -- -0.019423097435953676
	pesos_i(14472) := b"1111111111111111_1111111111111111_1111001111100101_0110010111010001"; -- -0.04728091860294562
	pesos_i(14473) := b"0000000000000000_0000000000000000_0000001100111001_1101000110110011"; -- 0.01260100008454003
	pesos_i(14474) := b"0000000000000000_0000000000000000_0010000101101100_1010100001001001"; -- 0.13056422969800707
	pesos_i(14475) := b"0000000000000000_0000000000000000_0000000001010010_0111110011000110"; -- 0.0012586578345341356
	pesos_i(14476) := b"0000000000000000_0000000000000000_0001111110100010_1101000111000011"; -- 0.12357817648520984
	pesos_i(14477) := b"0000000000000000_0000000000000000_0001111100010110_1011010111101001"; -- 0.12144028610314647
	pesos_i(14478) := b"1111111111111111_1111111111111111_1111001001100111_1110110011110010"; -- -0.053101721725394575
	pesos_i(14479) := b"1111111111111111_1111111111111111_1111010001001011_1111110111010011"; -- -0.045715461692289606
	pesos_i(14480) := b"1111111111111111_1111111111111111_1110111010011010_1001110011011100"; -- -0.0679532970247582
	pesos_i(14481) := b"1111111111111111_1111111111111111_1111001101000000_0101011011100000"; -- -0.04979950940368171
	pesos_i(14482) := b"0000000000000000_0000000000000000_0000101000001001_1011010010101101"; -- 0.03921059819905071
	pesos_i(14483) := b"0000000000000000_0000000000000000_0000111110000111_0101101110000001"; -- 0.06065914055692221
	pesos_i(14484) := b"0000000000000000_0000000000000000_0001000001001000_1101000100111010"; -- 0.06361110371834812
	pesos_i(14485) := b"1111111111111111_1111111111111111_1111001011010000_1010010001101010"; -- -0.05150387210178548
	pesos_i(14486) := b"1111111111111111_1111111111111111_1110111001000101_0111010011010110"; -- -0.06925267960193726
	pesos_i(14487) := b"1111111111111111_1111111111111111_1110110111101110_0010010001000100"; -- -0.07058499663592592
	pesos_i(14488) := b"1111111111111111_1111111111111111_1111110110101000_0111011111001000"; -- -0.009148133963368294
	pesos_i(14489) := b"0000000000000000_0000000000000000_0001011010010100_0101000100111100"; -- 0.08820064267201501
	pesos_i(14490) := b"1111111111111111_1111111111111111_1110111101001010_0001001110010001"; -- -0.06527593345980943
	pesos_i(14491) := b"0000000000000000_0000000000000000_0001000011100111_0110001110110110"; -- 0.0660307234356097
	pesos_i(14492) := b"0000000000000000_0000000000000000_0000111111100010_0111000111100011"; -- 0.06204902448939161
	pesos_i(14493) := b"1111111111111111_1111111111111111_1101101011111111_1100100010010110"; -- -0.14453455304858023
	pesos_i(14494) := b"1111111111111111_1111111111111111_1111110101001000_0010111010010100"; -- -0.010617340840314897
	pesos_i(14495) := b"0000000000000000_0000000000000000_0000101101000111_1010101010001101"; -- 0.044062289583072047
	pesos_i(14496) := b"1111111111111111_1111111111111111_1111001001011100_1010101111000101"; -- -0.05327345306997869
	pesos_i(14497) := b"1111111111111111_1111111111111111_1110010101011010_1000010101111111"; -- -0.10408750191766072
	pesos_i(14498) := b"1111111111111111_1111111111111111_1111100110000001_1001101111010110"; -- -0.025366077568255173
	pesos_i(14499) := b"1111111111111111_1111111111111111_1111111010101101_1111111100000100"; -- -0.005157529393410469
	pesos_i(14500) := b"1111111111111111_1111111111111111_1110111100101011_1100110101011010"; -- -0.06573788215603565
	pesos_i(14501) := b"0000000000000000_0000000000000000_0000001111110111_1010111100010001"; -- 0.015498105747034883
	pesos_i(14502) := b"0000000000000000_0000000000000000_0001011110000011_1101110110011000"; -- 0.09185585931892595
	pesos_i(14503) := b"1111111111111111_1111111111111111_1110111010010010_0100011100100000"; -- -0.06808047735306479
	pesos_i(14504) := b"1111111111111111_1111111111111111_1111011001110001_1111000110110010"; -- -0.03732385068386662
	pesos_i(14505) := b"0000000000000000_0000000000000000_0010000011001000_1011000000010100"; -- 0.1280622529170885
	pesos_i(14506) := b"0000000000000000_0000000000000000_0000110100110111_1010001100101111"; -- 0.0516302098418905
	pesos_i(14507) := b"0000000000000000_0000000000000000_0000011110111110_0110100101100010"; -- 0.03024920130931465
	pesos_i(14508) := b"0000000000000000_0000000000000000_0000100111110001_1111010000011100"; -- 0.038848168327951196
	pesos_i(14509) := b"0000000000000000_0000000000000000_0010010100011001_0100100001010011"; -- 0.14491703050772287
	pesos_i(14510) := b"0000000000000000_0000000000000000_0001101001000100_1101100111001001"; -- 0.10261307870317014
	pesos_i(14511) := b"0000000000000000_0000000000000000_0000111101101100_0010111110010001"; -- 0.06024453447886599
	pesos_i(14512) := b"1111111111111111_1111111111111111_1110010110011101_0011100110111101"; -- -0.10306967865359994
	pesos_i(14513) := b"0000000000000000_0000000000000000_0000011100011010_1011000111010000"; -- 0.02775107692748117
	pesos_i(14514) := b"1111111111111111_1111111111111111_1110111001110010_0110000101101001"; -- -0.06856719185967296
	pesos_i(14515) := b"0000000000000000_0000000000000000_0000100111101001_0110110011111110"; -- 0.0387180443680951
	pesos_i(14516) := b"1111111111111111_1111111111111111_1101100011011011_1010111001001010"; -- -0.15289793674807825
	pesos_i(14517) := b"1111111111111111_1111111111111111_1111011111010010_1101000011011000"; -- -0.03193945631102709
	pesos_i(14518) := b"0000000000000000_0000000000000000_0001001011000010_0010000101001011"; -- 0.0732746894438135
	pesos_i(14519) := b"1111111111111111_1111111111111111_1111011100100111_0111001101111101"; -- -0.03455427354894671
	pesos_i(14520) := b"0000000000000000_0000000000000000_0010010110111111_1000100101010010"; -- 0.14745386365935925
	pesos_i(14521) := b"1111111111111111_1111111111111111_1111101111100111_0000001010110110"; -- -0.016006308147562123
	pesos_i(14522) := b"1111111111111111_1111111111111111_1111001011101111_1010011000100010"; -- -0.05103074708466106
	pesos_i(14523) := b"1111111111111111_1111111111111111_1110011001111101_1111101100111010"; -- -0.09964017701244637
	pesos_i(14524) := b"1111111111111111_1111111111111111_1101101110010000_1010000110111011"; -- -0.14232434453523135
	pesos_i(14525) := b"0000000000000000_0000000000000000_0000001111111000_1000111000101000"; -- 0.015511402838683007
	pesos_i(14526) := b"1111111111111111_1111111111111111_1101110110101110_1110010111100101"; -- -0.13405001797094135
	pesos_i(14527) := b"0000000000000000_0000000000000000_0001010000111001_0101000101101001"; -- 0.0789996034076056
	pesos_i(14528) := b"0000000000000000_0000000000000000_0001100110100001_1101010100000010"; -- 0.10012561135224116
	pesos_i(14529) := b"0000000000000000_0000000000000000_0001101101000000_0011001101100100"; -- 0.1064483755329198
	pesos_i(14530) := b"0000000000000000_0000000000000000_0000110010010110_1111110011000101"; -- 0.049178884524737114
	pesos_i(14531) := b"1111111111111111_1111111111111111_1110001110100001_0001101101011111"; -- -0.11082295362999187
	pesos_i(14532) := b"1111111111111111_1111111111111111_1110011000100110_0011000001000001"; -- -0.10097978981472663
	pesos_i(14533) := b"1111111111111111_1111111111111111_1101110101000101_1101111100111000"; -- -0.1356525887541612
	pesos_i(14534) := b"1111111111111111_1111111111111111_1101011001001111_1111101011010011"; -- -0.16284210537317134
	pesos_i(14535) := b"0000000000000000_0000000000000000_0001111010011111_1100111100011010"; -- 0.11962599162267462
	pesos_i(14536) := b"0000000000000000_0000000000000000_0001010111100110_1101101000100110"; -- 0.08555377420317524
	pesos_i(14537) := b"0000000000000000_0000000000000000_0000111001010000_0000100000110001"; -- 0.055908691480105945
	pesos_i(14538) := b"1111111111111111_1111111111111111_1111001101110010_1000111101001100"; -- -0.049033207002328674
	pesos_i(14539) := b"1111111111111111_1111111111111111_1110000010100101_1000001100001110"; -- -0.12247448829558899
	pesos_i(14540) := b"1111111111111111_1111111111111111_1111010000110111_0010110110000101"; -- -0.04603305331239949
	pesos_i(14541) := b"1111111111111111_1111111111111111_1111101001010101_0100111100001110"; -- -0.022135790973290517
	pesos_i(14542) := b"1111111111111111_1111111111111111_1110100101010000_1111101011101110"; -- -0.08860809026386839
	pesos_i(14543) := b"1111111111111111_1111111111111111_1101111110110111_1011010001011001"; -- -0.1261031420683262
	pesos_i(14544) := b"0000000000000000_0000000000000000_0000001111100111_1010110010110111"; -- 0.015253824936690042
	pesos_i(14545) := b"0000000000000000_0000000000000000_0001000001000100_1101011101000101"; -- 0.06355042876514665
	pesos_i(14546) := b"1111111111111111_1111111111111111_1111000100100010_0000000010000011"; -- -0.058074920670957236
	pesos_i(14547) := b"1111111111111111_1111111111111111_1110000101000100_0100001001011000"; -- -0.12005219796782991
	pesos_i(14548) := b"1111111111111111_1111111111111111_1110100011111100_1100111011001010"; -- -0.08989245962534274
	pesos_i(14549) := b"1111111111111111_1111111111111111_1111010010101000_1110100010011110"; -- -0.04429765846505317
	pesos_i(14550) := b"1111111111111111_1111111111111111_1110011010100011_0011010110001100"; -- -0.09907212566726185
	pesos_i(14551) := b"1111111111111111_1111111111111111_1110010110111110_0101101011001111"; -- -0.10256416743620134
	pesos_i(14552) := b"1111111111111111_1111111111111111_1110000010100000_1111000110000101"; -- -0.1225441980462981
	pesos_i(14553) := b"0000000000000000_0000000000000000_0001000011101011_1110010011010001"; -- 0.06609945386630656
	pesos_i(14554) := b"1111111111111111_1111111111111111_1110000011111001_1001000111101000"; -- -0.12119186490725799
	pesos_i(14555) := b"1111111111111111_1111111111111111_1110011000110101_0011101101111101"; -- -0.10075023838692221
	pesos_i(14556) := b"0000000000000000_0000000000000000_0010001101001000_1111010100011011"; -- 0.13783199213269925
	pesos_i(14557) := b"0000000000000000_0000000000000000_0010000000010010_0000101011110110"; -- 0.1252753116362548
	pesos_i(14558) := b"0000000000000000_0000000000000000_0010000000100100_1111001101011010"; -- 0.12556382123629295
	pesos_i(14559) := b"1111111111111111_1111111111111111_1111101001110001_1110101000011011"; -- -0.021699303174343168
	pesos_i(14560) := b"1111111111111111_1111111111111111_1110101101100010_0110010111101000"; -- -0.08052981454174941
	pesos_i(14561) := b"0000000000000000_0000000000000000_0000000111100001_1000001110010000"; -- 0.007347319263745492
	pesos_i(14562) := b"1111111111111111_1111111111111111_1111110011111101_0010111111000111"; -- -0.011761678690825821
	pesos_i(14563) := b"0000000000000000_0000000000000000_0001001011011111_1001110100100010"; -- 0.0737245757075692
	pesos_i(14564) := b"1111111111111111_1111111111111111_1101111011101010_0011101100111100"; -- -0.12923841270098868
	pesos_i(14565) := b"1111111111111111_1111111111111111_1101101001010011_1010101011001101"; -- -0.14716083987673886
	pesos_i(14566) := b"1111111111111111_1111111111111111_1101101011111001_0000111111001111"; -- -0.14463711926175493
	pesos_i(14567) := b"1111111111111111_1111111111111111_1110001101011000_1101001100010110"; -- -0.1119258948499655
	pesos_i(14568) := b"0000000000000000_0000000000000000_0000011001110001_1011100001011100"; -- 0.02517273174134593
	pesos_i(14569) := b"1111111111111111_1111111111111111_1111111011010110_0010001011011010"; -- -0.004545041824355317
	pesos_i(14570) := b"1111111111111111_1111111111111111_1111000011001010_0111010101000100"; -- -0.059410735039790455
	pesos_i(14571) := b"0000000000000000_0000000000000000_0001110100111011_0111100001001111"; -- 0.11418868962171155
	pesos_i(14572) := b"0000000000000000_0000000000000000_0000110110010010_1111101000110100"; -- 0.05302394653736808
	pesos_i(14573) := b"0000000000000000_0000000000000000_0010000011101001_1100101101110011"; -- 0.12856742444058025
	pesos_i(14574) := b"1111111111111111_1111111111111111_1110011110100100_0101100110101011"; -- -0.09514846400219722
	pesos_i(14575) := b"1111111111111111_1111111111111111_1111110010010000_0111010110011101"; -- -0.013420724192320616
	pesos_i(14576) := b"0000000000000000_0000000000000000_0001000010101001_1110111100010110"; -- 0.0650929858730249
	pesos_i(14577) := b"0000000000000000_0000000000000000_0001110011100000_0010010100011101"; -- 0.11279518091467974
	pesos_i(14578) := b"1111111111111111_1111111111111111_1110111100001110_0000010010100011"; -- -0.06619235059071495
	pesos_i(14579) := b"1111111111111111_1111111111111111_1101111011000011_1111100111010010"; -- -0.12982214561244484
	pesos_i(14580) := b"0000000000000000_0000000000000000_0001100101001010_1000001011110000"; -- 0.09879320482770376
	pesos_i(14581) := b"1111111111111111_1111111111111111_1101110110110110_0011000011001100"; -- -0.1339387418274031
	pesos_i(14582) := b"0000000000000000_0000000000000000_0000011111001110_1001111001100010"; -- 0.030496500988537033
	pesos_i(14583) := b"1111111111111111_1111111111111111_1110010111110101_1101011111011011"; -- -0.10171748071877619
	pesos_i(14584) := b"0000000000000000_0000000000000000_0001101111010001_0110111100101010"; -- 0.10866446269721436
	pesos_i(14585) := b"1111111111111111_1111111111111111_1111101100011010_1100000010011100"; -- -0.019123041071335046
	pesos_i(14586) := b"1111111111111111_1111111111111111_1110101010111111_0011111010111101"; -- -0.08301933173172756
	pesos_i(14587) := b"0000000000000000_0000000000000000_0001011100101011_0010110000000111"; -- 0.0905025021468415
	pesos_i(14588) := b"0000000000000000_0000000000000000_0000000010100000_1110000100011110"; -- 0.0024548242835393404
	pesos_i(14589) := b"0000000000000000_0000000000000000_0001010100011011_0100110010001100"; -- 0.08244779979681863
	pesos_i(14590) := b"1111111111111111_1111111111111111_1110101111100000_1001010011000101"; -- -0.07860441393991796
	pesos_i(14591) := b"0000000000000000_0000000000000000_0000100101100101_1111111010111010"; -- 0.03671257057375727
	pesos_i(14592) := b"1111111111111111_1111111111111111_1111000110001101_0100000110001010"; -- -0.056438354423247204
	pesos_i(14593) := b"1111111111111111_1111111111111111_1101110011001100_0111011111000100"; -- -0.13750506836501405
	pesos_i(14594) := b"0000000000000000_0000000000000000_0001011100000101_0010010100111100"; -- 0.08992226326093526
	pesos_i(14595) := b"1111111111111111_1111111111111111_1110011100100001_0010100100010111"; -- -0.09715026088588366
	pesos_i(14596) := b"1111111111111111_1111111111111111_1111010110000011_1000101101010110"; -- -0.04096154357856714
	pesos_i(14597) := b"0000000000000000_0000000000000000_0001001110011011_1000011111100011"; -- 0.07659196170979864
	pesos_i(14598) := b"1111111111111111_1111111111111111_1110110101011100_0110001111111100"; -- -0.07280898190530642
	pesos_i(14599) := b"0000000000000000_0000000000000000_0000111110010010_0001100011100001"; -- 0.060823016183974614
	pesos_i(14600) := b"0000000000000000_0000000000000000_0001001111011101_0010001111011101"; -- 0.07759308004970653
	pesos_i(14601) := b"0000000000000000_0000000000000000_0001000001110110_1010011001111101"; -- 0.06431046069450759
	pesos_i(14602) := b"1111111111111111_1111111111111111_1110001011110100_1100011111010000"; -- -0.11345244570687113
	pesos_i(14603) := b"1111111111111111_1111111111111111_1110110010010000_1000001010111111"; -- -0.07591994121306414
	pesos_i(14604) := b"1111111111111111_1111111111111111_1111001111010111_1010001100001010"; -- -0.047490892514299166
	pesos_i(14605) := b"1111111111111111_1111111111111111_1111111011010100_1100101011101110"; -- -0.004565541241510654
	pesos_i(14606) := b"0000000000000000_0000000000000000_0010001011000111_1010000000101001"; -- 0.13585854530569563
	pesos_i(14607) := b"0000000000000000_0000000000000000_0001001001100101_1111110011101001"; -- 0.07186871230310249
	pesos_i(14608) := b"0000000000000000_0000000000000000_0000110001111000_1010100110011001"; -- 0.04871616343100621
	pesos_i(14609) := b"1111111111111111_1111111111111111_1111000001000110_1110000101001001"; -- -0.06141845663050674
	pesos_i(14610) := b"0000000000000000_0000000000000000_0000101000101100_1010100101111100"; -- 0.03974398879342932
	pesos_i(14611) := b"1111111111111111_1111111111111111_1111001011111000_0010111011011011"; -- -0.050900527608791116
	pesos_i(14612) := b"0000000000000000_0000000000000000_0010100011010010_0010001111110010"; -- 0.15945648812164057
	pesos_i(14613) := b"1111111111111111_1111111111111111_1101111010001100_1001000100111111"; -- -0.13066761214385844
	pesos_i(14614) := b"0000000000000000_0000000000000000_0001100111110010_0100000111111001"; -- 0.10135280927530531
	pesos_i(14615) := b"1111111111111111_1111111111111111_1110111101111101_1000000000101111"; -- -0.06449126105475406
	pesos_i(14616) := b"0000000000000000_0000000000000000_0001111010111011_1100111110111101"; -- 0.12005327569180703
	pesos_i(14617) := b"0000000000000000_0000000000000000_0000010000011010_1101101010000101"; -- 0.01603475327508159
	pesos_i(14618) := b"1111111111111111_1111111111111111_1110000100111001_0110100010100000"; -- -0.12021776291087756
	pesos_i(14619) := b"0000000000000000_0000000000000000_0000111110011110_1001111101101001"; -- 0.061014140181648205
	pesos_i(14620) := b"1111111111111111_1111111111111111_1111011001100010_1011110010111110"; -- -0.037555888811913005
	pesos_i(14621) := b"1111111111111111_1111111111111111_1110101110110101_1010010110001011"; -- -0.07925954202969465
	pesos_i(14622) := b"0000000000000000_0000000000000000_0000100000100101_1001100000111111"; -- 0.0318236497637898
	pesos_i(14623) := b"1111111111111111_1111111111111111_1111001011010111_1100001111110111"; -- -0.05139517995672668
	pesos_i(14624) := b"1111111111111111_1111111111111111_1111101110101000_1101011010101101"; -- -0.01695497784873754
	pesos_i(14625) := b"0000000000000000_0000000000000000_0000011110000110_1001000100110010"; -- 0.0293970821393957
	pesos_i(14626) := b"0000000000000000_0000000000000000_0010000111111110_1000101011111011"; -- 0.13279026639130112
	pesos_i(14627) := b"0000000000000000_0000000000000000_0010100010101001_1000111011101101"; -- 0.15883725448641003
	pesos_i(14628) := b"1111111111111111_1111111111111111_1111001000011101_0110100000100000"; -- -0.054238788718821034
	pesos_i(14629) := b"0000000000000000_0000000000000000_0001100101100100_1001100001100010"; -- 0.09919121167335936
	pesos_i(14630) := b"1111111111111111_1111111111111111_1110011111110010_0110100010111010"; -- -0.09395738085079645
	pesos_i(14631) := b"0000000000000000_0000000000000000_0001000001011110_0100010011000010"; -- 0.06393842453695091
	pesos_i(14632) := b"0000000000000000_0000000000000000_0010011101000111_1111101000011100"; -- 0.15344203159395392
	pesos_i(14633) := b"1111111111111111_1111111111111111_1110000011010110_0000010000011100"; -- -0.12173437417026962
	pesos_i(14634) := b"1111111111111111_1111111111111111_1101101011100110_1111001010101110"; -- -0.14491351370877992
	pesos_i(14635) := b"0000000000000000_0000000000000000_0000000011010100_1010001011011101"; -- 0.0032445707575072787
	pesos_i(14636) := b"1111111111111111_1111111111111111_1111100010011011_0100000001001110"; -- -0.028881054848148433
	pesos_i(14637) := b"0000000000000000_0000000000000000_0001010010110101_0100000010101000"; -- 0.08089069461857422
	pesos_i(14638) := b"0000000000000000_0000000000000000_0000100101100100_1101001010010000"; -- 0.03669467945057664
	pesos_i(14639) := b"1111111111111111_1111111111111111_1110111110010110_0111011110101000"; -- -0.06411029962773988
	pesos_i(14640) := b"1111111111111111_1111111111111111_1111000110001101_1001011110110011"; -- -0.056433218772259014
	pesos_i(14641) := b"0000000000000000_0000000000000000_0001100111110011_1101001101101101"; -- 0.10137673771700738
	pesos_i(14642) := b"0000000000000000_0000000000000000_0000001100001100_0010001010011010"; -- 0.011903917892482858
	pesos_i(14643) := b"0000000000000000_0000000000000000_0000000000101001_0000110000110011"; -- 0.0006263375112752496
	pesos_i(14644) := b"1111111111111111_1111111111111111_1111001011010011_0111010001110110"; -- -0.0514609538885702
	pesos_i(14645) := b"0000000000000000_0000000000000000_0000011101000110_1111000011110011"; -- 0.02842622689059666
	pesos_i(14646) := b"1111111111111111_1111111111111111_1111110001000100_0111110100101111"; -- -0.014579940754067254
	pesos_i(14647) := b"1111111111111111_1111111111111111_1111100110101011_0010111010010100"; -- -0.02473172083198974
	pesos_i(14648) := b"0000000000000000_0000000000000000_0001100100010111_0101000110100010"; -- 0.09801206787239378
	pesos_i(14649) := b"1111111111111111_1111111111111111_1110110010100111_0101101001011111"; -- -0.07557139570823097
	pesos_i(14650) := b"0000000000000000_0000000000000000_0010000010001110_1100001011000110"; -- 0.1271783574612893
	pesos_i(14651) := b"1111111111111111_1111111111111111_1110000111010011_0011000100111110"; -- -0.11787121035008503
	pesos_i(14652) := b"1111111111111111_1111111111111111_1110000110001011_0111110001010111"; -- -0.118965367070743
	pesos_i(14653) := b"0000000000000000_0000000000000000_0000101111101010_1111101100101101"; -- 0.04655427793352598
	pesos_i(14654) := b"0000000000000000_0000000000000000_0000101000100100_0000000011100001"; -- 0.03961186875265862
	pesos_i(14655) := b"0000000000000000_0000000000000000_0001111000000110_0001010101110111"; -- 0.11728033219596379
	pesos_i(14656) := b"0000000000000000_0000000000000000_0001011001110100_1001001100100001"; -- 0.08771628916503679
	pesos_i(14657) := b"1111111111111111_1111111111111111_1110111100100110_1111000101010101"; -- -0.06581203142640536
	pesos_i(14658) := b"1111111111111111_1111111111111111_1110100000101100_1011001011000111"; -- -0.09306795739219766
	pesos_i(14659) := b"0000000000000000_0000000000000000_0010010010101110_1101101110101010"; -- 0.14329312227191174
	pesos_i(14660) := b"0000000000000000_0000000000000000_0000101110001011_1101001011110110"; -- 0.045102296033332594
	pesos_i(14661) := b"1111111111111111_1111111111111111_1110001011011001_1000010110111101"; -- -0.11386837144919826
	pesos_i(14662) := b"1111111111111111_1111111111111111_1101110011011111_1001011010010110"; -- -0.13721331440489568
	pesos_i(14663) := b"1111111111111111_1111111111111111_1110100011111001_1111011100110111"; -- -0.08993582640109396
	pesos_i(14664) := b"1111111111111111_1111111111111111_1110101111101110_1101100000010100"; -- -0.07838677884193682
	pesos_i(14665) := b"0000000000000000_0000000000000000_0001011011011000_0100100010001000"; -- 0.08923772174769544
	pesos_i(14666) := b"1111111111111111_1111111111111111_1110000001010011_0000100110101000"; -- -0.12373294504639068
	pesos_i(14667) := b"0000000000000000_0000000000000000_0000001011110001_0010001001001010"; -- 0.011491912005284226
	pesos_i(14668) := b"0000000000000000_0000000000000000_0000011010011011_1011110101001001"; -- 0.025813894671370182
	pesos_i(14669) := b"0000000000000000_0000000000000000_0001001100110110_0101010101110000"; -- 0.07504781697859418
	pesos_i(14670) := b"1111111111111111_1111111111111111_1111001001111011_1001100110010100"; -- -0.052801515090664386
	pesos_i(14671) := b"1111111111111111_1111111111111111_1110001111110011_0011111110111010"; -- -0.10956956580700952
	pesos_i(14672) := b"1111111111111111_1111111111111111_1111011000111110_0001111011101110"; -- -0.03811461146128361
	pesos_i(14673) := b"1111111111111111_1111111111111111_1110100001010000_0110101010101101"; -- -0.09252293855490798
	pesos_i(14674) := b"0000000000000000_0000000000000000_0000101011011011_1001010000000000"; -- 0.04241299627633904
	pesos_i(14675) := b"1111111111111111_1111111111111111_1110010111011100_0001000101000100"; -- -0.10211078721784649
	pesos_i(14676) := b"0000000000000000_0000000000000000_0001111011001000_1011110101100111"; -- 0.12025054709975518
	pesos_i(14677) := b"1111111111111111_1111111111111111_1101101111011011_0101010011011100"; -- -0.14118451713425006
	pesos_i(14678) := b"1111111111111111_1111111111111111_1101111010001010_1011000000011110"; -- -0.1306962897347331
	pesos_i(14679) := b"1111111111111111_1111111111111111_1111100101001110_1101000110001000"; -- -0.026141075453515794
	pesos_i(14680) := b"1111111111111111_1111111111111111_1110110010111110_0100000111001001"; -- -0.07522190892313771
	pesos_i(14681) := b"1111111111111111_1111111111111111_1110111100101100_1110001110111110"; -- -0.06572128877579743
	pesos_i(14682) := b"0000000000000000_0000000000000000_0010001000100011_1101100010001110"; -- 0.1333594652004522
	pesos_i(14683) := b"0000000000000000_0000000000000000_0000111100101010_1101111100011100"; -- 0.05924791753058915
	pesos_i(14684) := b"0000000000000000_0000000000000000_0001100100110110_1100010111001000"; -- 0.09849201325311284
	pesos_i(14685) := b"0000000000000000_0000000000000000_0010000110110000_1000001000111001"; -- 0.13159955874420798
	pesos_i(14686) := b"1111111111111111_1111111111111111_1101011001010111_0101110100110010"; -- -0.1627294305630238
	pesos_i(14687) := b"0000000000000000_0000000000000000_0001001110011100_1100101100101011"; -- 0.0766112307562805
	pesos_i(14688) := b"0000000000000000_0000000000000000_0010000000111011_0001111010000010"; -- 0.1259020869801718
	pesos_i(14689) := b"1111111111111111_1111111111111111_1101111000010010_0000101111111101"; -- -0.13253712716675406
	pesos_i(14690) := b"0000000000000000_0000000000000000_0001110001101100_1000001001110110"; -- 0.11103072524776873
	pesos_i(14691) := b"1111111111111111_1111111111111111_1110011000110011_0010101111100111"; -- -0.10078168496444063
	pesos_i(14692) := b"1111111111111111_1111111111111111_1110011111100111_0001101101000110"; -- -0.09412984414475022
	pesos_i(14693) := b"0000000000000000_0000000000000000_0010010111100111_0011100011001100"; -- 0.14805941569647868
	pesos_i(14694) := b"1111111111111111_1111111111111111_1111000100010110_1000111111011001"; -- -0.05824948260021073
	pesos_i(14695) := b"1111111111111111_1111111111111111_1110100010011011_1001111011011111"; -- -0.09137541835162653
	pesos_i(14696) := b"0000000000000000_0000000000000000_0000100000000101_1100111111111111"; -- 0.031338691556425005
	pesos_i(14697) := b"0000000000000000_0000000000000000_0001111011000010_0011000100000111"; -- 0.12015062736382495
	pesos_i(14698) := b"1111111111111111_1111111111111111_1111100000110110_1100111001100000"; -- -0.030413724381291203
	pesos_i(14699) := b"1111111111111111_1111111111111111_1110100111010101_1011101100100010"; -- -0.08658247391491153
	pesos_i(14700) := b"1111111111111111_1111111111111111_1110000100010001_0110000001011000"; -- -0.12082860795741883
	pesos_i(14701) := b"1111111111111111_1111111111111111_1110111000011110_1111111001010100"; -- -0.06983957710418545
	pesos_i(14702) := b"1111111111111111_1111111111111111_1110000010111000_0011000011010100"; -- -0.12218947254256644
	pesos_i(14703) := b"1111111111111111_1111111111111111_1110110010011110_0011010101010000"; -- -0.07571093368001997
	pesos_i(14704) := b"1111111111111111_1111111111111111_1110001001110111_1000101011111101"; -- -0.11536341968784458
	pesos_i(14705) := b"1111111111111111_1111111111111111_1111111000101011_1010110110100101"; -- -0.007146022059315085
	pesos_i(14706) := b"1111111111111111_1111111111111111_1111011111001100_1000100001000111"; -- -0.032035334382774935
	pesos_i(14707) := b"0000000000000000_0000000000000000_0010010010000110_0001011011101101"; -- 0.1426710441945335
	pesos_i(14708) := b"0000000000000000_0000000000000000_0000001100010000_1100010100100110"; -- 0.011974641508795002
	pesos_i(14709) := b"0000000000000000_0000000000000000_0001100100011010_0000110110100111"; -- 0.09805379228914489
	pesos_i(14710) := b"1111111111111111_1111111111111111_1110011101000110_1100011110000001"; -- -0.09657624340545976
	pesos_i(14711) := b"1111111111111111_1111111111111111_1101110011010101_1011001000110111"; -- -0.13736425555057122
	pesos_i(14712) := b"1111111111111111_1111111111111111_1111100101010111_1000110110011011"; -- -0.026007794935829685
	pesos_i(14713) := b"0000000000000000_0000000000000000_0000110001011101_0011010110011101"; -- 0.0482972630330701
	pesos_i(14714) := b"0000000000000000_0000000000000000_0010110010000111_0010010000100111"; -- 0.17393709135413093
	pesos_i(14715) := b"1111111111111111_1111111111111111_1110010111011000_0100110001100000"; -- -0.1021682992252418
	pesos_i(14716) := b"0000000000000000_0000000000000000_0001110110010101_1100011011110010"; -- 0.11556666756376606
	pesos_i(14717) := b"1111111111111111_1111111111111111_1110110101101100_0010011010100111"; -- -0.07256849688824338
	pesos_i(14718) := b"0000000000000000_0000000000000000_0000111000100110_1000001001111001"; -- 0.05527511083140633
	pesos_i(14719) := b"0000000000000000_0000000000000000_0001011000000000_0001001010001010"; -- 0.08593860494938074
	pesos_i(14720) := b"1111111111111111_1111111111111111_1110010110001011_1010110111011001"; -- -0.10333741613428471
	pesos_i(14721) := b"0000000000000000_0000000000000000_0000101111001000_0111010111101111"; -- 0.046027537202256226
	pesos_i(14722) := b"0000000000000000_0000000000000000_0001110000100001_0011100111000110"; -- 0.10988198366737095
	pesos_i(14723) := b"0000000000000000_0000000000000000_0001101101010001_1101011000000010"; -- 0.1067174677933618
	pesos_i(14724) := b"1111111111111111_1111111111111111_1110001010100100_0000111111111001"; -- -0.11468410648063929
	pesos_i(14725) := b"0000000000000000_0000000000000000_0001010110011011_1011011000111100"; -- 0.08440722429644093
	pesos_i(14726) := b"0000000000000000_0000000000000000_0001111001000110_1111001001110111"; -- 0.11827006717176881
	pesos_i(14727) := b"0000000000000000_0000000000000000_0001000000000010_0011100000010000"; -- 0.06253385905984526
	pesos_i(14728) := b"0000000000000000_0000000000000000_0001101010100011_0010011100100001"; -- 0.10405201484223536
	pesos_i(14729) := b"1111111111111111_1111111111111111_1101101010110010_0110011000011101"; -- -0.14571534912051937
	pesos_i(14730) := b"1111111111111111_1111111111111111_1110011100110101_1111100101001101"; -- -0.09683267472300208
	pesos_i(14731) := b"1111111111111111_1111111111111111_1110000001110100_1110000110000110"; -- -0.12321653814880075
	pesos_i(14732) := b"1111111111111111_1111111111111111_1111010001111000_0101101110001101"; -- -0.04503848850475002
	pesos_i(14733) := b"0000000000000000_0000000000000000_0001110011101010_0101111000100010"; -- 0.11295116732425473
	pesos_i(14734) := b"0000000000000000_0000000000000000_0000000100011001_0001001000001100"; -- 0.004288795520067567
	pesos_i(14735) := b"0000000000000000_0000000000000000_0001011100100010_0001001011001110"; -- 0.090363669620937
	pesos_i(14736) := b"1111111111111111_1111111111111111_1110101111001011_0010011000010100"; -- -0.07893144611398656
	pesos_i(14737) := b"0000000000000000_0000000000000000_0010001010101101_0110011000111011"; -- 0.13545836384368595
	pesos_i(14738) := b"1111111111111111_1111111111111111_1110000101101110_1010001011000110"; -- -0.1194055812311487
	pesos_i(14739) := b"1111111111111111_1111111111111111_1101111101011110_0011000110111001"; -- -0.12746896003881983
	pesos_i(14740) := b"0000000000000000_0000000000000000_0000011111011011_0000111010000110"; -- 0.030686290475344755
	pesos_i(14741) := b"0000000000000000_0000000000000000_0001100101101101_0101011101010010"; -- 0.09932466275263296
	pesos_i(14742) := b"0000000000000000_0000000000000000_0001100101110000_0000010100001010"; -- 0.0993655348342641
	pesos_i(14743) := b"0000000000000000_0000000000000000_0001001110101000_1101000000110100"; -- 0.07679463639844801
	pesos_i(14744) := b"1111111111111111_1111111111111111_1111111101001010_0011101000110111"; -- -0.002773629638263482
	pesos_i(14745) := b"1111111111111111_1111111111111111_1110100010110111_0101100110101100"; -- -0.09095229675018429
	pesos_i(14746) := b"0000000000000000_0000000000000000_0001101011100110_0010000111001000"; -- 0.1050740351002321
	pesos_i(14747) := b"0000000000000000_0000000000000000_0001111110000001_1111100010000100"; -- 0.12307694642851015
	pesos_i(14748) := b"1111111111111111_1111111111111111_1111110001010011_1110000000010000"; -- -0.014345165455755433
	pesos_i(14749) := b"1111111111111111_1111111111111111_1111000001001010_1100100100000100"; -- -0.061358868104655094
	pesos_i(14750) := b"1111111111111111_1111111111111111_1110100011000011_0101001001000011"; -- -0.09076963288386498
	pesos_i(14751) := b"1111111111111111_1111111111111111_1111100101011010_1011010111110011"; -- -0.025959613948860517
	pesos_i(14752) := b"0000000000000000_0000000000000000_0000111010111001_0110000000101001"; -- 0.057516107650898006
	pesos_i(14753) := b"1111111111111111_1111111111111111_1110110000000110_0010100101100100"; -- -0.07803098023911993
	pesos_i(14754) := b"1111111111111111_1111111111111111_1111010010010101_1100010000100011"; -- -0.044589749822395906
	pesos_i(14755) := b"1111111111111111_1111111111111111_1110110110110000_0001110000101010"; -- -0.07153152444912259
	pesos_i(14756) := b"0000000000000000_0000000000000000_0001111100110100_1000100001111011"; -- 0.1218953420085736
	pesos_i(14757) := b"0000000000000000_0000000000000000_0001010100010110_0010001011100111"; -- 0.08236902381186262
	pesos_i(14758) := b"0000000000000000_0000000000000000_0001110011110111_0110010101010100"; -- 0.11314996050759733
	pesos_i(14759) := b"1111111111111111_1111111111111111_1110100001111111_0011110111100000"; -- -0.09180844586344306
	pesos_i(14760) := b"0000000000000000_0000000000000000_0010001110001011_1111000101100101"; -- 0.13885410993764558
	pesos_i(14761) := b"1111111111111111_1111111111111111_1111111010101110_0000100100111110"; -- -0.005156919730183237
	pesos_i(14762) := b"0000000000000000_0000000000000000_0000100101110110_1001001001000010"; -- 0.036965504820931035
	pesos_i(14763) := b"0000000000000000_0000000000000000_0001111100100111_0010011011001111"; -- 0.12169115604077402
	pesos_i(14764) := b"1111111111111111_1111111111111111_1101111101011000_0011001001010101"; -- -0.12756047663185668
	pesos_i(14765) := b"1111111111111111_1111111111111111_1110111001111101_1001110010100101"; -- -0.06839581459278765
	pesos_i(14766) := b"0000000000000000_0000000000000000_0000001001001100_1101110010110100"; -- 0.00898532295048471
	pesos_i(14767) := b"1111111111111111_1111111111111111_1111000100101100_1001000011001000"; -- -0.05791373372803787
	pesos_i(14768) := b"0000000000000000_0000000000000000_0001100000111011_1011011111001101"; -- 0.09466122385670112
	pesos_i(14769) := b"1111111111111111_1111111111111111_1101111011010101_0010001110101101"; -- -0.12956025138015187
	pesos_i(14770) := b"0000000000000000_0000000000000000_0001100011100100_0110101011011000"; -- 0.09723537224133144
	pesos_i(14771) := b"0000000000000000_0000000000000000_0001100111110111_1001101001110101"; -- 0.10143437736144557
	pesos_i(14772) := b"1111111111111111_1111111111111111_1111100011111101_1100001111110001"; -- -0.027377847377784294
	pesos_i(14773) := b"1111111111111111_1111111111111111_1110111011100100_0100000011110001"; -- -0.06682962537304125
	pesos_i(14774) := b"0000000000000000_0000000000000000_0000100110100011_0001011011111101"; -- 0.037644802860543086
	pesos_i(14775) := b"0000000000000000_0000000000000000_0000011010001010_0100110011101011"; -- 0.02554779751432597
	pesos_i(14776) := b"0000000000000000_0000000000000000_0000111011100110_1000001000011001"; -- 0.05820477594396353
	pesos_i(14777) := b"1111111111111111_1111111111111111_1101110001111101_1110111100101001"; -- -0.13870339642086016
	pesos_i(14778) := b"1111111111111111_1111111111111111_1101110010111100_1000010111001111"; -- -0.13774837208252683
	pesos_i(14779) := b"0000000000000000_0000000000000000_0010010110111100_0001011110111100"; -- 0.14740131705677897
	pesos_i(14780) := b"1111111111111111_1111111111111111_1111001110100011_0101011110110110"; -- -0.048288839327136186
	pesos_i(14781) := b"0000000000000000_0000000000000000_0000101111101000_1001010111001110"; -- 0.046517718008273
	pesos_i(14782) := b"0000000000000000_0000000000000000_0000011100100101_0110111101000101"; -- 0.027914957334270424
	pesos_i(14783) := b"0000000000000000_0000000000000000_0001110100011111_1100010011111001"; -- 0.11376601294834494
	pesos_i(14784) := b"0000000000000000_0000000000000000_0000000111011000_1101000011100110"; -- 0.007214599837698602
	pesos_i(14785) := b"0000000000000000_0000000000000000_0001001010101011_1100000100101111"; -- 0.0729332675685564
	pesos_i(14786) := b"1111111111111111_1111111111111111_1110110111000001_1010010101110001"; -- -0.07126394252602884
	pesos_i(14787) := b"1111111111111111_1111111111111111_1101111100011001_0100100111011100"; -- -0.12852037796702745
	pesos_i(14788) := b"0000000000000000_0000000000000000_0001001111011101_1111101001000101"; -- 0.07760585950734888
	pesos_i(14789) := b"1111111111111111_1111111111111111_1111011001011000_0100001100100001"; -- -0.03771572528252775
	pesos_i(14790) := b"1111111111111111_1111111111111111_1111111011101100_1010001001111101"; -- -0.004201740831675097
	pesos_i(14791) := b"1111111111111111_1111111111111111_1111001011010010_1001001111000101"; -- -0.051474346435361654
	pesos_i(14792) := b"1111111111111111_1111111111111111_1110001110111100_0101010001101101"; -- -0.11040756541000225
	pesos_i(14793) := b"1111111111111111_1111111111111111_1110101011010000_1101100100011100"; -- -0.08275073105325152
	pesos_i(14794) := b"0000000000000000_0000000000000000_0000111000101000_0011001100001000"; -- 0.05530089330707987
	pesos_i(14795) := b"0000000000000000_0000000000000000_0001110010000000_0110011000101001"; -- 0.11133421429712864
	pesos_i(14796) := b"1111111111111111_1111111111111111_1110101000001001_1111111011010101"; -- -0.08578498183626189
	pesos_i(14797) := b"1111111111111111_1111111111111111_1101110111001001_0011100001111001"; -- -0.13364836729227042
	pesos_i(14798) := b"1111111111111111_1111111111111111_1111000000011111_1101010001111100"; -- -0.06201431248620958
	pesos_i(14799) := b"0000000000000000_0000000000000000_0000010111010000_1010001110001111"; -- 0.022714826921356818
	pesos_i(14800) := b"1111111111111111_1111111111111111_1111110110111001_0000100001101001"; -- -0.00889537276374248
	pesos_i(14801) := b"0000000000000000_0000000000000000_0001100000110100_1100000011001110"; -- 0.09455494903794368
	pesos_i(14802) := b"1111111111111111_1111111111111111_1111110001011000_0001111001001001"; -- -0.014280421530962584
	pesos_i(14803) := b"1111111111111111_1111111111111111_1110110001100011_0100000100100100"; -- -0.0766104972277129
	pesos_i(14804) := b"1111111111111111_1111111111111111_1110010000111100_1011000011011110"; -- -0.10844893061778846
	pesos_i(14805) := b"1111111111111111_1111111111111111_1110011000110001_1110101100000000"; -- -0.10080081215676771
	pesos_i(14806) := b"1111111111111111_1111111111111111_1110101110011101_0000110010001001"; -- -0.07963487295895001
	pesos_i(14807) := b"1111111111111111_1111111111111111_1110101010100010_0110011001111100"; -- -0.08345946768302902
	pesos_i(14808) := b"0000000000000000_0000000000000000_0001000011010100_1101000111001011"; -- 0.06574736796348399
	pesos_i(14809) := b"1111111111111111_1111111111111111_1110010001001100_0010000001110011"; -- -0.10821339784102822
	pesos_i(14810) := b"1111111111111111_1111111111111111_1110011010110111_0101100111010101"; -- -0.09876478721702299
	pesos_i(14811) := b"0000000000000000_0000000000000000_0010010010001010_0011000101001010"; -- 0.14273365084993014
	pesos_i(14812) := b"0000000000000000_0000000000000000_0000011101110110_0100111111101100"; -- 0.029149050822245448
	pesos_i(14813) := b"1111111111111111_1111111111111111_1101101010000100_1111111000100111"; -- -0.14640819107881817
	pesos_i(14814) := b"1111111111111111_1111111111111111_1111001001100001_0001101000101100"; -- -0.053205837391300304
	pesos_i(14815) := b"1111111111111111_1111111111111111_1110110011101010_1111010100011010"; -- -0.07453983407846262
	pesos_i(14816) := b"1111111111111111_1111111111111111_1101101001101101_0011000001001110"; -- -0.1467714128878849
	pesos_i(14817) := b"1111111111111111_1111111111111111_1111011010010100_0000100000010101"; -- -0.03680371741449256
	pesos_i(14818) := b"0000000000000000_0000000000000000_0001001010001011_0000111111001000"; -- 0.07243441230303377
	pesos_i(14819) := b"1111111111111111_1111111111111111_1110001000011111_1011110011010001"; -- -0.11670322326888571
	pesos_i(14820) := b"0000000000000000_0000000000000000_0000110001000100_1110010101111111"; -- 0.04792627671803611
	pesos_i(14821) := b"0000000000000000_0000000000000000_0000111001011111_0110000101111001"; -- 0.05614289488790534
	pesos_i(14822) := b"0000000000000000_0000000000000000_0001000110000011_1001101110110001"; -- 0.06841443131304413
	pesos_i(14823) := b"0000000000000000_0000000000000000_0001100101010111_1001101001101111"; -- 0.09899296972180455
	pesos_i(14824) := b"1111111111111111_1111111111111111_1111101110000101_1010000000001001"; -- -0.01749229213331737
	pesos_i(14825) := b"1111111111111111_1111111111111111_1110100011110011_0001101110101010"; -- -0.09004046525242197
	pesos_i(14826) := b"0000000000000000_0000000000000000_0000000101010111_1100111110111110"; -- 0.005246147051899895
	pesos_i(14827) := b"0000000000000000_0000000000000000_0001111000111111_1001011111110010"; -- 0.11815786041105142
	pesos_i(14828) := b"1111111111111111_1111111111111111_1101110001010001_1101101110000101"; -- -0.13937595368315242
	pesos_i(14829) := b"1111111111111111_1111111111111111_1110100110101000_0110000001000111"; -- -0.0872745347879874
	pesos_i(14830) := b"0000000000000000_0000000000000000_0000001010000111_1100101100010011"; -- 0.009884540780039879
	pesos_i(14831) := b"1111111111111111_1111111111111111_1110100101110011_0111010000001111"; -- -0.08808207165131503
	pesos_i(14832) := b"0000000000000000_0000000000000000_0000010001010101_1101111000100111"; -- 0.016935238401966375
	pesos_i(14833) := b"1111111111111111_1111111111111111_1110100100111101_0001101111000111"; -- -0.08891130817139775
	pesos_i(14834) := b"1111111111111111_1111111111111111_1110010001101101_1001000010011000"; -- -0.10770317349767204
	pesos_i(14835) := b"0000000000000000_0000000000000000_0000110111111100_0111100110001010"; -- 0.05463370923594019
	pesos_i(14836) := b"1111111111111111_1111111111111111_1101110111110010_0111100010101111"; -- -0.1330189297135742
	pesos_i(14837) := b"1111111111111111_1111111111111111_1111110010100101_0011100110000011"; -- -0.013103871801484014
	pesos_i(14838) := b"1111111111111111_1111111111111111_1101101100000101_1110101011100001"; -- -0.1444409562107872
	pesos_i(14839) := b"1111111111111111_1111111111111111_1110111101110111_1110111100111100"; -- -0.06457619466667495
	pesos_i(14840) := b"0000000000000000_0000000000000000_0001110010100110_1000000011100111"; -- 0.11191564214032738
	pesos_i(14841) := b"0000000000000000_0000000000000000_0001101100011001_0110010101100001"; -- 0.10585626237400694
	pesos_i(14842) := b"0000000000000000_0000000000000000_0000001010000111_1110101000000110"; -- 0.00988638535976871
	pesos_i(14843) := b"0000000000000000_0000000000000000_0001011100110110_0101110001001011"; -- 0.09067322562722845
	pesos_i(14844) := b"1111111111111111_1111111111111111_1110110101111011_1101011001000001"; -- -0.07232914848061506
	pesos_i(14845) := b"0000000000000000_0000000000000000_0000000100001010_0001001100101111"; -- 0.004059981402991341
	pesos_i(14846) := b"0000000000000000_0000000000000000_0000011011011011_0010010110101100"; -- 0.026781420200050803
	pesos_i(14847) := b"1111111111111111_1111111111111111_1110100100001011_1001000110111000"; -- -0.08966721780924729
	pesos_i(14848) := b"0000000000000000_0000000000000000_0001101000010010_1011101000000011"; -- 0.10184824528192295
	pesos_i(14849) := b"1111111111111111_1111111111111111_1111100100110011_1110010111110000"; -- -0.02655184644333763
	pesos_i(14850) := b"1111111111111111_1111111111111111_1110001101001000_0111101100110100"; -- -0.11217527366032409
	pesos_i(14851) := b"0000000000000000_0000000000000000_0000111001000100_0011011100110000"; -- 0.055728386982073747
	pesos_i(14852) := b"1111111111111111_1111111111111111_1110001011000100_1100111110111010"; -- -0.1141843958361604
	pesos_i(14853) := b"1111111111111111_1111111111111111_1111111101010111_0111101101110100"; -- -0.0025713770445905493
	pesos_i(14854) := b"0000000000000000_0000000000000000_0000110010010111_1011100111011110"; -- 0.049190155785993596
	pesos_i(14855) := b"1111111111111111_1111111111111111_1110100101010111_1000101000011111"; -- -0.08850800258094078
	pesos_i(14856) := b"1111111111111111_1111111111111111_1110011110010001_1111011110011110"; -- -0.0954289665409992
	pesos_i(14857) := b"1111111111111111_1111111111111111_1110111110101100_0111110001011000"; -- -0.06377432671969427
	pesos_i(14858) := b"0000000000000000_0000000000000000_0001100100010111_0101000011011010"; -- 0.09801202116847446
	pesos_i(14859) := b"1111111111111111_1111111111111111_1110001000011101_0001000010011001"; -- -0.11674400593213244
	pesos_i(14860) := b"0000000000000000_0000000000000000_0000110100111111_1010111100100011"; -- 0.051752992634949535
	pesos_i(14861) := b"1111111111111111_1111111111111111_1101111011101100_1011011100110000"; -- -0.12920050704690647
	pesos_i(14862) := b"0000000000000000_0000000000000000_0001100011010001_0010011110111100"; -- 0.09694145528226851
	pesos_i(14863) := b"1111111111111111_1111111111111111_1110000011110011_1110100111111000"; -- -0.12127816868718702
	pesos_i(14864) := b"0000000000000000_0000000000000000_0001011000110010_1001000111101010"; -- 0.08670913655327286
	pesos_i(14865) := b"1111111111111111_1111111111111111_1111111000011011_0011101001010001"; -- -0.007397036834629951
	pesos_i(14866) := b"0000000000000000_0000000000000000_0000011011011010_1001100101011001"; -- 0.026773056137007777
	pesos_i(14867) := b"0000000000000000_0000000000000000_0000101011111110_0011111101011001"; -- 0.042942008264590374
	pesos_i(14868) := b"1111111111111111_1111111111111111_1101100110111001_1111000111110101"; -- -0.14950645221546757
	pesos_i(14869) := b"0000000000000000_0000000000000000_0010010100001110_0101100100011011"; -- 0.14475018423931135
	pesos_i(14870) := b"1111111111111111_1111111111111111_1110101101010110_1011010110110010"; -- -0.0807081642706156
	pesos_i(14871) := b"1111111111111111_1111111111111111_1110111111000111_0100100001000100"; -- -0.06336544358492407
	pesos_i(14872) := b"0000000000000000_0000000000000000_0000011000101110_0001000010001011"; -- 0.024140390227330607
	pesos_i(14873) := b"1111111111111111_1111111111111111_1101111001001110_1010010110010010"; -- -0.13161244565506935
	pesos_i(14874) := b"0000000000000000_0000000000000000_0001001110100011_0011011111111101"; -- 0.07670926967125113
	pesos_i(14875) := b"0000000000000000_0000000000000000_0010000101011011_0000010111110111"; -- 0.13029515538317657
	pesos_i(14876) := b"0000000000000000_0000000000000000_0001101111111101_1110111110000100"; -- 0.10934349989719669
	pesos_i(14877) := b"0000000000000000_0000000000000000_0000011110110110_1110000100001100"; -- 0.03013426349680581
	pesos_i(14878) := b"0000000000000000_0000000000000000_0001100011010010_1001000100000111"; -- 0.0969629900979602
	pesos_i(14879) := b"1111111111111111_1111111111111111_1101110101001110_0001001111100100"; -- -0.1355273787855174
	pesos_i(14880) := b"0000000000000000_0000000000000000_0000000111011000_1000110001011000"; -- 0.007210513639868191
	pesos_i(14881) := b"1111111111111111_1111111111111111_1111010010110011_1010101000101101"; -- -0.04413353347312099
	pesos_i(14882) := b"0000000000000000_0000000000000000_0001111111100001_1100000110110111"; -- 0.12453852375078057
	pesos_i(14883) := b"0000000000000000_0000000000000000_0000111000111000_0101001100110010"; -- 0.055546950917450225
	pesos_i(14884) := b"0000000000000000_0000000000000000_0000101110101000_0010100100010001"; -- 0.045534674418283114
	pesos_i(14885) := b"1111111111111111_1111111111111111_1111101110100110_0101111010111011"; -- -0.01699264467788095
	pesos_i(14886) := b"0000000000000000_0000000000000000_0001100010011110_1011010111010001"; -- 0.09617172572895387
	pesos_i(14887) := b"1111111111111111_1111111111111111_1110101000011011_1001000111011000"; -- -0.08551681962660722
	pesos_i(14888) := b"1111111111111111_1111111111111111_1111000000110100_0111111001110000"; -- -0.06169900675814854
	pesos_i(14889) := b"1111111111111111_1111111111111111_1110011010001010_1110111011011001"; -- -0.09944255062272356
	pesos_i(14890) := b"0000000000000000_0000000000000000_0010010011011010_0011111000101100"; -- 0.14395512171248126
	pesos_i(14891) := b"0000000000000000_0000000000000000_0001000111001111_1010011010000100"; -- 0.06957474453747493
	pesos_i(14892) := b"0000000000000000_0000000000000000_0001000010100100_0101111111110011"; -- 0.06500816039732986
	pesos_i(14893) := b"0000000000000000_0000000000000000_0010010101010000_0001101001001110"; -- 0.14575352102935918
	pesos_i(14894) := b"0000000000000000_0000000000000000_0000011001001011_1010000110010110"; -- 0.02459154055906631
	pesos_i(14895) := b"0000000000000000_0000000000000000_0001011111100111_0100010001010101"; -- 0.09337260318561338
	pesos_i(14896) := b"0000000000000000_0000000000000000_0001011101111010_0110000011101100"; -- 0.09171109935268885
	pesos_i(14897) := b"1111111111111111_1111111111111111_1110000111001101_1001110001111011"; -- -0.1179563712830396
	pesos_i(14898) := b"0000000000000000_0000000000000000_0000011010100110_1001101111000011"; -- 0.025979743002588995
	pesos_i(14899) := b"1111111111111111_1111111111111111_1101111111110101_1001110101000110"; -- -0.12515847247424763
	pesos_i(14900) := b"0000000000000000_0000000000000000_0000110101000010_1101111100111101"; -- 0.0518016361372422
	pesos_i(14901) := b"1111111111111111_1111111111111111_1111110011001100_1101101010101000"; -- -0.012499174014257874
	pesos_i(14902) := b"0000000000000000_0000000000000000_0000010011010110_1001100010101010"; -- 0.018899480327804648
	pesos_i(14903) := b"0000000000000000_0000000000000000_0001000111011111_1100001110001111"; -- 0.06982061621671229
	pesos_i(14904) := b"0000000000000000_0000000000000000_0000110111111101_0101110010011001"; -- 0.05464724299753788
	pesos_i(14905) := b"0000000000000000_0000000000000000_0000001110001001_1111010110011100"; -- 0.013823843503768106
	pesos_i(14906) := b"1111111111111111_1111111111111111_1110000111011101_1101111101101001"; -- -0.11770824142060338
	pesos_i(14907) := b"1111111111111111_1111111111111111_1101101001110101_1100000110001011"; -- -0.14664068564895413
	pesos_i(14908) := b"1111111111111111_1111111111111111_1101000111101001_1111110001101100"; -- -0.18002340667083502
	pesos_i(14909) := b"1111111111111111_1111111111111111_1111011011101001_0101000010010110"; -- -0.035502398966804315
	pesos_i(14910) := b"1111111111111111_1111111111111111_1111010011101011_0100000000110010"; -- -0.04328535830502939
	pesos_i(14911) := b"1111111111111111_1111111111111111_1111100001101111_1111011100111011"; -- -0.02954153839031817
	pesos_i(14912) := b"0000000000000000_0000000000000000_0010001011100011_1110010001010111"; -- 0.13628985533397858
	pesos_i(14913) := b"1111111111111111_1111111111111111_1110111010110010_0110000001101101"; -- -0.06759068806791058
	pesos_i(14914) := b"0000000000000000_0000000000000000_0001011101010000_0000101111101100"; -- 0.09106516383851998
	pesos_i(14915) := b"1111111111111111_1111111111111111_1111010011000111_1010001110010101"; -- -0.0438287507230357
	pesos_i(14916) := b"0000000000000000_0000000000000000_0001001010001001_1101101110110000"; -- 0.07241604855575179
	pesos_i(14917) := b"1111111111111111_1111111111111111_1110000000100001_0000111001110001"; -- -0.12449559920059092
	pesos_i(14918) := b"0000000000000000_0000000000000000_0001011110101110_1001110100111001"; -- 0.09250815058439196
	pesos_i(14919) := b"0000000000000000_0000000000000000_0000100100011001_0010101010001011"; -- 0.0355402554416869
	pesos_i(14920) := b"0000000000000000_0000000000000000_0000100101000111_0010010010110111"; -- 0.036241812422522036
	pesos_i(14921) := b"0000000000000000_0000000000000000_0001100101010100_0010001000111011"; -- 0.09894002865208468
	pesos_i(14922) := b"1111111111111111_1111111111111111_1101101110101011_1100011011111111"; -- -0.14191013607271266
	pesos_i(14923) := b"0000000000000000_0000000000000000_0000110001110011_0000110100000000"; -- 0.04863053563696339
	pesos_i(14924) := b"0000000000000000_0000000000000000_0001010100011000_0011011001101111"; -- 0.08240070552031047
	pesos_i(14925) := b"1111111111111111_1111111111111111_1111101001010110_0000101011001110"; -- -0.02212460014358429
	pesos_i(14926) := b"1111111111111111_1111111111111111_1111100010011111_1100001101011111"; -- -0.02881220761847749
	pesos_i(14927) := b"0000000000000000_0000000000000000_0001011000100110_1011110101111111"; -- 0.08652862892087523
	pesos_i(14928) := b"0000000000000000_0000000000000000_0000001101000010_0011010111001111"; -- 0.012729037394416463
	pesos_i(14929) := b"0000000000000000_0000000000000000_0000001011101011_0011011001011110"; -- 0.011401555941561708
	pesos_i(14930) := b"0000000000000000_0000000000000000_0000011111111111_1110110011111000"; -- 0.031248865629852445
	pesos_i(14931) := b"1111111111111111_1111111111111111_1111111001000010_1011010001001011"; -- -0.006794673677511769
	pesos_i(14932) := b"1111111111111111_1111111111111111_1101101100011000_1001101110010110"; -- -0.14415576532534066
	pesos_i(14933) := b"0000000000000000_0000000000000000_0000111000101001_0110111111110110"; -- 0.05531978380205064
	pesos_i(14934) := b"0000000000000000_0000000000000000_0001100100101001_0101011010000011"; -- 0.09828701685100025
	pesos_i(14935) := b"1111111111111111_1111111111111111_1110100011111111_0010111000010010"; -- -0.08985626275992306
	pesos_i(14936) := b"0000000000000000_0000000000000000_0000001100101110_1110110010111110"; -- 0.0124347651398539
	pesos_i(14937) := b"0000000000000000_0000000000000000_0001001100000000_0111000011111110"; -- 0.07422548495679139
	pesos_i(14938) := b"0000000000000000_0000000000000000_0001011111010001_1011010011011011"; -- 0.0930436167645685
	pesos_i(14939) := b"1111111111111111_1111111111111111_1111010010110011_1111010011000001"; -- -0.04412908823165248
	pesos_i(14940) := b"0000000000000000_0000000000000000_0010010000100101_0011010000101100"; -- 0.14119268478064095
	pesos_i(14941) := b"0000000000000000_0000000000000000_0000001000011100_0101011110000110"; -- 0.008244962878041705
	pesos_i(14942) := b"0000000000000000_0000000000000000_0000010011000111_1101010101111010"; -- 0.018674223262096654
	pesos_i(14943) := b"1111111111111111_1111111111111111_1111010101001001_0111101010110111"; -- -0.04184754396623715
	pesos_i(14944) := b"1111111111111111_1111111111111111_1111101000110111_0111000010000000"; -- -0.02259156106468098
	pesos_i(14945) := b"0000000000000000_0000000000000000_0001100111001000_1011100011111000"; -- 0.10071903280123369
	pesos_i(14946) := b"0000000000000000_0000000000000000_0000111101000101_1000001010111111"; -- 0.059654399464998994
	pesos_i(14947) := b"1111111111111111_1111111111111111_1111101010111011_0101111010100100"; -- -0.020578465477118824
	pesos_i(14948) := b"0000000000000000_0000000000000000_0001001110111001_0101000000101100"; -- 0.07704640462894537
	pesos_i(14949) := b"0000000000000000_0000000000000000_0001101001011010_0111100000100000"; -- 0.10294295111583386
	pesos_i(14950) := b"1111111111111111_1111111111111111_1111101010010001_1100010000100110"; -- -0.021213284112260717
	pesos_i(14951) := b"1111111111111111_1111111111111111_1110100110011111_0011111010111000"; -- -0.08741386415488007
	pesos_i(14952) := b"1111111111111111_1111111111111111_1111011100110110_0001101101110011"; -- -0.03433063940577198
	pesos_i(14953) := b"1111111111111111_1111111111111111_1101111000101101_0001011100011101"; -- -0.13212447682925085
	pesos_i(14954) := b"0000000000000000_0000000000000000_0000000101101001_1110101100010000"; -- 0.005522433616287964
	pesos_i(14955) := b"1111111111111111_1111111111111111_1111110011001011_1000111011011011"; -- -0.012518950949225604
	pesos_i(14956) := b"1111111111111111_1111111111111111_1110100110101000_1101011110101101"; -- -0.0872674181684624
	pesos_i(14957) := b"0000000000000000_0000000000000000_0000111100010111_0111100000000111"; -- 0.05895185639039578
	pesos_i(14958) := b"1111111111111111_1111111111111111_1101111010101110_0011100110010000"; -- -0.1301540396467361
	pesos_i(14959) := b"1111111111111111_1111111111111111_1101110111010010_0111100010001111"; -- -0.1335072185369412
	pesos_i(14960) := b"0000000000000000_0000000000000000_0000011100100100_0010110001011010"; -- 0.027895710025281652
	pesos_i(14961) := b"0000000000000000_0000000000000000_0001100011101001_1000111011000111"; -- 0.09731380806221374
	pesos_i(14962) := b"1111111111111111_1111111111111111_1111110000001011_1101100010111000"; -- -0.015444235911857507
	pesos_i(14963) := b"0000000000000000_0000000000000000_0000011100100010_1010001111010001"; -- 0.02787231296196298
	pesos_i(14964) := b"1111111111111111_1111111111111111_1110011100011000_1110111100011100"; -- -0.09727578696750228
	pesos_i(14965) := b"1111111111111111_1111111111111111_1111101111011000_1110000001110001"; -- -0.016221973703171008
	pesos_i(14966) := b"0000000000000000_0000000000000000_0000001001111100_0001001001000000"; -- 0.00970567752082624
	pesos_i(14967) := b"1111111111111111_1111111111111111_1110101010111101_1100010101001000"; -- -0.08304183001437702
	pesos_i(14968) := b"1111111111111111_1111111111111111_1111110101000000_1000101101101100"; -- -0.010733877356893786
	pesos_i(14969) := b"0000000000000000_0000000000000000_0000110110001101_1001110100111100"; -- 0.05294211126367163
	pesos_i(14970) := b"1111111111111111_1111111111111111_1110100011101110_0110101101111111"; -- -0.0901120008423648
	pesos_i(14971) := b"1111111111111111_1111111111111111_1101111110001001_1010111000010100"; -- -0.1268054201191692
	pesos_i(14972) := b"1111111111111111_1111111111111111_1110001011101101_0011101100111111"; -- -0.11356763558261472
	pesos_i(14973) := b"0000000000000000_0000000000000000_0010010010100110_0010111110000111"; -- 0.14316079178795982
	pesos_i(14974) := b"1111111111111111_1111111111111111_1111110001011100_0111101100001010"; -- -0.014213857712558125
	pesos_i(14975) := b"0000000000000000_0000000000000000_0001110100011101_1000001001000000"; -- 0.11373151837103788
	pesos_i(14976) := b"0000000000000000_0000000000000000_0001010001010110_1010101101000101"; -- 0.07944746430743516
	pesos_i(14977) := b"1111111111111111_1111111111111111_1111101011000000_1100001011111011"; -- -0.020496190717963818
	pesos_i(14978) := b"0000000000000000_0000000000000000_0001110000110011_1100111001000100"; -- 0.11016549265472401
	pesos_i(14979) := b"0000000000000000_0000000000000000_0001110001001000_0101010001101001"; -- 0.11047866414243329
	pesos_i(14980) := b"1111111111111111_1111111111111111_1111110010100001_0011100110000000"; -- -0.013164907628074103
	pesos_i(14981) := b"0000000000000000_0000000000000000_0010000111101111_1010010000010001"; -- 0.13256287973143557
	pesos_i(14982) := b"0000000000000000_0000000000000000_0001101110101101_1100000100100110"; -- 0.10812003306975344
	pesos_i(14983) := b"1111111111111111_1111111111111111_1101111001000100_1010110000011100"; -- -0.13176464385907058
	pesos_i(14984) := b"1111111111111111_1111111111111111_1110000010100000_0001111111010101"; -- -0.12255669645169645
	pesos_i(14985) := b"1111111111111111_1111111111111111_1110110100000110_1110011110110101"; -- -0.07411338637838853
	pesos_i(14986) := b"0000000000000000_0000000000000000_0001111010000010_0001110111111011"; -- 0.11917292947091052
	pesos_i(14987) := b"0000000000000000_0000000000000000_0000001001001110_0010100001011111"; -- 0.009005091762417417
	pesos_i(14988) := b"1111111111111111_1111111111111111_1111011001111000_1011110000101000"; -- -0.037220230212112924
	pesos_i(14989) := b"0000000000000000_0000000000000000_0000101000000111_0111001101110000"; -- 0.03917619212932052
	pesos_i(14990) := b"0000000000000000_0000000000000000_0001100011100110_0110101000101101"; -- 0.09726585009626906
	pesos_i(14991) := b"1111111111111111_1111111111111111_1111001100100111_1000010111100000"; -- -0.05017817774464611
	pesos_i(14992) := b"1111111111111111_1111111111111111_1110111110100100_0101101110100011"; -- -0.06389834653337273
	pesos_i(14993) := b"0000000000000000_0000000000000000_0001110011010111_1111110100101010"; -- 0.11267072948337999
	pesos_i(14994) := b"1111111111111111_1111111111111111_1101101000001111_1001110110011001"; -- -0.14819922470275165
	pesos_i(14995) := b"0000000000000000_0000000000000000_0001001011010001_0001110100011111"; -- 0.07350332255647997
	pesos_i(14996) := b"1111111111111111_1111111111111111_1111100001101001_1010011010110000"; -- -0.029637891687932637
	pesos_i(14997) := b"0000000000000000_0000000000000000_0001101111110010_0101111001000111"; -- 0.10916699629759316
	pesos_i(14998) := b"0000000000000000_0000000000000000_0000001011111011_1011101101010111"; -- 0.011653622434474901
	pesos_i(14999) := b"1111111111111111_1111111111111111_1110001001001001_0110111110101000"; -- -0.11606695326148453
	pesos_i(15000) := b"1111111111111111_1111111111111111_1110101110101100_1011010000110010"; -- -0.07939599788910337
	pesos_i(15001) := b"0000000000000000_0000000000000000_0001000100011100_0000111101110011"; -- 0.06683441701309221
	pesos_i(15002) := b"0000000000000000_0000000000000000_0000011010010001_1100110000011101"; -- 0.02566219059506469
	pesos_i(15003) := b"0000000000000000_0000000000000000_0000111110110111_1100110100001000"; -- 0.061398329189704975
	pesos_i(15004) := b"0000000000000000_0000000000000000_0001101101101111_1011010100111001"; -- 0.10717327729679346
	pesos_i(15005) := b"0000000000000000_0000000000000000_0000000100100000_0110011001111010"; -- 0.004400639439334419
	pesos_i(15006) := b"1111111111111111_1111111111111111_1110111100011011_1010101000000001"; -- -0.06598412973678881
	pesos_i(15007) := b"0000000000000000_0000000000000000_0001100010011111_0000100000110101"; -- 0.09617663674363754
	pesos_i(15008) := b"0000000000000000_0000000000000000_0000101001100011_1101011010011100"; -- 0.04058591184818789
	pesos_i(15009) := b"1111111111111111_1111111111111111_1111100000111011_0000011110011001"; -- -0.03034927867100404
	pesos_i(15010) := b"0000000000000000_0000000000000000_0000011000110100_0000000011110100"; -- 0.02423101391599212
	pesos_i(15011) := b"0000000000000000_0000000000000000_0000010000111101_1101000111111001"; -- 0.016568301538209887
	pesos_i(15012) := b"1111111111111111_1111111111111111_1101101110001111_1110001100110110"; -- -0.14233570027942063
	pesos_i(15013) := b"1111111111111111_1111111111111111_1110111101100011_1101111010011101"; -- -0.06488236104010918
	pesos_i(15014) := b"1111111111111111_1111111111111111_1101101100011010_0110101101010000"; -- -0.1441281252118408
	pesos_i(15015) := b"1111111111111111_1111111111111111_1110010100011011_0010100000110100"; -- -0.10505436644371242
	pesos_i(15016) := b"0000000000000000_0000000000000000_0000010010110110_1011100101100011"; -- 0.01841314950500087
	pesos_i(15017) := b"0000000000000000_0000000000000000_0001110001101011_1110111000001100"; -- 0.11102187919990464
	pesos_i(15018) := b"1111111111111111_1111111111111111_1110100111011110_0001001010001001"; -- -0.08645519402273795
	pesos_i(15019) := b"1111111111111111_1111111111111111_1111101011101110_0111100001110111"; -- -0.019798728018456585
	pesos_i(15020) := b"1111111111111111_1111111111111111_1111110001000010_0101010100001100"; -- -0.014612850694348933
	pesos_i(15021) := b"1111111111111111_1111111111111111_1110100101000010_0010001001111010"; -- -0.08883461498894164
	pesos_i(15022) := b"0000000000000000_0000000000000000_0001111010011101_1110101001101000"; -- 0.11959710158022453
	pesos_i(15023) := b"1111111111111111_1111111111111111_1110101001111111_1111011100011101"; -- -0.08398490457736671
	pesos_i(15024) := b"1111111111111111_1111111111111111_1111111011010110_0110110000000011"; -- -0.004540681141961174
	pesos_i(15025) := b"0000000000000000_0000000000000000_0001100001011010_1101111100011100"; -- 0.09513658939889981
	pesos_i(15026) := b"1111111111111111_1111111111111111_1111111100111110_0001010100001011"; -- -0.002958950923341289
	pesos_i(15027) := b"0000000000000000_0000000000000000_0000010111000000_1111100001110111"; -- 0.022475747259711687
	pesos_i(15028) := b"1111111111111111_1111111111111111_1110001010100101_0011000010010011"; -- -0.11466690463274609
	pesos_i(15029) := b"0000000000000000_0000000000000000_0001101101111101_0100111010001011"; -- 0.1073807800604878
	pesos_i(15030) := b"1111111111111111_1111111111111111_1110001001101100_0101101010010010"; -- -0.11553415235790421
	pesos_i(15031) := b"0000000000000000_0000000000000000_0000110000101010_0101100011111010"; -- 0.047521172563228034
	pesos_i(15032) := b"0000000000000000_0000000000000000_0001110010110110_1011000000001010"; -- 0.11216259237534537
	pesos_i(15033) := b"1111111111111111_1111111111111111_1111001000011000_0111010111100111"; -- -0.054314261576808895
	pesos_i(15034) := b"1111111111111111_1111111111111111_1110001101111101_1110011111101110"; -- -0.11136007735572062
	pesos_i(15035) := b"0000000000000000_0000000000000000_0010001011100010_1010000001000011"; -- 0.13627053863952737
	pesos_i(15036) := b"0000000000000000_0000000000000000_0010000001101110_1110000011101100"; -- 0.12669187323679534
	pesos_i(15037) := b"0000000000000000_0000000000000000_0001101101001000_1011011011101001"; -- 0.10657828521754086
	pesos_i(15038) := b"1111111111111111_1111111111111111_1111101111010010_1100010101000100"; -- -0.01631514626999679
	pesos_i(15039) := b"1111111111111111_1111111111111111_1111101000000010_1010111111101111"; -- -0.02339649593998415
	pesos_i(15040) := b"1111111111111111_1111111111111111_1111001100011011_1111010010010100"; -- -0.05035468477866962
	pesos_i(15041) := b"0000000000000000_0000000000000000_0000010100100100_1001110100011111"; -- 0.02008993158705423
	pesos_i(15042) := b"0000000000000000_0000000000000000_0001011110010000_0111100011111110"; -- 0.09204822722832058
	pesos_i(15043) := b"1111111111111111_1111111111111111_1111001010101001_0001110111110101"; -- -0.052106979171869676
	pesos_i(15044) := b"0000000000000000_0000000000000000_0001110111000100_0011110010000110"; -- 0.11627558022888154
	pesos_i(15045) := b"0000000000000000_0000000000000000_0010000111011101_1010101100100100"; -- 0.1322886430836357
	pesos_i(15046) := b"1111111111111111_1111111111111111_1101110011011000_1110010111000100"; -- -0.13731540638583203
	pesos_i(15047) := b"0000000000000000_0000000000000000_0000111000100100_1110010111101111"; -- 0.05525052156646692
	pesos_i(15048) := b"1111111111111111_1111111111111111_1111010000111100_0001001011101010"; -- -0.04595834530801569
	pesos_i(15049) := b"1111111111111111_1111111111111111_1110000100110011_1000111000011001"; -- -0.12030708213850798
	pesos_i(15050) := b"0000000000000000_0000000000000000_0001001101010111_1100100101010010"; -- 0.07555826418679289
	pesos_i(15051) := b"1111111111111111_1111111111111111_1110100111000101_1101100000010011"; -- -0.08682488954868466
	pesos_i(15052) := b"0000000000000000_0000000000000000_0010011110000011_1111110010000011"; -- 0.15435770218022385
	pesos_i(15053) := b"1111111111111111_1111111111111111_1110011001000110_0010001010000100"; -- -0.10049232754680713
	pesos_i(15054) := b"0000000000000000_0000000000000000_0000001001011011_1101110111000110"; -- 0.009214268491086287
	pesos_i(15055) := b"0000000000000000_0000000000000000_0000101100101101_1001111001010000"; -- 0.04366483175125808
	pesos_i(15056) := b"0000000000000000_0000000000000000_0001111101001110_1101111111100001"; -- 0.12229727987747376
	pesos_i(15057) := b"1111111111111111_1111111111111111_1101111100111010_0000110101000010"; -- -0.12802045009744206
	pesos_i(15058) := b"0000000000000000_0000000000000000_0001110101111000_0110110001010001"; -- 0.11511876088198861
	pesos_i(15059) := b"1111111111111111_1111111111111111_1110101101000110_1101101001000110"; -- -0.08095012454144704
	pesos_i(15060) := b"0000000000000000_0000000000000000_0000101111100100_0110110100110100"; -- 0.046454262904500776
	pesos_i(15061) := b"0000000000000000_0000000000000000_0001101111001110_1100100111001100"; -- 0.10862408850146595
	pesos_i(15062) := b"1111111111111111_1111111111111111_1101111000100110_0010110111001010"; -- -0.13222993677222192
	pesos_i(15063) := b"0000000000000000_0000000000000000_0000000000101111_1101100110111110"; -- 0.0007301416244896933
	pesos_i(15064) := b"0000000000000000_0000000000000000_0000111111100001_1101101010011110"; -- 0.06204000824753583
	pesos_i(15065) := b"1111111111111111_1111111111111111_1110001101100110_0111111000001011"; -- -0.11171734086183806
	pesos_i(15066) := b"0000000000000000_0000000000000000_0000111000101111_1001010010000000"; -- 0.05541351440728011
	pesos_i(15067) := b"1111111111111111_1111111111111111_1101111100100111_0111000000000110"; -- -0.12830448005213882
	pesos_i(15068) := b"1111111111111111_1111111111111111_1111110010000101_0100010001000010"; -- -0.013591512500426332
	pesos_i(15069) := b"0000000000000000_0000000000000000_0001100110100111_0001100000010010"; -- 0.10020590240991618
	pesos_i(15070) := b"1111111111111111_1111111111111111_1110000110101011_1001110000100001"; -- -0.11847519112056515
	pesos_i(15071) := b"1111111111111111_1111111111111111_1101111011100010_1001000111111000"; -- -0.12935531336882286
	pesos_i(15072) := b"0000000000000000_0000000000000000_0000101111011010_1000101011100101"; -- 0.046303444754384526
	pesos_i(15073) := b"1111111111111111_1111111111111111_1111111111001011_1101101100011010"; -- -0.0007956564653303085
	pesos_i(15074) := b"1111111111111111_1111111111111111_1111110000011101_0110000001100100"; -- -0.015176749748926195
	pesos_i(15075) := b"1111111111111111_1111111111111111_1111111011101001_1101100101100100"; -- -0.004244244613679014
	pesos_i(15076) := b"1111111111111111_1111111111111111_1101101011101110_0001011010001100"; -- -0.14480456433226271
	pesos_i(15077) := b"1111111111111111_1111111111111111_1110111010111100_1010111001101101"; -- -0.06743345115652714
	pesos_i(15078) := b"0000000000000000_0000000000000000_0000100101101101_1101000001001011"; -- 0.0368318731302531
	pesos_i(15079) := b"0000000000000000_0000000000000000_0001001000111101_1010101110000010"; -- 0.0712535089077489
	pesos_i(15080) := b"1111111111111111_1111111111111111_1110101101110001_0111110100111001"; -- -0.08029954301700819
	pesos_i(15081) := b"1111111111111111_1111111111111111_1110010001100100_1100111111100101"; -- -0.1078367296564381
	pesos_i(15082) := b"0000000000000000_0000000000000000_0000000000111010_0011011010101111"; -- 0.000888269218845742
	pesos_i(15083) := b"0000000000000000_0000000000000000_0010011000101110_1011101010110001"; -- 0.14915053200000958
	pesos_i(15084) := b"0000000000000000_0000000000000000_0001010101110010_1101110110100000"; -- 0.08378396173695812
	pesos_i(15085) := b"1111111111111111_1111111111111111_1110100001000011_0111000011011000"; -- -0.09272093508976134
	pesos_i(15086) := b"1111111111111111_1111111111111111_1111111100001110_0111100000101100"; -- -0.0036854641476601487
	pesos_i(15087) := b"0000000000000000_0000000000000000_0000010010111010_1100101011011010"; -- 0.01847522558806838
	pesos_i(15088) := b"1111111111111111_1111111111111111_1110100100010101_0100110000000111"; -- -0.08951878388480679
	pesos_i(15089) := b"0000000000000000_0000000000000000_0000111100011000_1100101101010111"; -- 0.05897208083310114
	pesos_i(15090) := b"1111111111111111_1111111111111111_1110001001101000_1010100011010101"; -- -0.11559052268266448
	pesos_i(15091) := b"1111111111111111_1111111111111111_1110011111011000_1111000111101001"; -- -0.09434593258310542
	pesos_i(15092) := b"1111111111111111_1111111111111111_1101101110001100_1100011110111011"; -- -0.14238311463302164
	pesos_i(15093) := b"0000000000000000_0000000000000000_0000011001100110_1110101000101010"; -- 0.02500785373972705
	pesos_i(15094) := b"1111111111111111_1111111111111111_1110010010111110_0110111001111000"; -- -0.1064692455196848
	pesos_i(15095) := b"1111111111111111_1111111111111111_1111111001011100_0011000100001001"; -- -0.006405768773479639
	pesos_i(15096) := b"0000000000000000_0000000000000000_0000000110101010_0010110011100110"; -- 0.0065029203251259675
	pesos_i(15097) := b"0000000000000000_0000000000000000_0010000110110100_0001100001111101"; -- 0.13165429155979103
	pesos_i(15098) := b"0000000000000000_0000000000000000_0001111111011011_1101101010100100"; -- 0.1244484568832454
	pesos_i(15099) := b"0000000000000000_0000000000000000_0000110111010001_0110101111011001"; -- 0.053976765139466296
	pesos_i(15100) := b"0000000000000000_0000000000000000_0000010111111111_0011000011100101"; -- 0.023425155654200287
	pesos_i(15101) := b"0000000000000000_0000000000000000_0000110011100101_1001011011110011"; -- 0.050378260061524516
	pesos_i(15102) := b"1111111111111111_1111111111111111_1111101101010101_0100111011010001"; -- -0.018229555174607455
	pesos_i(15103) := b"1111111111111111_1111111111111111_1110111011110000_0101100001000101"; -- -0.0666451294048169
	pesos_i(15104) := b"1111111111111111_1111111111111111_1111010001000101_1110110010110100"; -- -0.04580803505786501
	pesos_i(15105) := b"0000000000000000_0000000000000000_0000101011100000_0000101011101010"; -- 0.042481119274517434
	pesos_i(15106) := b"0000000000000000_0000000000000000_0000001011100011_0001110010110101"; -- 0.01127795613062135
	pesos_i(15107) := b"1111111111111111_1111111111111111_1111010111001000_1110110010101110"; -- -0.03990288491214867
	pesos_i(15108) := b"1111111111111111_1111111111111111_1101111011001111_0101100001010111"; -- -0.12964866528617625
	pesos_i(15109) := b"1111111111111111_1111111111111111_1101100110001100_0100011000001010"; -- -0.15020334484956815
	pesos_i(15110) := b"0000000000000000_0000000000000000_0010010110001101_1001110011110101"; -- 0.1466920945133511
	pesos_i(15111) := b"1111111111111111_1111111111111111_1101110101010000_0110010101110100"; -- -0.13549199990011188
	pesos_i(15112) := b"1111111111111111_1111111111111111_1111100110001011_0011110100100100"; -- -0.025219134156972366
	pesos_i(15113) := b"0000000000000000_0000000000000000_0000100000000000_1000010100100011"; -- 0.03125793554062693
	pesos_i(15114) := b"0000000000000000_0000000000000000_0000111110111000_1111001010100101"; -- 0.06141583001006027
	pesos_i(15115) := b"0000000000000000_0000000000000000_0000010011010011_1001000000110110"; -- 0.01885320014611304
	pesos_i(15116) := b"1111111111111111_1111111111111111_1111010001011101_1001011011100011"; -- -0.04544693906960556
	pesos_i(15117) := b"1111111111111111_1111111111111111_1110000011000011_1010100110110000"; -- -0.12201442185546703
	pesos_i(15118) := b"1111111111111111_1111111111111111_1111111101111111_1101000110101000"; -- -0.001955887251734705
	pesos_i(15119) := b"1111111111111111_1111111111111111_1111100000011011_0000101101011111"; -- -0.030837334845292722
	pesos_i(15120) := b"0000000000000000_0000000000000000_0010001001011010_0001100010111101"; -- 0.13418726563965147
	pesos_i(15121) := b"0000000000000000_0000000000000000_0000010111101100_1011010000100001"; -- 0.023143060697617353
	pesos_i(15122) := b"1111111111111111_1111111111111111_1111101000001010_1000010111100010"; -- -0.023276932102765092
	pesos_i(15123) := b"1111111111111111_1111111111111111_1111100010100011_1001111110101101"; -- -0.028753300004559623
	pesos_i(15124) := b"1111111111111111_1111111111111111_1111100101100111_0010001111011001"; -- -0.025769958025974805
	pesos_i(15125) := b"1111111111111111_1111111111111111_1111010001100110_0011010111110000"; -- -0.04531538859895726
	pesos_i(15126) := b"0000000000000000_0000000000000000_0000100010000011_0010001001111110"; -- 0.03325095728279655
	pesos_i(15127) := b"1111111111111111_1111111111111111_1111101001000010_1111111001101010"; -- -0.022415255769835253
	pesos_i(15128) := b"0000000000000000_0000000000000000_0001110101000000_1101001000100001"; -- 0.1142703370972597
	pesos_i(15129) := b"0000000000000000_0000000000000000_0001111110000001_0111101010000101"; -- 0.1230694366161011
	pesos_i(15130) := b"0000000000000000_0000000000000000_0001000100010110_1101011000011110"; -- 0.06675470569404755
	pesos_i(15131) := b"0000000000000000_0000000000000000_0001001110111010_1100000110001001"; -- 0.07706842024781425
	pesos_i(15132) := b"1111111111111111_1111111111111111_1111001000001011_1101001101111000"; -- -0.054507048717184564
	pesos_i(15133) := b"1111111111111111_1111111111111111_1111011011110010_0011100011000000"; -- -0.03536649042421043
	pesos_i(15134) := b"0000000000000000_0000000000000000_0001110011010110_0010001100101100"; -- 0.11264247717900643
	pesos_i(15135) := b"0000000000000000_0000000000000000_0001000110010010_1001001100010010"; -- 0.0686427992928376
	pesos_i(15136) := b"1111111111111111_1111111111111111_1110101000001111_0100010110111100"; -- -0.08570446165402726
	pesos_i(15137) := b"0000000000000000_0000000000000000_0000110000010010_1000111011111110"; -- 0.04715818117317693
	pesos_i(15138) := b"0000000000000000_0000000000000000_0001101110111000_1100100000000011"; -- 0.10828828887074032
	pesos_i(15139) := b"0000000000000000_0000000000000000_0001011000101011_1000011110000100"; -- 0.08660170519336405
	pesos_i(15140) := b"0000000000000000_0000000000000000_0000111001000110_0101010000011011"; -- 0.05576062825639474
	pesos_i(15141) := b"1111111111111111_1111111111111111_1111001000010101_1111010011010110"; -- -0.05435247212614948
	pesos_i(15142) := b"0000000000000000_0000000000000000_0000011101011001_1110110111000111"; -- 0.028715954919219293
	pesos_i(15143) := b"1111111111111111_1111111111111111_1111011111010011_1010011010110011"; -- -0.03192670938414332
	pesos_i(15144) := b"0000000000000000_0000000000000000_0000010111111100_0110001100110010"; -- 0.0233823772389836
	pesos_i(15145) := b"0000000000000000_0000000000000000_0001101010101001_0000110110110011"; -- 0.10414205192589793
	pesos_i(15146) := b"1111111111111111_1111111111111111_1110111101001100_1110011111100010"; -- -0.06523276064884699
	pesos_i(15147) := b"0000000000000000_0000000000000000_0000100101011100_1000101111111000"; -- 0.03656840140334504
	pesos_i(15148) := b"0000000000000000_0000000000000000_0000010111110111_1011110110000011"; -- 0.02331146667146667
	pesos_i(15149) := b"0000000000000000_0000000000000000_0010000000001010_0011110011001110"; -- 0.12515621207223193
	pesos_i(15150) := b"0000000000000000_0000000000000000_0010000100001000_0101000110101101"; -- 0.1290331885255858
	pesos_i(15151) := b"1111111111111111_1111111111111111_1110000010001001_0100101110100000"; -- -0.12290503824890343
	pesos_i(15152) := b"0000000000000000_0000000000000000_0000001111011100_0111110000010101"; -- 0.01508307937283441
	pesos_i(15153) := b"0000000000000000_0000000000000000_0001101101000110_1011100110110011"; -- 0.10654793370275835
	pesos_i(15154) := b"1111111111111111_1111111111111111_1111001011010001_0110110100001111"; -- -0.051491912590229144
	pesos_i(15155) := b"1111111111111111_1111111111111111_1101111100110100_1110110110110111"; -- -0.1280986239512371
	pesos_i(15156) := b"0000000000000000_0000000000000000_0001100000001010_1110000101101011"; -- 0.09391602380792818
	pesos_i(15157) := b"0000000000000000_0000000000000000_0000100111000101_0100000100101111"; -- 0.03816611676242979
	pesos_i(15158) := b"1111111111111111_1111111111111111_1110111110101110_0100110111111100"; -- -0.06374657248970142
	pesos_i(15159) := b"1111111111111111_1111111111111111_1111010100111011_1011110011110000"; -- -0.042057219788316245
	pesos_i(15160) := b"1111111111111111_1111111111111111_1111100000111001_1100011010010010"; -- -0.030368413279302824
	pesos_i(15161) := b"1111111111111111_1111111111111111_1101100111110001_1010100111111001"; -- -0.1486562507555555
	pesos_i(15162) := b"1111111111111111_1111111111111111_1111110001001000_1000111000110011"; -- -0.014517891338320904
	pesos_i(15163) := b"1111111111111111_1111111111111111_1110011100111110_1001110101000001"; -- -0.09670083205154814
	pesos_i(15164) := b"0000000000000000_0000000000000000_0001011000101100_1001001100010110"; -- 0.08661765377945903
	pesos_i(15165) := b"1111111111111111_1111111111111111_1111011111101100_1000000000111110"; -- -0.03154753198060686
	pesos_i(15166) := b"0000000000000000_0000000000000000_0001000101110101_1011000001011110"; -- 0.06820204055392899
	pesos_i(15167) := b"0000000000000000_0000000000000000_0010010110101101_0100010010010100"; -- 0.147175108141742
	pesos_i(15168) := b"0000000000000000_0000000000000000_0001000010000010_0101110011001101"; -- 0.06448917391212004
	pesos_i(15169) := b"1111111111111111_1111111111111111_1111111100101010_1111111011101100"; -- -0.0032501862604972643
	pesos_i(15170) := b"0000000000000000_0000000000000000_0010000100010111_0001101000001110"; -- 0.129258755177848
	pesos_i(15171) := b"0000000000000000_0000000000000000_0001110111011011_0110011001111100"; -- 0.1166290333514398
	pesos_i(15172) := b"1111111111111111_1111111111111111_1111111000000110_1011101100001110"; -- -0.007709797917375856
	pesos_i(15173) := b"1111111111111111_1111111111111111_1110010111000101_1001110110001110"; -- -0.10245337749411343
	pesos_i(15174) := b"0000000000000000_0000000000000000_0001111100110100_0000011101111011"; -- 0.12188765288303485
	pesos_i(15175) := b"1111111111111111_1111111111111111_1101101110011100_1010010011010001"; -- -0.14214105510494007
	pesos_i(15176) := b"0000000000000000_0000000000000000_0001011011101011_0000010000110110"; -- 0.08952356633661049
	pesos_i(15177) := b"1111111111111111_1111111111111111_1110001000001110_1000011111101011"; -- -0.1169657754982085
	pesos_i(15178) := b"1111111111111111_1111111111111111_1111001000011000_1100001011100001"; -- -0.05430967339047776
	pesos_i(15179) := b"1111111111111111_1111111111111111_1110110011110100_0011011010100000"; -- -0.0743985994971965
	pesos_i(15180) := b"0000000000000000_0000000000000000_0001011110000100_1010000110111010"; -- 0.09186754984574053
	pesos_i(15181) := b"0000000000000000_0000000000000000_0010001010011001_0010100011001011"; -- 0.13514952625594398
	pesos_i(15182) := b"1111111111111111_1111111111111111_1111101010110111_0011011011000100"; -- -0.02064187733083597
	pesos_i(15183) := b"1111111111111111_1111111111111111_1111001110011111_1110100101100010"; -- -0.048341191807188495
	pesos_i(15184) := b"0000000000000000_0000000000000000_0010100101111001_0010000101101011"; -- 0.16200455525370352
	pesos_i(15185) := b"1111111111111111_1111111111111111_1111011001011111_1111110100001011"; -- -0.037597832510114164
	pesos_i(15186) := b"1111111111111111_1111111111111111_1110010000011000_0101111110111111"; -- -0.10900308219994755
	pesos_i(15187) := b"1111111111111111_1111111111111111_1110100110110000_1011010010110011"; -- -0.0871474325396704
	pesos_i(15188) := b"1111111111111111_1111111111111111_1111011010000110_1101001000001100"; -- -0.037005302552438994
	pesos_i(15189) := b"0000000000000000_0000000000000000_0001111000000001_0101011101100011"; -- 0.11720796750803221
	pesos_i(15190) := b"0000000000000000_0000000000000000_0001010000000100_1110010001000111"; -- 0.07819964147381891
	pesos_i(15191) := b"0000000000000000_0000000000000000_0001011101000000_1000101000101110"; -- 0.09082854869802795
	pesos_i(15192) := b"1111111111111111_1111111111111111_1111011000101011_1110011100100010"; -- -0.03839259558583267
	pesos_i(15193) := b"1111111111111111_1111111111111111_1111101010011111_1111011000110001"; -- -0.02099667842892934
	pesos_i(15194) := b"1111111111111111_1111111111111111_1111001001101100_0001000111101101"; -- -0.053038482224897106
	pesos_i(15195) := b"0000000000000000_0000000000000000_0001011100101110_0101001100011110"; -- 0.09055060835343963
	pesos_i(15196) := b"0000000000000000_0000000000000000_0000001111101000_0110000111110101"; -- 0.015264627710447325
	pesos_i(15197) := b"1111111111111111_1111111111111111_1111100111001001_0111110111111000"; -- -0.024269225038560382
	pesos_i(15198) := b"1111111111111111_1111111111111111_1110010100001001_1100100000011011"; -- -0.10531949365851642
	pesos_i(15199) := b"0000000000000000_0000000000000000_0010000110010011_1000100100011101"; -- 0.1311574645075317
	pesos_i(15200) := b"1111111111111111_1111111111111111_1111001011010110_1111110001101100"; -- -0.051407073542165276
	pesos_i(15201) := b"0000000000000000_0000000000000000_0001000000001010_0101010010110011"; -- 0.06265763635852471
	pesos_i(15202) := b"1111111111111111_1111111111111111_1111100011010111_0111000001101011"; -- -0.02796265982829319
	pesos_i(15203) := b"0000000000000000_0000000000000000_0001111010101111_0111000100010100"; -- 0.11986452817197878
	pesos_i(15204) := b"1111111111111111_1111111111111111_1101111101111110_1111010001000100"; -- -0.12696908316440836
	pesos_i(15205) := b"1111111111111111_1111111111111111_1101100010111011_0001111011010010"; -- -0.15339476944666505
	pesos_i(15206) := b"1111111111111111_1111111111111111_1111100000111000_1011010011110001"; -- -0.03038472277983417
	pesos_i(15207) := b"0000000000000000_0000000000000000_0010001100001101_0101101110011011"; -- 0.1369225743797766
	pesos_i(15208) := b"1111111111111111_1111111111111111_1111110000111011_1011110010100011"; -- -0.01471348792089394
	pesos_i(15209) := b"1111111111111111_1111111111111111_1110100000010011_1111011101101010"; -- -0.0934453360178056
	pesos_i(15210) := b"1111111111111111_1111111111111111_1111011100000101_1110100100110100"; -- -0.035066055956151754
	pesos_i(15211) := b"0000000000000000_0000000000000000_0001011110001011_0011100110110101"; -- 0.09196816130182349
	pesos_i(15212) := b"0000000000000000_0000000000000000_0001101101010110_1001001111110000"; -- 0.1067898236119679
	pesos_i(15213) := b"1111111111111111_1111111111111111_1111111001011010_0000110011011100"; -- -0.006438442485296509
	pesos_i(15214) := b"0000000000000000_0000000000000000_0000100100001101_1001010101100011"; -- 0.03536351840129967
	pesos_i(15215) := b"0000000000000000_0000000000000000_0010000100110111_0011111111111001"; -- 0.1297492963733901
	pesos_i(15216) := b"1111111111111111_1111111111111111_1110101001111011_1110010001000010"; -- -0.08404706364334139
	pesos_i(15217) := b"0000000000000000_0000000000000000_0001000111001100_1111101000011010"; -- 0.06953395012612963
	pesos_i(15218) := b"1111111111111111_1111111111111111_1111111011101001_1110001101111111"; -- -0.004243642281391061
	pesos_i(15219) := b"1111111111111111_1111111111111111_1110001010110111_0000010100011101"; -- -0.11439483674303995
	pesos_i(15220) := b"0000000000000000_0000000000000000_0001111100101011_0001100101101110"; -- 0.12175139360056307
	pesos_i(15221) := b"0000000000000000_0000000000000000_0000001011011010_0101001001100001"; -- 0.011143826103820748
	pesos_i(15222) := b"1111111111111111_1111111111111111_1110111010011101_1001010000101011"; -- -0.06790803862317205
	pesos_i(15223) := b"1111111111111111_1111111111111111_1101110101110010_0011101001101111"; -- -0.13497576518357485
	pesos_i(15224) := b"1111111111111111_1111111111111111_1101110110101100_0010100100010000"; -- -0.1340917907931986
	pesos_i(15225) := b"0000000000000000_0000000000000000_0010000001000001_1101010011011010"; -- 0.12600450833052257
	pesos_i(15226) := b"0000000000000000_0000000000000000_0001001111100010_1111100101101011"; -- 0.07768210281386577
	pesos_i(15227) := b"0000000000000000_0000000000000000_0000011100100110_1111010100111010"; -- 0.02793820061615288
	pesos_i(15228) := b"1111111111111111_1111111111111111_1111101010111100_1010011101111111"; -- -0.02055886407902009
	pesos_i(15229) := b"1111111111111111_1111111111111111_1110110100001111_0001000000011011"; -- -0.0739889082383261
	pesos_i(15230) := b"0000000000000000_0000000000000000_0000100001110011_1001101010011100"; -- 0.033013976202981174
	pesos_i(15231) := b"0000000000000000_0000000000000000_0001001010101000_1011111010101001"; -- 0.07288734079601547
	pesos_i(15232) := b"1111111111111111_1111111111111111_1101111111011101_1110011101110110"; -- -0.1255202614359468
	pesos_i(15233) := b"0000000000000000_0000000000000000_0001110001001000_1000100000011000"; -- 0.11048174452887306
	pesos_i(15234) := b"0000000000000000_0000000000000000_0000001110010101_0000001111101100"; -- 0.013992543382581449
	pesos_i(15235) := b"0000000000000000_0000000000000000_0001010000011010_1111011001110000"; -- 0.07853641734999012
	pesos_i(15236) := b"0000000000000000_0000000000000000_0000111010010111_0000010111000111"; -- 0.05699192148665938
	pesos_i(15237) := b"1111111111111111_1111111111111111_1111111010010100_0111000011011010"; -- -0.005547472752290501
	pesos_i(15238) := b"0000000000000000_0000000000000000_0001100000000100_0100011001110101"; -- 0.09381523461117794
	pesos_i(15239) := b"1111111111111111_1111111111111111_1101100111110110_0100101001101000"; -- -0.1485856529288302
	pesos_i(15240) := b"0000000000000000_0000000000000000_0000110101011010_0110000101000110"; -- 0.05216033894608829
	pesos_i(15241) := b"0000000000000000_0000000000000000_0000101110101010_1110000100110001"; -- 0.04557616669265777
	pesos_i(15242) := b"1111111111111111_1111111111111111_1111001001110111_0110100100101101"; -- -0.05286543523504154
	pesos_i(15243) := b"0000000000000000_0000000000000000_0000110110001111_1111011101111111"; -- 0.052978008829784394
	pesos_i(15244) := b"0000000000000000_0000000000000000_0000111001100111_0001100101111011"; -- 0.05626067392008442
	pesos_i(15245) := b"1111111111111111_1111111111111111_1110011101011101_0100010101011001"; -- -0.09623304920213376
	pesos_i(15246) := b"1111111111111111_1111111111111111_1111110011100000_1000101010011110"; -- -0.01219876892573988
	pesos_i(15247) := b"1111111111111111_1111111111111111_1111110000010111_0001000111000110"; -- -0.015272988585698961
	pesos_i(15248) := b"0000000000000000_0000000000000000_0001011000100011_0111000101001110"; -- 0.0864783110843961
	pesos_i(15249) := b"1111111111111111_1111111111111111_1111101010000001_1011011101110000"; -- -0.021458182509276304
	pesos_i(15250) := b"1111111111111111_1111111111111111_1110000100000111_0010100101000010"; -- -0.12098447922170942
	pesos_i(15251) := b"1111111111111111_1111111111111111_1111001111111101_0000011100101011"; -- -0.04692034906110008
	pesos_i(15252) := b"0000000000000000_0000000000000000_0001011000010010_0011111100011110"; -- 0.08621592030211435
	pesos_i(15253) := b"0000000000000000_0000000000000000_0010000010010011_0011011100011101"; -- 0.12724632694174262
	pesos_i(15254) := b"0000000000000000_0000000000000000_0001110011011001_0110100111010111"; -- 0.11269246575748057
	pesos_i(15255) := b"1111111111111111_1111111111111111_1101101000100001_1100000011100011"; -- -0.1479224630820666
	pesos_i(15256) := b"1111111111111111_1111111111111111_1111010101001011_0001111001011010"; -- -0.04182253182030285
	pesos_i(15257) := b"0000000000000000_0000000000000000_0001111001100011_1101000001100111"; -- 0.11871054184858827
	pesos_i(15258) := b"0000000000000000_0000000000000000_0000011010111100_0001000110000000"; -- 0.026307195512566463
	pesos_i(15259) := b"0000000000000000_0000000000000000_0010001011100110_1010100010110010"; -- 0.13633207656479573
	pesos_i(15260) := b"0000000000000000_0000000000000000_0001110100110100_0111000011111111"; -- 0.1140814421773146
	pesos_i(15261) := b"1111111111111111_1111111111111111_1110011000111010_0010000010101000"; -- -0.10067554382176357
	pesos_i(15262) := b"1111111111111111_1111111111111111_1111000110110010_0110100010111100"; -- -0.05587144299912981
	pesos_i(15263) := b"1111111111111111_1111111111111111_1110010000000000_0011110110000010"; -- -0.10937133380051012
	pesos_i(15264) := b"1111111111111111_1111111111111111_1110011011001011_1010000110010111"; -- -0.0984553343135663
	pesos_i(15265) := b"1111111111111111_1111111111111111_1111101000001100_0000110000001000"; -- -0.023253677355835552
	pesos_i(15266) := b"1111111111111111_1111111111111111_1111111000010011_0010010111101110"; -- -0.007520322225956618
	pesos_i(15267) := b"1111111111111111_1111111111111111_1111111010010001_0100011111001011"; -- -0.005595696341598926
	pesos_i(15268) := b"0000000000000000_0000000000000000_0001000111110111_0000110100000010"; -- 0.07017594611640397
	pesos_i(15269) := b"1111111111111111_1111111111111111_1110100011101011_1010011100101001"; -- -0.09015422094456177
	pesos_i(15270) := b"1111111111111111_1111111111111111_1111101001100000_1100111000111010"; -- -0.021960364196266638
	pesos_i(15271) := b"0000000000000000_0000000000000000_0010011101110000_1001000110110001"; -- 0.15406141828018843
	pesos_i(15272) := b"1111111111111111_1111111111111111_1111000110100100_1000010011000111"; -- -0.056083394453814286
	pesos_i(15273) := b"1111111111111111_1111111111111111_1111110110010000_0010011101011010"; -- -0.009519138759921483
	pesos_i(15274) := b"0000000000000000_0000000000000000_0001001100001101_0100100001011111"; -- 0.07442142797888131
	pesos_i(15275) := b"1111111111111111_1111111111111111_1110010011111010_0010110001110111"; -- -0.10555765249821335
	pesos_i(15276) := b"1111111111111111_1111111111111111_1111101011000011_1101010000110010"; -- -0.020449388352786667
	pesos_i(15277) := b"1111111111111111_1111111111111111_1110001011111110_0001111100000111"; -- -0.113309918246891
	pesos_i(15278) := b"1111111111111111_1111111111111111_1110101011000000_1011000110011011"; -- -0.08299722635729265
	pesos_i(15279) := b"1111111111111111_1111111111111111_1110000101110100_1101010010001000"; -- -0.11931106257543643
	pesos_i(15280) := b"0000000000000000_0000000000000000_0000000100001101_1011110010110010"; -- 0.004115861414976117
	pesos_i(15281) := b"1111111111111111_1111111111111111_1101111011001100_0110010110011100"; -- -0.12969365058816165
	pesos_i(15282) := b"0000000000000000_0000000000000000_0000010101100110_0011100011000110"; -- 0.021091030346189445
	pesos_i(15283) := b"0000000000000000_0000000000000000_0010010110000101_1100110000001110"; -- 0.1465728316590369
	pesos_i(15284) := b"1111111111111111_1111111111111111_1111110110110100_1111000010001000"; -- -0.008957831122675954
	pesos_i(15285) := b"1111111111111111_1111111111111111_1111010011100110_0000101101010101"; -- -0.04336480310306524
	pesos_i(15286) := b"0000000000000000_0000000000000000_0001101000101100_1110010111001010"; -- 0.10224758330360001
	pesos_i(15287) := b"1111111111111111_1111111111111111_1110101101111011_0011011001111101"; -- -0.08015117115654845
	pesos_i(15288) := b"1111111111111111_1111111111111111_1111011001000100_0010010100110101"; -- -0.038022684656571215
	pesos_i(15289) := b"0000000000000000_0000000000000000_0010010101010010_1011110110000011"; -- 0.14579376642099504
	pesos_i(15290) := b"0000000000000000_0000000000000000_0000011001101000_1110000010111001"; -- 0.025037808550298274
	pesos_i(15291) := b"1111111111111111_1111111111111111_1110011001101111_1000010010000100"; -- -0.09986087589632477
	pesos_i(15292) := b"0000000000000000_0000000000000000_0001000100111100_0101110010110100"; -- 0.06732730294262036
	pesos_i(15293) := b"1111111111111111_1111111111111111_1111011100100001_0011011111100011"; -- -0.034649378826236824
	pesos_i(15294) := b"1111111111111111_1111111111111111_1110011111011011_0011011110101110"; -- -0.09431125638988713
	pesos_i(15295) := b"1111111111111111_1111111111111111_1110101011101100_1110100100010111"; -- -0.08232253265997466
	pesos_i(15296) := b"1111111111111111_1111111111111111_1110000010100111_1000011110010011"; -- -0.12244370134672082
	pesos_i(15297) := b"0000000000000000_0000000000000000_0000010010100111_1011000000110010"; -- 0.01818371975811062
	pesos_i(15298) := b"1111111111111111_1111111111111111_1110111100000001_0011011110100011"; -- -0.06638767504694636
	pesos_i(15299) := b"1111111111111111_1111111111111111_1110111111010011_1100100101100110"; -- -0.06317464128653921
	pesos_i(15300) := b"1111111111111111_1111111111111111_1110000110010001_0010100111110001"; -- -0.11887872569991546
	pesos_i(15301) := b"1111111111111111_1111111111111111_1110101001010001_1101110101100001"; -- -0.0846883428779772
	pesos_i(15302) := b"0000000000000000_0000000000000000_0001110000110110_0101001101101001"; -- 0.11020394632183765
	pesos_i(15303) := b"0000000000000000_0000000000000000_0001111110011110_0101010110010111"; -- 0.12350974011507974
	pesos_i(15304) := b"1111111111111111_1111111111111111_1110110000111000_0001001010110101"; -- -0.07726939276856219
	pesos_i(15305) := b"0000000000000000_0000000000000000_0000011111011011_1011111100111100"; -- 0.03069682318540076
	pesos_i(15306) := b"1111111111111111_1111111111111111_1111110100011001_0101110111001100"; -- -0.011331689536215491
	pesos_i(15307) := b"1111111111111111_1111111111111111_1101111111010011_0001010111010000"; -- -0.12568534543425405
	pesos_i(15308) := b"0000000000000000_0000000000000000_0000100101101100_1100010100111001"; -- 0.03681595455598547
	pesos_i(15309) := b"0000000000000000_0000000000000000_0000011001011110_0110101111010000"; -- 0.024878252213708475
	pesos_i(15310) := b"0000000000000000_0000000000000000_0000001111110011_1011111011110001"; -- 0.015438016630466856
	pesos_i(15311) := b"1111111111111111_1111111111111111_1111001110111110_0000011000110110"; -- -0.04788170985685195
	pesos_i(15312) := b"0000000000000000_0000000000000000_0000100110011111_1000101100111000"; -- 0.03759069562958422
	pesos_i(15313) := b"1111111111111111_1111111111111111_1111001110010111_0111101111110000"; -- -0.04846978564846632
	pesos_i(15314) := b"0000000000000000_0000000000000000_0000000001100011_1110001111011001"; -- 0.0015242009597008321
	pesos_i(15315) := b"1111111111111111_1111111111111111_1110000000111000_0101011000001000"; -- -0.12414037987958049
	pesos_i(15316) := b"0000000000000000_0000000000000000_0000100000111110_0011111100100100"; -- 0.03219980839052795
	pesos_i(15317) := b"1111111111111111_1111111111111111_1110111110001011_1100100000001100"; -- -0.06427335454638126
	pesos_i(15318) := b"0000000000000000_0000000000000000_0001000011100000_1000010000001000"; -- 0.06592583849214262
	pesos_i(15319) := b"0000000000000000_0000000000000000_0001011111010011_0110100001101011"; -- 0.09306957837505395
	pesos_i(15320) := b"1111111111111111_1111111111111111_1110001111111111_1110001110011001"; -- -0.10937669295586633
	pesos_i(15321) := b"1111111111111111_1111111111111111_1111101001011110_0111101011101110"; -- -0.021995846609178596
	pesos_i(15322) := b"0000000000000000_0000000000000000_0000011100011100_1110100111101010"; -- 0.02778493853502306
	pesos_i(15323) := b"0000000000000000_0000000000000000_0000111000100001_1001111100110000"; -- 0.0552005283576168
	pesos_i(15324) := b"0000000000000000_0000000000000000_0001100010000100_1101100111100100"; -- 0.09577714740993831
	pesos_i(15325) := b"0000000000000000_0000000000000000_0001101101011010_0100101010000001"; -- 0.10684648172408555
	pesos_i(15326) := b"0000000000000000_0000000000000000_0001001111110110_0100010100000100"; -- 0.07797652584030142
	pesos_i(15327) := b"0000000000000000_0000000000000000_0001101111100001_0101000110000011"; -- 0.1089068360897429
	pesos_i(15328) := b"0000000000000000_0000000000000000_0001001001100001_1100010000110101"; -- 0.07180429749308757
	pesos_i(15329) := b"1111111111111111_1111111111111111_1101011001101111_1011000110101000"; -- -0.16235818539174252
	pesos_i(15330) := b"1111111111111111_1111111111111111_1111001010110100_0111010011001100"; -- -0.051933956430987506
	pesos_i(15331) := b"1111111111111111_1111111111111111_1110100111100000_0111000100000011"; -- -0.0864190452175587
	pesos_i(15332) := b"0000000000000000_0000000000000000_0001001101011101_1111011000010101"; -- 0.07565248505014466
	pesos_i(15333) := b"0000000000000000_0000000000000000_0000011011110101_0001101010111010"; -- 0.027177496247075456
	pesos_i(15334) := b"0000000000000000_0000000000000000_0001001100010111_0111110100111010"; -- 0.07457716625725797
	pesos_i(15335) := b"1111111111111111_1111111111111111_1111100111111010_0001101010010100"; -- -0.0235274685644898
	pesos_i(15336) := b"1111111111111111_1111111111111111_1111001110001010_0101110010011011"; -- -0.048670017488691396
	pesos_i(15337) := b"0000000000000000_0000000000000000_0001111101100000_1010001110101011"; -- 0.1225683491300506
	pesos_i(15338) := b"0000000000000000_0000000000000000_0010001011000111_0111011001011110"; -- 0.1358560542931223
	pesos_i(15339) := b"0000000000000000_0000000000000000_0001101001101011_0001001010110001"; -- 0.1031963045812931
	pesos_i(15340) := b"0000000000000000_0000000000000000_0001001010011000_0010001010100011"; -- 0.07263390042358672
	pesos_i(15341) := b"1111111111111111_1111111111111111_1110000111010111_0001000100100111"; -- -0.11781208810744209
	pesos_i(15342) := b"0000000000000000_0000000000000000_0000001011001111_1101010100101010"; -- 0.010983774997181929
	pesos_i(15343) := b"1111111111111111_1111111111111111_1101100000100000_1011000001011010"; -- -0.15575120744250057
	pesos_i(15344) := b"0000000000000000_0000000000000000_0001100110011110_1100110000101000"; -- 0.10007930744554584
	pesos_i(15345) := b"1111111111111111_1111111111111111_1111101101110000_0010011110001000"; -- -0.01781990942092052
	pesos_i(15346) := b"0000000000000000_0000000000000000_0000111000101011_0110010100100100"; -- 0.05534965636576925
	pesos_i(15347) := b"1111111111111111_1111111111111111_1101101100101110_0010010010001100"; -- -0.14382716727423736
	pesos_i(15348) := b"0000000000000000_0000000000000000_0000010101011111_1100100111110000"; -- 0.020992871357851564
	pesos_i(15349) := b"1111111111111111_1111111111111111_1110100110011110_0100000000000110"; -- -0.08742904530375281
	pesos_i(15350) := b"1111111111111111_1111111111111111_1110100011000110_1100110010110001"; -- -0.09071655915988827
	pesos_i(15351) := b"1111111111111111_1111111111111111_1101100110110110_1001001011000100"; -- -0.14955790237735658
	pesos_i(15352) := b"0000000000000000_0000000000000000_0001000000101110_0010001000001101"; -- 0.06320393385275588
	pesos_i(15353) := b"0000000000000000_0000000000000000_0001001011000010_0101011010000010"; -- 0.07327786132928593
	pesos_i(15354) := b"1111111111111111_1111111111111111_1111011000100010_0111101111100111"; -- -0.038536316086368816
	pesos_i(15355) := b"1111111111111111_1111111111111111_1110010111110010_1001111011100111"; -- -0.10176665180073662
	pesos_i(15356) := b"1111111111111111_1111111111111111_1111011001110100_0101110100010001"; -- -0.037286933330723256
	pesos_i(15357) := b"0000000000000000_0000000000000000_0001010110000000_1101011010110110"; -- 0.08399717287873341
	pesos_i(15358) := b"1111111111111111_1111111111111111_1101100110000101_1001111110001010"; -- -0.150304821895053
	pesos_i(15359) := b"0000000000000000_0000000000000000_0000011001000001_1101110010011010"; -- 0.024442470098428263
	pesos_i(15360) := b"1111111111111111_1111111111111111_1111000101100110_1101000010111000"; -- -0.05702491302039206
	pesos_i(15361) := b"0000000000000000_0000000000000000_0000111000011010_0111011011101000"; -- 0.055091315789154174
	pesos_i(15362) := b"0000000000000000_0000000000000000_0001010110000101_0010110101000100"; -- 0.08406336698932072
	pesos_i(15363) := b"1111111111111111_1111111111111111_1111101110111000_0011101101100111"; -- -0.016720092179712865
	pesos_i(15364) := b"0000000000000000_0000000000000000_0000111111110001_1101010100000100"; -- 0.06228381483917926
	pesos_i(15365) := b"0000000000000000_0000000000000000_0010001001101100_1011111110000110"; -- 0.13447186480912837
	pesos_i(15366) := b"0000000000000000_0000000000000000_0000001101011101_0000000101001111"; -- 0.013137895269188028
	pesos_i(15367) := b"0000000000000000_0000000000000000_0000100110001111_0111100000100100"; -- 0.03734541780295184
	pesos_i(15368) := b"1111111111111111_1111111111111111_1110010001100010_1100111111110110"; -- -0.10786724322583376
	pesos_i(15369) := b"0000000000000000_0000000000000000_0000101111110011_0110000011100010"; -- 0.04668241038221733
	pesos_i(15370) := b"1111111111111111_1111111111111111_1111100100101101_1110010100111011"; -- -0.02664344136371683
	pesos_i(15371) := b"1111111111111111_1111111111111111_1110000010000000_1000110011100010"; -- -0.12303847766843776
	pesos_i(15372) := b"1111111111111111_1111111111111111_1111001110111011_1010011110101111"; -- -0.04791786171496439
	pesos_i(15373) := b"0000000000000000_0000000000000000_0010010000111011_0101011001001110"; -- 0.14153041270917022
	pesos_i(15374) := b"0000000000000000_0000000000000000_0010001011010010_0100111011111000"; -- 0.13602155266180993
	pesos_i(15375) := b"0000000000000000_0000000000000000_0010000000011101_1100010100110000"; -- 0.12545425817376382
	pesos_i(15376) := b"0000000000000000_0000000000000000_0010011000001101_1101010000111010"; -- 0.14864851387270953
	pesos_i(15377) := b"0000000000000000_0000000000000000_0000111100110110_0100110010100010"; -- 0.05942229234255098
	pesos_i(15378) := b"1111111111111111_1111111111111111_1110111001000000_1011000001111001"; -- -0.06932541894235048
	pesos_i(15379) := b"0000000000000000_0000000000000000_0001011000110100_1111111010001110"; -- 0.08674612976391387
	pesos_i(15380) := b"0000000000000000_0000000000000000_0000000011011111_0101100010011111"; -- 0.0034079922211915892
	pesos_i(15381) := b"0000000000000000_0000000000000000_0001001000000101_1010000000101011"; -- 0.07039834064335355
	pesos_i(15382) := b"1111111111111111_1111111111111111_1101100110111010_1001001000000000"; -- -0.14949691299508494
	pesos_i(15383) := b"0000000000000000_0000000000000000_0001110111011110_0010010110111110"; -- 0.11667095082025424
	pesos_i(15384) := b"1111111111111111_1111111111111111_1110100001011001_1010110111000101"; -- -0.09238161033828357
	pesos_i(15385) := b"1111111111111111_1111111111111111_1111010101111010_1011100011100010"; -- -0.041096157940338135
	pesos_i(15386) := b"1111111111111111_1111111111111111_1111100000110101_1001011110100011"; -- -0.030432245895820983
	pesos_i(15387) := b"1111111111111111_1111111111111111_1110110001100011_1000101101011100"; -- -0.07660607351625338
	pesos_i(15388) := b"1111111111111111_1111111111111111_1111101100100110_1010111100110100"; -- -0.018940972993908872
	pesos_i(15389) := b"0000000000000000_0000000000000000_0001011111100011_1010111100100000"; -- 0.0933179332687808
	pesos_i(15390) := b"1111111111111111_1111111111111111_1101110110101010_1100001110110111"; -- -0.1341130902305681
	pesos_i(15391) := b"0000000000000000_0000000000000000_0000010101001011_1010110010011110"; -- 0.02068594801333601
	pesos_i(15392) := b"1111111111111111_1111111111111111_1110111101000111_1001101000010011"; -- -0.06531369248529748
	pesos_i(15393) := b"0000000000000000_0000000000000000_0000111110110001_1111001101100001"; -- 0.061309062291397716
	pesos_i(15394) := b"0000000000000000_0000000000000000_0010100001001100_1001000110110011"; -- 0.1574183522204029
	pesos_i(15395) := b"1111111111111111_1111111111111111_1111011010011100_0101100001110101"; -- -0.036676856381770914
	pesos_i(15396) := b"1111111111111111_1111111111111111_1101110111100000_0111001010011010"; -- -0.13329395049481654
	pesos_i(15397) := b"1111111111111111_1111111111111111_1110000110101100_0100100101110101"; -- -0.11846485996219183
	pesos_i(15398) := b"1111111111111111_1111111111111111_1111111010110001_0110010110101111"; -- -0.005105633406623713
	pesos_i(15399) := b"1111111111111111_1111111111111111_1110110010010001_0010001101011010"; -- -0.07591036840223808
	pesos_i(15400) := b"0000000000000000_0000000000000000_0001110111001110_0011011100100111"; -- 0.1164278479593184
	pesos_i(15401) := b"0000000000000000_0000000000000000_0000111001001000_1000010011011000"; -- 0.055794051018828235
	pesos_i(15402) := b"0000000000000000_0000000000000000_0001101110011111_1001001010000001"; -- 0.1079036298858133
	pesos_i(15403) := b"1111111111111111_1111111111111111_1110011100011010_1011101110111011"; -- -0.09724833178836563
	pesos_i(15404) := b"0000000000000000_0000000000000000_0010001101111010_0110001110110011"; -- 0.1385862647502611
	pesos_i(15405) := b"1111111111111111_1111111111111111_1111100000111101_1001010011100110"; -- -0.03031033879354494
	pesos_i(15406) := b"0000000000000000_0000000000000000_0000001001100101_0100110111100111"; -- 0.009358281085955041
	pesos_i(15407) := b"0000000000000000_0000000000000000_0010001001101001_0000000101001100"; -- 0.13441475009973353
	pesos_i(15408) := b"1111111111111111_1111111111111111_1101111001010100_0101111011101001"; -- -0.1315251045417763
	pesos_i(15409) := b"0000000000000000_0000000000000000_0000101111010010_1101011000101010"; -- 0.04618586093883695
	pesos_i(15410) := b"0000000000000000_0000000000000000_0001011001101000_0011101100100011"; -- 0.0875279389589487
	pesos_i(15411) := b"0000000000000000_0000000000000000_0001110110010001_0001001001100001"; -- 0.11549486988106787
	pesos_i(15412) := b"0000000000000000_0000000000000000_0000010000011001_0101110001001101"; -- 0.01601197132516946
	pesos_i(15413) := b"1111111111111111_1111111111111111_1110110001110011_0000100000111001"; -- -0.07636974909700399
	pesos_i(15414) := b"0000000000000000_0000000000000000_0000101100111000_1111011001100011"; -- 0.043837927884358266
	pesos_i(15415) := b"0000000000000000_0000000000000000_0000001111111100_0011100101100111"; -- 0.015567386316768022
	pesos_i(15416) := b"0000000000000000_0000000000000000_0010011011000000_1110000101010000"; -- 0.1513806171772706
	pesos_i(15417) := b"0000000000000000_0000000000000000_0001101100100101_0011110001000100"; -- 0.10603691734822404
	pesos_i(15418) := b"1111111111111111_1111111111111111_1111100101011000_1010110010110111"; -- -0.025990682060542943
	pesos_i(15419) := b"0000000000000000_0000000000000000_0010000110111111_0001100101100011"; -- 0.13182219194016995
	pesos_i(15420) := b"1111111111111111_1111111111111111_1110110000001010_0001100101010000"; -- -0.07797090337330954
	pesos_i(15421) := b"1111111111111111_1111111111111111_1110100011011000_1000101001110101"; -- -0.09044584878567784
	pesos_i(15422) := b"0000000000000000_0000000000000000_0001000100000010_1000111100000111"; -- 0.06644529272110673
	pesos_i(15423) := b"1111111111111111_1111111111111111_1110011100100011_0010100111100011"; -- -0.0971196957929365
	pesos_i(15424) := b"0000000000000000_0000000000000000_0001101011000001_1001111101111000"; -- 0.10451695144204506
	pesos_i(15425) := b"1111111111111111_1111111111111111_1110010111000101_0010110111001101"; -- -0.10246003859642182
	pesos_i(15426) := b"0000000000000000_0000000000000000_0001100111001111_1111101101110101"; -- 0.10082980729011168
	pesos_i(15427) := b"0000000000000000_0000000000000000_0010000011001000_0100001000110110"; -- 0.1280557041791831
	pesos_i(15428) := b"1111111111111111_1111111111111111_1101101110111111_0100110101000000"; -- -0.14161221682158817
	pesos_i(15429) := b"0000000000000000_0000000000000000_0000111100100111_0010110000001100"; -- 0.05919146825303312
	pesos_i(15430) := b"1111111111111111_1111111111111111_1110101101000001_0100010000111101"; -- -0.08103536149615735
	pesos_i(15431) := b"0000000000000000_0000000000000000_0001000010000111_1011101100111100"; -- 0.06457109660125614
	pesos_i(15432) := b"0000000000000000_0000000000000000_0010000101011000_1100100111010110"; -- 0.1302610538724256
	pesos_i(15433) := b"0000000000000000_0000000000000000_0000011110101100_1101111000001000"; -- 0.029981495783733665
	pesos_i(15434) := b"1111111111111111_1111111111111111_1101011110111010_0011110100001000"; -- -0.15731447751745267
	pesos_i(15435) := b"0000000000000000_0000000000000000_0000111111001000_1011000011101110"; -- 0.061656053530020134
	pesos_i(15436) := b"1111111111111111_1111111111111111_1111100001000000_1000101010111101"; -- -0.03026516811974238
	pesos_i(15437) := b"1111111111111111_1111111111111111_1110100101100010_1101000010010011"; -- -0.08833595656805768
	pesos_i(15438) := b"0000000000000000_0000000000000000_0010011011000110_0010110101111101"; -- 0.15146145161362196
	pesos_i(15439) := b"1111111111111111_1111111111111111_1111101001011100_0010000100101100"; -- -0.0220317142711628
	pesos_i(15440) := b"0000000000000000_0000000000000000_0000000101110010_1011000101101111"; -- 0.0056563278230903884
	pesos_i(15441) := b"1111111111111111_1111111111111111_1110000111110011_0111111100111110"; -- -0.11737828012815696
	pesos_i(15442) := b"0000000000000000_0000000000000000_0000011011011011_1011101010101111"; -- 0.026790301975921967
	pesos_i(15443) := b"0000000000000000_0000000000000000_0001001011011010_1110010110000000"; -- 0.07365259519612455
	pesos_i(15444) := b"1111111111111111_1111111111111111_1101111111000101_1111111000110101"; -- -0.12588511661771437
	pesos_i(15445) := b"1111111111111111_1111111111111111_1110110100011010_0100001101011010"; -- -0.07381800703429749
	pesos_i(15446) := b"1111111111111111_1111111111111111_1101100000110000_1111011001001101"; -- -0.15550289744642345
	pesos_i(15447) := b"1111111111111111_1111111111111111_1110110011000001_0001001000101011"; -- -0.07517897092731056
	pesos_i(15448) := b"0000000000000000_0000000000000000_0001011101101000_1001110110000001"; -- 0.09144005192346932
	pesos_i(15449) := b"0000000000000000_0000000000000000_0001101111110010_0110110100111100"; -- 0.10916788778491858
	pesos_i(15450) := b"1111111111111111_1111111111111111_1111111000011110_0110010011100010"; -- -0.007348723348877714
	pesos_i(15451) := b"1111111111111111_1111111111111111_1110010110011011_0110001101110101"; -- -0.10309770968938368
	pesos_i(15452) := b"1111111111111111_1111111111111111_1110011001001101_1110110110111100"; -- -0.10037340314623892
	pesos_i(15453) := b"1111111111111111_1111111111111111_1111100111100011_0000110111000110"; -- -0.02387918384387779
	pesos_i(15454) := b"1111111111111111_1111111111111111_1111000011101111_0001101011000010"; -- -0.05885155454509593
	pesos_i(15455) := b"0000000000000000_0000000000000000_0001010111111110_0001001111100110"; -- 0.08590816852138793
	pesos_i(15456) := b"1111111111111111_1111111111111111_1110100111010110_0001100011100101"; -- -0.08657688539462244
	pesos_i(15457) := b"1111111111111111_1111111111111111_1110001101100100_0111010111110011"; -- -0.1117483408167873
	pesos_i(15458) := b"0000000000000000_0000000000000000_0010001101000110_0111111111101101"; -- 0.1377944902341521
	pesos_i(15459) := b"1111111111111111_1111111111111111_1111000001110011_1000001010111010"; -- -0.06073744735859943
	pesos_i(15460) := b"0000000000000000_0000000000000000_0001011100101001_0101101001000000"; -- 0.09047473973927694
	pesos_i(15461) := b"0000000000000000_0000000000000000_0001001100010101_0001011000101101"; -- 0.07454050643341001
	pesos_i(15462) := b"1111111111111111_1111111111111111_1111011100011011_0001000111001001"; -- -0.03474320257013297
	pesos_i(15463) := b"0000000000000000_0000000000000000_0000111001110111_0010101010011111"; -- 0.056505836328382505
	pesos_i(15464) := b"0000000000000000_0000000000000000_0000010101111101_0101101010100110"; -- 0.021444001762967825
	pesos_i(15465) := b"0000000000000000_0000000000000000_0001001110100110_0111001000100000"; -- 0.07675851145666202
	pesos_i(15466) := b"1111111111111111_1111111111111111_1111011101010010_0011101111010100"; -- -0.033901463166188556
	pesos_i(15467) := b"1111111111111111_1111111111111111_1110001110011000_1010001101011101"; -- -0.11095217695768876
	pesos_i(15468) := b"1111111111111111_1111111111111111_1111110100101000_0001100100010100"; -- -0.011106903706982314
	pesos_i(15469) := b"1111111111111111_1111111111111111_1110010010000110_0000011001101111"; -- -0.10732993870867387
	pesos_i(15470) := b"0000000000000000_0000000000000000_0010010000100111_0000100101100010"; -- 0.14122065203131437
	pesos_i(15471) := b"1111111111111111_1111111111111111_1110001101010000_1011010000010011"; -- -0.11204981362204808
	pesos_i(15472) := b"0000000000000000_0000000000000000_0001001111011111_0011110100010001"; -- 0.07762509975241604
	pesos_i(15473) := b"1111111111111111_1111111111111111_1101111101011001_0111000000011011"; -- -0.12754153572452098
	pesos_i(15474) := b"0000000000000000_0000000000000000_0001000110010011_1100111101111110"; -- 0.06866165951536154
	pesos_i(15475) := b"1111111111111111_1111111111111111_1111110101111011_1100101011110100"; -- -0.009829821914505099
	pesos_i(15476) := b"0000000000000000_0000000000000000_0001001110101101_1100110010110110"; -- 0.07687072222516778
	pesos_i(15477) := b"0000000000000000_0000000000000000_0001111001010110_1101101011111000"; -- 0.11851280748856537
	pesos_i(15478) := b"1111111111111111_1111111111111111_1110100101101011_0101111100110000"; -- -0.0882053858462033
	pesos_i(15479) := b"0000000000000000_0000000000000000_0001011110010101_0000011101110110"; -- 0.09211775435666822
	pesos_i(15480) := b"0000000000000000_0000000000000000_0001100011101010_1110100011111110"; -- 0.09733444406234801
	pesos_i(15481) := b"1111111111111111_1111111111111111_1110100001110010_1100110010010000"; -- -0.09199830525318299
	pesos_i(15482) := b"1111111111111111_1111111111111111_1111011000001011_0001100000000100"; -- -0.03889322193883459
	pesos_i(15483) := b"1111111111111111_1111111111111111_1110110001101010_1000010111111111"; -- -0.07649958148967015
	pesos_i(15484) := b"0000000000000000_0000000000000000_0010010100011001_0100001000110100"; -- 0.14491666582492507
	pesos_i(15485) := b"1111111111111111_1111111111111111_1111101101110000_0000111000101100"; -- -0.017821420800517962
	pesos_i(15486) := b"1111111111111111_1111111111111111_1111110000001101_1001110101011101"; -- -0.015417256069787921
	pesos_i(15487) := b"1111111111111111_1111111111111111_1111010010001101_0011100010111110"; -- -0.044720128756588005
	pesos_i(15488) := b"0000000000000000_0000000000000000_0000001001010110_0001010010111000"; -- 0.009125990780292777
	pesos_i(15489) := b"1111111111111111_1111111111111111_1110011101101011_0011101001110101"; -- -0.0960200753204707
	pesos_i(15490) := b"0000000000000000_0000000000000000_0001111001100001_0010111110101110"; -- 0.11867044435996828
	pesos_i(15491) := b"0000000000000000_0000000000000000_0001101011010111_1110000000001001"; -- 0.10485649315267229
	pesos_i(15492) := b"0000000000000000_0000000000000000_0010000101100010_1010011110001000"; -- 0.13041159707653135
	pesos_i(15493) := b"1111111111111111_1111111111111111_1101100110001010_1001010000101001"; -- -0.15022920602156328
	pesos_i(15494) := b"1111111111111111_1111111111111111_1110111111101010_1101001111100001"; -- -0.06282306448957402
	pesos_i(15495) := b"1111111111111111_1111111111111111_1110000110011110_1110001100001101"; -- -0.11866932796269258
	pesos_i(15496) := b"0000000000000000_0000000000000000_0010011110001001_1101110100011100"; -- 0.15444738327971544
	pesos_i(15497) := b"0000000000000000_0000000000000000_0000011110000100_0101101111110000"; -- 0.029363390041891646
	pesos_i(15498) := b"0000000000000000_0000000000000000_0001001001001000_1010000001000011"; -- 0.07142068520902561
	pesos_i(15499) := b"0000000000000000_0000000000000000_0001011011101101_1011101100000111"; -- 0.0895649806236459
	pesos_i(15500) := b"1111111111111111_1111111111111111_1110100000110110_0011111110011000"; -- -0.09292223496488071
	pesos_i(15501) := b"0000000000000000_0000000000000000_0010010011100111_1110000000010100"; -- 0.1441631362678124
	pesos_i(15502) := b"0000000000000000_0000000000000000_0000000101010000_0101111111111110"; -- 0.00513267462550687
	pesos_i(15503) := b"0000000000000000_0000000000000000_0000110011011100_0001001001101011"; -- 0.050233031348594526
	pesos_i(15504) := b"1111111111111111_1111111111111111_1111100110101000_0010001111111001"; -- -0.02477812934638108
	pesos_i(15505) := b"1111111111111111_1111111111111111_1110101001100000_1111100101100001"; -- -0.08445779206158945
	pesos_i(15506) := b"0000000000000000_0000000000000000_0001010010100010_0001000010100010"; -- 0.08059791533611546
	pesos_i(15507) := b"1111111111111111_1111111111111111_1111001010000100_0000010111110000"; -- -0.05267298593912441
	pesos_i(15508) := b"0000000000000000_0000000000000000_0001110010001100_1100011001010001"; -- 0.11152305093325943
	pesos_i(15509) := b"1111111111111111_1111111111111111_1111011001110010_0011111100111110"; -- -0.03731922852476707
	pesos_i(15510) := b"0000000000000000_0000000000000000_0001101010010011_0100011001010011"; -- 0.10380973362594756
	pesos_i(15511) := b"0000000000000000_0000000000000000_0010001011000000_0001001100011000"; -- 0.13574332567930525
	pesos_i(15512) := b"0000000000000000_0000000000000000_0001101101000110_0011011000001101"; -- 0.10654008693239442
	pesos_i(15513) := b"0000000000000000_0000000000000000_0001001001011101_1011001110001000"; -- 0.07174226826939209
	pesos_i(15514) := b"0000000000000000_0000000000000000_0010010100001010_0101101001000101"; -- 0.14468921840957236
	pesos_i(15515) := b"0000000000000000_0000000000000000_0000001000011100_0110000111100111"; -- 0.008245581567477487
	pesos_i(15516) := b"1111111111111111_1111111111111111_1110011010110101_1010110110101010"; -- -0.09879030791939816
	pesos_i(15517) := b"0000000000000000_0000000000000000_0001001010110101_1111100000001110"; -- 0.0730891259501571
	pesos_i(15518) := b"0000000000000000_0000000000000000_0001111100010011_1001000001110001"; -- 0.12139227645892131
	pesos_i(15519) := b"0000000000000000_0000000000000000_0000100010000101_0101000101110000"; -- 0.03328427299784622
	pesos_i(15520) := b"0000000000000000_0000000000000000_0010001101001110_0100000000000000"; -- 0.13791275018683521
	pesos_i(15521) := b"1111111111111111_1111111111111111_1111110101101010_0101010001111010"; -- -0.010096283060156593
	pesos_i(15522) := b"0000000000000000_0000000000000000_0001010111101101_0110001111110011"; -- 0.08565354038440479
	pesos_i(15523) := b"0000000000000000_0000000000000000_0001111000000110_1001100001001011"; -- 0.11728813013935
	pesos_i(15524) := b"0000000000000000_0000000000000000_0000101100011000_0000110001000110"; -- 0.043335692548924075
	pesos_i(15525) := b"1111111111111111_1111111111111111_1111111000100100_0111000001011111"; -- -0.007256485771354488
	pesos_i(15526) := b"0000000000000000_0000000000000000_0000111101011000_0111011110001000"; -- 0.059943648144321515
	pesos_i(15527) := b"1111111111111111_1111111111111111_1110110010101111_1011111011000100"; -- -0.07544334149463167
	pesos_i(15528) := b"0000000000000000_0000000000000000_0010000100110000_1100000101100100"; -- 0.12965019894730895
	pesos_i(15529) := b"1111111111111111_1111111111111111_1111100110011000_1010000100110001"; -- -0.02501480625351089
	pesos_i(15530) := b"1111111111111111_1111111111111111_1110010100111101_1010001001110101"; -- -0.10452828064520238
	pesos_i(15531) := b"1111111111111111_1111111111111111_1101111100100101_1101111011001100"; -- -0.1283283950683804
	pesos_i(15532) := b"1111111111111111_1111111111111111_1110010111010100_0111010111101101"; -- -0.10222685788812365
	pesos_i(15533) := b"1111111111111111_1111111111111111_1111111111010110_1111010000110000"; -- -0.0006263143873450892
	pesos_i(15534) := b"0000000000000000_0000000000000000_0000111000110010_0111111110011011"; -- 0.055458045283071
	pesos_i(15535) := b"1111111111111111_1111111111111111_1110010001011010_0101011100111111"; -- -0.10799650880554258
	pesos_i(15536) := b"1111111111111111_1111111111111111_1111111011010111_0000011110000011"; -- -0.004531412689507341
	pesos_i(15537) := b"0000000000000000_0000000000000000_0010010101001110_1010011100011010"; -- 0.14573139555627024
	pesos_i(15538) := b"1111111111111111_1111111111111111_1111000010110101_1010001001101100"; -- -0.059728478049451535
	pesos_i(15539) := b"0000000000000000_0000000000000000_0010010011010100_0001111000101110"; -- 0.14386166206451703
	pesos_i(15540) := b"1111111111111111_1111111111111111_1111011100000000_1010011010010001"; -- -0.035146321935548994
	pesos_i(15541) := b"0000000000000000_0000000000000000_0001100111101011_0110101111101110"; -- 0.10124849845593252
	pesos_i(15542) := b"1111111111111111_1111111111111111_1110010110011101_1101001010011110"; -- -0.10306056625755813
	pesos_i(15543) := b"0000000000000000_0000000000000000_0001000010010001_0101000111010111"; -- 0.06471740254030361
	pesos_i(15544) := b"1111111111111111_1111111111111111_1110101100100000_0011010001100100"; -- -0.08153984598712362
	pesos_i(15545) := b"0000000000000000_0000000000000000_0000001100010010_0011000011000010"; -- 0.011996314363761437
	pesos_i(15546) := b"0000000000000000_0000000000000000_0001110110100010_0000001000110010"; -- 0.11575330468684575
	pesos_i(15547) := b"1111111111111111_1111111111111111_1101110101010001_0010101110011001"; -- -0.13548018949556276
	pesos_i(15548) := b"1111111111111111_1111111111111111_1110100110101000_0111010111110101"; -- -0.08727324271471541
	pesos_i(15549) := b"0000000000000000_0000000000000000_0001110101100000_1111100101111100"; -- 0.11476096421714492
	pesos_i(15550) := b"0000000000000000_0000000000000000_0000000110100110_0011010010011001"; -- 0.006442343950521994
	pesos_i(15551) := b"0000000000000000_0000000000000000_0010010010001110_1010011011111111"; -- 0.14280170171401632
	pesos_i(15552) := b"0000000000000000_0000000000000000_0010000101000110_0010000110010010"; -- 0.12997636612850613
	pesos_i(15553) := b"1111111111111111_1111111111111111_1110101101101110_0001100001011000"; -- -0.08035133212806539
	pesos_i(15554) := b"0000000000000000_0000000000000000_0000100000110101_1110010001010000"; -- 0.03207232432905424
	pesos_i(15555) := b"0000000000000000_0000000000000000_0001101111010110_1010001010011110"; -- 0.1087438236056228
	pesos_i(15556) := b"0000000000000000_0000000000000000_0001101111011101_0010110011011111"; -- 0.10884361687883315
	pesos_i(15557) := b"0000000000000000_0000000000000000_0000101101000010_1110101110110011"; -- 0.043989878806015605
	pesos_i(15558) := b"1111111111111111_1111111111111111_1101111101100000_1000001001110001"; -- -0.12743363143353956
	pesos_i(15559) := b"1111111111111111_1111111111111111_1110011101101011_0110100111101100"; -- -0.09601724604095294
	pesos_i(15560) := b"0000000000000000_0000000000000000_0010010000011000_1011111110110000"; -- 0.1410026365031272
	pesos_i(15561) := b"1111111111111111_1111111111111111_1110010000000110_1101110010111001"; -- -0.10927029122205688
	pesos_i(15562) := b"0000000000000000_0000000000000000_0001001110011000_0101011001011100"; -- 0.07654323339871971
	pesos_i(15563) := b"1111111111111111_1111111111111111_1111101100010011_1001111111111110"; -- -0.019231796776971864
	pesos_i(15564) := b"0000000000000000_0000000000000000_0001100011001010_0000010101010001"; -- 0.09683259231603975
	pesos_i(15565) := b"0000000000000000_0000000000000000_0000000010100011_0000010110110000"; -- 0.0024875215170346104
	pesos_i(15566) := b"0000000000000000_0000000000000000_0010100001001111_1111010010010011"; -- 0.1574700220149149
	pesos_i(15567) := b"1111111111111111_1111111111111111_1110010111000010_1000011101100001"; -- -0.1025004756696327
	pesos_i(15568) := b"1111111111111111_1111111111111111_1111100111111010_1110101010101000"; -- -0.023515066151212245
	pesos_i(15569) := b"1111111111111111_1111111111111111_1110111000100011_1011011000000111"; -- -0.06976759266518041
	pesos_i(15570) := b"0000000000000000_0000000000000000_0000110100000001_0101101000101101"; -- 0.0508018837908721
	pesos_i(15571) := b"1111111111111111_1111111111111111_1110100000101101_1110000111100000"; -- -0.09304989127562856
	pesos_i(15572) := b"1111111111111111_1111111111111111_1111110000000000_1000100011100111"; -- -0.015616840078913815
	pesos_i(15573) := b"0000000000000000_0000000000000000_0001011100111111_1010110111101110"; -- 0.09081542084124071
	pesos_i(15574) := b"1111111111111111_1111111111111111_1111101111111111_1001001111010101"; -- -0.015631447204794837
	pesos_i(15575) := b"0000000000000000_0000000000000000_0000001011100000_1101100001110011"; -- 0.011243370126074601
	pesos_i(15576) := b"0000000000000000_0000000000000000_0000101101001000_1111110000000001"; -- 0.04408240332245799
	pesos_i(15577) := b"1111111111111111_1111111111111111_1110011011111010_0111100101011000"; -- -0.09774057016709053
	pesos_i(15578) := b"0000000000000000_0000000000000000_0000101000000110_1100011000001100"; -- 0.03916585717461207
	pesos_i(15579) := b"1111111111111111_1111111111111111_1111010110111101_0101110110011110"; -- -0.04007925889837406
	pesos_i(15580) := b"1111111111111111_1111111111111111_1101111010110001_1110010011111000"; -- -0.13009804684831475
	pesos_i(15581) := b"1111111111111111_1111111111111111_1110011110001001_0100010000010110"; -- -0.09556173758400802
	pesos_i(15582) := b"0000000000000000_0000000000000000_0001000000111000_1011011110011010"; -- 0.06336543562852885
	pesos_i(15583) := b"0000000000000000_0000000000000000_0010001110100100_1110101010010001"; -- 0.13923517254095336
	pesos_i(15584) := b"1111111111111111_1111111111111111_1111110100110000_1010010010101000"; -- -0.010976513960204265
	pesos_i(15585) := b"0000000000000000_0000000000000000_0000010100101110_0011100101010000"; -- 0.020236570435926842
	pesos_i(15586) := b"1111111111111111_1111111111111111_1110110001111010_1011001111010001"; -- -0.07625270979499377
	pesos_i(15587) := b"0000000000000000_0000000000000000_0001110110101110_1011100111100100"; -- 0.11594735918531553
	pesos_i(15588) := b"0000000000000000_0000000000000000_0001000010101111_1000001000111001"; -- 0.06517804989499063
	pesos_i(15589) := b"0000000000000000_0000000000000000_0001111010000110_0000100000011111"; -- 0.1192326618308219
	pesos_i(15590) := b"1111111111111111_1111111111111111_1101010101011011_0011011101011100"; -- -0.16657690051241353
	pesos_i(15591) := b"1111111111111111_1111111111111111_1110001010110000_0000100000011001"; -- -0.11450147040278238
	pesos_i(15592) := b"0000000000000000_0000000000000000_0010010100100011_0111010010011000"; -- 0.14507225704028162
	pesos_i(15593) := b"1111111111111111_1111111111111111_1111001110110011_1010001011010110"; -- -0.048040221071222605
	pesos_i(15594) := b"1111111111111111_1111111111111111_1110001110100000_1010101110000110"; -- -0.110829620187047
	pesos_i(15595) := b"0000000000000000_0000000000000000_0010001010100110_0100110010100001"; -- 0.13535002636858265
	pesos_i(15596) := b"1111111111111111_1111111111111111_1110110010010000_1100111110110101"; -- -0.07591535405325885
	pesos_i(15597) := b"1111111111111111_1111111111111111_1111001011001100_0001000100101011"; -- -0.05157368384251917
	pesos_i(15598) := b"0000000000000000_0000000000000000_0001011100001010_0110100010100111"; -- 0.0900025756610477
	pesos_i(15599) := b"1111111111111111_1111111111111111_1111001110110100_1010010110000001"; -- -0.0480248032153593
	pesos_i(15600) := b"1111111111111111_1111111111111111_1110011000111001_1110010111101011"; -- -0.10067904482098525
	pesos_i(15601) := b"0000000000000000_0000000000000000_0000010101110010_0101100110111011"; -- 0.021276100318031343
	pesos_i(15602) := b"0000000000000000_0000000000000000_0000101100010110_0100010000001000"; -- 0.043308498278647356
	pesos_i(15603) := b"0000000000000000_0000000000000000_0001001100000110_0010110100110100"; -- 0.07431299699610752
	pesos_i(15604) := b"0000000000000000_0000000000000000_0010000000111001_1000000101000010"; -- 0.1258774553363524
	pesos_i(15605) := b"0000000000000000_0000000000000000_0000100010010101_0110100000011111"; -- 0.03352976573862496
	pesos_i(15606) := b"1111111111111111_1111111111111111_1111011100011011_0010010110110010"; -- -0.034742015876465436
	pesos_i(15607) := b"1111111111111111_1111111111111111_1110110001111000_1100000000111110"; -- -0.0762824868580548
	pesos_i(15608) := b"0000000000000000_0000000000000000_0001010100000010_0000101101111101"; -- 0.08206245239451822
	pesos_i(15609) := b"1111111111111111_1111111111111111_1110011111100110_1111101111111101"; -- -0.09413170880171097
	pesos_i(15610) := b"1111111111111111_1111111111111111_1110000000011110_1001101111000111"; -- -0.124532951221434
	pesos_i(15611) := b"1111111111111111_1111111111111111_1110100100111010_1011001010110011"; -- -0.08894808891488648
	pesos_i(15612) := b"1111111111111111_1111111111111111_1110001100001011_1110101000110011"; -- -0.1130994438870314
	pesos_i(15613) := b"1111111111111111_1111111111111111_1111010011010000_0011001001011010"; -- -0.04369817062226487
	pesos_i(15614) := b"1111111111111111_1111111111111111_1110101001000101_1100001101000110"; -- -0.08487300441984535
	pesos_i(15615) := b"0000000000000000_0000000000000000_0000101100000101_0010010000100101"; -- 0.043047198387402
	pesos_i(15616) := b"1111111111111111_1111111111111111_1110010110100011_1111110010101000"; -- -0.10296650787754541
	pesos_i(15617) := b"1111111111111111_1111111111111111_1111000011101111_1001010000111011"; -- -0.05884431408387914
	pesos_i(15618) := b"0000000000000000_0000000000000000_0000000110010110_1111100000001111"; -- 0.006209853845044751
	pesos_i(15619) := b"0000000000000000_0000000000000000_0000111001010101_0101101010010011"; -- 0.055989895820081494
	pesos_i(15620) := b"1111111111111111_1111111111111111_1111001001100010_0110001000101001"; -- -0.053186287967024626
	pesos_i(15621) := b"0000000000000000_0000000000000000_0000110100000011_1111011000010011"; -- 0.050841693556570484
	pesos_i(15622) := b"0000000000000000_0000000000000000_0001011000110001_1001001010010000"; -- 0.086693916512551
	pesos_i(15623) := b"1111111111111111_1111111111111111_1101111000101001_1001100011100001"; -- -0.13217777729823843
	pesos_i(15624) := b"1111111111111111_1111111111111111_1110101000010110_0000010100011011"; -- -0.08560150244564953
	pesos_i(15625) := b"0000000000000000_0000000000000000_0001111101110011_1110100100010001"; -- 0.12286240261308973
	pesos_i(15626) := b"1111111111111111_1111111111111111_1110101101110110_0110010101000010"; -- -0.08022467749570662
	pesos_i(15627) := b"1111111111111111_1111111111111111_1111001111000011_0010001000001111"; -- -0.04780375611959745
	pesos_i(15628) := b"1111111111111111_1111111111111111_1101101100111010_0100011110010001"; -- -0.14364197454088581
	pesos_i(15629) := b"1111111111111111_1111111111111111_1110110001010000_1011000100010111"; -- -0.07689374159569076
	pesos_i(15630) := b"1111111111111111_1111111111111111_1111010111011100_1001110010110110"; -- -0.03960247559932296
	pesos_i(15631) := b"1111111111111111_1111111111111111_1110111001001100_1001000001110100"; -- -0.06914422200571765
	pesos_i(15632) := b"1111111111111111_1111111111111111_1110111011001101_0010110111111110"; -- -0.06718170684239924
	pesos_i(15633) := b"1111111111111111_1111111111111111_1110010010100000_0101001001001101"; -- -0.10692868827165421
	pesos_i(15634) := b"1111111111111111_1111111111111111_1111011001010010_0100010110111100"; -- -0.037807122905990816
	pesos_i(15635) := b"0000000000000000_0000000000000000_0001011101011000_1111111100001000"; -- 0.09120172442441273
	pesos_i(15636) := b"0000000000000000_0000000000000000_0001111001111010_1111101100101010"; -- 0.11906404274307736
	pesos_i(15637) := b"1111111111111111_1111111111111111_1111100001000100_1000101110100101"; -- -0.030204078824909546
	pesos_i(15638) := b"1111111111111111_1111111111111111_1111100101100101_0100101000100100"; -- -0.025798193118567767
	pesos_i(15639) := b"1111111111111111_1111111111111111_1111001101001001_0001111000011100"; -- -0.04966556378106556
	pesos_i(15640) := b"1111111111111111_1111111111111111_1110001110110110_0010010000000011"; -- -0.11050200391468504
	pesos_i(15641) := b"1111111111111111_1111111111111111_1110111111111100_1110010001111011"; -- -0.06254741657734586
	pesos_i(15642) := b"1111111111111111_1111111111111111_1110101101010101_1110101010010001"; -- -0.08072027175117455
	pesos_i(15643) := b"0000000000000000_0000000000000000_0001110010101100_0101111011001001"; -- 0.11200516146947435
	pesos_i(15644) := b"0000000000000000_0000000000000000_0010000101010110_0101001111100111"; -- 0.1302235067705361
	pesos_i(15645) := b"0000000000000000_0000000000000000_0001100110111111_0000110011111111"; -- 0.10057145335839177
	pesos_i(15646) := b"1111111111111111_1111111111111111_1110100100100010_1001011011101000"; -- -0.08931595648333364
	pesos_i(15647) := b"0000000000000000_0000000000000000_0000011000110110_1010000010001001"; -- 0.024271043267845193
	pesos_i(15648) := b"1111111111111111_1111111111111111_1111101100000100_1001100010000110"; -- -0.019461123670657315
	pesos_i(15649) := b"1111111111111111_1111111111111111_1110110010100101_0011001000000000"; -- -0.07560431961396431
	pesos_i(15650) := b"1111111111111111_1111111111111111_1110111001111010_1100000001011011"; -- -0.06843946245716859
	pesos_i(15651) := b"1111111111111111_1111111111111111_1101101111100000_0010110101010100"; -- -0.14111057936735627
	pesos_i(15652) := b"1111111111111111_1111111111111111_1101111110101001_1001011111000100"; -- -0.12631846865328766
	pesos_i(15653) := b"1111111111111111_1111111111111111_1101101110011001_1011011111101010"; -- -0.14218569306987588
	pesos_i(15654) := b"1111111111111111_1111111111111111_1101100001111000_1001001101000101"; -- -0.15441016738615712
	pesos_i(15655) := b"1111111111111111_1111111111111111_1111110011001011_0111100101000001"; -- -0.012520238638096934
	pesos_i(15656) := b"1111111111111111_1111111111111111_1111001011010101_1011010110111100"; -- -0.05142654574319775
	pesos_i(15657) := b"0000000000000000_0000000000000000_0001010010100101_0011010011110000"; -- 0.0806458555056468
	pesos_i(15658) := b"1111111111111111_1111111111111111_1111000011111110_1100010110010101"; -- -0.058612490689681294
	pesos_i(15659) := b"1111111111111111_1111111111111111_1110101101100111_1101101011111110"; -- -0.08044654182685156
	pesos_i(15660) := b"1111111111111111_1111111111111111_1110010111111000_1011111111010100"; -- -0.10167313652274249
	pesos_i(15661) := b"1111111111111111_1111111111111111_1110100010011101_1010011001111101"; -- -0.09134444669107272
	pesos_i(15662) := b"0000000000000000_0000000000000000_0001010000110010_0001001000011001"; -- 0.07888901809444335
	pesos_i(15663) := b"0000000000000000_0000000000000000_0001101110100110_1111100111010110"; -- 0.10801660041218131
	pesos_i(15664) := b"0000000000000000_0000000000000000_0010001111001011_1010010001101000"; -- 0.13982608346588643
	pesos_i(15665) := b"0000000000000000_0000000000000000_0000011101100010_0001001001110100"; -- 0.02884021118521021
	pesos_i(15666) := b"1111111111111111_1111111111111111_1101111010001011_1000101110011011"; -- -0.13068320721802262
	pesos_i(15667) := b"1111111111111111_1111111111111111_1110001110011110_1100001000001101"; -- -0.11085879506749145
	pesos_i(15668) := b"0000000000000000_0000000000000000_0000110011010010_1111011000100000"; -- 0.05009401593231947
	pesos_i(15669) := b"1111111111111111_1111111111111111_1110110111101001_1110100001011111"; -- -0.07064960175849559
	pesos_i(15670) := b"0000000000000000_0000000000000000_0000011110000101_0101100000110011"; -- 0.029378426141109356
	pesos_i(15671) := b"1111111111111111_1111111111111111_1110100001011010_0000111000111000"; -- -0.09237586156640017
	pesos_i(15672) := b"0000000000000000_0000000000000000_0000000010001110_0101001011011101"; -- 0.0021716871122968735
	pesos_i(15673) := b"1111111111111111_1111111111111111_1101101010101001_1110011000101100"; -- -0.1458450452842811
	pesos_i(15674) := b"1111111111111111_1111111111111111_1111000011011110_1101011001000010"; -- -0.05909977803182875
	pesos_i(15675) := b"1111111111111111_1111111111111111_1111100010000001_0110010100010010"; -- -0.02927559185293686
	pesos_i(15676) := b"1111111111111111_1111111111111111_1111010110010000_1010000010110001"; -- -0.04076190636156088
	pesos_i(15677) := b"1111111111111111_1111111111111111_1111111111100011_0100000001100100"; -- -0.0004386668489192294
	pesos_i(15678) := b"1111111111111111_1111111111111111_1110000010110111_1110100110010000"; -- -0.12219372017191793
	pesos_i(15679) := b"0000000000000000_0000000000000000_0001001101001110_1001110001011000"; -- 0.07541825441241282
	pesos_i(15680) := b"1111111111111111_1111111111111111_1111001101001110_1010001111010001"; -- -0.04958130014909354
	pesos_i(15681) := b"0000000000000000_0000000000000000_0000011011111000_1101101011110101"; -- 0.027234730616732795
	pesos_i(15682) := b"1111111111111111_1111111111111111_1110110010101101_1010000101010011"; -- -0.07547561384324658
	pesos_i(15683) := b"1111111111111111_1111111111111111_1111000000011100_0011001101000110"; -- -0.06206969776798549
	pesos_i(15684) := b"1111111111111111_1111111111111111_1111101011011110_1100110100111110"; -- -0.020037815388651598
	pesos_i(15685) := b"0000000000000000_0000000000000000_0001100101100111_0100110111101010"; -- 0.09923254938337606
	pesos_i(15686) := b"0000000000000000_0000000000000000_0001001101110101_0111000001101110"; -- 0.07601072961812062
	pesos_i(15687) := b"0000000000000000_0000000000000000_0001011011101000_1000110111001011"; -- 0.08948599061222766
	pesos_i(15688) := b"1111111111111111_1111111111111111_1111110001000111_1100111000010100"; -- -0.014529342861833053
	pesos_i(15689) := b"1111111111111111_1111111111111111_1110101011011011_0010110001110010"; -- -0.08259317614672708
	pesos_i(15690) := b"1111111111111111_1111111111111111_1110110011000111_1110110000101010"; -- -0.07507442459938383
	pesos_i(15691) := b"1111111111111111_1111111111111111_1101110110000111_0110011010101110"; -- -0.13465269336470664
	pesos_i(15692) := b"0000000000000000_0000000000000000_0001000110001001_0010000101011100"; -- 0.06849869251721293
	pesos_i(15693) := b"0000000000000000_0000000000000000_0001111110001001_0110011100010111"; -- 0.12319034863447485
	pesos_i(15694) := b"0000000000000000_0000000000000000_0001101111101010_1011011100111011"; -- 0.10905022794047918
	pesos_i(15695) := b"1111111111111111_1111111111111111_1110110100110001_0011110000101010"; -- -0.07346748320780637
	pesos_i(15696) := b"1111111111111111_1111111111111111_1101110010100010_1010000001100001"; -- -0.13814351676597558
	pesos_i(15697) := b"0000000000000000_0000000000000000_0001100000111010_1010110010000001"; -- 0.0946452917170625
	pesos_i(15698) := b"1111111111111111_1111111111111111_1111111111110010_0100100111011010"; -- -0.00020922106826555043
	pesos_i(15699) := b"1111111111111111_1111111111111111_1111011101001110_1011111111111011"; -- -0.03395462157026445
	pesos_i(15700) := b"1111111111111111_1111111111111111_1111011111010000_0110011010101101"; -- -0.03197630200073993
	pesos_i(15701) := b"0000000000000000_0000000000000000_0001011101000110_0001101011010000"; -- 0.09091346327310736
	pesos_i(15702) := b"1111111111111111_1111111111111111_1110000110000110_0110111010000011"; -- -0.11904248523497536
	pesos_i(15703) := b"0000000000000000_0000000000000000_0000000000010001_1100100010011100"; -- 0.00027135673335222166
	pesos_i(15704) := b"0000000000000000_0000000000000000_0001010001110100_1110000100100110"; -- 0.07990843933990327
	pesos_i(15705) := b"0000000000000000_0000000000000000_0001000100011100_0010100000111011"; -- 0.06683589408101558
	pesos_i(15706) := b"1111111111111111_1111111111111111_1111011101101101_0100110110110000"; -- -0.033488411387122004
	pesos_i(15707) := b"1111111111111111_1111111111111111_1111011111011001_0100100011101001"; -- -0.031840746960246816
	pesos_i(15708) := b"0000000000000000_0000000000000000_0010010101001110_1000110000100010"; -- 0.1457297881850176
	pesos_i(15709) := b"1111111111111111_1111111111111111_1111010100000111_1110110110000000"; -- -0.042847782431625944
	pesos_i(15710) := b"0000000000000000_0000000000000000_0001011100111111_0000010111010111"; -- 0.09080540183818754
	pesos_i(15711) := b"0000000000000000_0000000000000000_0000000110010011_0101010110110001"; -- 0.006154399704466894
	pesos_i(15712) := b"1111111111111111_1111111111111111_1110001011101111_1001011001011001"; -- -0.11353168795561773
	pesos_i(15713) := b"1111111111111111_1111111111111111_1111101000010110_0011110010010101"; -- -0.02309819565397403
	pesos_i(15714) := b"1111111111111111_1111111111111111_1111001000110100_0000111100110010"; -- -0.053893137318398135
	pesos_i(15715) := b"1111111111111111_1111111111111111_1111001001010110_0000001010011101"; -- -0.05337508832595687
	pesos_i(15716) := b"1111111111111111_1111111111111111_1110101001001000_0100010101010001"; -- -0.08483473559537939
	pesos_i(15717) := b"1111111111111111_1111111111111111_1111110111101111_0010101001000010"; -- -0.008069380715871698
	pesos_i(15718) := b"1111111111111111_1111111111111111_1111000111110001_0101000101001111"; -- -0.05491153552594936
	pesos_i(15719) := b"1111111111111111_1111111111111111_1111100100100011_1100010001011011"; -- -0.02679798857277785
	pesos_i(15720) := b"0000000000000000_0000000000000000_0010001000010111_0001100101111110"; -- 0.13316497156976803
	pesos_i(15721) := b"1111111111111111_1111111111111111_1111100111101111_1111111111001011"; -- -0.023681653067471782
	pesos_i(15722) := b"0000000000000000_0000000000000000_0000100010110100_1101100101010111"; -- 0.03400953644344673
	pesos_i(15723) := b"1111111111111111_1111111111111111_1101100101100101_1100111100000000"; -- -0.15079027408985105
	pesos_i(15724) := b"1111111111111111_1111111111111111_1110101000001110_0100110001100100"; -- -0.08571932377629851
	pesos_i(15725) := b"1111111111111111_1111111111111111_1111110010001001_0110101000001011"; -- -0.013528225241471624
	pesos_i(15726) := b"0000000000000000_0000000000000000_0001110100110101_1000010101101101"; -- 0.1140979187253911
	pesos_i(15727) := b"0000000000000000_0000000000000000_0001110011100110_1000000001110111"; -- 0.11289217856587616
	pesos_i(15728) := b"1111111111111111_1111111111111111_1110101111111100_1001000011101010"; -- -0.07817739757260127
	pesos_i(15729) := b"0000000000000000_0000000000000000_0000100110110110_1101110010010111"; -- 0.037946497859461366
	pesos_i(15730) := b"1111111111111111_1111111111111111_1110100111101101_0010111001011110"; -- -0.08622465322375816
	pesos_i(15731) := b"1111111111111111_1111111111111111_1110000010101111_1101011001111001"; -- -0.1223169282945371
	pesos_i(15732) := b"1111111111111111_1111111111111111_1101110000111111_1011110110011100"; -- -0.1396523947754529
	pesos_i(15733) := b"1111111111111111_1111111111111111_1110110110011111_1110111000010000"; -- -0.07177841294137519
	pesos_i(15734) := b"0000000000000000_0000000000000000_0000011101101100_1101110100100001"; -- 0.02900487941250684
	pesos_i(15735) := b"1111111111111111_1111111111111111_1101110001010111_0111111011011010"; -- -0.13928992429649642
	pesos_i(15736) := b"1111111111111111_1111111111111111_1110010000000101_0011101011010000"; -- -0.10929520063401944
	pesos_i(15737) := b"1111111111111111_1111111111111111_1110011011011100_1011100001010100"; -- -0.0981945795758235
	pesos_i(15738) := b"1111111111111111_1111111111111111_1111000101010110_0010110111111011"; -- -0.05727875350273204
	pesos_i(15739) := b"1111111111111111_1111111111111111_1101111101001111_0010000101011110"; -- -0.1276988167937032
	pesos_i(15740) := b"1111111111111111_1111111111111111_1111110111000011_0111110101110100"; -- -0.008735808573396814
	pesos_i(15741) := b"0000000000000000_0000000000000000_0010010000100010_0001000011101001"; -- 0.1411448067136008
	pesos_i(15742) := b"1111111111111111_1111111111111111_1110000100001000_1110111101110111"; -- -0.12095740638167875
	pesos_i(15743) := b"1111111111111111_1111111111111111_1111000110001011_0000000100100011"; -- -0.056472710475406245
	pesos_i(15744) := b"0000000000000000_0000000000000000_0001000111110110_1101110010110001"; -- 0.07017306635057322
	pesos_i(15745) := b"1111111111111111_1111111111111111_1111100001001010_1111101001010000"; -- -0.030105929826566243
	pesos_i(15746) := b"0000000000000000_0000000000000000_0010110001101000_1110110010101011"; -- 0.1734760206207126
	pesos_i(15747) := b"0000000000000000_0000000000000000_0000011100110010_0010001000011000"; -- 0.028108721707206394
	pesos_i(15748) := b"0000000000000000_0000000000000000_0000100101000011_1100010011000001"; -- 0.03619031635039261
	pesos_i(15749) := b"1111111111111111_1111111111111111_1110111011001100_1010111011010100"; -- -0.06718928652520302
	pesos_i(15750) := b"1111111111111111_1111111111111111_1111000010101101_1110011000010000"; -- -0.0598465166425129
	pesos_i(15751) := b"0000000000000000_0000000000000000_0001111010111011_0101010011101110"; -- 0.1200459558247836
	pesos_i(15752) := b"1111111111111111_1111111111111111_1110100100000000_1010011101001001"; -- -0.08983377908524989
	pesos_i(15753) := b"1111111111111111_1111111111111111_1110001110110010_0110100101100111"; -- -0.11055890315832365
	pesos_i(15754) := b"1111111111111111_1111111111111111_1111110000111100_0110111001110100"; -- -0.014702889119619025
	pesos_i(15755) := b"0000000000000000_0000000000000000_0000111101000100_1100110110001011"; -- 0.05964359897508264
	pesos_i(15756) := b"1111111111111111_1111111111111111_1110100000111110_1001010000111110"; -- -0.09279511919629546
	pesos_i(15757) := b"0000000000000000_0000000000000000_0000110011110011_0101010001111101"; -- 0.0505879215598322
	pesos_i(15758) := b"0000000000000000_0000000000000000_0010001111011111_1100111100001000"; -- 0.1401337998839673
	pesos_i(15759) := b"1111111111111111_1111111111111111_1111001000110010_1101001111100110"; -- -0.05391193042294744
	pesos_i(15760) := b"0000000000000000_0000000000000000_0001011111011001_1000111000001110"; -- 0.09316337429641296
	pesos_i(15761) := b"0000000000000000_0000000000000000_0000101100011100_1011010010111000"; -- 0.043406767877149297
	pesos_i(15762) := b"0000000000000000_0000000000000000_0010010001111101_0110110011110110"; -- 0.142538843137672
	pesos_i(15763) := b"1111111111111111_1111111111111111_1111110000001100_0101001110110001"; -- -0.015436906250515438
	pesos_i(15764) := b"1111111111111111_1111111111111111_1111100101100010_0111000000001001"; -- -0.02584171092685654
	pesos_i(15765) := b"0000000000000000_0000000000000000_0000000100100010_0001110001101001"; -- 0.004426742230031552
	pesos_i(15766) := b"1111111111111111_1111111111111111_1111101010111010_1011111010110100"; -- -0.020587998555664032
	pesos_i(15767) := b"0000000000000000_0000000000000000_0000101101000000_0100100000001011"; -- 0.04394960666384673
	pesos_i(15768) := b"1111111111111111_1111111111111111_1110000101010110_0000010000111001"; -- -0.11978124234950904
	pesos_i(15769) := b"0000000000000000_0000000000000000_0001011111110111_0100101011100010"; -- 0.09361713436632008
	pesos_i(15770) := b"0000000000000000_0000000000000000_0000110010011100_1011001100100100"; -- 0.04926604860698197
	pesos_i(15771) := b"0000000000000000_0000000000000000_0001001010001111_0111000000100010"; -- 0.07250119053360399
	pesos_i(15772) := b"1111111111111111_1111111111111111_1110011010000111_0110100100101101"; -- -0.09949629452993348
	pesos_i(15773) := b"0000000000000000_0000000000000000_0000001010011000_0110111100010011"; -- 0.010138456413010496
	pesos_i(15774) := b"1111111111111111_1111111111111111_1111100000100101_1011001001111101"; -- -0.03067478608284233
	pesos_i(15775) := b"0000000000000000_0000000000000000_0001001110011010_1001011101101001"; -- 0.07657762834060956
	pesos_i(15776) := b"0000000000000000_0000000000000000_0000100011011011_1101011010010001"; -- 0.03460446388488601
	pesos_i(15777) := b"0000000000000000_0000000000000000_0000101110111000_1001011011101011"; -- 0.045785362681264416
	pesos_i(15778) := b"0000000000000000_0000000000000000_0001000100100100_0000001101010101"; -- 0.06695576512296945
	pesos_i(15779) := b"1111111111111111_1111111111111111_1110000001110110_1011010100001101"; -- -0.1231886715170797
	pesos_i(15780) := b"1111111111111111_1111111111111111_1110111000111110_0010111111001110"; -- -0.06936360558495822
	pesos_i(15781) := b"0000000000000000_0000000000000000_0010011011001011_1000111011010101"; -- 0.15154354757155006
	pesos_i(15782) := b"1111111111111111_1111111111111111_1111001110011010_0110101000001111"; -- -0.04842507483387504
	pesos_i(15783) := b"1111111111111111_1111111111111111_1111100110000110_0010001110111100"; -- -0.025296942261083685
	pesos_i(15784) := b"0000000000000000_0000000000000000_0010001111111110_1001001110011000"; -- 0.14060327980371576
	pesos_i(15785) := b"1111111111111111_1111111111111111_1111101101011101_1111010110000001"; -- -0.01809754950692387
	pesos_i(15786) := b"0000000000000000_0000000000000000_0001111001110100_1111001101010111"; -- 0.1189720237755135
	pesos_i(15787) := b"1111111111111111_1111111111111111_1111100011100000_0000110000101011"; -- -0.02783130600902947
	pesos_i(15788) := b"0000000000000000_0000000000000000_0010000100111100_0100111110011010"; -- 0.1298265220716643
	pesos_i(15789) := b"0000000000000000_0000000000000000_0000101110000011_1000010111001011"; -- 0.04497562604792009
	pesos_i(15790) := b"0000000000000000_0000000000000000_0000010100100100_1101110001101100"; -- 0.02009370468249822
	pesos_i(15791) := b"0000000000000000_0000000000000000_0000111101000000_1111011010001011"; -- 0.05958500754149759
	pesos_i(15792) := b"1111111111111111_1111111111111111_1111100000100011_0111010001111111"; -- -0.030708998600820128
	pesos_i(15793) := b"0000000000000000_0000000000000000_0000100000000011_0000101111100000"; -- 0.031296484077487606
	pesos_i(15794) := b"1111111111111111_1111111111111111_1110110110111101_1111011100100110"; -- -0.07132010762698211
	pesos_i(15795) := b"1111111111111111_1111111111111111_1111110000001101_1110011010101011"; -- -0.015412886866192405
	pesos_i(15796) := b"1111111111111111_1111111111111111_1110111011010101_0110000000011000"; -- -0.06705665020749005
	pesos_i(15797) := b"0000000000000000_0000000000000000_0000000100000100_1111100101000111"; -- 0.003982143355265321
	pesos_i(15798) := b"1111111111111111_1111111111111111_1111110010100111_1001010111101111"; -- -0.013067845552289232
	pesos_i(15799) := b"0000000000000000_0000000000000000_0000011011111101_0011010001100001"; -- 0.027301095619574393
	pesos_i(15800) := b"1111111111111111_1111111111111111_1110110010001111_0101011111011101"; -- -0.0759377560089468
	pesos_i(15801) := b"0000000000000000_0000000000000000_0001010110011100_1101001010011011"; -- 0.0844241742521834
	pesos_i(15802) := b"0000000000000000_0000000000000000_0001010111001111_1110110101011000"; -- 0.08520396611866153
	pesos_i(15803) := b"1111111111111111_1111111111111111_1111010110110011_0010010101001000"; -- -0.04023520469285672
	pesos_i(15804) := b"1111111111111111_1111111111111111_1110000111001111_0100000000110000"; -- -0.11793135485738836
	pesos_i(15805) := b"1111111111111111_1111111111111111_1110000010101110_1001111000011000"; -- -0.12233554760740857
	pesos_i(15806) := b"0000000000000000_0000000000000000_0000001101010101_1010111111111001"; -- 0.013026235953834075
	pesos_i(15807) := b"0000000000000000_0000000000000000_0001000001110110_0000101011010111"; -- 0.06430118320797133
	pesos_i(15808) := b"1111111111111111_1111111111111111_1110000110010010_0000110111110101"; -- -0.11886513496412324
	pesos_i(15809) := b"0000000000000000_0000000000000000_0001111000111011_1101011100011010"; -- 0.11810058950707497
	pesos_i(15810) := b"0000000000000000_0000000000000000_0000111001100100_1101100111100000"; -- 0.05622636525452945
	pesos_i(15811) := b"0000000000000000_0000000000000000_0010000011001001_0111101000100010"; -- 0.1280742961904068
	pesos_i(15812) := b"1111111111111111_1111111111111111_1111011111011101_1111110001110110"; -- -0.03176900986244448
	pesos_i(15813) := b"1111111111111111_1111111111111111_1111100010111011_1000110010111100"; -- -0.028388218103666214
	pesos_i(15814) := b"0000000000000000_0000000000000000_0001100010001000_1100100011101101"; -- 0.0958371713693721
	pesos_i(15815) := b"0000000000000000_0000000000000000_0000100001100101_1100001110010100"; -- 0.03280279502389527
	pesos_i(15816) := b"0000000000000000_0000000000000000_0001110001000011_1100011101101111"; -- 0.11040922593817051
	pesos_i(15817) := b"0000000000000000_0000000000000000_0001011011000011_1100010010010011"; -- 0.08892468066112974
	pesos_i(15818) := b"1111111111111111_1111111111111111_1111110100001101_0001111111100101"; -- -0.01151848478922661
	pesos_i(15819) := b"0000000000000000_0000000000000000_0001111010001000_0001011001110010"; -- 0.11926403324093517
	pesos_i(15820) := b"1111111111111111_1111111111111111_1110001111011100_0100100001100100"; -- -0.10992000149603748
	pesos_i(15821) := b"0000000000000000_0000000000000000_0000011000001111_0000110000010111"; -- 0.023667102549087257
	pesos_i(15822) := b"0000000000000000_0000000000000000_0010001001111011_0111100000010100"; -- 0.13469648833825612
	pesos_i(15823) := b"1111111111111111_1111111111111111_1110000001111100_1011010110111111"; -- -0.1230970771919814
	pesos_i(15824) := b"0000000000000000_0000000000000000_0001111101010100_0111011110000001"; -- 0.12238261125722279
	pesos_i(15825) := b"1111111111111111_1111111111111111_1111110010011011_1100111101100010"; -- -0.013247526749726263
	pesos_i(15826) := b"1111111111111111_1111111111111111_1110001011011001_0001111110101010"; -- -0.11387445544383022
	pesos_i(15827) := b"1111111111111111_1111111111111111_1101010011110001_1101000010100011"; -- -0.16818519615563754
	pesos_i(15828) := b"0000000000000000_0000000000000000_0000011100100101_0001001101001100"; -- 0.02790947536064249
	pesos_i(15829) := b"0000000000000000_0000000000000000_0001010001100000_1110101111001101"; -- 0.07960389845565102
	pesos_i(15830) := b"1111111111111111_1111111111111111_1110101010100010_1110010001010011"; -- -0.0834519669531359
	pesos_i(15831) := b"0000000000000000_0000000000000000_0001001110000100_1100110001011101"; -- 0.07624509111225519
	pesos_i(15832) := b"1111111111111111_1111111111111111_1111101011011110_0010111111010000"; -- -0.020047198992953125
	pesos_i(15833) := b"1111111111111111_1111111111111111_1111011001010010_1110101010110110"; -- -0.03779728954792086
	pesos_i(15834) := b"0000000000000000_0000000000000000_0001010101100111_0001101010011011"; -- 0.08360449112801734
	pesos_i(15835) := b"1111111111111111_1111111111111111_1111110010100111_1100001100110101"; -- -0.013065146991761756
	pesos_i(15836) := b"1111111111111111_1111111111111111_1110000111010111_1001101000101000"; -- -0.11780392195097819
	pesos_i(15837) := b"1111111111111111_1111111111111111_1110010000111000_1011110101011000"; -- -0.1085092219384428
	pesos_i(15838) := b"1111111111111111_1111111111111111_1110000010011001_1110111100111001"; -- -0.12265114651898786
	pesos_i(15839) := b"0000000000000000_0000000000000000_0000100100110101_0011011111011011"; -- 0.035968295089931435
	pesos_i(15840) := b"0000000000000000_0000000000000000_0000010101110011_1000110100000010"; -- 0.02129441536679341
	pesos_i(15841) := b"1111111111111111_1111111111111111_1110110110100101_0111011111100101"; -- -0.07169390362504775
	pesos_i(15842) := b"1111111111111111_1111111111111111_1110100001000001_1011001001010110"; -- -0.09274754911471973
	pesos_i(15843) := b"1111111111111111_1111111111111111_1110100001100110_0011001100111010"; -- -0.092190550166493
	pesos_i(15844) := b"0000000000000000_0000000000000000_0000000001110100_1000111000111000"; -- 0.0017784964911983427
	pesos_i(15845) := b"1111111111111111_1111111111111111_1101111100000010_1110001011001011"; -- -0.12886221442587753
	pesos_i(15846) := b"0000000000000000_0000000000000000_0010101010010111_0001110110010111"; -- 0.166368340793469
	pesos_i(15847) := b"0000000000000000_0000000000000000_0000111111101010_0011101111001000"; -- 0.06216786983306981
	pesos_i(15848) := b"1111111111111111_1111111111111111_1101110001000011_0000111100011010"; -- -0.13960176109509492
	pesos_i(15849) := b"0000000000000000_0000000000000000_0001101111110011_0101011011110010"; -- 0.10918181815297398
	pesos_i(15850) := b"0000000000000000_0000000000000000_0001111010001010_0000101011110010"; -- 0.11929386530703144
	pesos_i(15851) := b"0000000000000000_0000000000000000_0000010111000010_1100000000101101"; -- 0.022502909539972075
	pesos_i(15852) := b"0000000000000000_0000000000000000_0001011110100110_1100101110101010"; -- 0.092388848269023
	pesos_i(15853) := b"1111111111111111_1111111111111111_1101110010100010_0011101010100000"; -- -0.1381495819435529
	pesos_i(15854) := b"1111111111111111_1111111111111111_1111110001010001_0110011010000011"; -- -0.014382927923668581
	pesos_i(15855) := b"0000000000000000_0000000000000000_0001110100001010_0010000001110000"; -- 0.11343577132684474
	pesos_i(15856) := b"1111111111111111_1111111111111111_1110000000000111_1010001100100000"; -- -0.12488346555237072
	pesos_i(15857) := b"1111111111111111_1111111111111111_1110000001001010_1111111001110010"; -- -0.12385568337256495
	pesos_i(15858) := b"1111111111111111_1111111111111111_1111101111110000_1111010010010000"; -- -0.01585456363188115
	pesos_i(15859) := b"0000000000000000_0000000000000000_0000010101011101_1010010011010101"; -- 0.02096014206003576
	pesos_i(15860) := b"0000000000000000_0000000000000000_0000110111101000_1001111010001110"; -- 0.05433073962635417
	pesos_i(15861) := b"0000000000000000_0000000000000000_0010110000011111_0001101101000000"; -- 0.17234964673548625
	pesos_i(15862) := b"0000000000000000_0000000000000000_0001100101011000_0100100001111100"; -- 0.09900334374715257
	pesos_i(15863) := b"1111111111111111_1111111111111111_1110100011001011_0101111100000001"; -- -0.09064680324157037
	pesos_i(15864) := b"1111111111111111_1111111111111111_1101101000100001_0110101000000101"; -- -0.1479276407913947
	pesos_i(15865) := b"1111111111111111_1111111111111111_1101101111111100_1011001010011001"; -- -0.14067538994706436
	pesos_i(15866) := b"1111111111111111_1111111111111111_1111011010000011_1100111101100011"; -- -0.03705123741866127
	pesos_i(15867) := b"0000000000000000_0000000000000000_0010000100101001_0000011111100111"; -- 0.12953233136687398
	pesos_i(15868) := b"0000000000000000_0000000000000000_0000011000000010_0100011011101001"; -- 0.023472244140051564
	pesos_i(15869) := b"0000000000000000_0000000000000000_0010001110111110_1010011100100101"; -- 0.13962788254812603
	pesos_i(15870) := b"1111111111111111_1111111111111111_1110001001010010_1010000101011000"; -- -0.1159266623832612
	pesos_i(15871) := b"1111111111111111_1111111111111111_1110101101101101_1010001101001000"; -- -0.08035830958397797
	pesos_i(15872) := b"1111111111111111_1111111111111111_1101111000101100_1001100011110011"; -- -0.13213199676039442
	pesos_i(15873) := b"1111111111111111_1111111111111111_1111110111010111_0010111000011101"; -- -0.00843536176840339
	pesos_i(15874) := b"0000000000000000_0000000000000000_0010110011000110_1010011011000010"; -- 0.17490617975694817
	pesos_i(15875) := b"0000000000000000_0000000000000000_0000111000101101_1111001011000000"; -- 0.055388614526883394
	pesos_i(15876) := b"0000000000000000_0000000000000000_0001010011010011_0111110110100010"; -- 0.0813520928780076
	pesos_i(15877) := b"0000000000000000_0000000000000000_0001101111111001_0000110101001100"; -- 0.10926898103168442
	pesos_i(15878) := b"1111111111111111_1111111111111111_1111000000110111_0011001100011000"; -- -0.06165772119041596
	pesos_i(15879) := b"1111111111111111_1111111111111111_1111010100101011_0100000100100000"; -- -0.04230874024483804
	pesos_i(15880) := b"1111111111111111_1111111111111111_1110011000111101_0001101100100011"; -- -0.10063009638934914
	pesos_i(15881) := b"1111111111111111_1111111111111111_1110001101011101_0001111000011000"; -- -0.11186038886446593
	pesos_i(15882) := b"0000000000000000_0000000000000000_0000010000001100_0011100001011100"; -- 0.01581146485098663
	pesos_i(15883) := b"1111111111111111_1111111111111111_1110101001111011_1001001101110111"; -- -0.0840518793260301
	pesos_i(15884) := b"1111111111111111_1111111111111111_1110110110001100_0010001111111101"; -- -0.07208037448565173
	pesos_i(15885) := b"0000000000000000_0000000000000000_0010011100001010_0000110001101010"; -- 0.15249707779324803
	pesos_i(15886) := b"0000000000000000_0000000000000000_0010011001011100_1100101011110100"; -- 0.14985340548699563
	pesos_i(15887) := b"0000000000000000_0000000000000000_0001111001101001_1100000001111000"; -- 0.11880114477276875
	pesos_i(15888) := b"0000000000000000_0000000000000000_0001010001011000_1101100110110010"; -- 0.0794807490031473
	pesos_i(15889) := b"1111111111111111_1111111111111111_1110000000000101_1111110001101001"; -- -0.12490866113082391
	pesos_i(15890) := b"0000000000000000_0000000000000000_0010101010101110_1101000001100110"; -- 0.1667299508688062
	pesos_i(15891) := b"1111111111111111_1111111111111111_1110001011000111_1000001110001001"; -- -0.11414316097422775
	pesos_i(15892) := b"1111111111111111_1111111111111111_1110000100101000_1110111000110111"; -- -0.12046919982678973
	pesos_i(15893) := b"1111111111111111_1111111111111111_1110001011100010_1010010001100101"; -- -0.11372921509184168
	pesos_i(15894) := b"1111111111111111_1111111111111111_1111010100000110_0100001101011100"; -- -0.04287318244063877
	pesos_i(15895) := b"1111111111111111_1111111111111111_1101111011110101_1101011010010101"; -- -0.12906130654133588
	pesos_i(15896) := b"0000000000000000_0000000000000000_0000011010100101_1001110000001010"; -- 0.025964500932056326
	pesos_i(15897) := b"1111111111111111_1111111111111111_1110011011000011_0111100100101000"; -- -0.09857981467431298
	pesos_i(15898) := b"0000000000000000_0000000000000000_0000111000110000_1011011111100101"; -- 0.05543088289138413
	pesos_i(15899) := b"1111111111111111_1111111111111111_1111111101101011_1010100011110001"; -- -0.002263489958501805
	pesos_i(15900) := b"1111111111111111_1111111111111111_1101101111010011_1011001111001001"; -- -0.14130092946870176
	pesos_i(15901) := b"1111111111111111_1111111111111111_1101111110000101_1000111100110011"; -- -0.1268682956733031
	pesos_i(15902) := b"1111111111111111_1111111111111111_1110010000100010_1010100000011110"; -- -0.10884618067116839
	pesos_i(15903) := b"1111111111111111_1111111111111111_1111110100010100_1101111011011101"; -- -0.011400290602973115
	pesos_i(15904) := b"1111111111111111_1111111111111111_1111001011011011_1101110000010000"; -- -0.05133270854541833
	pesos_i(15905) := b"0000000000000000_0000000000000000_0000111001011110_0101111010010100"; -- 0.056127463499628036
	pesos_i(15906) := b"1111111111111111_1111111111111111_1110100010111000_0000011100101110"; -- -0.09094195487796725
	pesos_i(15907) := b"1111111111111111_1111111111111111_1111111011011110_1001011001011001"; -- -0.004416087507698645
	pesos_i(15908) := b"1111111111111111_1111111111111111_1110011000110111_0011011001000110"; -- -0.10072003160551858
	pesos_i(15909) := b"0000000000000000_0000000000000000_0000000101110101_0111100001101110"; -- 0.005698706445075492
	pesos_i(15910) := b"0000000000000000_0000000000000000_0000100111010110_1001101110100011"; -- 0.03843090748939078
	pesos_i(15911) := b"0000000000000000_0000000000000000_0000011010010001_1101001100110110"; -- 0.025662613682920738
	pesos_i(15912) := b"1111111111111111_1111111111111111_1110110110101100_1000000111101000"; -- -0.07158649517327435
	pesos_i(15913) := b"0000000000000000_0000000000000000_0000110001110011_0110101111000111"; -- 0.048636184833840794
	pesos_i(15914) := b"1111111111111111_1111111111111111_1110110101010000_0101010110010010"; -- -0.07299294640764817
	pesos_i(15915) := b"0000000000000000_0000000000000000_0000001001001100_0111111101001000"; -- 0.00897975456254145
	pesos_i(15916) := b"1111111111111111_1111111111111111_1110100011110110_1010111011111001"; -- -0.08998590875372996
	pesos_i(15917) := b"1111111111111111_1111111111111111_1110101101010110_1001000010001001"; -- -0.0807103792687704
	pesos_i(15918) := b"0000000000000000_0000000000000000_0000010010011101_1101110100110001"; -- 0.018033813897126112
	pesos_i(15919) := b"0000000000000000_0000000000000000_0010100111010000_1101000110111100"; -- 0.16334257915635803
	pesos_i(15920) := b"0000000000000000_0000000000000000_0001111000011101_1000001111111011"; -- 0.11763787147510439
	pesos_i(15921) := b"0000000000000000_0000000000000000_0001110001000110_1010001000110000"; -- 0.11045278224952812
	pesos_i(15922) := b"1111111111111111_1111111111111111_1110011011000100_1011100101011101"; -- -0.0985607287164079
	pesos_i(15923) := b"1111111111111111_1111111111111111_1101110001111011_1111100100100011"; -- -0.13873331928401503
	pesos_i(15924) := b"1111111111111111_1111111111111111_1110010000010110_0000011101010110"; -- -0.10903886938757214
	pesos_i(15925) := b"0000000000000000_0000000000000000_0000100011011010_0000011110111111"; -- 0.03457687780439111
	pesos_i(15926) := b"0000000000000000_0000000000000000_0010000010110111_1001011101111010"; -- 0.12780138706853794
	pesos_i(15927) := b"1111111111111111_1111111111111111_1101110011110000_1001111101010111"; -- -0.13695339333700082
	pesos_i(15928) := b"1111111111111111_1111111111111111_1111110000010010_0100111101111100"; -- -0.015345604195908307
	pesos_i(15929) := b"0000000000000000_0000000000000000_0010010101000000_1000010001101010"; -- 0.14551570509696912
	pesos_i(15930) := b"1111111111111111_1111111111111111_1111001110011000_0101110101010111"; -- -0.04845635059492579
	pesos_i(15931) := b"0000000000000000_0000000000000000_0001010010001110_1001001101111000"; -- 0.08030053777608108
	pesos_i(15932) := b"1111111111111111_1111111111111111_1110001101101110_1011011110111010"; -- -0.11159183221291982
	pesos_i(15933) := b"0000000000000000_0000000000000000_0001011101001011_0000101101011011"; -- 0.09098883611598349
	pesos_i(15934) := b"1111111111111111_1111111111111111_1101111001100001_1110010010000111"; -- -0.13131877614291113
	pesos_i(15935) := b"1111111111111111_1111111111111111_1111010011011010_0010010000110101"; -- -0.04354642593273099
	pesos_i(15936) := b"1111111111111111_1111111111111111_1111111011011100_0110100011101001"; -- -0.004449313327212487
	pesos_i(15937) := b"1111111111111111_1111111111111111_1111110000100000_1001110111100010"; -- -0.015127308211167836
	pesos_i(15938) := b"1111111111111111_1111111111111111_1111111010001001_0001110011000010"; -- -0.005720331717621798
	pesos_i(15939) := b"0000000000000000_0000000000000000_0000111100111010_1110111000010000"; -- 0.059492949292357065
	pesos_i(15940) := b"0000000000000000_0000000000000000_0000000100011000_1011101000011000"; -- 0.004283553046238796
	pesos_i(15941) := b"0000000000000000_0000000000000000_0000000100110101_0000100010110111"; -- 0.004715485303001428
	pesos_i(15942) := b"0000000000000000_0000000000000000_0001011101011110_1000110010110111"; -- 0.0912864633618231
	pesos_i(15943) := b"0000000000000000_0000000000000000_0001000010010001_1110111101101000"; -- 0.06472679421631256
	pesos_i(15944) := b"1111111111111111_1111111111111111_1110110111000011_0011001110001100"; -- -0.07124021364756031
	pesos_i(15945) := b"0000000000000000_0000000000000000_0000111100100110_1000010100110101"; -- 0.059181523682624866
	pesos_i(15946) := b"0000000000000000_0000000000000000_0010101100110101_1001110100010110"; -- 0.16878682890445781
	pesos_i(15947) := b"1111111111111111_1111111111111111_1101110111001100_1001010100101001"; -- -0.13359706632354035
	pesos_i(15948) := b"1111111111111111_1111111111111111_1110100110001010_0011110110011100"; -- -0.08773436486603983
	pesos_i(15949) := b"1111111111111111_1111111111111111_1101101011100001_1110100010110111"; -- -0.14499040154711845
	pesos_i(15950) := b"1111111111111111_1111111111111111_1110100110000000_0100011010101011"; -- -0.0878864127530228
	pesos_i(15951) := b"0000000000000000_0000000000000000_0000011101011000_0101101000001010"; -- 0.0286918900992865
	pesos_i(15952) := b"0000000000000000_0000000000000000_0010000010000011_1101111101011111"; -- 0.12701221532957307
	pesos_i(15953) := b"1111111111111111_1111111111111111_1110111010010100_1110001110001101"; -- -0.06804063623738371
	pesos_i(15954) := b"0000000000000000_0000000000000000_0001000101001110_1000111001101000"; -- 0.06760492369042317
	pesos_i(15955) := b"1111111111111111_1111111111111111_1110010001000101_0110000011100000"; -- -0.10831636936912208
	pesos_i(15956) := b"1111111111111111_1111111111111111_1111000000110101_1100101110011001"; -- -0.061679148738034505
	pesos_i(15957) := b"0000000000000000_0000000000000000_0000101010111101_0101100100001010"; -- 0.04195171829563081
	pesos_i(15958) := b"0000000000000000_0000000000000000_0000110100001011_1001110000111010"; -- 0.05095840848619743
	pesos_i(15959) := b"1111111111111111_1111111111111111_1111111011100100_0011100001000010"; -- -0.004330142858006185
	pesos_i(15960) := b"1111111111111111_1111111111111111_1110100111110101_0110010011101101"; -- -0.08609933109858586
	pesos_i(15961) := b"0000000000000000_0000000000000000_0000101011010111_1100111100101000"; -- 0.04235548714706392
	pesos_i(15962) := b"0000000000000000_0000000000000000_0010000000101111_1110001001101110"; -- 0.12573065938676417
	pesos_i(15963) := b"0000000000000000_0000000000000000_0000001100101111_0100001010100100"; -- 0.012439885105860938
	pesos_i(15964) := b"1111111111111111_1111111111111111_1111111011001011_1100000001010000"; -- -0.004703503002506545
	pesos_i(15965) := b"0000000000000000_0000000000000000_0000011011000100_1001001011010010"; -- 0.02643697376042538
	pesos_i(15966) := b"0000000000000000_0000000000000000_0010000110000010_0001001111011110"; -- 0.1308910767343391
	pesos_i(15967) := b"1111111111111111_1111111111111111_1110010110110011_0000010001110010"; -- -0.10273716181926872
	pesos_i(15968) := b"1111111111111111_1111111111111111_1111011111001111_1110001100110110"; -- -0.03198413788411644
	pesos_i(15969) := b"1111111111111111_1111111111111111_1101111110100000_1111100000100110"; -- -0.1264500528403091
	pesos_i(15970) := b"0000000000000000_0000000000000000_0001001001111010_0101001101101011"; -- 0.07217904425273987
	pesos_i(15971) := b"1111111111111111_1111111111111111_1111001111010010_1001010000111101"; -- -0.04756806858436572
	pesos_i(15972) := b"0000000000000000_0000000000000000_0010000000011010_1010111100101011"; -- 0.12540716924389342
	pesos_i(15973) := b"0000000000000000_0000000000000000_0000110101010101_0111100010110001"; -- 0.05208544091728327
	pesos_i(15974) := b"1111111111111111_1111111111111111_1110010110011001_0001101001110111"; -- -0.10313257790322884
	pesos_i(15975) := b"1111111111111111_1111111111111111_1110101000000010_1111000111110010"; -- -0.08589256125106444
	pesos_i(15976) := b"0000000000000000_0000000000000000_0001100011101111_1101011100000011"; -- 0.09740966624871066
	pesos_i(15977) := b"0000000000000000_0000000000000000_0001100111010001_0000110001101100"; -- 0.10084607736609573
	pesos_i(15978) := b"1111111111111111_1111111111111111_1101110110001111_1101011100001100"; -- -0.13452392536384133
	pesos_i(15979) := b"1111111111111111_1111111111111111_1110101001010010_0001101000110000"; -- -0.08468471841421614
	pesos_i(15980) := b"0000000000000000_0000000000000000_0001101000100011_0110101011010010"; -- 0.10210292457753754
	pesos_i(15981) := b"1111111111111111_1111111111111111_1111101111010111_1001101010010010"; -- -0.016241397251255108
	pesos_i(15982) := b"1111111111111111_1111111111111111_1111110100001000_1111001111101000"; -- -0.01158214173433405
	pesos_i(15983) := b"0000000000000000_0000000000000000_0001111010001010_1011000101100110"; -- 0.11930378675341556
	pesos_i(15984) := b"1111111111111111_1111111111111111_1111100101111000_0001110010111100"; -- -0.025510982589881572
	pesos_i(15985) := b"0000000000000000_0000000000000000_0001011001110010_0110101000100000"; -- 0.08768332755369926
	pesos_i(15986) := b"0000000000000000_0000000000000000_0010001001011010_0110000100110110"; -- 0.13419158531559816
	pesos_i(15987) := b"0000000000000000_0000000000000000_0000011000011010_0000110100100001"; -- 0.023835011101410012
	pesos_i(15988) := b"0000000000000000_0000000000000000_0001000000000110_1100000010111111"; -- 0.0626030412763702
	pesos_i(15989) := b"1111111111111111_1111111111111111_1111100101101111_0010000011110111"; -- -0.025648059613346753
	pesos_i(15990) := b"0000000000000000_0000000000000000_0000111101111000_1110110011110101"; -- 0.060438928377619903
	pesos_i(15991) := b"1111111111111111_1111111111111111_1111010111101011_1111000000100001"; -- -0.039368621726767805
	pesos_i(15992) := b"1111111111111111_1111111111111111_1111010010001001_0001101110101000"; -- -0.04478289736563715
	pesos_i(15993) := b"0000000000000000_0000000000000000_0000101110100100_0111011010111001"; -- 0.045478267918524745
	pesos_i(15994) := b"0000000000000000_0000000000000000_0000111110000010_0001001000110000"; -- 0.06057847673329904
	pesos_i(15995) := b"1111111111111111_1111111111111111_1110001110111111_0011100100101000"; -- -0.11036341450889793
	pesos_i(15996) := b"0000000000000000_0000000000000000_0001011000110010_1001110111110001"; -- 0.08670985356102072
	pesos_i(15997) := b"0000000000000000_0000000000000000_0000000110010101_0101111101110001"; -- 0.006185498261955568
	pesos_i(15998) := b"1111111111111111_1111111111111111_1111111101100000_1010011110100010"; -- -0.0024314144494713636
	pesos_i(15999) := b"1111111111111111_1111111111111111_1110001010011010_1100111010110011"; -- -0.1148253261890759
	pesos_i(16000) := b"1111111111111111_1111111111111111_1111100101011101_1011000010001111"; -- -0.025914158877943273
	pesos_i(16001) := b"1111111111111111_1111111111111111_1110010111101110_1111110101011110"; -- -0.10182205629208037
	pesos_i(16002) := b"0000000000000000_0000000000000000_0010111001111110_1100000011101000"; -- 0.18162160554284384
	pesos_i(16003) := b"0000000000000000_0000000000000000_0001001000000101_0010010110010010"; -- 0.07039103325599749
	pesos_i(16004) := b"1111111111111111_1111111111111111_1101110011000110_1110000010101101"; -- -0.13759036806060967
	pesos_i(16005) := b"0000000000000000_0000000000000000_0000110100010101_1000101010101100"; -- 0.05110994996771928
	pesos_i(16006) := b"1111111111111111_1111111111111111_1111010010001011_0000000111110110"; -- -0.04475391152871983
	pesos_i(16007) := b"1111111111111111_1111111111111111_1111101110111101_1101110001101100"; -- -0.01663420065546847
	pesos_i(16008) := b"0000000000000000_0000000000000000_0000100110001111_0010010010100011"; -- 0.037340440500266234
	pesos_i(16009) := b"0000000000000000_0000000000000000_0010010110110001_0100010011001011"; -- 0.1472361559712018
	pesos_i(16010) := b"0000000000000000_0000000000000000_0010011001011010_0001001111000111"; -- 0.14981196988300088
	pesos_i(16011) := b"1111111111111111_1111111111111111_1111010110101111_0011000001011011"; -- -0.04029557971999987
	pesos_i(16012) := b"0000000000000000_0000000000000000_0000011110010000_0001000111001010"; -- 0.029542076028868543
	pesos_i(16013) := b"1111111111111111_1111111111111111_1111101000101101_1110010011100010"; -- -0.02273721210867721
	pesos_i(16014) := b"1111111111111111_1111111111111111_1110110000001010_0100011010010001"; -- -0.07796820591161699
	pesos_i(16015) := b"1111111111111111_1111111111111111_1111111111000111_1010111110101010"; -- -0.0008592806190859654
	pesos_i(16016) := b"0000000000000000_0000000000000000_0001100100000111_0110011010010100"; -- 0.09776917567439233
	pesos_i(16017) := b"0000000000000000_0000000000000000_0000010110101010_1001001100111010"; -- 0.022134019479556375
	pesos_i(16018) := b"1111111111111111_1111111111111111_1111111011110101_0100101011011001"; -- -0.004069635464049725
	pesos_i(16019) := b"0000000000000000_0000000000000000_0001010111110111_0101000000011101"; -- 0.08580494602870119
	pesos_i(16020) := b"1111111111111111_1111111111111111_1110001110110111_0101101010100000"; -- -0.11048349001394608
	pesos_i(16021) := b"1111111111111111_1111111111111111_1111110001101011_1001101000010100"; -- -0.013983125736842456
	pesos_i(16022) := b"1111111111111111_1111111111111111_1111001010111110_0101100000111000"; -- -0.05178307176567389
	pesos_i(16023) := b"1111111111111111_1111111111111111_1111101000110101_0001110101111101"; -- -0.022627026548407172
	pesos_i(16024) := b"0000000000000000_0000000000000000_0001110111010000_1110011011111111"; -- 0.11646884665528427
	pesos_i(16025) := b"0000000000000000_0000000000000000_0000010000011011_1101000101110110"; -- 0.016049472099271992
	pesos_i(16026) := b"1111111111111111_1111111111111111_1110010101010100_0111110011001011"; -- -0.10417957350456657
	pesos_i(16027) := b"1111111111111111_1111111111111111_1101101000010010_1011101001010000"; -- -0.1481517366986948
	pesos_i(16028) := b"0000000000000000_0000000000000000_0000001110001000_0000011011010111"; -- 0.01379435297152064
	pesos_i(16029) := b"1111111111111111_1111111111111111_1110001011010101_0011101100001011"; -- -0.11393385871374959
	pesos_i(16030) := b"1111111111111111_1111111111111111_1111000100110011_0101100000110100"; -- -0.05781029442859459
	pesos_i(16031) := b"1111111111111111_1111111111111111_1110001001001111_0000000001101000"; -- -0.11598203156239058
	pesos_i(16032) := b"1111111111111111_1111111111111111_1111000001011100_0101000010011101"; -- -0.06109138658482336
	pesos_i(16033) := b"0000000000000000_0000000000000000_0001010101100111_0111101010010100"; -- 0.08361021143662362
	pesos_i(16034) := b"0000000000000000_0000000000000000_0001010111001000_0110101000011110"; -- 0.08508933284375043
	pesos_i(16035) := b"0000000000000000_0000000000000000_0001110110111110_0001101010110111"; -- 0.11618201216622807
	pesos_i(16036) := b"1111111111111111_1111111111111111_1111010100111101_0111000100110001"; -- -0.04203121715329076
	pesos_i(16037) := b"1111111111111111_1111111111111111_1110010100101111_0000100010111100"; -- -0.10475106637873854
	pesos_i(16038) := b"1111111111111111_1111111111111111_1101101100110110_0110101000010010"; -- -0.14370095303029642
	pesos_i(16039) := b"1111111111111111_1111111111111111_1110010101011010_0101100010010111"; -- -0.10409017851035446
	pesos_i(16040) := b"1111111111111111_1111111111111111_1111111010100111_1001111110100010"; -- -0.005254767318616789
	pesos_i(16041) := b"0000000000000000_0000000000000000_0001110000000000_1010111110110111"; -- 0.10938547345041853
	pesos_i(16042) := b"1111111111111111_1111111111111111_1111111100011111_0111010000001111"; -- -0.0034263100060671035
	pesos_i(16043) := b"1111111111111111_1111111111111111_1101011111000100_1101000110110110"; -- -0.15715302752224428
	pesos_i(16044) := b"1111111111111111_1111111111111111_1110000000000000_0111110110010010"; -- -0.12499251535688655
	pesos_i(16045) := b"1111111111111111_1111111111111111_1111100011001010_0000111110000000"; -- -0.0281668006815624
	pesos_i(16046) := b"0000000000000000_0000000000000000_0001011001011100_0010100100011101"; -- 0.08734375913190583
	pesos_i(16047) := b"1111111111111111_1111111111111111_1111101001010000_0110100010101100"; -- -0.022210557956001877
	pesos_i(16048) := b"1111111111111111_1111111111111111_1111111011000000_1000011010001001"; -- -0.004874793591864758
	pesos_i(16049) := b"1111111111111111_1111111111111111_1110110100100100_1000010001010100"; -- -0.07366154628260947
	pesos_i(16050) := b"0000000000000000_0000000000000000_0001000111011001_0101100110000000"; -- 0.069722741922141
	pesos_i(16051) := b"0000000000000000_0000000000000000_0001100101010111_1000011000101011"; -- 0.09899176175922823
	pesos_i(16052) := b"1111111111111111_1111111111111111_1101101011111001_0011010110011100"; -- -0.14463486605993553
	pesos_i(16053) := b"1111111111111111_1111111111111111_1111001011101101_1100000100000001"; -- -0.05105966299001762
	pesos_i(16054) := b"1111111111111111_1111111111111111_1111110010110011_0101100110100100"; -- -0.012888333745826189
	pesos_i(16055) := b"1111111111111111_1111111111111111_1111111110001100_1011001011011100"; -- -0.0017593586882055274
	pesos_i(16056) := b"0000000000000000_0000000000000000_0010000011101010_0101111100111100"; -- 0.12857623305436466
	pesos_i(16057) := b"0000000000000000_0000000000000000_0001101110110010_0000000010000101"; -- 0.10818484547924938
	pesos_i(16058) := b"0000000000000000_0000000000000000_0000110011101000_1101001100001011"; -- 0.0504276181025442
	pesos_i(16059) := b"1111111111111111_1111111111111111_1110000100101000_1110100000000001"; -- -0.12046956983132573
	pesos_i(16060) := b"0000000000000000_0000000000000000_0001110100111110_1001101111010100"; -- 0.11423658294931105
	pesos_i(16061) := b"0000000000000000_0000000000000000_0000001011001111_1111001001001100"; -- 0.010985511344926504
	pesos_i(16062) := b"1111111111111111_1111111111111111_1110101010000101_0110000010111111"; -- -0.08390231458444429
	pesos_i(16063) := b"1111111111111111_1111111111111111_1101110101110101_1011100110101011"; -- -0.1349224049690937
	pesos_i(16064) := b"1111111111111111_1111111111111111_1110001011101011_1101111100101110"; -- -0.11358838200646469
	pesos_i(16065) := b"1111111111111111_1111111111111111_1110110111000110_0110000100010011"; -- -0.07119172357798978
	pesos_i(16066) := b"1111111111111111_1111111111111111_1111101001000101_1000001001100010"; -- -0.022376872239817585
	pesos_i(16067) := b"1111111111111111_1111111111111111_1110001101000101_1011000001010101"; -- -0.1122178833167098
	pesos_i(16068) := b"0000000000000000_0000000000000000_0000110001100100_0011100101100110"; -- 0.048404300175886775
	pesos_i(16069) := b"1111111111111111_1111111111111111_1111011011010001_1010100110111011"; -- -0.03586329625702176
	pesos_i(16070) := b"1111111111111111_1111111111111111_1101111100000100_1010001101111000"; -- -0.12883547128608092
	pesos_i(16071) := b"0000000000000000_0000000000000000_0010000010010001_1111111000000101"; -- 0.1272276650541761
	pesos_i(16072) := b"1111111111111111_1111111111111111_1101111101010011_1011100011001000"; -- -0.12762875668505286
	pesos_i(16073) := b"1111111111111111_1111111111111111_1111100010001010_0010101011010110"; -- -0.02914173380530087
	pesos_i(16074) := b"0000000000000000_0000000000000000_0010101001111011_1011101010111111"; -- 0.16595046196365348
	pesos_i(16075) := b"1111111111111111_1111111111111111_1110010101101101_0101110111010010"; -- -0.10379994986301042
	pesos_i(16076) := b"0000000000000000_0000000000000000_0001110100000111_1011000001000100"; -- 0.11339856777910778
	pesos_i(16077) := b"0000000000000000_0000000000000000_0001110010101111_1010111100110111"; -- 0.11205573168585334
	pesos_i(16078) := b"1111111111111111_1111111111111111_1110001000011100_1001101110001010"; -- -0.11675098314345791
	pesos_i(16079) := b"1111111111111111_1111111111111111_1110110110101100_1100111110110111"; -- -0.07158185748875687
	pesos_i(16080) := b"0000000000000000_0000000000000000_0000110110101000_0110100100110000"; -- 0.053350996147229386
	pesos_i(16081) := b"1111111111111111_1111111111111111_1111100011001110_1011110110000110"; -- -0.028095392989611598
	pesos_i(16082) := b"1111111111111111_1111111111111111_1110101001010000_0001100000011010"; -- -0.08471536031632466
	pesos_i(16083) := b"1111111111111111_1111111111111111_1111010001011101_1111111111011110"; -- -0.04544068163946916
	pesos_i(16084) := b"1111111111111111_1111111111111111_1111010001111001_0101111111101001"; -- -0.045022969837891495
	pesos_i(16085) := b"1111111111111111_1111111111111111_1111111111000111_0111101000111010"; -- -0.0008624656226691128
	pesos_i(16086) := b"0000000000000000_0000000000000000_0001111111110111_0010000111001101"; -- 0.12486468554133637
	pesos_i(16087) := b"0000000000000000_0000000000000000_0000110111111010_1110010100010000"; -- 0.05460960056375827
	pesos_i(16088) := b"1111111111111111_1111111111111111_1111111100000110_0110000010011000"; -- -0.0038089397299221855
	pesos_i(16089) := b"1111111111111111_1111111111111111_1110011110001010_0000110100010000"; -- -0.09554975858458424
	pesos_i(16090) := b"0000000000000000_0000000000000000_0000011101110011_0101111000011011"; -- 0.029104119810164295
	pesos_i(16091) := b"1111111111111111_1111111111111111_1110000001011001_1100110101100101"; -- -0.12362972524402714
	pesos_i(16092) := b"1111111111111111_1111111111111111_1110110110100110_1110001100100010"; -- -0.07167225287992234
	pesos_i(16093) := b"0000000000000000_0000000000000000_0010001111110001_1000011101010010"; -- 0.14040418398748308
	pesos_i(16094) := b"1111111111111111_1111111111111111_1110000100110001_1101110001101011"; -- -0.12033293146643893
	pesos_i(16095) := b"1111111111111111_1111111111111111_1101111101001000_1011110100101111"; -- -0.12779634097241852
	pesos_i(16096) := b"1111111111111111_1111111111111111_1111010100100001_1000000101001001"; -- -0.042457503990340754
	pesos_i(16097) := b"0000000000000000_0000000000000000_0000111000111010_1100100110001011"; -- 0.055584522600106163
	pesos_i(16098) := b"0000000000000000_0000000000000000_0000101101110000_1100100110101111"; -- 0.04468975571221327
	pesos_i(16099) := b"1111111111111111_1111111111111111_1111111101001000_0100011011101000"; -- -0.002803390789855138
	pesos_i(16100) := b"0000000000000000_0000000000000000_0000101010101001_0110000010110101"; -- 0.041646999650671195
	pesos_i(16101) := b"0000000000000000_0000000000000000_0000111010100110_0110011001111010"; -- 0.05722656713627449
	pesos_i(16102) := b"0000000000000000_0000000000000000_0000010100101110_1101100100100111"; -- 0.020246097629355857
	pesos_i(16103) := b"0000000000000000_0000000000000000_0010000111000101_0001101001110110"; -- 0.13191380859925425
	pesos_i(16104) := b"0000000000000000_0000000000000000_0000100001001101_1010010001010001"; -- 0.03243472074004312
	pesos_i(16105) := b"1111111111111111_1111111111111111_1101111111100000_1000101110010001"; -- -0.12547996232829953
	pesos_i(16106) := b"1111111111111111_1111111111111111_1101100110100000_1011010000110101"; -- -0.14989160254011427
	pesos_i(16107) := b"0000000000000000_0000000000000000_0010010110010101_1011011001010001"; -- 0.1468156764954205
	pesos_i(16108) := b"1111111111111111_1111111111111111_1111110101001110_0100011100010010"; -- -0.01052432838477123
	pesos_i(16109) := b"0000000000000000_0000000000000000_0000010110000010_1011000100110100"; -- 0.021525454790716297
	pesos_i(16110) := b"0000000000000000_0000000000000000_0000010101010111_0001010010111100"; -- 0.020860000555063145
	pesos_i(16111) := b"1111111111111111_1111111111111111_1111101111011101_1111111000101001"; -- -0.01614390853490617
	pesos_i(16112) := b"1111111111111111_1111111111111111_1101111011001101_1011101100111000"; -- -0.12967328916875417
	pesos_i(16113) := b"1111111111111111_1111111111111111_1101110111010001_1100000110100001"; -- -0.1335181218254681
	pesos_i(16114) := b"0000000000000000_0000000000000000_0000011011011100_0000100010101010"; -- 0.026794950059264733
	pesos_i(16115) := b"1111111111111111_1111111111111111_1111010111000111_0001110000100010"; -- -0.039930574096553456
	pesos_i(16116) := b"0000000000000000_0000000000000000_0001011101100110_0011110100001100"; -- 0.09140378525070636
	pesos_i(16117) := b"1111111111111111_1111111111111111_1111111010100111_1111110101010011"; -- -0.005249182847477219
	pesos_i(16118) := b"1111111111111111_1111111111111111_1101111001100001_1111101011010010"; -- -0.1313174473778313
	pesos_i(16119) := b"0000000000000000_0000000000000000_0010010101101101_0101000011000101"; -- 0.14619927232927138
	pesos_i(16120) := b"0000000000000000_0000000000000000_0001000011111101_1011101100001110"; -- 0.06637162287312869
	pesos_i(16121) := b"1111111111111111_1111111111111111_1110001111110100_1000000110100111"; -- -0.10955037768489415
	pesos_i(16122) := b"1111111111111111_1111111111111111_1111001011001011_1010011111100011"; -- -0.05157995891587382
	pesos_i(16123) := b"1111111111111111_1111111111111111_1110010110111001_1110011001111001"; -- -0.10263213677730464
	pesos_i(16124) := b"0000000000000000_0000000000000000_0001001110011110_1100101100111001"; -- 0.07664175176883349
	pesos_i(16125) := b"1111111111111111_1111111111111111_1111101110100110_0000101011010111"; -- -0.016997644979906017
	pesos_i(16126) := b"1111111111111111_1111111111111111_1111011110000000_0111011110111111"; -- -0.03319598766097681
	pesos_i(16127) := b"0000000000000000_0000000000000000_0000001110111101_0100101110101100"; -- 0.014607171444644006
	pesos_i(16128) := b"0000000000000000_0000000000000000_0001100001100111_1011110110101110"; -- 0.09533296105176711
	pesos_i(16129) := b"1111111111111111_1111111111111111_1110010010000111_0110000011110001"; -- -0.10730928531822227
	pesos_i(16130) := b"0000000000000000_0000000000000000_0001101110011001_1101001101010100"; -- 0.10781594093119139
	pesos_i(16131) := b"1111111111111111_1111111111111111_1110110111000011_1011001111010010"; -- -0.07123256805728027
	pesos_i(16132) := b"0000000000000000_0000000000000000_0001110100000000_1100101000000000"; -- 0.11329329003582995
	pesos_i(16133) := b"0000000000000000_0000000000000000_0000001011011101_0010001100000000"; -- 0.01118677844485717
	pesos_i(16134) := b"0000000000000000_0000000000000000_0001001100010010_1111100011010001"; -- 0.07450823871785436
	pesos_i(16135) := b"1111111111111111_1111111111111111_1110111010011111_0000110000010011"; -- -0.06788563276049925
	pesos_i(16136) := b"1111111111111111_1111111111111111_1111011001010000_0010101010000010"; -- -0.03783926316167305
	pesos_i(16137) := b"0000000000000000_0000000000000000_0010011110000011_0111011101010100"; -- 0.15434976381255175
	pesos_i(16138) := b"0000000000000000_0000000000000000_0000010000010011_1000100100101011"; -- 0.01592309295252135
	pesos_i(16139) := b"0000000000000000_0000000000000000_0010000011101101_0101010010110101"; -- 0.12862138202852064
	pesos_i(16140) := b"0000000000000000_0000000000000000_0001101111001101_0110111010011101"; -- 0.10860339490820144
	pesos_i(16141) := b"1111111111111111_1111111111111111_1110001110101101_1111110000100010"; -- -0.11062645116286587
	pesos_i(16142) := b"0000000000000000_0000000000000000_0000000110100111_0011110100101101"; -- 0.006458114108265622
	pesos_i(16143) := b"0000000000000000_0000000000000000_0010001010111001_0000011100100010"; -- 0.13563580104856932
	pesos_i(16144) := b"0000000000000000_0000000000000000_0000101110011011_0110101001011001"; -- 0.0453402010421414
	pesos_i(16145) := b"0000000000000000_0000000000000000_0000011010110101_0010010100000010"; -- 0.026201546570464425
	pesos_i(16146) := b"0000000000000000_0000000000000000_0001011110110110_1100000111000111"; -- 0.09263239962745791
	pesos_i(16147) := b"1111111111111111_1111111111111111_1110100111111001_1010101000100010"; -- -0.08603417081788277
	pesos_i(16148) := b"1111111111111111_1111111111111111_1111010000001001_1001101010111010"; -- -0.04672844843581406
	pesos_i(16149) := b"0000000000000000_0000000000000000_0010101000100011_0111101110101000"; -- 0.16460392806895477
	pesos_i(16150) := b"0000000000000000_0000000000000000_0001001011011001_1011110011111010"; -- 0.0736349211246181
	pesos_i(16151) := b"1111111111111111_1111111111111111_1111111000111101_0001011010010110"; -- -0.0068803676001850675
	pesos_i(16152) := b"1111111111111111_1111111111111111_1110000010000000_0100110000110000"; -- -0.12304233381265842
	pesos_i(16153) := b"0000000000000000_0000000000000000_0001010001110110_0011110011101101"; -- 0.07992916853011287
	pesos_i(16154) := b"0000000000000000_0000000000000000_0000010111011000_1111001100011100"; -- 0.022841638875898893
	pesos_i(16155) := b"1111111111111111_1111111111111111_1101100101011110_0010110101110001"; -- -0.1509067152941591
	pesos_i(16156) := b"1111111111111111_1111111111111111_1111101000001001_1011011000111100"; -- -0.02328930896208642
	pesos_i(16157) := b"0000000000000000_0000000000000000_0001011110011100_0001101001111001"; -- 0.09222569909286125
	pesos_i(16158) := b"1111111111111111_1111111111111111_1110001111000110_1111000111000100"; -- -0.11024559933661222
	pesos_i(16159) := b"0000000000000000_0000000000000000_0000010110000101_0001110111111011"; -- 0.021562456021061105
	pesos_i(16160) := b"1111111111111111_1111111111111111_1111010101010111_0010101101010110"; -- -0.04163865242167872
	pesos_i(16161) := b"0000000000000000_0000000000000000_0010000010010000_1011101011010110"; -- 0.12720840181578183
	pesos_i(16162) := b"1111111111111111_1111111111111111_1110000011110001_0010110111110110"; -- -0.12131989237913741
	pesos_i(16163) := b"1111111111111111_1111111111111111_1111010011101000_1000100111101101"; -- -0.04332674000806373
	pesos_i(16164) := b"0000000000000000_0000000000000000_0000010111011010_0101111100011101"; -- 0.022863335155543573
	pesos_i(16165) := b"1111111111111111_1111111111111111_1101101110011001_1110001100100000"; -- -0.14218311745551226
	pesos_i(16166) := b"1111111111111111_1111111111111111_1111101010110110_1011100011010111"; -- -0.020649383044339453
	pesos_i(16167) := b"1111111111111111_1111111111111111_1111010001110111_1001101011000111"; -- -0.045049978609670846
	pesos_i(16168) := b"0000000000000000_0000000000000000_0001000100101111_1110100010010101"; -- 0.0671372760773262
	pesos_i(16169) := b"1111111111111111_1111111111111111_1110111110100000_0100110011101100"; -- -0.06396025895554051
	pesos_i(16170) := b"0000000000000000_0000000000000000_0001110011010001_1011101110101101"; -- 0.11257527330417964
	pesos_i(16171) := b"1111111111111111_1111111111111111_1101111100100100_0011010111101001"; -- -0.12835372028437933
	pesos_i(16172) := b"0000000000000000_0000000000000000_0001001000111101_0001001010010111"; -- 0.07124439408478006
	pesos_i(16173) := b"0000000000000000_0000000000000000_0000001010001011_0000010011001011"; -- 0.009933757288525724
	pesos_i(16174) := b"1111111111111111_1111111111111111_1110000111101100_1100101110100110"; -- -0.11748053736170173
	pesos_i(16175) := b"1111111111111111_1111111111111111_1111011011110100_0011100110001110"; -- -0.03533592503924057
	pesos_i(16176) := b"1111111111111111_1111111111111111_1110111000001101_0101001000001011"; -- -0.07010924560831482
	pesos_i(16177) := b"0000000000000000_0000000000000000_0001000001100100_1111111101100000"; -- 0.06404110053220068
	pesos_i(16178) := b"1111111111111111_1111111111111111_1101110100011111_1111111100010011"; -- -0.1362305239596933
	pesos_i(16179) := b"0000000000000000_0000000000000000_0000110111011011_0100011100011000"; -- 0.05412716233200668
	pesos_i(16180) := b"0000000000000000_0000000000000000_0010000110111000_1101001100100111"; -- 0.13172645281936
	pesos_i(16181) := b"1111111111111111_1111111111111111_1110101111110000_0111100110101110"; -- -0.07836188790309814
	pesos_i(16182) := b"1111111111111111_1111111111111111_1110010011011000_0110101010111101"; -- -0.10607273955933294
	pesos_i(16183) := b"0000000000000000_0000000000000000_0010011101111011_1100000010010011"; -- 0.15423205946750226
	pesos_i(16184) := b"0000000000000000_0000000000000000_0001000000010100_0010010101110101"; -- 0.06280740842995518
	pesos_i(16185) := b"1111111111111111_1111111111111111_1101011110110100_0110011111010000"; -- -0.15740348025825907
	pesos_i(16186) := b"1111111111111111_1111111111111111_1111010100110111_1110011110111011"; -- -0.04211570442045168
	pesos_i(16187) := b"0000000000000000_0000000000000000_0001101110110100_0110000100101011"; -- 0.10822112369501356
	pesos_i(16188) := b"0000000000000000_0000000000000000_0010000110110011_0101101110101010"; -- 0.13164303681552264
	pesos_i(16189) := b"0000000000000000_0000000000000000_0010011011111001_0110000011101101"; -- 0.152242715669686
	pesos_i(16190) := b"1111111111111111_1111111111111111_1111010010111100_1010010011011100"; -- -0.043996521283348265
	pesos_i(16191) := b"1111111111111111_1111111111111111_1110001001000010_1111000011101010"; -- -0.11616606022041644
	pesos_i(16192) := b"0000000000000000_0000000000000000_0000010000110111_0001100101000001"; -- 0.016465738538075123
	pesos_i(16193) := b"0000000000000000_0000000000000000_0010000110000100_1100010101000010"; -- 0.13093216765181837
	pesos_i(16194) := b"0000000000000000_0000000000000000_0001011000110101_0111100110111001"; -- 0.08675347106742598
	pesos_i(16195) := b"0000000000000000_0000000000000000_0000101010001101_0010001110001111"; -- 0.041216108754603444
	pesos_i(16196) := b"1111111111111111_1111111111111111_1111001010100000_0010000001110111"; -- -0.05224415867785193
	pesos_i(16197) := b"0000000000000000_0000000000000000_0010001001101001_0111101100100111"; -- 0.13442201336503198
	pesos_i(16198) := b"0000000000000000_0000000000000000_0001001000101000_0000110001110001"; -- 0.07092359319006838
	pesos_i(16199) := b"0000000000000000_0000000000000000_0001111110110111_0110100010110011"; -- 0.12389234884338177
	pesos_i(16200) := b"0000000000000000_0000000000000000_0001100001100001_0011111001000111"; -- 0.09523381463368302
	pesos_i(16201) := b"1111111111111111_1111111111111111_1110001000101101_1101001110011001"; -- -0.11648824228186029
	pesos_i(16202) := b"0000000000000000_0000000000000000_0001110101001000_1011111001011111"; -- 0.11439122989469913
	pesos_i(16203) := b"1111111111111111_1111111111111111_1110000000111001_1011100011001011"; -- -0.12411923458279671
	pesos_i(16204) := b"1111111111111111_1111111111111111_1101101100000011_0100011100001000"; -- -0.14448123978898103
	pesos_i(16205) := b"0000000000000000_0000000000000000_0001111111101111_1000011100011110"; -- 0.12474865416008844
	pesos_i(16206) := b"1111111111111111_1111111111111111_1111111110000011_0000010000001010"; -- -0.0019071079551881212
	pesos_i(16207) := b"0000000000000000_0000000000000000_0000101111001101_1101100110011011"; -- 0.046109772124024596
	pesos_i(16208) := b"0000000000000000_0000000000000000_0001111011111111_1101101001100010"; -- 0.12109150773091715
	pesos_i(16209) := b"0000000000000000_0000000000000000_0000001111100101_1100101000100000"; -- 0.015225060231161044
	pesos_i(16210) := b"1111111111111111_1111111111111111_1110101001000101_0001001100110100"; -- -0.08488349894350265
	pesos_i(16211) := b"1111111111111111_1111111111111111_1111111000101011_0111010111001111"; -- -0.007149350140013532
	pesos_i(16212) := b"1111111111111111_1111111111111111_1101100010110101_0100110100110001"; -- -0.15348355832073593
	pesos_i(16213) := b"1111111111111111_1111111111111111_1101100010001000_0110101110010110"; -- -0.15416839207580188
	pesos_i(16214) := b"0000000000000000_0000000000000000_0001000001110001_1000001001011101"; -- 0.06423201345448237
	pesos_i(16215) := b"1111111111111111_1111111111111111_1110001010000010_1010010110001100"; -- -0.11519399008645116
	pesos_i(16216) := b"1111111111111111_1111111111111111_1101110111110110_0111100111110010"; -- -0.13295781927488737
	pesos_i(16217) := b"0000000000000000_0000000000000000_0010100101010101_1000100010011101"; -- 0.16146138984700142
	pesos_i(16218) := b"1111111111111111_1111111111111111_1101111001000010_1110100000000110"; -- -0.13179159025688586
	pesos_i(16219) := b"0000000000000000_0000000000000000_0010001111101101_1010000000010101"; -- 0.14034462472125234
	pesos_i(16220) := b"0000000000000000_0000000000000000_0001001010010000_0101111111111011"; -- 0.07251548640762642
	pesos_i(16221) := b"0000000000000000_0000000000000000_0000000011010010_0100010111101010"; -- 0.0032085129714036565
	pesos_i(16222) := b"1111111111111111_1111111111111111_1111111110000010_1010100101000010"; -- -0.0019125188057756892
	pesos_i(16223) := b"0000000000000000_0000000000000000_0000110011011001_0101101001110000"; -- 0.05019154766950921
	pesos_i(16224) := b"1111111111111111_1111111111111111_1111110011100011_1011011111011111"; -- -0.012150295405704569
	pesos_i(16225) := b"0000000000000000_0000000000000000_0001000001011001_1110101100111111"; -- 0.06387205390954354
	pesos_i(16226) := b"0000000000000000_0000000000000000_0001010001000001_0110001000101011"; -- 0.07912267261672648
	pesos_i(16227) := b"1111111111111111_1111111111111111_1110110111110101_0010111111001100"; -- -0.07047749786059895
	pesos_i(16228) := b"1111111111111111_1111111111111111_1110001110100000_0110000000110000"; -- -0.11083411050939448
	pesos_i(16229) := b"0000000000000000_0000000000000000_0010000111110010_0000011111000100"; -- 0.13259933981238084
	pesos_i(16230) := b"1111111111111111_1111111111111111_1101110111111111_1111000001100001"; -- -0.13281343112385782
	pesos_i(16231) := b"0000000000000000_0000000000000000_0000010001111011_1000101000100100"; -- 0.017510064853598968
	pesos_i(16232) := b"1111111111111111_1111111111111111_1111100000001101_0000111000111100"; -- -0.031050787208566313
	pesos_i(16233) := b"1111111111111111_1111111111111111_1111110000110001_1001010100000011"; -- -0.014868437480602181
	pesos_i(16234) := b"0000000000000000_0000000000000000_0000010100011011_0010011101010010"; -- 0.01994558095460453
	pesos_i(16235) := b"1111111111111111_1111111111111111_1101111001000110_1100101110101110"; -- -0.13173224440340833
	pesos_i(16236) := b"1111111111111111_1111111111111111_1110101110100111_0110000101110101"; -- -0.07947722324215371
	pesos_i(16237) := b"1111111111111111_1111111111111111_1110001011000100_0100100101100001"; -- -0.11419240372200691
	pesos_i(16238) := b"1111111111111111_1111111111111111_1111110110111111_1001001101001110"; -- -0.008795541191535841
	pesos_i(16239) := b"1111111111111111_1111111111111111_1110011001110000_0010110011001000"; -- -0.09985084655458429
	pesos_i(16240) := b"1111111111111111_1111111111111111_1111000111001100_1011101111111001"; -- -0.05546975307562655
	pesos_i(16241) := b"0000000000000000_0000000000000000_0001000101011011_0111111011011111"; -- 0.06780236189641276
	pesos_i(16242) := b"1111111111111111_1111111111111111_1111011100100011_0010010101110100"; -- -0.03461996000572974
	pesos_i(16243) := b"0000000000000000_0000000000000000_0000111000110001_0101010011111001"; -- 0.05544024534197937
	pesos_i(16244) := b"0000000000000000_0000000000000000_0000010100001110_0111100100100111"; -- 0.019752094381985833
	pesos_i(16245) := b"1111111111111111_1111111111111111_1111000000111010_1000100110111011"; -- -0.06160678083335263
	pesos_i(16246) := b"1111111111111111_1111111111111111_1101100001101101_1110100011110001"; -- -0.15457290756661038
	pesos_i(16247) := b"0000000000000000_0000000000000000_0010001010011110_0011101001111110"; -- 0.1352268751653936
	pesos_i(16248) := b"0000000000000000_0000000000000000_0001101100100010_1100011011011011"; -- 0.10599940163956047
	pesos_i(16249) := b"1111111111111111_1111111111111111_1101111011011001_0111110110011010"; -- -0.12949385635324207
	pesos_i(16250) := b"1111111111111111_1111111111111111_1111011000000001_1011111101000111"; -- -0.03903584026444716
	pesos_i(16251) := b"1111111111111111_1111111111111111_1110111111010111_0000000101111000"; -- -0.06312552291315794
	pesos_i(16252) := b"0000000000000000_0000000000000000_0001010101100001_1001101101100000"; -- 0.08352061361954334
	pesos_i(16253) := b"0000000000000000_0000000000000000_0010010111001011_0000110111011101"; -- 0.14762961037954409
	pesos_i(16254) := b"1111111111111111_1111111111111111_1101111010100101_0111001110111101"; -- -0.13028790130224627
	pesos_i(16255) := b"1111111111111111_1111111111111111_1101110100001111_0101000000000011"; -- -0.1364850990876458
	pesos_i(16256) := b"0000000000000000_0000000000000000_0000110011101100_0011111010101110"; -- 0.05047981016134725
	pesos_i(16257) := b"1111111111111111_1111111111111111_1111011010011000_1100110010010001"; -- -0.03673097092977251
	pesos_i(16258) := b"0000000000000000_0000000000000000_0010100101100111_1100000001110101"; -- 0.16173937656453533
	pesos_i(16259) := b"1111111111111111_1111111111111111_1110011011010101_1101010010100100"; -- -0.09829970355606299
	pesos_i(16260) := b"1111111111111111_1111111111111111_1111100000011110_1100000011100101"; -- -0.030780738927422516
	pesos_i(16261) := b"0000000000000000_0000000000000000_0000011010010110_0001011111111000"; -- 0.025727747042449293
	pesos_i(16262) := b"0000000000000000_0000000000000000_0010001011101111_1111110111000010"; -- 0.13647447572135168
	pesos_i(16263) := b"1111111111111111_1111111111111111_1111110111111001_1100011010111011"; -- -0.007907466171983662
	pesos_i(16264) := b"1111111111111111_1111111111111111_1110110110100101_0001010101000110"; -- -0.0716997818761117
	pesos_i(16265) := b"1111111111111111_1111111111111111_1111111111000100_0010000011010100"; -- -0.0009135706681728254
	pesos_i(16266) := b"0000000000000000_0000000000000000_0001101000100101_1110001001011110"; -- 0.10214056771336444
	pesos_i(16267) := b"0000000000000000_0000000000000000_0000001011101011_1000000011001101"; -- 0.011405992576447697
	pesos_i(16268) := b"1111111111111111_1111111111111111_1110011111100011_0111011001011000"; -- -0.09418545100585492
	pesos_i(16269) := b"1111111111111111_1111111111111111_1111111100010101_1110101101011101"; -- -0.0035717866733177904
	pesos_i(16270) := b"0000000000000000_0000000000000000_0000001010101000_0101110001001010"; -- 0.010381477347043888
	pesos_i(16271) := b"0000000000000000_0000000000000000_0000111011001111_0110111000110101"; -- 0.05785263814309682
	pesos_i(16272) := b"0000000000000000_0000000000000000_0000010010111101_1001100101001101"; -- 0.018518048660226983
	pesos_i(16273) := b"1111111111111111_1111111111111111_1101110100111111_0101001001110111"; -- -0.13575253111499155
	pesos_i(16274) := b"0000000000000000_0000000000000000_0000000011010101_1010010000011100"; -- 0.0032599036766873908
	pesos_i(16275) := b"1111111111111111_1111111111111111_1110000010011101_1010010010110000"; -- -0.12259455388037396
	pesos_i(16276) := b"0000000000000000_0000000000000000_0000100011001100_0100001011110000"; -- 0.034366782696268076
	pesos_i(16277) := b"0000000000000000_0000000000000000_0001110101001101_1101000011000100"; -- 0.11446862015043101
	pesos_i(16278) := b"1111111111111111_1111111111111111_1110010101001000_0101111010101111"; -- -0.10436447366424234
	pesos_i(16279) := b"1111111111111111_1111111111111111_1111101101101101_0100110100010111"; -- -0.0178634470829147
	pesos_i(16280) := b"1111111111111111_1111111111111111_1110100101110011_1100111100100100"; -- -0.08807664276292544
	pesos_i(16281) := b"0000000000000000_0000000000000000_0000000101110011_0101111001101000"; -- 0.0056666377394607136
	pesos_i(16282) := b"1111111111111111_1111111111111111_1110101011010000_0100011111000111"; -- -0.08275939371604299
	pesos_i(16283) := b"1111111111111111_1111111111111111_1110010101100111_1010011100011110"; -- -0.10388713381871606
	pesos_i(16284) := b"0000000000000000_0000000000000000_0010000001001101_1110100100101101"; -- 0.12618882513609145
	pesos_i(16285) := b"1111111111111111_1111111111111111_1101110011110101_1110110101000000"; -- -0.13687245538726067
	pesos_i(16286) := b"1111111111111111_1111111111111111_1110100100110000_1101100000011111"; -- -0.08909844634912009
	pesos_i(16287) := b"0000000000000000_0000000000000000_0010000110100010_1000001010011111"; -- 0.13138595941430573
	pesos_i(16288) := b"0000000000000000_0000000000000000_0001000001011000_0001001110101000"; -- 0.0638439450193851
	pesos_i(16289) := b"0000000000000000_0000000000000000_0001101001010100_0111100011010011"; -- 0.10285144007786517
	pesos_i(16290) := b"1111111111111111_1111111111111111_1110110111100110_1110110011001101"; -- -0.07069511414965847
	pesos_i(16291) := b"0000000000000000_0000000000000000_0000100111101111_1000001101100011"; -- 0.038810931881461376
	pesos_i(16292) := b"0000000000000000_0000000000000000_0010000011010101_0010001000111100"; -- 0.12825216251889124
	pesos_i(16293) := b"0000000000000000_0000000000000000_0000111001110110_0100011001010001"; -- 0.05649222836078101
	pesos_i(16294) := b"0000000000000000_0000000000000000_0000101010000100_1011011001110110"; -- 0.04108753568957073
	pesos_i(16295) := b"0000000000000000_0000000000000000_0010010111100000_1101100011100111"; -- 0.14796214721284354
	pesos_i(16296) := b"1111111111111111_1111111111111111_1110011100101100_0100100100100010"; -- -0.09698050412646195
	pesos_i(16297) := b"0000000000000000_0000000000000000_0000100101011011_0000000000010000"; -- 0.036544803589505716
	pesos_i(16298) := b"0000000000000000_0000000000000000_0000111010110111_1110001110110000"; -- 0.0574934295648742
	pesos_i(16299) := b"0000000000000000_0000000000000000_0001100110101110_1001110010111100"; -- 0.10032062133499912
	pesos_i(16300) := b"1111111111111111_1111111111111111_1110010101001101_1000111001100000"; -- -0.10428533692945881
	pesos_i(16301) := b"1111111111111111_1111111111111111_1110110010010111_0111010000101001"; -- -0.07581399926053996
	pesos_i(16302) := b"1111111111111111_1111111111111111_1111001111111011_0101011010001101"; -- -0.04694613520424062
	pesos_i(16303) := b"0000000000000000_0000000000000000_0000110000100011_0100001000001100"; -- 0.04741299425116185
	pesos_i(16304) := b"0000000000000000_0000000000000000_0000111110011000_1100000011010110"; -- 0.06092457993281221
	pesos_i(16305) := b"0000000000000000_0000000000000000_0001110010000111_1001101011110110"; -- 0.11144417282509704
	pesos_i(16306) := b"1111111111111111_1111111111111111_1111100010010100_1101000100001010"; -- -0.02897923955168839
	pesos_i(16307) := b"1111111111111111_1111111111111111_1111000011101101_1000011100000101"; -- -0.05887561929158031
	pesos_i(16308) := b"0000000000000000_0000000000000000_0000111100001100_0011100010100001"; -- 0.058780230855603174
	pesos_i(16309) := b"0000000000000000_0000000000000000_0000011101110001_1000110111011111"; -- 0.029076449320999107
	pesos_i(16310) := b"1111111111111111_1111111111111111_1110110101000110_1100010101110101"; -- -0.07313886551433099
	pesos_i(16311) := b"0000000000000000_0000000000000000_0010001101010110_0101000010111000"; -- 0.13803581701631032
	pesos_i(16312) := b"0000000000000000_0000000000000000_0000001101011100_0001000011101001"; -- 0.01312356647903392
	pesos_i(16313) := b"1111111111111111_1111111111111111_1110010111101010_1100001111110111"; -- -0.10188651299372715
	pesos_i(16314) := b"0000000000000000_0000000000000000_0010011011110100_1011010110110100"; -- 0.15217147480882887
	pesos_i(16315) := b"0000000000000000_0000000000000000_0001010011001010_0100000011111110"; -- 0.08121114915692655
	pesos_i(16316) := b"0000000000000000_0000000000000000_0001011001010111_1011100110110111"; -- 0.08727608420813947
	pesos_i(16317) := b"1111111111111111_1111111111111111_1110111110100001_1111111100010011"; -- -0.06393438140992774
	pesos_i(16318) := b"0000000000000000_0000000000000000_0001101101000011_0001110000110010"; -- 0.10649276933525831
	pesos_i(16319) := b"0000000000000000_0000000000000000_0010010101110000_1000000000101010"; -- 0.1462478734827656
	pesos_i(16320) := b"0000000000000000_0000000000000000_0001110110100001_0110011000111111"; -- 0.11574400946315792
	pesos_i(16321) := b"1111111111111111_1111111111111111_1101100101100010_1100011000001101"; -- -0.1508365839247948
	pesos_i(16322) := b"1111111111111111_1111111111111111_1111000100010101_1010110101010110"; -- -0.05826298382403514
	pesos_i(16323) := b"1111111111111111_1111111111111111_1101100001110011_1100001001111111"; -- -0.15448364650110308
	pesos_i(16324) := b"0000000000000000_0000000000000000_0010000101110000_1111101110100001"; -- 0.1306302327184921
	pesos_i(16325) := b"1111111111111111_1111111111111111_1110100011000001_0111110010100100"; -- -0.09079762447186178
	pesos_i(16326) := b"0000000000000000_0000000000000000_0001111111110010_1110100001110000"; -- 0.12480023136367292
	pesos_i(16327) := b"1111111111111111_1111111111111111_1111100100100101_1010101010101010"; -- -0.026769002469807866
	pesos_i(16328) := b"0000000000000000_0000000000000000_0000101011011010_0001100001011110"; -- 0.042390368307225285
	pesos_i(16329) := b"1111111111111111_1111111111111111_1111111010100101_0101001101100010"; -- -0.005289829686622613
	pesos_i(16330) := b"1111111111111111_1111111111111111_1110101011111101_1010000010100011"; -- -0.08206745166348003
	pesos_i(16331) := b"0000000000000000_0000000000000000_0000011011100111_0001101010011000"; -- 0.026963865367485698
	pesos_i(16332) := b"0000000000000000_0000000000000000_0000100101001010_0110011101010000"; -- 0.03629155834029741
	pesos_i(16333) := b"1111111111111111_1111111111111111_1101110001101101_1001011011101110"; -- -0.13895279596024748
	pesos_i(16334) := b"0000000000000000_0000000000000000_0000011011001101_0101110100110011"; -- 0.026571106783336254
	pesos_i(16335) := b"1111111111111111_1111111111111111_1111010001010011_0100011100001100"; -- -0.04560428583768775
	pesos_i(16336) := b"1111111111111111_1111111111111111_1111000101111001_1100000001110101"; -- -0.056735965195800715
	pesos_i(16337) := b"0000000000000000_0000000000000000_0000011010110011_1010000001101011"; -- 0.026178384996854764
	pesos_i(16338) := b"0000000000000000_0000000000000000_0000100001101101_1110111010101001"; -- 0.032927433348952886
	pesos_i(16339) := b"0000000000000000_0000000000000000_0010000001111011_1100011010111100"; -- 0.12688867652762395
	pesos_i(16340) := b"1111111111111111_1111111111111111_1111111100011110_0010110111000011"; -- -0.0034457587819284666
	pesos_i(16341) := b"0000000000000000_0000000000000000_0001100101101110_0000101100010001"; -- 0.09933537636201993
	pesos_i(16342) := b"1111111111111111_1111111111111111_1111101010101100_1001100010011000"; -- -0.020803892891114374
	pesos_i(16343) := b"0000000000000000_0000000000000000_0001001010001111_0010001010101000"; -- 0.07249657256553363
	pesos_i(16344) := b"0000000000000000_0000000000000000_0000110101000000_1011101010010111"; -- 0.051768934064708304
	pesos_i(16345) := b"1111111111111111_1111111111111111_1110100100001110_1011001100101000"; -- -0.08961944837003079
	pesos_i(16346) := b"1111111111111111_1111111111111111_1110111111000101_1101101000011100"; -- -0.06338726812221597
	pesos_i(16347) := b"1111111111111111_1111111111111111_1110111011010111_1110001111100100"; -- -0.0670182770858524
	pesos_i(16348) := b"1111111111111111_1111111111111111_1111101110101110_0100010100111001"; -- -0.016872094771825472
	pesos_i(16349) := b"1111111111111111_1111111111111111_1111101010101001_1000000011100111"; -- -0.02085108153239553
	pesos_i(16350) := b"1111111111111111_1111111111111111_1110001011011001_1101100001101011"; -- -0.11386344324042336
	pesos_i(16351) := b"1111111111111111_1111111111111111_1101101011001111_0101000011011000"; -- -0.145274112053198
	pesos_i(16352) := b"1111111111111111_1111111111111111_1111101111111011_1011011100100010"; -- -0.015690378397035826
	pesos_i(16353) := b"0000000000000000_0000000000000000_0000011101011010_1011111110101100"; -- 0.0287284656090128
	pesos_i(16354) := b"0000000000000000_0000000000000000_0001011010000011_0001001100100001"; -- 0.08793754153420472
	pesos_i(16355) := b"0000000000000000_0000000000000000_0000001001111000_0001101010110101"; -- 0.009645146550089414
	pesos_i(16356) := b"1111111111111111_1111111111111111_1110111110111111_0010110010010010"; -- -0.06348916475674031
	pesos_i(16357) := b"1111111111111111_1111111111111111_1101100010101011_0110111110010101"; -- -0.1536340962794287
	pesos_i(16358) := b"0000000000000000_0000000000000000_0001110010100101_0010010101000111"; -- 0.11189492219742549
	pesos_i(16359) := b"0000000000000000_0000000000000000_0001000000000001_1000011111101100"; -- 0.06252336046023352
	pesos_i(16360) := b"0000000000000000_0000000000000000_0000100011110100_0100111100001011"; -- 0.03497785592261722
	pesos_i(16361) := b"1111111111111111_1111111111111111_1110100010111110_1010100010110001"; -- -0.09084077530637318
	pesos_i(16362) := b"0000000000000000_0000000000000000_0001010101000101_1100110010101010"; -- 0.08309630533120096
	pesos_i(16363) := b"1111111111111111_1111111111111111_1111011011011001_0011110000101001"; -- -0.035747756993491524
	pesos_i(16364) := b"1111111111111111_1111111111111111_1110111001100100_0000110110101111"; -- -0.06878580549315672
	pesos_i(16365) := b"0000000000000000_0000000000000000_0001101010110110_1001110010110001"; -- 0.10434893921877945
	pesos_i(16366) := b"1111111111111111_1111111111111111_1111000101110001_0000100000000111"; -- -0.05686902846309237
	pesos_i(16367) := b"1111111111111111_1111111111111111_1110011101110101_0110110110111000"; -- -0.09586443197531272
	pesos_i(16368) := b"0000000000000000_0000000000000000_0000010101011111_1010011111001011"; -- 0.020990836222371287
	pesos_i(16369) := b"0000000000000000_0000000000000000_0000111010111100_1001010001101011"; -- 0.05756499881163861
	pesos_i(16370) := b"0000000000000000_0000000000000000_0001111000000000_0111111001011001"; -- 0.1171950310080407
	pesos_i(16371) := b"1111111111111111_1111111111111111_1110000110101101_0110000010011010"; -- -0.1184482216523543
	pesos_i(16372) := b"0000000000000000_0000000000000000_0001100111101011_0111100001100001"; -- 0.10124924059113041
	pesos_i(16373) := b"0000000000000000_0000000000000000_0001010000101011_1101111011011001"; -- 0.07879441071352465
	pesos_i(16374) := b"0000000000000000_0000000000000000_0010001101101111_0110110001000001"; -- 0.13841892809728884
	pesos_i(16375) := b"0000000000000000_0000000000000000_0001110001111111_0011001011110011"; -- 0.11131590311728566
	pesos_i(16376) := b"0000000000000000_0000000000000000_0010011000011011_1001100010110110"; -- 0.14885858962101506
	pesos_i(16377) := b"0000000000000000_0000000000000000_0001001011011101_0010110111111110"; -- 0.07368743368970365
	pesos_i(16378) := b"0000000000000000_0000000000000000_0010000100100011_1110000010101000"; -- 0.1294536980580039
	pesos_i(16379) := b"0000000000000000_0000000000000000_0001100011001001_1100111000111001"; -- 0.09682930834472378
	pesos_i(16380) := b"0000000000000000_0000000000000000_0000001000110011_1110101010010110"; -- 0.008604680641061417
	pesos_i(16381) := b"1111111111111111_1111111111111111_1111011111001010_1101000000110010"; -- -0.032061565174104634
	pesos_i(16382) := b"0000000000000000_0000000000000000_0010010101000111_1100001011111111"; -- 0.14562624680588318
	pesos_i(16383) := b"1111111111111111_1111111111111111_1110101011010100_0111010001011001"; -- -0.08269570192554171
	pesos_i(16384) := b"1111111111111111_1111111111111111_1110000011001100_1101110101001011"; -- -0.12187401705509204
	pesos_i(16385) := b"0000000000000000_0000000000000000_0010000000111011_1010100111100000"; -- 0.12591039396460288
	pesos_i(16386) := b"1111111111111111_1111111111111111_1111001001001010_0000110001110101"; -- -0.053557607117034785
	pesos_i(16387) := b"0000000000000000_0000000000000000_0010011011110111_1101000101101110"; -- 0.1522189038922654
	pesos_i(16388) := b"0000000000000000_0000000000000000_0001010110101100_1011101000000101"; -- 0.08466684933429836
	pesos_i(16389) := b"0000000000000000_0000000000000000_0000001111010111_1001110010001001"; -- 0.015008719794843244
	pesos_i(16390) := b"1111111111111111_1111111111111111_1111011100011000_0100100001000110"; -- -0.03478573128045215
	pesos_i(16391) := b"1111111111111111_1111111111111111_1111100010100100_1110010010000100"; -- -0.028733937889337615
	pesos_i(16392) := b"0000000000000000_0000000000000000_0010000001000110_1001111000001101"; -- 0.12607753580006287
	pesos_i(16393) := b"0000000000000000_0000000000000000_0001111000101011_1010010101110100"; -- 0.11785348960279193
	pesos_i(16394) := b"0000000000000000_0000000000000000_0001101000001011_0101100001110110"; -- 0.10173561930925595
	pesos_i(16395) := b"1111111111111111_1111111111111111_1110111111100011_1110011110100001"; -- -0.06292869868887366
	pesos_i(16396) := b"0000000000000000_0000000000000000_0001011101001010_0110101111100100"; -- 0.09097933107226408
	pesos_i(16397) := b"0000000000000000_0000000000000000_0000100001100111_1010001000000001"; -- 0.032831311550682515
	pesos_i(16398) := b"0000000000000000_0000000000000000_0000110111001000_1001100100000101"; -- 0.05384212842950066
	pesos_i(16399) := b"0000000000000000_0000000000000000_0001111110001011_1001101000001010"; -- 0.12322390301925049
	pesos_i(16400) := b"1111111111111111_1111111111111111_1111000010000100_1010001000111111"; -- -0.06047616933074833
	pesos_i(16401) := b"1111111111111111_1111111111111111_1110110110101111_1000010101110101"; -- -0.07154050730044796
	pesos_i(16402) := b"0000000000000000_0000000000000000_0000000110010111_0101110011011000"; -- 0.0062158609588506076
	pesos_i(16403) := b"0000000000000000_0000000000000000_0000111110110001_0001110000100110"; -- 0.06129623354295596
	pesos_i(16404) := b"1111111111111111_1111111111111111_1111100011010010_0100110100110010"; -- -0.028041053017071438
	pesos_i(16405) := b"1111111111111111_1111111111111111_1111110100110111_0000000101011011"; -- -0.010879435751179544
	pesos_i(16406) := b"1111111111111111_1111111111111111_1111011011001001_0101100000000000"; -- -0.03599023818001874
	pesos_i(16407) := b"1111111111111111_1111111111111111_1101111000010010_1111000111010110"; -- -0.13252342729575456
	pesos_i(16408) := b"0000000000000000_0000000000000000_0000101111101100_1101011010100011"; -- 0.0465826175683667
	pesos_i(16409) := b"1111111111111111_1111111111111111_1110001010101111_0101000111000010"; -- -0.11451233885298748
	pesos_i(16410) := b"0000000000000000_0000000000000000_0000000111110101_1000110000110111"; -- 0.007653010875279052
	pesos_i(16411) := b"1111111111111111_1111111111111111_1111100100000001_1011100001011100"; -- -0.027317502615425062
	pesos_i(16412) := b"0000000000000000_0000000000000000_0010010001100100_0100110010110011"; -- 0.14215545062838564
	pesos_i(16413) := b"1111111111111111_1111111111111111_1110000110001110_1111000001011001"; -- -0.1189126760288403
	pesos_i(16414) := b"1111111111111111_1111111111111111_1111010001010010_0101101000101100"; -- -0.0456184047048558
	pesos_i(16415) := b"0000000000000000_0000000000000000_0000111000100101_0111101011101011"; -- 0.055259401607940704
	pesos_i(16416) := b"0000000000000000_0000000000000000_0001110110101101_1011101001100011"; -- 0.11593213001998141
	pesos_i(16417) := b"1111111111111111_1111111111111111_1110000010111010_0110101100000111"; -- -0.12215548589844913
	pesos_i(16418) := b"1111111111111111_1111111111111111_1101101101001001_1110011110010001"; -- -0.14340355593177231
	pesos_i(16419) := b"1111111111111111_1111111111111111_1110110111010110_0010110011110010"; -- -0.07095069017984357
	pesos_i(16420) := b"1111111111111111_1111111111111111_1110000010010010_1000011000101111"; -- -0.1227642187546695
	pesos_i(16421) := b"0000000000000000_0000000000000000_0000011011010111_0100101011110001"; -- 0.026722606419541127
	pesos_i(16422) := b"0000000000000000_0000000000000000_0000001101001010_0010110010010100"; -- 0.012850557468173996
	pesos_i(16423) := b"1111111111111111_1111111111111111_1111010100010000_0001101110011101"; -- -0.042722963441979886
	pesos_i(16424) := b"0000000000000000_0000000000000000_0001001100100100_0110100011101001"; -- 0.07477431961819815
	pesos_i(16425) := b"1111111111111111_1111111111111111_1110001011101001_0100101010110110"; -- -0.11362774905672386
	pesos_i(16426) := b"0000000000000000_0000000000000000_0000101001111101_1010011001001001"; -- 0.04097976000792911
	pesos_i(16427) := b"0000000000000000_0000000000000000_0000011101101000_1011111100101010"; -- 0.028942058368511908
	pesos_i(16428) := b"1111111111111111_1111111111111111_1110010010000111_1000001100000000"; -- -0.10730725525275907
	pesos_i(16429) := b"1111111111111111_1111111111111111_1111000110101011_1011111101000000"; -- -0.055973097613217726
	pesos_i(16430) := b"0000000000000000_0000000000000000_0001110100001101_1001100100011010"; -- 0.1134887398481137
	pesos_i(16431) := b"1111111111111111_1111111111111111_1111101100110100_1001011110110010"; -- -0.01872875121935733
	pesos_i(16432) := b"0000000000000000_0000000000000000_0010011110110011_1011001000001000"; -- 0.1550856848121211
	pesos_i(16433) := b"0000000000000000_0000000000000000_0010001111000111_1001101101100110"; -- 0.1397645114591176
	pesos_i(16434) := b"1111111111111111_1111111111111111_1111001011100111_1101100100111010"; -- -0.05114977202208439
	pesos_i(16435) := b"0000000000000000_0000000000000000_0001100110111110_1110111100101000"; -- 0.10056967462912594
	pesos_i(16436) := b"0000000000000000_0000000000000000_0001111111000100_1001011000010100"; -- 0.12409341808832597
	pesos_i(16437) := b"1111111111111111_1111111111111111_1110001101011101_0111101011111110"; -- -0.111854851818005
	pesos_i(16438) := b"1111111111111111_1111111111111111_1110011001000010_0000101001001001"; -- -0.10055480695005145
	pesos_i(16439) := b"0000000000000000_0000000000000000_0000010101011010_1101010011111110"; -- 0.020917236366688442
	pesos_i(16440) := b"0000000000000000_0000000000000000_0000000000101001_1000101001111001"; -- 0.0006338640676260015
	pesos_i(16441) := b"1111111111111111_1111111111111111_1110011111000010_1110010011100000"; -- -0.09468240299178897
	pesos_i(16442) := b"1111111111111111_1111111111111111_1110011110111101_1010111111101000"; -- -0.09476185399880244
	pesos_i(16443) := b"1111111111111111_1111111111111111_1110010110111100_0001100010000011"; -- -0.10259863670703805
	pesos_i(16444) := b"0000000000000000_0000000000000000_0000000010010110_0011101011110110"; -- 0.0022923326285793208
	pesos_i(16445) := b"0000000000000000_0000000000000000_0010101100011110_1000011001101001"; -- 0.16843452522779592
	pesos_i(16446) := b"1111111111111111_1111111111111111_1111011111110001_1100111101110010"; -- -0.03146651723660717
	pesos_i(16447) := b"0000000000000000_0000000000000000_0001110110000001_0100100111011100"; -- 0.11525403607926078
	pesos_i(16448) := b"0000000000000000_0000000000000000_0010000111010101_1011101100000000"; -- 0.13216751806466845
	pesos_i(16449) := b"1111111111111111_1111111111111111_1111000111001010_0001011111101111"; -- -0.05551004813086992
	pesos_i(16450) := b"1111111111111111_1111111111111111_1101101000001011_1001111000001011"; -- -0.14826023319252163
	pesos_i(16451) := b"0000000000000000_0000000000000000_0001001011111100_0011011011001010"; -- 0.07416098048783591
	pesos_i(16452) := b"1111111111111111_1111111111111111_1101101100111011_0010000110010001"; -- -0.1436289806677527
	pesos_i(16453) := b"0000000000000000_0000000000000000_0000111100000100_1011001101101010"; -- 0.05866547913815189
	pesos_i(16454) := b"1111111111111111_1111111111111111_1111011000011010_1011101101101010"; -- -0.03865460074631138
	pesos_i(16455) := b"1111111111111111_1111111111111111_1110000010010111_1110000100010100"; -- -0.12268250725820148
	pesos_i(16456) := b"1111111111111111_1111111111111111_1111001111100111_0111011011010011"; -- -0.047249387202093304
	pesos_i(16457) := b"0000000000000000_0000000000000000_0001010010111100_1000110110001011"; -- 0.08100208885783079
	pesos_i(16458) := b"1111111111111111_1111111111111111_1110101110111111_1001000000101100"; -- -0.07910822804785382
	pesos_i(16459) := b"1111111111111111_1111111111111111_1110111010101111_1111011000111101"; -- -0.06762753490101606
	pesos_i(16460) := b"1111111111111111_1111111111111111_1110111001000100_0110010101000010"; -- -0.06926886688770743
	pesos_i(16461) := b"0000000000000000_0000000000000000_0000111011100000_0101010111001100"; -- 0.05811058272943634
	pesos_i(16462) := b"1111111111111111_1111111111111111_1111000111100100_1111100010100111"; -- -0.05509992516004518
	pesos_i(16463) := b"0000000000000000_0000000000000000_0010000010010111_0011101001111110"; -- 0.12730756357461864
	pesos_i(16464) := b"0000000000000000_0000000000000000_0000111001101001_1110010111011111"; -- 0.056303374217371076
	pesos_i(16465) := b"0000000000000000_0000000000000000_0010011001010000_1000000110001001"; -- 0.14966592411568735
	pesos_i(16466) := b"0000000000000000_0000000000000000_0010001101110001_1101010111110111"; -- 0.138455746558602
	pesos_i(16467) := b"1111111111111111_1111111111111111_1110000100100110_1110100001111011"; -- -0.12050005917207846
	pesos_i(16468) := b"1111111111111111_1111111111111111_1110101100100001_1110011101010101"; -- -0.08151392148218435
	pesos_i(16469) := b"0000000000000000_0000000000000000_0000010001001100_0101000100111000"; -- 0.016789508951022727
	pesos_i(16470) := b"1111111111111111_1111111111111111_1110000001010000_0110010001101010"; -- -0.1237733117125269
	pesos_i(16471) := b"0000000000000000_0000000000000000_0000100110110000_0000100111111110"; -- 0.0378423925387495
	pesos_i(16472) := b"0000000000000000_0000000000000000_0001010001001110_1001001000011011"; -- 0.07932389414809686
	pesos_i(16473) := b"1111111111111111_1111111111111111_1110011110000011_0001010011000110"; -- -0.09565611053435927
	pesos_i(16474) := b"0000000000000000_0000000000000000_0001011011100000_1001110000100100"; -- 0.08936477555976559
	pesos_i(16475) := b"0000000000000000_0000000000000000_0001001110100001_1111100000011000"; -- 0.07669020263159122
	pesos_i(16476) := b"1111111111111111_1111111111111111_1111011001110011_1100001010100001"; -- -0.03729613842352622
	pesos_i(16477) := b"1111111111111111_1111111111111111_1111000010000100_1101111010011011"; -- -0.06047257156441061
	pesos_i(16478) := b"1111111111111111_1111111111111111_1111110010100110_1011000110001001"; -- -0.01308145907433637
	pesos_i(16479) := b"0000000000000000_0000000000000000_0001111011011110_1000101000001000"; -- 0.1205831785301528
	pesos_i(16480) := b"1111111111111111_1111111111111111_1110101111110010_0000101011110000"; -- -0.07833797109836142
	pesos_i(16481) := b"1111111111111111_1111111111111111_1111110010101101_0101011000101111"; -- -0.012980092479323097
	pesos_i(16482) := b"0000000000000000_0000000000000000_0000011001100010_0001101010111110"; -- 0.024934455309650484
	pesos_i(16483) := b"1111111111111111_1111111111111111_1110101100111000_1011101010100000"; -- -0.08116563400969
	pesos_i(16484) := b"1111111111111111_1111111111111111_1111111000001010_0100100001111101"; -- -0.007655591483482777
	pesos_i(16485) := b"1111111111111111_1111111111111111_1111011110110010_1101110100010101"; -- -0.032427007986049666
	pesos_i(16486) := b"1111111111111111_1111111111111111_1110100101110010_1110001000011110"; -- -0.08809077049374626
	pesos_i(16487) := b"1111111111111111_1111111111111111_1110100100010100_1011001011100111"; -- -0.08952791077864493
	pesos_i(16488) := b"0000000000000000_0000000000000000_0010001000010000_1111110001000100"; -- 0.13307167674213155
	pesos_i(16489) := b"0000000000000000_0000000000000000_0001110101001000_1011001101111011"; -- 0.11439058057236232
	pesos_i(16490) := b"0000000000000000_0000000000000000_0001100000011101_0110110000101010"; -- 0.09419895190257628
	pesos_i(16491) := b"0000000000000000_0000000000000000_0001010001010110_0000010101110010"; -- 0.07943758043276677
	pesos_i(16492) := b"1111111111111111_1111111111111111_1111101101110010_1110111001111110"; -- -0.017777532852775703
	pesos_i(16493) := b"0000000000000000_0000000000000000_0000100001000011_0110010110101010"; -- 0.032278398461088986
	pesos_i(16494) := b"1111111111111111_1111111111111111_1110110001100010_1001111100111111"; -- -0.07662014682910204
	pesos_i(16495) := b"0000000000000000_0000000000000000_0000100101111100_1001111110000101"; -- 0.03705784805553125
	pesos_i(16496) := b"0000000000000000_0000000000000000_0000001010001000_1101111110010010"; -- 0.009901021080753443
	pesos_i(16497) := b"1111111111111111_1111111111111111_1101011111100000_1111001111010110"; -- -0.15672374750687915
	pesos_i(16498) := b"1111111111111111_1111111111111111_1110100101010011_1110110100011101"; -- -0.08856313741488417
	pesos_i(16499) := b"1111111111111111_1111111111111111_1101100011001011_0111000011010101"; -- -0.15314574048354915
	pesos_i(16500) := b"0000000000000000_0000000000000000_0000011010011000_0100111111110011"; -- 0.025761601224312106
	pesos_i(16501) := b"1111111111111111_1111111111111111_1101111111010011_1100100001000010"; -- -0.12567470909613226
	pesos_i(16502) := b"0000000000000000_0000000000000000_0000000111110011_0111001000111011"; -- 0.007620944352965608
	pesos_i(16503) := b"0000000000000000_0000000000000000_0000100001010100_1011011101000101"; -- 0.03254266189627683
	pesos_i(16504) := b"1111111111111111_1111111111111111_1111100010101110_0111110001111110"; -- -0.028587550403772734
	pesos_i(16505) := b"0000000000000000_0000000000000000_0001110010000000_1100011111111110"; -- 0.11134004540953957
	pesos_i(16506) := b"0000000000000000_0000000000000000_0001001100000010_1011100101000000"; -- 0.07426030931245235
	pesos_i(16507) := b"1111111111111111_1111111111111111_1111000110101100_1000001010111011"; -- -0.055961446090137534
	pesos_i(16508) := b"0000000000000000_0000000000000000_0001010000101101_0011111101111011"; -- 0.07881542928831142
	pesos_i(16509) := b"0000000000000000_0000000000000000_0010000011110100_0010010111101100"; -- 0.12872540483656436
	pesos_i(16510) := b"1111111111111111_1111111111111111_1111100000100011_0110111101000010"; -- -0.030709310804422376
	pesos_i(16511) := b"1111111111111111_1111111111111111_1111110100100110_0011011001100111"; -- -0.011135673403533549
	pesos_i(16512) := b"0000000000000000_0000000000000000_0000001001001010_1010101001100001"; -- 0.008951805810678065
	pesos_i(16513) := b"1111111111111111_1111111111111111_1111011110101111_0010011010011101"; -- -0.032483660281325655
	pesos_i(16514) := b"0000000000000000_0000000000000000_0001100001101011_0000001100101001"; -- 0.09538287867329273
	pesos_i(16515) := b"0000000000000000_0000000000000000_0010010110000011_0011001100100010"; -- 0.14653319913805243
	pesos_i(16516) := b"0000000000000000_0000000000000000_0000110000111101_0001011000110010"; -- 0.04780710916114401
	pesos_i(16517) := b"0000000000000000_0000000000000000_0001100000100100_1111011101010001"; -- 0.09431405772527877
	pesos_i(16518) := b"1111111111111111_1111111111111111_1110010011111100_1010111101100011"; -- -0.1055193312565093
	pesos_i(16519) := b"0000000000000000_0000000000000000_0000010010011100_1000011001000000"; -- 0.01801337303069122
	pesos_i(16520) := b"0000000000000000_0000000000000000_0001111010010000_0100010000101100"; -- 0.11938882888918759
	pesos_i(16521) := b"1111111111111111_1111111111111111_1111001010001110_0000010001101111"; -- -0.052520487584578904
	pesos_i(16522) := b"1111111111111111_1111111111111111_1111011100001110_1001110000100001"; -- -0.03493332095587575
	pesos_i(16523) := b"0000000000000000_0000000000000000_0000011100100001_1110101001001010"; -- 0.027861254836272196
	pesos_i(16524) := b"0000000000000000_0000000000000000_0001001100011111_0111010010110111"; -- 0.07469872921822042
	pesos_i(16525) := b"1111111111111111_1111111111111111_1111110111100110_1110110101110001"; -- -0.008195075820555378
	pesos_i(16526) := b"0000000000000000_0000000000000000_0010011110101000_0101100010001000"; -- 0.15491250334112183
	pesos_i(16527) := b"1111111111111111_1111111111111111_1111111011100010_0100110011101110"; -- -0.00435942828333195
	pesos_i(16528) := b"1111111111111111_1111111111111111_1101111000011110_0111100110011011"; -- -0.13234748807171637
	pesos_i(16529) := b"0000000000000000_0000000000000000_0001010111011011_1100010110011000"; -- 0.0853847022397815
	pesos_i(16530) := b"0000000000000000_0000000000000000_0001010101000010_1100011101000101"; -- 0.08305020753508849
	pesos_i(16531) := b"0000000000000000_0000000000000000_0001010111101001_0001011001000100"; -- 0.08558787497080976
	pesos_i(16532) := b"1111111111111111_1111111111111111_1110111010010000_1100001111110011"; -- -0.06810355478474106
	pesos_i(16533) := b"0000000000000000_0000000000000000_0000000111010111_1101101010111101"; -- 0.007199927397305195
	pesos_i(16534) := b"1111111111111111_1111111111111111_1111001010111110_0010000101011001"; -- -0.05178634231759164
	pesos_i(16535) := b"1111111111111111_1111111111111111_1111111110000101_1111000111001000"; -- -0.0018624196664419692
	pesos_i(16536) := b"0000000000000000_0000000000000000_0010011111010111_1110110101000011"; -- 0.15563853149928208
	pesos_i(16537) := b"1111111111111111_1111111111111111_1110101111100101_1011000011000010"; -- -0.07852645178463546
	pesos_i(16538) := b"0000000000000000_0000000000000000_0001010101011011_0001001100010001"; -- 0.08342093614499212
	pesos_i(16539) := b"1111111111111111_1111111111111111_1111110101110111_1011110000110001"; -- -0.009891737115399174
	pesos_i(16540) := b"0000000000000000_0000000000000000_0000001111001010_1000000011111111"; -- 0.014808714138297626
	pesos_i(16541) := b"1111111111111111_1111111111111111_1101111001100111_1011110100011111"; -- -0.1312295722171385
	pesos_i(16542) := b"1111111111111111_1111111111111111_1110111011111010_0001110110110001"; -- -0.06649603292410847
	pesos_i(16543) := b"0000000000000000_0000000000000000_0001111100011110_1111001001001010"; -- 0.12156595533579964
	pesos_i(16544) := b"0000000000000000_0000000000000000_0001101001100101_0001010001001100"; -- 0.10310484739105223
	pesos_i(16545) := b"0000000000000000_0000000000000000_0010001111110111_1011100110111001"; -- 0.14049874083169528
	pesos_i(16546) := b"0000000000000000_0000000000000000_0000111011111111_1100110011001010"; -- 0.05859069755645005
	pesos_i(16547) := b"0000000000000000_0000000000000000_0001110000001111_0111011001101100"; -- 0.10961094034642634
	pesos_i(16548) := b"1111111111111111_1111111111111111_1111111100011101_1101100001000100"; -- -0.0034508545734727876
	pesos_i(16549) := b"1111111111111111_1111111111111111_1111100101110001_1110100110100100"; -- -0.025605580801567454
	pesos_i(16550) := b"0000000000000000_0000000000000000_0000110110000000_0111011000101011"; -- 0.05274141824647413
	pesos_i(16551) := b"0000000000000000_0000000000000000_0001100000011011_1010010100101000"; -- 0.09417183136386172
	pesos_i(16552) := b"0000000000000000_0000000000000000_0001011010010111_1010110110101100"; -- 0.08825192869162987
	pesos_i(16553) := b"0000000000000000_0000000000000000_0001101100110000_0101000111000110"; -- 0.10620604596576964
	pesos_i(16554) := b"1111111111111111_1111111111111111_1110110010000001_1111000110111101"; -- -0.0761422075033188
	pesos_i(16555) := b"0000000000000000_0000000000000000_0010001000010111_1110011000001100"; -- 0.13317716410065591
	pesos_i(16556) := b"1111111111111111_1111111111111111_1111001011000001_0100000100100100"; -- -0.05173867100185079
	pesos_i(16557) := b"0000000000000000_0000000000000000_0000111111110111_0011000010001011"; -- 0.06236556422154187
	pesos_i(16558) := b"0000000000000000_0000000000000000_0001011010001001_0101010111111000"; -- 0.08803307819417162
	pesos_i(16559) := b"1111111111111111_1111111111111111_1111110100101001_1001110110101101"; -- -0.011083741339130251
	pesos_i(16560) := b"1111111111111111_1111111111111111_1110101001110101_0100011010111101"; -- -0.08414800526044178
	pesos_i(16561) := b"0000000000000000_0000000000000000_0001010001101101_0111010101111010"; -- 0.0797952101413627
	pesos_i(16562) := b"0000000000000000_0000000000000000_0000000001101011_0010011011101011"; -- 0.0016350100584820815
	pesos_i(16563) := b"0000000000000000_0000000000000000_0000011001011011_1100101000010111"; -- 0.0248380953298739
	pesos_i(16564) := b"0000000000000000_0000000000000000_0000101101100001_1001100101101010"; -- 0.04445799671565839
	pesos_i(16565) := b"0000000000000000_0000000000000000_0000110011010000_0010001100101101"; -- 0.05005092479576497
	pesos_i(16566) := b"0000000000000000_0000000000000000_0001110000111101_1000101101011101"; -- 0.1103140928596361
	pesos_i(16567) := b"1111111111111111_1111111111111111_1110001111101011_0011011110110011"; -- -0.10969211468809188
	pesos_i(16568) := b"1111111111111111_1111111111111111_1110001001100111_1011100110001110"; -- -0.11560478487134361
	pesos_i(16569) := b"1111111111111111_1111111111111111_1111000111011100_0110101101011111"; -- -0.05523041663700978
	pesos_i(16570) := b"1111111111111111_1111111111111111_1101110111001010_1011101111011011"; -- -0.13362527758535797
	pesos_i(16571) := b"1111111111111111_1111111111111111_1111000001001000_0000010001001001"; -- -0.06140111177150397
	pesos_i(16572) := b"0000000000000000_0000000000000000_0000111011111001_0101110110101101"; -- 0.05849252207958135
	pesos_i(16573) := b"0000000000000000_0000000000000000_0000100010110000_1001111010010110"; -- 0.033944999418064205
	pesos_i(16574) := b"1111111111111111_1111111111111111_1110010011001101_1111011111000001"; -- -0.10623218095352717
	pesos_i(16575) := b"1111111111111111_1111111111111111_1110101010001000_1000001100000100"; -- -0.08385449543618598
	pesos_i(16576) := b"1111111111111111_1111111111111111_1101111100001111_1001101101101111"; -- -0.1286681034944667
	pesos_i(16577) := b"0000000000000000_0000000000000000_0001010110100001_1011110001001010"; -- 0.08449913791767322
	pesos_i(16578) := b"1111111111111111_1111111111111111_1110010101111110_1001000110011100"; -- -0.1035374635726661
	pesos_i(16579) := b"0000000000000000_0000000000000000_0001001100101110_1000000110011111"; -- 0.07492838041592041
	pesos_i(16580) := b"1111111111111111_1111111111111111_1110010111000110_0100011100101101"; -- -0.10244326735222616
	pesos_i(16581) := b"0000000000000000_0000000000000000_0000111011101100_0110001010000010"; -- 0.058294445691348624
	pesos_i(16582) := b"0000000000000000_0000000000000000_0001101111001100_0001011100101000"; -- 0.10858292325528986
	pesos_i(16583) := b"1111111111111111_1111111111111111_1101111001111110_0000101001110110"; -- -0.13088926906830886
	pesos_i(16584) := b"0000000000000000_0000000000000000_0000001101111100_1000100000101001"; -- 0.013618955729194639
	pesos_i(16585) := b"1111111111111111_1111111111111111_1111110000001101_0010110110001100"; -- -0.015423920843697203
	pesos_i(16586) := b"1111111111111111_1111111111111111_1111001111000011_0010100001110001"; -- -0.04780337563520218
	pesos_i(16587) := b"1111111111111111_1111111111111111_1110111011011011_0101000101000111"; -- -0.06696598069824772
	pesos_i(16588) := b"1111111111111111_1111111111111111_1101110011010010_0001001001010000"; -- -0.13741956280572315
	pesos_i(16589) := b"1111111111111111_1111111111111111_1111111111111010_0111011111110101"; -- -8.440283900771336e-05
	pesos_i(16590) := b"1111111111111111_1111111111111111_1111110110001111_1110011010110101"; -- -0.009522991988980838
	pesos_i(16591) := b"0000000000000000_0000000000000000_0000001111010110_0010101000010100"; -- 0.01498663883265419
	pesos_i(16592) := b"0000000000000000_0000000000000000_0010010000011110_0001110111001001"; -- 0.14108453900806295
	pesos_i(16593) := b"0000000000000000_0000000000000000_0000101010110111_0101000001110000"; -- 0.041859652772205526
	pesos_i(16594) := b"1111111111111111_1111111111111111_1110010100010101_1110101100100101"; -- -0.1051342997353098
	pesos_i(16595) := b"1111111111111111_1111111111111111_1101110001111001_1100010110010000"; -- -0.13876691097325122
	pesos_i(16596) := b"0000000000000000_0000000000000000_0001000100101110_0010101001111110"; -- 0.0671106870857825
	pesos_i(16597) := b"0000000000000000_0000000000000000_0001010100011001_0110101101111110"; -- 0.08241912672504026
	pesos_i(16598) := b"1111111111111111_1111111111111111_1111000011101111_1001011101111110"; -- -0.058844119844420416
	pesos_i(16599) := b"1111111111111111_1111111111111111_1101110010110011_0001011110110101"; -- -0.1378922637976879
	pesos_i(16600) := b"1111111111111111_1111111111111111_1110011011110111_0001010001000111"; -- -0.09779237048538408
	pesos_i(16601) := b"0000000000000000_0000000000000000_0000111111010011_1110101111111001"; -- 0.06182741953511684
	pesos_i(16602) := b"0000000000000000_0000000000000000_0010000001000110_0010110011100001"; -- 0.12607079021864118
	pesos_i(16603) := b"1111111111111111_1111111111111111_1111100100100010_1100110111100011"; -- -0.02681267929218331
	pesos_i(16604) := b"0000000000000000_0000000000000000_0001111101010111_0001001000001111"; -- 0.12242234099348095
	pesos_i(16605) := b"0000000000000000_0000000000000000_0001001100000011_1001100101111010"; -- 0.0742736743751958
	pesos_i(16606) := b"0000000000000000_0000000000000000_0010010101101101_0101101001000011"; -- 0.14619983801291078
	pesos_i(16607) := b"1111111111111111_1111111111111111_1111010001000011_1100001001111101"; -- -0.04584106876058541
	pesos_i(16608) := b"1111111111111111_1111111111111111_1110000101111110_1100001101001010"; -- -0.11915950232666335
	pesos_i(16609) := b"0000000000000000_0000000000000000_0001011011010010_0101001001111110"; -- 0.08914676253178473
	pesos_i(16610) := b"0000000000000000_0000000000000000_0001011010100011_0100001101011000"; -- 0.08842869667430306
	pesos_i(16611) := b"0000000000000000_0000000000000000_0000111110101100_1111100001100000"; -- 0.06123306593378517
	pesos_i(16612) := b"0000000000000000_0000000000000000_0001010111010000_1001110010010101"; -- 0.08521441107243978
	pesos_i(16613) := b"1111111111111111_1111111111111111_1111100001000100_1101011000110001"; -- -0.03019963563013639
	pesos_i(16614) := b"0000000000000000_0000000000000000_0010001101000000_0000000111100011"; -- 0.13769542491529482
	pesos_i(16615) := b"1111111111111111_1111111111111111_1110000101111001_0111001001110110"; -- -0.11924061419228173
	pesos_i(16616) := b"1111111111111111_1111111111111111_1110111100111001_0101000100000110"; -- -0.06553166960674717
	pesos_i(16617) := b"1111111111111111_1111111111111111_1101111010100111_0101100011000111"; -- -0.13025899079842118
	pesos_i(16618) := b"1111111111111111_1111111111111111_1111100000111100_1010110110100101"; -- -0.03032412267105981
	pesos_i(16619) := b"0000000000000000_0000000000000000_0000100111000110_1111000110100000"; -- 0.03819189223706566
	pesos_i(16620) := b"1111111111111111_1111111111111111_1110100100101000_1110111100011000"; -- -0.08921914737517789
	pesos_i(16621) := b"0000000000000000_0000000000000000_0001000001010111_1111011000011010"; -- 0.06384218350713441
	pesos_i(16622) := b"1111111111111111_1111111111111111_1101111111001010_1100010100101101"; -- -0.12581222208677456
	pesos_i(16623) := b"0000000000000000_0000000000000000_0000101111111000_0000000101111110"; -- 0.0467530186511631
	pesos_i(16624) := b"1111111111111111_1111111111111111_1110011111111010_0000111000110101"; -- -0.09384070592417172
	pesos_i(16625) := b"1111111111111111_1111111111111111_1101111101000001_1011100011101000"; -- -0.12790340743410664
	pesos_i(16626) := b"1111111111111111_1111111111111111_1110011011001010_0100110001000111"; -- -0.09847567808630225
	pesos_i(16627) := b"1111111111111111_1111111111111111_1101111100100101_1010011010010000"; -- -0.1283317469006575
	pesos_i(16628) := b"0000000000000000_0000000000000000_0001010010001010_0100000101010111"; -- 0.08023460746029668
	pesos_i(16629) := b"1111111111111111_1111111111111111_1110001011001010_0111001110011111"; -- -0.11409833315954443
	pesos_i(16630) := b"0000000000000000_0000000000000000_0000011111000000_0111110001001000"; -- 0.03028084524000876
	pesos_i(16631) := b"0000000000000000_0000000000000000_0010010101000001_1010011001010000"; -- 0.14553298432720685
	pesos_i(16632) := b"0000000000000000_0000000000000000_0000010111001011_0001101110101010"; -- 0.022630433150909447
	pesos_i(16633) := b"1111111111111111_1111111111111111_1111111010101000_0100010111101111"; -- -0.005244855059880464
	pesos_i(16634) := b"1111111111111111_1111111111111111_1111101011011111_0000111110000101"; -- -0.020033864897450238
	pesos_i(16635) := b"1111111111111111_1111111111111111_1111001001101011_0001001011011000"; -- -0.05305368635030951
	pesos_i(16636) := b"0000000000000000_0000000000000000_0000110000010100_0101111111110010"; -- 0.04718589455993841
	pesos_i(16637) := b"1111111111111111_1111111111111111_1111100010100010_1100101111011001"; -- -0.028765925988933214
	pesos_i(16638) := b"1111111111111111_1111111111111111_1111000100011010_1001001101011000"; -- -0.05818823920435211
	pesos_i(16639) := b"0000000000000000_0000000000000000_0010000010000001_1101100101100000"; -- 0.1269813403944699
	pesos_i(16640) := b"0000000000000000_0000000000000000_0000001110010001_0111100110000111"; -- 0.013938518122361705
	pesos_i(16641) := b"0000000000000000_0000000000000000_0001100110000111_0001101111101110"; -- 0.09971785117600349
	pesos_i(16642) := b"1111111111111111_1111111111111111_1110101101110000_0101000110001111"; -- -0.0803174042606179
	pesos_i(16643) := b"0000000000000000_0000000000000000_0000111111001010_0100010100001101"; -- 0.0616801410435471
	pesos_i(16644) := b"1111111111111111_1111111111111111_1110101010101111_1000110000100011"; -- -0.08325885915763274
	pesos_i(16645) := b"1111111111111111_1111111111111111_1111111101100001_0101110111111011"; -- -0.0024205458777468453
	pesos_i(16646) := b"0000000000000000_0000000000000000_0001100000011011_0001110100000000"; -- 0.09416371595329448
	pesos_i(16647) := b"0000000000000000_0000000000000000_0010010111011100_0111001110110011"; -- 0.1478950798814405
	pesos_i(16648) := b"0000000000000000_0000000000000000_0000011010010000_1101101000011001"; -- 0.025647765187038755
	pesos_i(16649) := b"0000000000000000_0000000000000000_0000010100010010_1111110010001101"; -- 0.01982096134944849
	pesos_i(16650) := b"0000000000000000_0000000000000000_0001100010000000_1101101000010111"; -- 0.0957161242122128
	pesos_i(16651) := b"1111111111111111_1111111111111111_1111001000110111_1011011111010111"; -- -0.05383730881819231
	pesos_i(16652) := b"1111111111111111_1111111111111111_1111111001100110_1010100000101110"; -- -0.006246079181317853
	pesos_i(16653) := b"1111111111111111_1111111111111111_1110010001111111_1101111110001101"; -- -0.1074238091109676
	pesos_i(16654) := b"0000000000000000_0000000000000000_0000001110010111_0001000010010110"; -- 0.014023815680041013
	pesos_i(16655) := b"1111111111111111_1111111111111111_1110110101110111_1001011000111000"; -- -0.07239400025957995
	pesos_i(16656) := b"1111111111111111_1111111111111111_1110011101100101_1100101110100111"; -- -0.09610297362277731
	pesos_i(16657) := b"0000000000000000_0000000000000000_0001010110001101_1011110001001001"; -- 0.0841939619943664
	pesos_i(16658) := b"0000000000000000_0000000000000000_0001101011010111_1011100011000111"; -- 0.10485415316564824
	pesos_i(16659) := b"0000000000000000_0000000000000000_0001101101111101_0111100010100101"; -- 0.10738328953467188
	pesos_i(16660) := b"1111111111111111_1111111111111111_1110011010111000_0110000101110010"; -- -0.09874907463662438
	pesos_i(16661) := b"1111111111111111_1111111111111111_1111001110001101_0110001111110111"; -- -0.048623802269152146
	pesos_i(16662) := b"0000000000000000_0000000000000000_0000010010001110_0101000100000100"; -- 0.01779657699308362
	pesos_i(16663) := b"0000000000000000_0000000000000000_0000011110010010_1000001011101110"; -- 0.029579337175990966
	pesos_i(16664) := b"1111111111111111_1111111111111111_1111100100000101_0110010101011100"; -- -0.027261414623218176
	pesos_i(16665) := b"0000000000000000_0000000000000000_0001010001001010_1101000010101100"; -- 0.07926658809694699
	pesos_i(16666) := b"0000000000000000_0000000000000000_0010010001101111_1111110010111111"; -- 0.14233379051767475
	pesos_i(16667) := b"1111111111111111_1111111111111111_1111101010101001_1110100111100010"; -- -0.02084482404556332
	pesos_i(16668) := b"0000000000000000_0000000000000000_0000001111101011_1101101000101111"; -- 0.015317570291230766
	pesos_i(16669) := b"1111111111111111_1111111111111111_1101100111010111_1011011001000000"; -- -0.1490522473575045
	pesos_i(16670) := b"0000000000000000_0000000000000000_0010000000101011_0101011110100100"; -- 0.1256613517196701
	pesos_i(16671) := b"1111111111111111_1111111111111111_1111000011000101_1101000101000011"; -- -0.059481545655017176
	pesos_i(16672) := b"0000000000000000_0000000000000000_0000101011001100_1100101000010000"; -- 0.04218733684295077
	pesos_i(16673) := b"0000000000000000_0000000000000000_0001011001110010_0011111111011100"; -- 0.08768080818152965
	pesos_i(16674) := b"1111111111111111_1111111111111111_1110101010001101_1011100100100110"; -- -0.0837749750499343
	pesos_i(16675) := b"0000000000000000_0000000000000000_0000101010010000_1110111010001110"; -- 0.041273984666679184
	pesos_i(16676) := b"1111111111111111_1111111111111111_1101111100010111_1101110111100101"; -- -0.12854207181321328
	pesos_i(16677) := b"0000000000000000_0000000000000000_0001111010000100_1001011010100000"; -- 0.11921063819479369
	pesos_i(16678) := b"1111111111111111_1111111111111111_1110100101000000_0111101001000001"; -- -0.08885990065216373
	pesos_i(16679) := b"1111111111111111_1111111111111111_1111001000111100_1100010111111101"; -- -0.05376017165604605
	pesos_i(16680) := b"0000000000000000_0000000000000000_0000100011011001_1110100101000011"; -- 0.03457506080301115
	pesos_i(16681) := b"0000000000000000_0000000000000000_0000110101110110_1111101101111111"; -- 0.05259677749270661
	pesos_i(16682) := b"0000000000000000_0000000000000000_0000110100011110_1100000110010100"; -- 0.05125055174987395
	pesos_i(16683) := b"0000000000000000_0000000000000000_0010010001000001_1111101000111110"; -- 0.1416317368418296
	pesos_i(16684) := b"0000000000000000_0000000000000000_0000001100000111_0111101001000101"; -- 0.011832849240818259
	pesos_i(16685) := b"1111111111111111_1111111111111111_1111001011100001_1101001110011100"; -- -0.051241659490746994
	pesos_i(16686) := b"1111111111111111_1111111111111111_1101101100101000_1000010111100010"; -- -0.14391291829439176
	pesos_i(16687) := b"1111111111111111_1111111111111111_1110001100010100_1000010000101111"; -- -0.11296819535477429
	pesos_i(16688) := b"1111111111111111_1111111111111111_1101110000100000_0111111101000001"; -- -0.14012913393565513
	pesos_i(16689) := b"1111111111111111_1111111111111111_1110000110101111_0001101110001011"; -- -0.11842182015639598
	pesos_i(16690) := b"1111111111111111_1111111111111111_1111001111101111_1001001001000010"; -- -0.04712568167918407
	pesos_i(16691) := b"0000000000000000_0000000000000000_0001011111101111_0110110011011000"; -- 0.09349708824445949
	pesos_i(16692) := b"1111111111111111_1111111111111111_1111000000010010_1100010001010110"; -- -0.0622136392386782
	pesos_i(16693) := b"1111111111111111_1111111111111111_1111011111110011_1010101000110111"; -- -0.03143821855692268
	pesos_i(16694) := b"1111111111111111_1111111111111111_1110011010001001_1101001011011000"; -- -0.09945947852857291
	pesos_i(16695) := b"1111111111111111_1111111111111111_1110001001010010_0110111010000010"; -- -0.11592969243308089
	pesos_i(16696) := b"0000000000000000_0000000000000000_0000110111101000_1101010101110010"; -- 0.054334011353668436
	pesos_i(16697) := b"0000000000000000_0000000000000000_0001000100010111_1101010111000101"; -- 0.0667699437099632
	pesos_i(16698) := b"0000000000000000_0000000000000000_0001100011010100_1010011010100001"; -- 0.09699479509750282
	pesos_i(16699) := b"1111111111111111_1111111111111111_1110101100000101_0010010010000111"; -- -0.08195277895444847
	pesos_i(16700) := b"1111111111111111_1111111111111111_1111000001110010_1110011110100010"; -- -0.060746691619813116
	pesos_i(16701) := b"0000000000000000_0000000000000000_0010011110100100_0000010011001001"; -- 0.15484647665803739
	pesos_i(16702) := b"0000000000000000_0000000000000000_0000110111101011_1111100101010111"; -- 0.05438192734854685
	pesos_i(16703) := b"0000000000000000_0000000000000000_0000111010101100_0010100011100111"; -- 0.05731444979815562
	pesos_i(16704) := b"0000000000000000_0000000000000000_0001101010010101_0000110011011010"; -- 0.10383682550223677
	pesos_i(16705) := b"1111111111111111_1111111111111111_1110001010111101_1001011101110010"; -- -0.1142945620646501
	pesos_i(16706) := b"1111111111111111_1111111111111111_1110111111111010_0001100100100100"; -- -0.0625900542153351
	pesos_i(16707) := b"1111111111111111_1111111111111111_1110101001010100_0000011000110101"; -- -0.08465539182186473
	pesos_i(16708) := b"1111111111111111_1111111111111111_1111100100001101_1101110000110101"; -- -0.02713226029802798
	pesos_i(16709) := b"0000000000000000_0000000000000000_0000100010110011_0101101000011000"; -- 0.03398669317600765
	pesos_i(16710) := b"0000000000000000_0000000000000000_0001001010101101_0100110110111110"; -- 0.07295690439104553
	pesos_i(16711) := b"1111111111111111_1111111111111111_1110001010000100_1010111100110101"; -- -0.11516289675939517
	pesos_i(16712) := b"0000000000000000_0000000000000000_0000111000100001_1110011111001000"; -- 0.055204855270658104
	pesos_i(16713) := b"0000000000000000_0000000000000000_0010001000101101_1111010000100011"; -- 0.13351369728535228
	pesos_i(16714) := b"0000000000000000_0000000000000000_0010001011111011_0111100110010101"; -- 0.1366497030074261
	pesos_i(16715) := b"0000000000000000_0000000000000000_0000010010111111_0100100101011110"; -- 0.01854380164271165
	pesos_i(16716) := b"1111111111111111_1111111111111111_1110111001011110_1100010001010100"; -- -0.06886647182140052
	pesos_i(16717) := b"1111111111111111_1111111111111111_1110011101100001_0100011111000010"; -- -0.09617187030582815
	pesos_i(16718) := b"1111111111111111_1111111111111111_1111011111011111_0100011000110000"; -- -0.03174935660017558
	pesos_i(16719) := b"0000000000000000_0000000000000000_0001111110011111_1110110110000010"; -- 0.12353405394308338
	pesos_i(16720) := b"0000000000000000_0000000000000000_0000001011001111_1110111110100011"; -- 0.01098535273810412
	pesos_i(16721) := b"0000000000000000_0000000000000000_0000100000011011_0001001000000001"; -- 0.031663060437128916
	pesos_i(16722) := b"0000000000000000_0000000000000000_0000110111110111_1111010011011110"; -- 0.054564766122990924
	pesos_i(16723) := b"1111111111111111_1111111111111111_1110011000001100_1010101100110100"; -- -0.10136919010415806
	pesos_i(16724) := b"0000000000000000_0000000000000000_0001010111001000_0011000011010110"; -- 0.08508591867274623
	pesos_i(16725) := b"0000000000000000_0000000000000000_0000101011010001_0000000001011010"; -- 0.042251607901390396
	pesos_i(16726) := b"1111111111111111_1111111111111111_1111000110000110_0010110110110111"; -- -0.05654634739155916
	pesos_i(16727) := b"1111111111111111_1111111111111111_1110101001000011_0110000000000110"; -- -0.08490943779829732
	pesos_i(16728) := b"1111111111111111_1111111111111111_1111101110010010_1110010010010001"; -- -0.0172898432671064
	pesos_i(16729) := b"1111111111111111_1111111111111111_1110110001100011_0011001000001000"; -- -0.07661139787982146
	pesos_i(16730) := b"0000000000000000_0000000000000000_0001011111100001_1010100000001001"; -- 0.09328699321530368
	pesos_i(16731) := b"0000000000000000_0000000000000000_0010011010000100_0000011110000100"; -- 0.15045210820927532
	pesos_i(16732) := b"1111111111111111_1111111111111111_1110001001110110_0100001101101000"; -- -0.11538294525079089
	pesos_i(16733) := b"1111111111111111_1111111111111111_1111010111110011_1100111001101000"; -- -0.039248561384004496
	pesos_i(16734) := b"0000000000000000_0000000000000000_0001011000101101_0111011010011110"; -- 0.0866312156034602
	pesos_i(16735) := b"1111111111111111_1111111111111111_1111011111010011_0100101000010011"; -- -0.03193223026398289
	pesos_i(16736) := b"0000000000000000_0000000000000000_0000001010111011_0111010001000010"; -- 0.010672823123393837
	pesos_i(16737) := b"0000000000000000_0000000000000000_0000000010010111_1011011000111100"; -- 0.002314939237999537
	pesos_i(16738) := b"1111111111111111_1111111111111111_1101111100010111_0101000010111111"; -- -0.12855048512159414
	pesos_i(16739) := b"0000000000000000_0000000000000000_0001011001110011_1101011000100110"; -- 0.08770502506756653
	pesos_i(16740) := b"1111111111111111_1111111111111111_1111100010111011_0111110000100000"; -- -0.028389207987520156
	pesos_i(16741) := b"1111111111111111_1111111111111111_1110000010100110_0000110000111001"; -- -0.12246631248524671
	pesos_i(16742) := b"0000000000000000_0000000000000000_0000110011111110_1010010111100111"; -- 0.050760621005646406
	pesos_i(16743) := b"0000000000000000_0000000000000000_0000001111011010_1001000011000100"; -- 0.015053794627444092
	pesos_i(16744) := b"1111111111111111_1111111111111111_1111000001111000_1011100111100101"; -- -0.06065786509839104
	pesos_i(16745) := b"1111111111111111_1111111111111111_1110000111100101_0011000101001001"; -- -0.11759654979278311
	pesos_i(16746) := b"1111111111111111_1111111111111111_1111100011110110_0011010100011110"; -- -0.02749317189441285
	pesos_i(16747) := b"0000000000000000_0000000000000000_0001010000111001_0010100110000101"; -- 0.07899722581955086
	pesos_i(16748) := b"1111111111111111_1111111111111111_1101100110111010_1110011000010011"; -- -0.14949190166759277
	pesos_i(16749) := b"0000000000000000_0000000000000000_0000010001110101_1100111010001000"; -- 0.01742258852200491
	pesos_i(16750) := b"0000000000000000_0000000000000000_0000000000001110_0110101110110001"; -- 0.00022004191857747895
	pesos_i(16751) := b"1111111111111111_1111111111111111_1111101011101000_0111101000010000"; -- -0.0198901854403685
	pesos_i(16752) := b"1111111111111111_1111111111111111_1111001111101100_0011001010101000"; -- -0.04717715640539689
	pesos_i(16753) := b"0000000000000000_0000000000000000_0001111001100110_0111000111110110"; -- 0.11875068919881507
	pesos_i(16754) := b"1111111111111111_1111111111111111_1101110010111110_0100001011101100"; -- -0.13772184114881172
	pesos_i(16755) := b"1111111111111111_1111111111111111_1111100001010110_1100010110011111"; -- -0.029925964939693746
	pesos_i(16756) := b"1111111111111111_1111111111111111_1101111111111010_0010010000101101"; -- -0.12508939647640216
	pesos_i(16757) := b"1111111111111111_1111111111111111_1111000100111111_1001010000010100"; -- -0.057623620109461766
	pesos_i(16758) := b"1111111111111111_1111111111111111_1111111001110010_0100100110010010"; -- -0.0060686129040827125
	pesos_i(16759) := b"0000000000000000_0000000000000000_0000011101100010_1111000110101101"; -- 0.02885351642787132
	pesos_i(16760) := b"1111111111111111_1111111111111111_1110110011011100_0110111010001100"; -- -0.07476147719812411
	pesos_i(16761) := b"1111111111111111_1111111111111111_1110111000111101_0010011010100100"; -- -0.06937941065221061
	pesos_i(16762) := b"0000000000000000_0000000000000000_0000011101101010_0111011001010111"; -- 0.028968235155879634
	pesos_i(16763) := b"0000000000000000_0000000000000000_0010000001101011_0001101011011110"; -- 0.1266342917712983
	pesos_i(16764) := b"1111111111111111_1111111111111111_1110011000000100_0001111111011100"; -- -0.10149956593600623
	pesos_i(16765) := b"0000000000000000_0000000000000000_0000000010100011_0100011111000101"; -- 0.002491460364506781
	pesos_i(16766) := b"1111111111111111_1111111111111111_1111011101111010_0101110110100011"; -- -0.033289096518786546
	pesos_i(16767) := b"1111111111111111_1111111111111111_1110000000110010_1011101001001000"; -- -0.12422595736026247
	pesos_i(16768) := b"0000000000000000_0000000000000000_0010010010001110_1011110110101110"; -- 0.14280305377739608
	pesos_i(16769) := b"0000000000000000_0000000000000000_0000001101110111_0100000111110010"; -- 0.013538476454005221
	pesos_i(16770) := b"0000000000000000_0000000000000000_0001000000011110_0110000100101100"; -- 0.06296355555586287
	pesos_i(16771) := b"1111111111111111_1111111111111111_1110011110011101_1011011101000001"; -- -0.09524969737605624
	pesos_i(16772) := b"0000000000000000_0000000000000000_0001001110000101_1101011100100010"; -- 0.0762609917594397
	pesos_i(16773) := b"0000000000000000_0000000000000000_0010000111101101_0000010101000100"; -- 0.13252289686273688
	pesos_i(16774) := b"0000000000000000_0000000000000000_0010010100111011_0111010111010001"; -- 0.14543854105317522
	pesos_i(16775) := b"1111111111111111_1111111111111111_1111101011001011_1111000110010010"; -- -0.020325567208037985
	pesos_i(16776) := b"0000000000000000_0000000000000000_0000000111001001_1011011101001010"; -- 0.00698419143471517
	pesos_i(16777) := b"0000000000000000_0000000000000000_0010001110010001_1111010001100100"; -- 0.13894584131440918
	pesos_i(16778) := b"1111111111111111_1111111111111111_1111011010011001_0001011111001110"; -- -0.03672648640485824
	pesos_i(16779) := b"1111111111111111_1111111111111111_1110100001001110_0111111010110110"; -- -0.0925522619042066
	pesos_i(16780) := b"0000000000000000_0000000000000000_0001000111000101_1110101000100100"; -- 0.06942618734622041
	pesos_i(16781) := b"0000000000000000_0000000000000000_0000000100101101_0011100010100110"; -- 0.0045962719161416745
	pesos_i(16782) := b"1111111111111111_1111111111111111_1101101101100000_1110110011100111"; -- -0.1430522857774825
	pesos_i(16783) := b"0000000000000000_0000000000000000_0001111100000101_0111110000111101"; -- 0.12117744913308343
	pesos_i(16784) := b"0000000000000000_0000000000000000_0001001101001011_1101010110000110"; -- 0.07537588623579433
	pesos_i(16785) := b"1111111111111111_1111111111111111_1110100100011101_0111000111010011"; -- -0.08939446061587167
	pesos_i(16786) := b"1111111111111111_1111111111111111_1110001101111100_1111011110100001"; -- -0.11137440029853442
	pesos_i(16787) := b"1111111111111111_1111111111111111_1101101100001111_1001011011111010"; -- -0.144293369227393
	pesos_i(16788) := b"0000000000000000_0000000000000000_0001001100100100_1110011100101001"; -- 0.07478184459363128
	pesos_i(16789) := b"0000000000000000_0000000000000000_0001001000011001_0111001100101001"; -- 0.07070083369322376
	pesos_i(16790) := b"1111111111111111_1111111111111111_1111010101111001_1110110001101000"; -- -0.04110834557520032
	pesos_i(16791) := b"1111111111111111_1111111111111111_1110111101101110_1110100111010101"; -- -0.06471384580025549
	pesos_i(16792) := b"1111111111111111_1111111111111111_1111001100101011_0101001101101101"; -- -0.05012014943455583
	pesos_i(16793) := b"0000000000000000_0000000000000000_0000101010001101_0111010000101100"; -- 0.04122091358180004
	pesos_i(16794) := b"1111111111111111_1111111111111111_1110101110010110_1111011010101000"; -- -0.07972772977274499
	pesos_i(16795) := b"0000000000000000_0000000000000000_0000011000000101_1110100100011111"; -- 0.023527688996650864
	pesos_i(16796) := b"0000000000000000_0000000000000000_0001101110010101_1010000101111000"; -- 0.10775193391497413
	pesos_i(16797) := b"1111111111111111_1111111111111111_1110101001010001_0100100010111010"; -- -0.08469720335920736
	pesos_i(16798) := b"0000000000000000_0000000000000000_0001001101000001_1110101101000001"; -- 0.07522459344592823
	pesos_i(16799) := b"0000000000000000_0000000000000000_0001110111111010_1000011110001100"; -- 0.1171040265430849
	pesos_i(16800) := b"1111111111111111_1111111111111111_1110000001100001_1110010010011110"; -- -0.1235062708406582
	pesos_i(16801) := b"0000000000000000_0000000000000000_0001001010101110_0100101010001000"; -- 0.07297197175052494
	pesos_i(16802) := b"1111111111111111_1111111111111111_1110101000001101_0010111000010011"; -- -0.08573638954040279
	pesos_i(16803) := b"1111111111111111_1111111111111111_1111101000000001_1111101110111101"; -- -0.023407236424431193
	pesos_i(16804) := b"0000000000000000_0000000000000000_0000000010000011_1110011110111110"; -- 0.002012714270234442
	pesos_i(16805) := b"0000000000000000_0000000000000000_0010000010101100_0100101111110100"; -- 0.12762903884998292
	pesos_i(16806) := b"0000000000000000_0000000000000000_0001000100010010_0011101101000111"; -- 0.06668444143603876
	pesos_i(16807) := b"1111111111111111_1111111111111111_1101101010110100_0110000000001110"; -- -0.14568519266187052
	pesos_i(16808) := b"1111111111111111_1111111111111111_1111001010101110_0111010011001001"; -- -0.05202550982315749
	pesos_i(16809) := b"1111111111111111_1111111111111111_1111000000011111_1000111100111111"; -- -0.062018439427317
	pesos_i(16810) := b"0000000000000000_0000000000000000_0010001110100100_1000000000100110"; -- 0.13922882953463567
	pesos_i(16811) := b"1111111111111111_1111111111111111_1101111000101110_0101010001000100"; -- -0.13210557319334568
	pesos_i(16812) := b"1111111111111111_1111111111111111_1101101010111111_1010000001000111"; -- -0.1455135180756449
	pesos_i(16813) := b"0000000000000000_0000000000000000_0001111101100110_1101101010101001"; -- 0.12266317959729224
	pesos_i(16814) := b"0000000000000000_0000000000000000_0010000000111111_1011100001000101"; -- 0.12597228699150168
	pesos_i(16815) := b"1111111111111111_1111111111111111_1110010111000100_1011000010011111"; -- -0.10246749998774801
	pesos_i(16816) := b"1111111111111111_1111111111111111_1110000000101011_0001010001011111"; -- -0.12434265796940676
	pesos_i(16817) := b"1111111111111111_1111111111111111_1110001010100010_1011100011111110"; -- -0.1147045497214576
	pesos_i(16818) := b"1111111111111111_1111111111111111_1110101001101110_0011000111110110"; -- -0.0842560553722108
	pesos_i(16819) := b"0000000000000000_0000000000000000_0001100011111010_0110010110101000"; -- 0.09757075645402057
	pesos_i(16820) := b"0000000000000000_0000000000000000_0000010111100110_1110110001010010"; -- 0.023054857240532477
	pesos_i(16821) := b"1111111111111111_1111111111111111_1111011111100001_0011110001000111"; -- -0.031719429595662464
	pesos_i(16822) := b"0000000000000000_0000000000000000_0001101111100100_0101101101010001"; -- 0.10895319675300032
	pesos_i(16823) := b"1111111111111111_1111111111111111_1111110010101001_1001111000010111"; -- -0.013036841851761407
	pesos_i(16824) := b"1111111111111111_1111111111111111_1101111110010001_1100000011010011"; -- -0.12668223247458632
	pesos_i(16825) := b"0000000000000000_0000000000000000_0001011000011011_1100000110010111"; -- 0.08636102614256465
	pesos_i(16826) := b"0000000000000000_0000000000000000_0000011001110000_0011111000111101"; -- 0.02515019400599065
	pesos_i(16827) := b"1111111111111111_1111111111111111_1111011111100111_0001011001100010"; -- -0.031630135575315764
	pesos_i(16828) := b"0000000000000000_0000000000000000_0000010101001001_1011100101011011"; -- 0.020656189558601226
	pesos_i(16829) := b"0000000000000000_0000000000000000_0000001100101001_1010100011100011"; -- 0.012354426836908612
	pesos_i(16830) := b"0000000000000000_0000000000000000_0010010101011100_1110101001111001"; -- 0.14594903420982389
	pesos_i(16831) := b"0000000000000000_0000000000000000_0000000110011110_1010110010101101"; -- 0.006327431059457497
	pesos_i(16832) := b"1111111111111111_1111111111111111_1110101000001001_0110101010011100"; -- -0.08579381643627303
	pesos_i(16833) := b"0000000000000000_0000000000000000_0000111110100000_1001001110011001"; -- 0.061043953768204956
	pesos_i(16834) := b"0000000000000000_0000000000000000_0001111000001000_1001101001000101"; -- 0.11731876545736415
	pesos_i(16835) := b"1111111111111111_1111111111111111_1110101111100011_1101001100010001"; -- -0.07855492444365944
	pesos_i(16836) := b"1111111111111111_1111111111111111_1110011111011111_1010001110000101"; -- -0.09424379346633581
	pesos_i(16837) := b"0000000000000000_0000000000000000_0000010010010000_0010001110010011"; -- 0.017824385898246906
	pesos_i(16838) := b"0000000000000000_0000000000000000_0000010011000011_1000111111001010"; -- 0.018609034452555823
	pesos_i(16839) := b"0000000000000000_0000000000000000_0001011111110111_0011110010101110"; -- 0.09361628773493663
	pesos_i(16840) := b"0000000000000000_0000000000000000_0001001111111000_0001000110111111"; -- 0.0780039874108931
	pesos_i(16841) := b"0000000000000000_0000000000000000_0000100000110100_0111110001111100"; -- 0.03205087683720155
	pesos_i(16842) := b"1111111111111111_1111111111111111_1111001000000010_0100010100110110"; -- -0.0546528570493533
	pesos_i(16843) := b"1111111111111111_1111111111111111_1110011101011110_1010111101101111"; -- -0.09621146708080199
	pesos_i(16844) := b"0000000000000000_0000000000000000_0000001011011111_0000110000110101"; -- 0.011215937495888341
	pesos_i(16845) := b"0000000000000000_0000000000000000_0001011111000100_0100101110100100"; -- 0.09283898127526492
	pesos_i(16846) := b"1111111111111111_1111111111111111_1110101100111110_0001011000111111"; -- -0.08108387908674786
	pesos_i(16847) := b"1111111111111111_1111111111111111_1111011010001010_1110011101100111"; -- -0.03694299434160009
	pesos_i(16848) := b"1111111111111111_1111111111111111_1111001001010110_0011110111000010"; -- -0.05337156301580399
	pesos_i(16849) := b"0000000000000000_0000000000000000_0000101011101001_0111001110011001"; -- 0.04262468811102447
	pesos_i(16850) := b"0000000000000000_0000000000000000_0010010000100000_0101111000110001"; -- 0.1411188954315163
	pesos_i(16851) := b"0000000000000000_0000000000000000_0010010011101110_1011000100000010"; -- 0.1442671423547615
	pesos_i(16852) := b"1111111111111111_1111111111111111_1111111011001010_0010101100111100"; -- -0.004727647735382684
	pesos_i(16853) := b"1111111111111111_1111111111111111_1101110101101101_1010000100011001"; -- -0.13504593984303756
	pesos_i(16854) := b"1111111111111111_1111111111111111_1111001101010100_0000111011001010"; -- -0.049498630111550215
	pesos_i(16855) := b"1111111111111111_1111111111111111_1110001010100101_0111010111000110"; -- -0.11466278002372461
	pesos_i(16856) := b"1111111111111111_1111111111111111_1101100111101010_0111010101100111"; -- -0.14876619565583085
	pesos_i(16857) := b"1111111111111111_1111111111111111_1111100100000111_0000101100010011"; -- -0.027236278364706712
	pesos_i(16858) := b"1111111111111111_1111111111111111_1101101011111001_0111101000100001"; -- -0.1446307820964019
	pesos_i(16859) := b"0000000000000000_0000000000000000_0000001001100001_1011100010101010"; -- 0.009303609285211439
	pesos_i(16860) := b"0000000000000000_0000000000000000_0000001100111011_0011111001000001"; -- 0.012622729234070405
	pesos_i(16861) := b"1111111111111111_1111111111111111_1101100011000100_1101100100101000"; -- -0.15324633387477768
	pesos_i(16862) := b"1111111111111111_1111111111111111_1101100010001011_1101011101100011"; -- -0.15411619033354904
	pesos_i(16863) := b"0000000000000000_0000000000000000_0001001100100001_1100110111111101"; -- 0.07473456782239034
	pesos_i(16864) := b"0000000000000000_0000000000000000_0000111110101010_0011111001010100"; -- 0.06119145909397131
	pesos_i(16865) := b"1111111111111111_1111111111111111_1110111101100111_1001000110100111"; -- -0.06482591311297731
	pesos_i(16866) := b"1111111111111111_1111111111111111_1110010010010000_0111010111100101"; -- -0.10717070729670827
	pesos_i(16867) := b"0000000000000000_0000000000000000_0001101110111010_1100011100110110"; -- 0.10831875858407164
	pesos_i(16868) := b"0000000000000000_0000000000000000_0001110101110010_0101111010011001"; -- 0.11502639052622089
	pesos_i(16869) := b"1111111111111111_1111111111111111_1111100000111100_0101011011111110"; -- -0.030329287486226025
	pesos_i(16870) := b"0000000000000000_0000000000000000_0000101110010011_1001010001001000"; -- 0.04522063020313478
	pesos_i(16871) := b"0000000000000000_0000000000000000_0001101110000100_1010101101111100"; -- 0.10749313137890858
	pesos_i(16872) := b"1111111111111111_1111111111111111_1111111101101101_0101100111100000"; -- -0.002237684969451148
	pesos_i(16873) := b"0000000000000000_0000000000000000_0000000101110000_0111110001000110"; -- 0.0056226416979867945
	pesos_i(16874) := b"0000000000000000_0000000000000000_0001000011100110_0001110110001101"; -- 0.06601128281938118
	pesos_i(16875) := b"0000000000000000_0000000000000000_0010011010000100_0100111110000001"; -- 0.1504563990040259
	pesos_i(16876) := b"1111111111111111_1111111111111111_1101101011000101_0000100000111101"; -- -0.14543102763092255
	pesos_i(16877) := b"0000000000000000_0000000000000000_0001101000011011_0100110010111010"; -- 0.10197906049076406
	pesos_i(16878) := b"1111111111111111_1111111111111111_1111010001111001_0100110000111000"; -- -0.04502414360251986
	pesos_i(16879) := b"0000000000000000_0000000000000000_0001000100000001_0001110110111101"; -- 0.06642328141287941
	pesos_i(16880) := b"1111111111111111_1111111111111111_1111011000010001_1100001010101111"; -- -0.038791496585922104
	pesos_i(16881) := b"0000000000000000_0000000000000000_0000001010010001_0110100001100101"; -- 0.010031246735903363
	pesos_i(16882) := b"1111111111111111_1111111111111111_1110111000100000_1010011001010100"; -- -0.06981430484293065
	pesos_i(16883) := b"0000000000000000_0000000000000000_0000111000010011_0010110101100111"; -- 0.054980123217581604
	pesos_i(16884) := b"1111111111111111_1111111111111111_1110110101000000_1011111101010111"; -- -0.07323078276510908
	pesos_i(16885) := b"0000000000000000_0000000000000000_0001110110111010_0010100000111011"; -- 0.11612178270055498
	pesos_i(16886) := b"0000000000000000_0000000000000000_0001001011011111_1001101100110011"; -- 0.07372446053064642
	pesos_i(16887) := b"1111111111111111_1111111111111111_1110111011100000_0110010111011101"; -- -0.06688845979636372
	pesos_i(16888) := b"1111111111111111_1111111111111111_1101110000010000_1101010110001001"; -- -0.14036813164067183
	pesos_i(16889) := b"1111111111111111_1111111111111111_1101100111100111_1110001101110101"; -- -0.148805412310816
	pesos_i(16890) := b"1111111111111111_1111111111111111_1110011111101101_0011010011001000"; -- -0.09403677106675398
	pesos_i(16891) := b"1111111111111111_1111111111111111_1111101001011101_0101011110011101"; -- -0.022013210536810254
	pesos_i(16892) := b"0000000000000000_0000000000000000_0001010111010000_1111110100101001"; -- 0.08522016771674958
	pesos_i(16893) := b"1111111111111111_1111111111111111_1101111001010100_1100000101011101"; -- -0.13151923629616638
	pesos_i(16894) := b"1111111111111111_1111111111111111_1111111001011110_0110111001101100"; -- -0.006371592282294613
	pesos_i(16895) := b"1111111111111111_1111111111111111_1111110010001100_1001111010010001"; -- -0.013479318251277152
	pesos_i(16896) := b"1111111111111111_1111111111111111_1111100000010111_1101111000101010"; -- -0.030885805874057804
	pesos_i(16897) := b"0000000000000000_0000000000000000_0001101100001001_1000100011000101"; -- 0.10561423131211796
	pesos_i(16898) := b"1111111111111111_1111111111111111_1111011100110110_0101111101001110"; -- -0.03432659485719753
	pesos_i(16899) := b"0000000000000000_0000000000000000_0010010000100101_0010100000000101"; -- 0.14119196057398203
	pesos_i(16900) := b"0000000000000000_0000000000000000_0010010000001010_0001010000100000"; -- 0.14077878752543582
	pesos_i(16901) := b"0000000000000000_0000000000000000_0001001000000001_0101100001110001"; -- 0.07033303036573223
	pesos_i(16902) := b"0000000000000000_0000000000000000_0000100110000100_1111001000110001"; -- 0.03718484582697407
	pesos_i(16903) := b"1111111111111111_1111111111111111_1110000100111001_0011101111011000"; -- -0.12022043209044246
	pesos_i(16904) := b"0000000000000000_0000000000000000_0001010011001001_0001101001011000"; -- 0.08119358677470986
	pesos_i(16905) := b"1111111111111111_1111111111111111_1111001001100000_0100110001101011"; -- -0.05321810133628594
	pesos_i(16906) := b"0000000000000000_0000000000000000_0000110010001110_1001101110110111"; -- 0.04905102938880027
	pesos_i(16907) := b"0000000000000000_0000000000000000_0000111000110011_0101101100100100"; -- 0.05547113073860155
	pesos_i(16908) := b"0000000000000000_0000000000000000_0000001000111111_0001100110101011"; -- 0.008775333689709263
	pesos_i(16909) := b"1111111111111111_1111111111111111_1111001001010011_1011000111010001"; -- -0.05341042186339291
	pesos_i(16910) := b"1111111111111111_1111111111111111_1111111000100110_1100010000110111"; -- -0.007220970698279144
	pesos_i(16911) := b"1111111111111111_1111111111111111_1111101011011000_0011111000110100"; -- -0.02013789404188431
	pesos_i(16912) := b"0000000000000000_0000000000000000_0001011110110110_0011111101111101"; -- 0.09262463376677925
	pesos_i(16913) := b"1111111111111111_1111111111111111_1110001010111001_1101110011000111"; -- -0.11435146476903917
	pesos_i(16914) := b"0000000000000000_0000000000000000_0001101001010101_0011011111010010"; -- 0.10286282426144731
	pesos_i(16915) := b"1111111111111111_1111111111111111_1110000011000010_0010101110110010"; -- -0.1220371905730089
	pesos_i(16916) := b"0000000000000000_0000000000000000_0010000110101000_0101100100110000"; -- 0.13147504246451686
	pesos_i(16917) := b"1111111111111111_1111111111111111_1101111011000001_0001011010110101"; -- -0.12986620018928796
	pesos_i(16918) := b"1111111111111111_1111111111111111_1110101000111011_1101101011000000"; -- -0.08502419287693654
	pesos_i(16919) := b"0000000000000000_0000000000000000_0000110101000110_0011110001011011"; -- 0.051852962626676886
	pesos_i(16920) := b"0000000000000000_0000000000000000_0001100110000010_1011101001010100"; -- 0.09965099857498384
	pesos_i(16921) := b"0000000000000000_0000000000000000_0000100110011111_0000011100100010"; -- 0.03758282270959106
	pesos_i(16922) := b"0000000000000000_0000000000000000_0001110101001111_1101010011011001"; -- 0.11449938114763751
	pesos_i(16923) := b"1111111111111111_1111111111111111_1111010001101000_0111111101001001"; -- -0.0452804991273404
	pesos_i(16924) := b"0000000000000000_0000000000000000_0000101110110100_1110110100101010"; -- 0.045729468114909605
	pesos_i(16925) := b"1111111111111111_1111111111111111_1110010001010100_0100010011101011"; -- -0.10808915393426569
	pesos_i(16926) := b"0000000000000000_0000000000000000_0000001101100000_0111010001110011"; -- 0.013190534645588054
	pesos_i(16927) := b"0000000000000000_0000000000000000_0001101111010100_1001110000101110"; -- 0.10871292230377438
	pesos_i(16928) := b"1111111111111111_1111111111111111_1110110100111101_0111110100010000"; -- -0.07328050955521431
	pesos_i(16929) := b"0000000000000000_0000000000000000_0010010010000010_1100011101001111"; -- 0.1426205222706437
	pesos_i(16930) := b"1111111111111111_1111111111111111_1111111001000010_0100100100110101"; -- -0.006801056376991616
	pesos_i(16931) := b"1111111111111111_1111111111111111_1101100001110111_1001101001010111"; -- -0.15442500463255174
	pesos_i(16932) := b"0000000000000000_0000000000000000_0001011001101110_1100101010011011"; -- 0.08762804304767378
	pesos_i(16933) := b"0000000000000000_0000000000000000_0001011010111111_1000001000001101"; -- 0.08885968038842897
	pesos_i(16934) := b"1111111111111111_1111111111111111_1110110000111000_0010111100110110"; -- -0.07726769381811853
	pesos_i(16935) := b"0000000000000000_0000000000000000_0010000100001101_1010111001101000"; -- 0.1291150095920106
	pesos_i(16936) := b"1111111111111111_1111111111111111_1111100100001111_0000000100111011"; -- -0.027114794731017012
	pesos_i(16937) := b"0000000000000000_0000000000000000_0000011000011110_0111010101100010"; -- 0.023902260228638336
	pesos_i(16938) := b"1111111111111111_1111111111111111_1110100000101100_0001110100000010"; -- -0.09307688434045072
	pesos_i(16939) := b"1111111111111111_1111111111111111_1110010000011111_1011011111000011"; -- -0.10889102450972689
	pesos_i(16940) := b"1111111111111111_1111111111111111_1111100100000110_1111101001001100"; -- -0.027237278311186632
	pesos_i(16941) := b"0000000000000000_0000000000000000_0000001010010100_1010011101000110"; -- 0.010080770991837263
	pesos_i(16942) := b"1111111111111111_1111111111111111_1101110010001001_0110100100110010"; -- -0.13852827587173766
	pesos_i(16943) := b"0000000000000000_0000000000000000_0010010011010110_1001110100000010"; -- 0.14389973935512243
	pesos_i(16944) := b"0000000000000000_0000000000000000_0010001011001110_0111001010001110"; -- 0.13596263853749724
	pesos_i(16945) := b"1111111111111111_1111111111111111_1110110100110101_1101101001000011"; -- -0.07339702486424175
	pesos_i(16946) := b"1111111111111111_1111111111111111_1111010000100110_0101110010001110"; -- -0.04628964921069993
	pesos_i(16947) := b"0000000000000000_0000000000000000_0001010001010010_1110100101010100"; -- 0.07939012816439152
	pesos_i(16948) := b"0000000000000000_0000000000000000_0001001110001100_1101010010001111"; -- 0.07636765003262393
	pesos_i(16949) := b"1111111111111111_1111111111111111_1110101101100110_0000001101110001"; -- -0.08047464847888425
	pesos_i(16950) := b"0000000000000000_0000000000000000_0010000010010101_1001101100011100"; -- 0.12728280475648593
	pesos_i(16951) := b"0000000000000000_0000000000000000_0000101000111010_1001011011011110"; -- 0.03995650225397717
	pesos_i(16952) := b"1111111111111111_1111111111111111_1110001010011101_1001100000110011"; -- -0.11478279837039516
	pesos_i(16953) := b"1111111111111111_1111111111111111_1101110011100101_0000011110011001"; -- -0.13713028435272076
	pesos_i(16954) := b"0000000000000000_0000000000000000_0000011000000100_0000011100010110"; -- 0.023498957480833037
	pesos_i(16955) := b"1111111111111111_1111111111111111_1111000101100011_0100110011111001"; -- -0.05707854199101851
	pesos_i(16956) := b"1111111111111111_1111111111111111_1111001000101000_0011111101101110"; -- -0.05407336781630332
	pesos_i(16957) := b"0000000000000000_0000000000000000_0000010000101000_1010000011111011"; -- 0.01624494663814575
	pesos_i(16958) := b"0000000000000000_0000000000000000_0010001100101101_0101000011011111"; -- 0.13741021587883556
	pesos_i(16959) := b"0000000000000000_0000000000000000_0000100010111011_0000001100000110"; -- 0.03410357370115574
	pesos_i(16960) := b"1111111111111111_1111111111111111_1101101110000101_0101010001011011"; -- -0.1424968030324929
	pesos_i(16961) := b"1111111111111111_1111111111111111_1110101011100100_0111001000000110"; -- -0.0824516997315355
	pesos_i(16962) := b"1111111111111111_1111111111111111_1111011000010000_1111110011001010"; -- -0.03880329197800103
	pesos_i(16963) := b"0000000000000000_0000000000000000_0001101100101001_0000111100101000"; -- 0.10609526379248167
	pesos_i(16964) := b"1111111111111111_1111111111111111_1111110111101011_0010100010110101"; -- -0.008130508290123573
	pesos_i(16965) := b"0000000000000000_0000000000000000_0000101010001100_0000100011000111"; -- 0.041199253609865774
	pesos_i(16966) := b"1111111111111111_1111111111111111_1110011110100100_1001111010001000"; -- -0.09514435948475665
	pesos_i(16967) := b"0000000000000000_0000000000000000_0000001101000010_0011111101010111"; -- 0.01272960550269451
	pesos_i(16968) := b"0000000000000000_0000000000000000_0001110001101010_0110001100010110"; -- 0.11099833771931182
	pesos_i(16969) := b"1111111111111111_1111111111111111_1111111010011000_0110011001101110"; -- -0.005487058822103148
	pesos_i(16970) := b"1111111111111111_1111111111111111_1110100101000100_0011001011110100"; -- -0.0888031153645112
	pesos_i(16971) := b"1111111111111111_1111111111111111_1110010001101110_1101110111101011"; -- -0.10768330585042071
	pesos_i(16972) := b"0000000000000000_0000000000000000_0010011001110101_1110010001001000"; -- 0.15023638485037277
	pesos_i(16973) := b"1111111111111111_1111111111111111_1111000101010001_1011000101011010"; -- -0.05734721700576558
	pesos_i(16974) := b"1111111111111111_1111111111111111_1101101000111010_1011000000111110"; -- -0.14754198548876551
	pesos_i(16975) := b"1111111111111111_1111111111111111_1110110110111000_1011011100100110"; -- -0.07140021634913948
	pesos_i(16976) := b"1111111111111111_1111111111111111_1111010111011110_0100101100011110"; -- -0.03957682139977003
	pesos_i(16977) := b"1111111111111111_1111111111111111_1101111111001000_0110110010010110"; -- -0.1258480199496623
	pesos_i(16978) := b"1111111111111111_1111111111111111_1110110111001010_1011110000100100"; -- -0.07112526055210186
	pesos_i(16979) := b"0000000000000000_0000000000000000_0000110011111001_0000011010010011"; -- 0.050674830282481986
	pesos_i(16980) := b"1111111111111111_1111111111111111_1111111010011010_1100110110100001"; -- -0.005450390108977156
	pesos_i(16981) := b"1111111111111111_1111111111111111_1110111001101011_0111010001111101"; -- -0.0686728663268224
	pesos_i(16982) := b"0000000000000000_0000000000000000_0001001001110101_1100010010101100"; -- 0.07210950093313787
	pesos_i(16983) := b"1111111111111111_1111111111111111_1110101101110110_0011000001110101"; -- -0.0802278245206881
	pesos_i(16984) := b"0000000000000000_0000000000000000_0000101001001111_1010111000100100"; -- 0.04027832388191692
	pesos_i(16985) := b"0000000000000000_0000000000000000_0001110111111100_0000111010110110"; -- 0.11712734170363552
	pesos_i(16986) := b"0000000000000000_0000000000000000_0000011010101100_0001001011001111"; -- 0.026063132881625796
	pesos_i(16987) := b"1111111111111111_1111111111111111_1110011101001011_1100001101111100"; -- -0.09650018911681751
	pesos_i(16988) := b"1111111111111111_1111111111111111_1110010011101110_1110011010110000"; -- -0.10572965814170296
	pesos_i(16989) := b"1111111111111111_1111111111111111_1111001001011100_0010001100110011"; -- -0.05328159327777476
	pesos_i(16990) := b"0000000000000000_0000000000000000_0000000100001100_1111100000011100"; -- 0.004104143958925162
	pesos_i(16991) := b"1111111111111111_1111111111111111_1110001001111100_0001101001001101"; -- -0.11529384239804555
	pesos_i(16992) := b"1111111111111111_1111111111111111_1110000111001011_0101000000110101"; -- -0.1179914351756431
	pesos_i(16993) := b"0000000000000000_0000000000000000_0000110011100000_0111111010100101"; -- 0.05030051738203364
	pesos_i(16994) := b"0000000000000000_0000000000000000_0010010011010101_0111111101010010"; -- 0.1438827110419901
	pesos_i(16995) := b"0000000000000000_0000000000000000_0000110100010110_0100100000000110"; -- 0.051121236190247374
	pesos_i(16996) := b"1111111111111111_1111111111111111_1111111111001000_0000010101010100"; -- -0.0008541746057652582
	pesos_i(16997) := b"0000000000000000_0000000000000000_0000001111001011_0111000111001110"; -- 0.01482306751875029
	pesos_i(16998) := b"1111111111111111_1111111111111111_1111110111110001_0111010110010101"; -- -0.008034373402832876
	pesos_i(16999) := b"1111111111111111_1111111111111111_1111000100001110_1111001110100101"; -- -0.058365604633160546
	pesos_i(17000) := b"0000000000000000_0000000000000000_0010001000101011_1101110110110110"; -- 0.1334818430067662
	pesos_i(17001) := b"1111111111111111_1111111111111111_1111010000111001_0011011101010101"; -- -0.04600195091991978
	pesos_i(17002) := b"0000000000000000_0000000000000000_0000110010010111_1000111001100000"; -- 0.0491875633021439
	pesos_i(17003) := b"0000000000000000_0000000000000000_0010001100000001_0110010011111110"; -- 0.13674002828756324
	pesos_i(17004) := b"1111111111111111_1111111111111111_1110010111011011_0110011010000000"; -- -0.10212096563660635
	pesos_i(17005) := b"0000000000000000_0000000000000000_0001001111111111_0000010000100111"; -- 0.07810998878597067
	pesos_i(17006) := b"0000000000000000_0000000000000000_0001100001101101_1100101111110101"; -- 0.09542536475205078
	pesos_i(17007) := b"1111111111111111_1111111111111111_1110101101111010_0100011010010111"; -- -0.08016547029693305
	pesos_i(17008) := b"1111111111111111_1111111111111111_1111111011110100_0100010001101010"; -- -0.004085277737935361
	pesos_i(17009) := b"1111111111111111_1111111111111111_1110000110001000_1011110111011101"; -- -0.11900723800284262
	pesos_i(17010) := b"0000000000000000_0000000000000000_0001011001101110_1010011000100011"; -- 0.08762586940364125
	pesos_i(17011) := b"1111111111111111_1111111111111111_1111011010011111_1110010111000101"; -- -0.036622657114895714
	pesos_i(17012) := b"0000000000000000_0000000000000000_0000110000010100_0101110111000011"; -- 0.047185764377825797
	pesos_i(17013) := b"0000000000000000_0000000000000000_0010000010111100_1010000100010110"; -- 0.12787825373409095
	pesos_i(17014) := b"1111111111111111_1111111111111111_1111010001110100_0000000110101001"; -- -0.045104881631190794
	pesos_i(17015) := b"1111111111111111_1111111111111111_1110010111011100_0000110101011111"; -- -0.10211101951327808
	pesos_i(17016) := b"1111111111111111_1111111111111111_1111111111100000_1110011100110111"; -- -0.0004744997172832566
	pesos_i(17017) := b"0000000000000000_0000000000000000_0001110010110001_1001000011001110"; -- 0.11208443678463305
	pesos_i(17018) := b"0000000000000000_0000000000000000_0000111110011100_0011001011111010"; -- 0.06097715945147442
	pesos_i(17019) := b"0000000000000000_0000000000000000_0000001010100101_0101001101010001"; -- 0.010335166334993382
	pesos_i(17020) := b"0000000000000000_0000000000000000_0001100011011111_0101000010101111"; -- 0.09715751918969773
	pesos_i(17021) := b"0000000000000000_0000000000000000_0001101100101010_1100101101000110"; -- 0.10612173521489775
	pesos_i(17022) := b"0000000000000000_0000000000000000_0001010010001110_1000000110100010"; -- 0.08029947486728495
	pesos_i(17023) := b"0000000000000000_0000000000000000_0000101001100100_1011010010110110"; -- 0.040599150120069254
	pesos_i(17024) := b"0000000000000000_0000000000000000_0000000001100001_0000110001000011"; -- 0.001480833454372974
	pesos_i(17025) := b"1111111111111111_1111111111111111_1110010001000000_0110110010111101"; -- -0.10839195612417775
	pesos_i(17026) := b"0000000000000000_0000000000000000_0001111011001000_0010101011000110"; -- 0.12024180740838372
	pesos_i(17027) := b"1111111111111111_1111111111111111_1110111100000101_1010010011000011"; -- -0.06632013542299223
	pesos_i(17028) := b"1111111111111111_1111111111111111_1101111100101011_1111101001001010"; -- -0.12823520377265504
	pesos_i(17029) := b"0000000000000000_0000000000000000_0010000001010011_1010100101001001"; -- 0.1262765696860417
	pesos_i(17030) := b"0000000000000000_0000000000000000_0001011110110110_0100010110100111"; -- 0.09262500120824563
	pesos_i(17031) := b"0000000000000000_0000000000000000_0001101110111001_1010110001100001"; -- 0.10830190047615584
	pesos_i(17032) := b"0000000000000000_0000000000000000_0001111011010110_0011100000001000"; -- 0.12045622064443429
	pesos_i(17033) := b"0000000000000000_0000000000000000_0001000010100001_1001110000011110"; -- 0.06496597031231184
	pesos_i(17034) := b"0000000000000000_0000000000000000_0000001000010100_1010011011101000"; -- 0.008127624170683419
	pesos_i(17035) := b"1111111111111111_1111111111111111_1110001101011101_1100111010110000"; -- -0.1118498630311688
	pesos_i(17036) := b"0000000000000000_0000000000000000_0010011111100011_1101001100011011"; -- 0.15582007809086101
	pesos_i(17037) := b"0000000000000000_0000000000000000_0001011101010111_1001100110001110"; -- 0.09118041732146472
	pesos_i(17038) := b"0000000000000000_0000000000000000_0010000100110111_1000100101000001"; -- 0.1297536644719778
	pesos_i(17039) := b"0000000000000000_0000000000000000_0001011000010001_1001000000000011"; -- 0.08620548308583843
	pesos_i(17040) := b"0000000000000000_0000000000000000_0000110000001111_0110101111011010"; -- 0.04711031019006714
	pesos_i(17041) := b"0000000000000000_0000000000000000_0000011101111110_1110110110011010"; -- 0.029280519611176423
	pesos_i(17042) := b"1111111111111111_1111111111111111_1111100101011110_0100011100100100"; -- -0.02590518350757798
	pesos_i(17043) := b"0000000000000000_0000000000000000_0000000000100101_0110110101000001"; -- 0.0005710872194766993
	pesos_i(17044) := b"0000000000000000_0000000000000000_0001010101101110_0111110110010011"; -- 0.08371720166998224
	pesos_i(17045) := b"0000000000000000_0000000000000000_0010001111100110_1100001010101011"; -- 0.1402398745198617
	pesos_i(17046) := b"0000000000000000_0000000000000000_0001110111100110_0001000001001110"; -- 0.11679174323217391
	pesos_i(17047) := b"1111111111111111_1111111111111111_1110110000110111_0010111101010000"; -- -0.07728294646149121
	pesos_i(17048) := b"0000000000000000_0000000000000000_0001101010000010_1110001101110100"; -- 0.10355969993033877
	pesos_i(17049) := b"0000000000000000_0000000000000000_0001111111001000_1100010100111100"; -- 0.1241572639706973
	pesos_i(17050) := b"0000000000000000_0000000000000000_0000011001111110_0100111010000100"; -- 0.02536478734630325
	pesos_i(17051) := b"1111111111111111_1111111111111111_1110000011011100_1010111101111110"; -- -0.12163260630050364
	pesos_i(17052) := b"0000000000000000_0000000000000000_0000111010000001_1111001101000001"; -- 0.056670382894487566
	pesos_i(17053) := b"1111111111111111_1111111111111111_1111001110011100_1100110100110111"; -- -0.04838864703310093
	pesos_i(17054) := b"0000000000000000_0000000000000000_0001011110100111_1000110101001011"; -- 0.09240038957231657
	pesos_i(17055) := b"0000000000000000_0000000000000000_0000101010111011_1110100111001101"; -- 0.04192982921511724
	pesos_i(17056) := b"0000000000000000_0000000000000000_0001100111001011_0110110101110110"; -- 0.10076030853396477
	pesos_i(17057) := b"1111111111111111_1111111111111111_1111100101001001_0111100111011101"; -- -0.026222594829512707
	pesos_i(17058) := b"1111111111111111_1111111111111111_1110001000100010_1011100111000000"; -- -0.1166576296932819
	pesos_i(17059) := b"0000000000000000_0000000000000000_0010010101110001_0101111101110111"; -- 0.14626118332006033
	pesos_i(17060) := b"0000000000000000_0000000000000000_0010010010000101_0001111101011001"; -- 0.14265628752469153
	pesos_i(17061) := b"1111111111111111_1111111111111111_1101100110001000_0101100110011101"; -- -0.1502632132797404
	pesos_i(17062) := b"0000000000000000_0000000000000000_0000010010011101_0111011001000010"; -- 0.01802767849253764
	pesos_i(17063) := b"0000000000000000_0000000000000000_0001111000000000_0111110100101100"; -- 0.11719496077751006
	pesos_i(17064) := b"1111111111111111_1111111111111111_1110111001000001_0100001101000000"; -- -0.06931667027870421
	pesos_i(17065) := b"1111111111111111_1111111111111111_1101011111000110_1000011111110110"; -- -0.1571269058145396
	pesos_i(17066) := b"1111111111111111_1111111111111111_1110100100111001_1010111000010110"; -- -0.088963622776783
	pesos_i(17067) := b"1111111111111111_1111111111111111_1111110010010001_0110000100011010"; -- -0.013406687993103244
	pesos_i(17068) := b"1111111111111111_1111111111111111_1101110010010011_0010111110000010"; -- -0.13837912642522776
	pesos_i(17069) := b"1111111111111111_1111111111111111_1110101011011000_0111010100100101"; -- -0.08263461916701288
	pesos_i(17070) := b"1111111111111111_1111111111111111_1110101101111000_0011011001010010"; -- -0.08019695764681065
	pesos_i(17071) := b"0000000000000000_0000000000000000_0000001011110001_0010100011000010"; -- 0.011492297491315263
	pesos_i(17072) := b"0000000000000000_0000000000000000_0000001100011111_0000000101011101"; -- 0.01219185362768964
	pesos_i(17073) := b"1111111111111111_1111111111111111_1101100101101011_1101110100110100"; -- -0.15069787489871064
	pesos_i(17074) := b"1111111111111111_1111111111111111_1101110011001111_1110000000000111"; -- -0.13745307767133527
	pesos_i(17075) := b"1111111111111111_1111111111111111_1111011000011011_1000100111001100"; -- -0.0386422994182959
	pesos_i(17076) := b"1111111111111111_1111111111111111_1101110011100110_0011111000000100"; -- -0.1371117820868374
	pesos_i(17077) := b"0000000000000000_0000000000000000_0001110100010100_0001001100100010"; -- 0.11358756616295378
	pesos_i(17078) := b"0000000000000000_0000000000000000_0000001010111110_0100000000010000"; -- 0.010715488277095632
	pesos_i(17079) := b"1111111111111111_1111111111111111_1111101010111111_1000111110111100"; -- -0.020514503983980265
	pesos_i(17080) := b"1111111111111111_1111111111111111_1110111100101101_0101000110001111"; -- -0.06571474312387049
	pesos_i(17081) := b"1111111111111111_1111111111111111_1110011111000001_0010100010110111"; -- -0.09470887690063187
	pesos_i(17082) := b"0000000000000000_0000000000000000_0000011101111011_0101011010100011"; -- 0.029225745011266305
	pesos_i(17083) := b"1111111111111111_1111111111111111_1101110111111101_0100010000011000"; -- -0.1328542177330785
	pesos_i(17084) := b"0000000000000000_0000000000000000_0001110110110011_1010101110100100"; -- 0.1160228037612287
	pesos_i(17085) := b"0000000000000000_0000000000000000_0001010101111100_0111110110001100"; -- 0.0839308230578097
	pesos_i(17086) := b"1111111111111111_1111111111111111_1111111110001100_1100111100011010"; -- -0.0017576752815718264
	pesos_i(17087) := b"1111111111111111_1111111111111111_1110001010000001_0111001010001110"; -- -0.11521228830600122
	pesos_i(17088) := b"1111111111111111_1111111111111111_1111111000010110_1000011101001101"; -- -0.00746874218059821
	pesos_i(17089) := b"1111111111111111_1111111111111111_1110011101000000_0101001001010010"; -- -0.09667478092053344
	pesos_i(17090) := b"0000000000000000_0000000000000000_0000001000011000_1110011101100101"; -- 0.008192503027201802
	pesos_i(17091) := b"1111111111111111_1111111111111111_1111011101110010_1010011100001000"; -- -0.03340679210804212
	pesos_i(17092) := b"0000000000000000_0000000000000000_0000000110000001_1101001010110010"; -- 0.005887192247626204
	pesos_i(17093) := b"0000000000000000_0000000000000000_0000001111000101_1001110111010101"; -- 0.014734139061927944
	pesos_i(17094) := b"1111111111111111_1111111111111111_1110101010100001_1011011111110100"; -- -0.08346987059688687
	pesos_i(17095) := b"1111111111111111_1111111111111111_1111110110110011_1101001011111010"; -- -0.008974851621360776
	pesos_i(17096) := b"1111111111111111_1111111111111111_1111011100101011_0100010101101001"; -- -0.0344959848542817
	pesos_i(17097) := b"1111111111111111_1111111111111111_1101111011001100_0100101101010000"; -- -0.12969521809359302
	pesos_i(17098) := b"1111111111111111_1111111111111111_1111101011100100_0110110011010100"; -- -0.019952009437375406
	pesos_i(17099) := b"1111111111111111_1111111111111111_1110100010111110_0110111111100110"; -- -0.09084416035784523
	pesos_i(17100) := b"1111111111111111_1111111111111111_1111011100001111_0111101011101010"; -- -0.034920041817527024
	pesos_i(17101) := b"1111111111111111_1111111111111111_1101101111100101_1101110010101001"; -- -0.14102383491618023
	pesos_i(17102) := b"1111111111111111_1111111111111111_1111110001111001_1111100111001101"; -- -0.013763797346809716
	pesos_i(17103) := b"0000000000000000_0000000000000000_0001111101001110_1011000101101011"; -- 0.12229451037802082
	pesos_i(17104) := b"1111111111111111_1111111111111111_1101110110101010_1010001011101101"; -- -0.134115044761612
	pesos_i(17105) := b"1111111111111111_1111111111111111_1111000000011110_0011111111001000"; -- -0.062038434669066424
	pesos_i(17106) := b"1111111111111111_1111111111111111_1111011011000101_1100111110100011"; -- -0.0360441423344604
	pesos_i(17107) := b"1111111111111111_1111111111111111_1101111110000111_0110110111010011"; -- -0.126839767446967
	pesos_i(17108) := b"1111111111111111_1111111111111111_1111010010100111_0000111011001100"; -- -0.044325900368422565
	pesos_i(17109) := b"0000000000000000_0000000000000000_0000011010111001_0110010100101100"; -- 0.026266406267689987
	pesos_i(17110) := b"0000000000000000_0000000000000000_0000111110110010_1111111010110100"; -- 0.06132499598812648
	pesos_i(17111) := b"0000000000000000_0000000000000000_0010000011111001_1101111001100101"; -- 0.12881269420627628
	pesos_i(17112) := b"0000000000000000_0000000000000000_0001000101101101_0110000100010000"; -- 0.06807524338365453
	pesos_i(17113) := b"0000000000000000_0000000000000000_0000101100001011_1001110110110011"; -- 0.04314599626256026
	pesos_i(17114) := b"1111111111111111_1111111111111111_1110100111011100_0100110001101011"; -- -0.08648226148358566
	pesos_i(17115) := b"0000000000000000_0000000000000000_0000100101111010_0010011101101011"; -- 0.03702017180425966
	pesos_i(17116) := b"1111111111111111_1111111111111111_1111101011110111_1001111100001111"; -- -0.019659098536687486
	pesos_i(17117) := b"0000000000000000_0000000000000000_0000101011001101_1110000101110110"; -- 0.0422039903267735
	pesos_i(17118) := b"1111111111111111_1111111111111111_1110110111100101_1000010101000001"; -- -0.07071654474982288
	pesos_i(17119) := b"1111111111111111_1111111111111111_1110100011101000_0010111000111110"; -- -0.09020720469960218
	pesos_i(17120) := b"1111111111111111_1111111111111111_1110000100011011_1110101011100111"; -- -0.12066776137024861
	pesos_i(17121) := b"0000000000000000_0000000000000000_0010000111011001_0110111011011000"; -- 0.13222401413620194
	pesos_i(17122) := b"0000000000000000_0000000000000000_0001000100011001_0111101010000000"; -- 0.06679502130235691
	pesos_i(17123) := b"1111111111111111_1111111111111111_1111100001010111_1101110000101111"; -- -0.029909361325027677
	pesos_i(17124) := b"0000000000000000_0000000000000000_0000101101111101_0100111111011100"; -- 0.04488085856325107
	pesos_i(17125) := b"1111111111111111_1111111111111111_1111111001101010_1001000001011010"; -- -0.006186464229175379
	pesos_i(17126) := b"1111111111111111_1111111111111111_1101101100000111_0010010100010000"; -- -0.14442222939035815
	pesos_i(17127) := b"0000000000000000_0000000000000000_0000101010010000_1011000010111011"; -- 0.041270299696196264
	pesos_i(17128) := b"0000000000000000_0000000000000000_0001001011111001_0011101110101110"; -- 0.0741154957445332
	pesos_i(17129) := b"1111111111111111_1111111111111111_1111001100111111_1101111110111010"; -- -0.04980661118468717
	pesos_i(17130) := b"1111111111111111_1111111111111111_1111001100000100_1101011010001000"; -- -0.05070742789026127
	pesos_i(17131) := b"1111111111111111_1111111111111111_1111001111100110_0011110001011011"; -- -0.04726813097961252
	pesos_i(17132) := b"1111111111111111_1111111111111111_1110100010101110_1011100000001111"; -- -0.09108399999762501
	pesos_i(17133) := b"1111111111111111_1111111111111111_1111101111010010_1001110100101011"; -- -0.016317536445223494
	pesos_i(17134) := b"1111111111111111_1111111111111111_1101110011100001_0111101101001110"; -- -0.13718442289922772
	pesos_i(17135) := b"1111111111111111_1111111111111111_1110100110110100_1011011111101111"; -- -0.08708620474766571
	pesos_i(17136) := b"0000000000000000_0000000000000000_0001000111110010_0110010101100001"; -- 0.07010491970215318
	pesos_i(17137) := b"0000000000000000_0000000000000000_0000110001101010_1001101001100010"; -- 0.048501633506812546
	pesos_i(17138) := b"0000000000000000_0000000000000000_0010001100101111_1000101111001111"; -- 0.13744424635425487
	pesos_i(17139) := b"1111111111111111_1111111111111111_1111111101110011_0011111101101000"; -- -0.0021477099564934377
	pesos_i(17140) := b"0000000000000000_0000000000000000_0000000001000100_1110100101011110"; -- 0.001051507394598441
	pesos_i(17141) := b"0000000000000000_0000000000000000_0001011001011001_1111101111110101"; -- 0.08731054997314353
	pesos_i(17142) := b"0000000000000000_0000000000000000_0001011100011100_0011101100000010"; -- 0.09027451313316642
	pesos_i(17143) := b"0000000000000000_0000000000000000_0001100000110010_1011010101011000"; -- 0.09452374829489414
	pesos_i(17144) := b"1111111111111111_1111111111111111_1110111110110001_0001110100001111"; -- -0.06370371227074006
	pesos_i(17145) := b"1111111111111111_1111111111111111_1110100011110000_1101110110111111"; -- -0.09007467363740508
	pesos_i(17146) := b"0000000000000000_0000000000000000_0001001001111011_0011101000101111"; -- 0.07219279909243274
	pesos_i(17147) := b"1111111111111111_1111111111111111_1111100001101111_0100111100010010"; -- -0.02955156140372518
	pesos_i(17148) := b"1111111111111111_1111111111111111_1101110001011100_1101110110111101"; -- -0.1392079747436822
	pesos_i(17149) := b"0000000000000000_0000000000000000_0000111010100110_1110001010101101"; -- 0.0572339699304333
	pesos_i(17150) := b"0000000000000000_0000000000000000_0001101010100100_1011000010010001"; -- 0.10407546563078869
	pesos_i(17151) := b"1111111111111111_1111111111111111_1111110011100010_1101101101011100"; -- -0.012163438750905038
	pesos_i(17152) := b"0000000000000000_0000000000000000_0001010111111110_1010000110011110"; -- 0.08591661545861265
	pesos_i(17153) := b"0000000000000000_0000000000000000_0001010000000101_0110001101010111"; -- 0.07820721502736926
	pesos_i(17154) := b"0000000000000000_0000000000000000_0000010111011000_0111010001011101"; -- 0.022834084129919368
	pesos_i(17155) := b"1111111111111111_1111111111111111_1111000111110101_1001011000110111"; -- -0.054846393209583816
	pesos_i(17156) := b"1111111111111111_1111111111111111_1111111000100000_0011110010111111"; -- -0.007320597958877086
	pesos_i(17157) := b"0000000000000000_0000000000000000_0010010101000011_1110110000101001"; -- 0.14556766515069136
	pesos_i(17158) := b"0000000000000000_0000000000000000_0010000100011110_0110001101101100"; -- 0.12936993976298136
	pesos_i(17159) := b"0000000000000000_0000000000000000_0000110011010010_0101000000000011"; -- 0.05008411482134842
	pesos_i(17160) := b"1111111111111111_1111111111111111_1101111011001011_1111010010100110"; -- -0.129700383628683
	pesos_i(17161) := b"1111111111111111_1111111111111111_1111111000111001_0001010000100001"; -- -0.006941549341670932
	pesos_i(17162) := b"0000000000000000_0000000000000000_0001101110011011_1011110011110110"; -- 0.10784512517618085
	pesos_i(17163) := b"0000000000000000_0000000000000000_0000011101000000_1101000011111001"; -- 0.028332768312028706
	pesos_i(17164) := b"1111111111111111_1111111111111111_1110110101011001_1010010100000110"; -- -0.07285088163673091
	pesos_i(17165) := b"0000000000000000_0000000000000000_0010011011110111_1001001101011010"; -- 0.1522152036405213
	pesos_i(17166) := b"0000000000000000_0000000000000000_0001001000101101_0010101011001110"; -- 0.07100169694035056
	pesos_i(17167) := b"0000000000000000_0000000000000000_0001010011101010_0111001101010010"; -- 0.08170243038107448
	pesos_i(17168) := b"0000000000000000_0000000000000000_0001110100001001_0100000110010010"; -- 0.11342248734484664
	pesos_i(17169) := b"1111111111111111_1111111111111111_1110011010101001_1110110101011100"; -- -0.09896961692178748
	pesos_i(17170) := b"0000000000000000_0000000000000000_0010011101011010_1110101001110111"; -- 0.1537310163017156
	pesos_i(17171) := b"0000000000000000_0000000000000000_0001111100110010_1101010001101001"; -- 0.12186935018632804
	pesos_i(17172) := b"0000000000000000_0000000000000000_0010000000010100_0001010000110011"; -- 0.12530637967212716
	pesos_i(17173) := b"1111111111111111_1111111111111111_1111010010010111_1100001100110110"; -- -0.04455928737590646
	pesos_i(17174) := b"1111111111111111_1111111111111111_1110000111100110_1011110011001110"; -- -0.11757297477316633
	pesos_i(17175) := b"1111111111111111_1111111111111111_1111010111100110_0001010010111001"; -- -0.03945799330482609
	pesos_i(17176) := b"1111111111111111_1111111111111111_1110010111111010_0001000010100100"; -- -0.10165306089158437
	pesos_i(17177) := b"0000000000000000_0000000000000000_0000010001111101_0110110100011101"; -- 0.017538852241387043
	pesos_i(17178) := b"1111111111111111_1111111111111111_1110111001101001_1010011000001010"; -- -0.06870043036616122
	pesos_i(17179) := b"0000000000000000_0000000000000000_0001111100010011_1001000110001100"; -- 0.12139234217344091
	pesos_i(17180) := b"0000000000000000_0000000000000000_0000001010011010_1100110001110101"; -- 0.010174540213962746
	pesos_i(17181) := b"1111111111111111_1111111111111111_1111110011010000_1001000111001111"; -- -0.012442481053714973
	pesos_i(17182) := b"1111111111111111_1111111111111111_1110110111110100_1011011000101000"; -- -0.07048474808264585
	pesos_i(17183) := b"0000000000000000_0000000000000000_0001011011011111_0010111000000010"; -- 0.08934295222395314
	pesos_i(17184) := b"0000000000000000_0000000000000000_0000011110111110_1100001111100100"; -- 0.030254596017679315
	pesos_i(17185) := b"0000000000000000_0000000000000000_0001100100001101_1110010110101010"; -- 0.09786830335112635
	pesos_i(17186) := b"1111111111111111_1111111111111111_1101100101000001_0110100001000110"; -- -0.1513457135907991
	pesos_i(17187) := b"1111111111111111_1111111111111111_1110011001000001_1001001000010110"; -- -0.10056197134124123
	pesos_i(17188) := b"1111111111111111_1111111111111111_1111011001111011_0011001100000110"; -- -0.03718262764192375
	pesos_i(17189) := b"1111111111111111_1111111111111111_1110011011101101_1101111000010100"; -- -0.0979329300539904
	pesos_i(17190) := b"1111111111111111_1111111111111111_1111101010000110_0010101111011100"; -- -0.021390207970409657
	pesos_i(17191) := b"0000000000000000_0000000000000000_0001011101001010_1010101010001111"; -- 0.090983066503851
	pesos_i(17192) := b"1111111111111111_1111111111111111_1110100101001101_0101010111111001"; -- -0.08866369887731208
	pesos_i(17193) := b"1111111111111111_1111111111111111_1110011100100000_0010100010101000"; -- -0.09716554537862485
	pesos_i(17194) := b"1111111111111111_1111111111111111_1111101001100000_1110001011110110"; -- -0.021959128227728133
	pesos_i(17195) := b"0000000000000000_0000000000000000_0010010000110000_1111011000111000"; -- 0.1413720976619192
	pesos_i(17196) := b"1111111111111111_1111111111111111_1110100001001000_1000111010001010"; -- -0.09264287117797596
	pesos_i(17197) := b"0000000000000000_0000000000000000_0001011011011001_1010011110110011"; -- 0.08925865282867998
	pesos_i(17198) := b"0000000000000000_0000000000000000_0001100100100100_1101001001100110"; -- 0.09821810721840073
	pesos_i(17199) := b"0000000000000000_0000000000000000_0000100000011011_1011111011100011"; -- 0.0316733650911018
	pesos_i(17200) := b"0000000000000000_0000000000000000_0000100000010011_0010111101011010"; -- 0.03154273934272983
	pesos_i(17201) := b"0000000000000000_0000000000000000_0001101000011100_0011011101010111"; -- 0.1019930446398123
	pesos_i(17202) := b"0000000000000000_0000000000000000_0001001101001001_1011001111000100"; -- 0.07534335638228395
	pesos_i(17203) := b"0000000000000000_0000000000000000_0010101001110101_0111000101001110"; -- 0.1658545317858055
	pesos_i(17204) := b"1111111111111111_1111111111111111_1110100110010001_1110000111000111"; -- -0.08761776826291304
	pesos_i(17205) := b"1111111111111111_1111111111111111_1110100001111100_0010001100010011"; -- -0.09185581961065935
	pesos_i(17206) := b"0000000000000000_0000000000000000_0001011110101111_1111011110101001"; -- 0.09252879979448096
	pesos_i(17207) := b"0000000000000000_0000000000000000_0000101001100110_1110001100010111"; -- 0.040632432047454675
	pesos_i(17208) := b"1111111111111111_1111111111111111_1110111100100101_0010011111001111"; -- -0.06583930197746975
	pesos_i(17209) := b"1111111111111111_1111111111111111_1111111010110011_0100111000010011"; -- -0.005076523147373372
	pesos_i(17210) := b"1111111111111111_1111111111111111_1111111011011010_0111010101001001"; -- -0.004479093210603666
	pesos_i(17211) := b"0000000000000000_0000000000000000_0001110000100001_1000001110010100"; -- 0.10988638268044033
	pesos_i(17212) := b"1111111111111111_1111111111111111_1110001111000001_0001011000101001"; -- -0.11033498280236387
	pesos_i(17213) := b"0000000000000000_0000000000000000_0001000100001011_1111001101010111"; -- 0.06658860075947758
	pesos_i(17214) := b"1111111111111111_1111111111111111_1110001111101110_0010111111101010"; -- -0.10964680239002837
	pesos_i(17215) := b"0000000000000000_0000000000000000_0010000110000111_1111001110001000"; -- 0.1309807021401603
	pesos_i(17216) := b"1111111111111111_1111111111111111_1110100101011001_0111000101010110"; -- -0.08847896233965177
	pesos_i(17217) := b"1111111111111111_1111111111111111_1101101010000110_0011100111100110"; -- -0.1463893711428132
	pesos_i(17218) := b"1111111111111111_1111111111111111_1111001110011100_1011001010101010"; -- -0.048390229622228345
	pesos_i(17219) := b"1111111111111111_1111111111111111_1111110100001110_0110100100101011"; -- -0.011498858393308088
	pesos_i(17220) := b"0000000000000000_0000000000000000_0000100011111011_0100101010000110"; -- 0.0350843980541957
	pesos_i(17221) := b"0000000000000000_0000000000000000_0000001000110001_1010010101000000"; -- 0.008570030386896589
	pesos_i(17222) := b"1111111111111111_1111111111111111_1111011101111011_1100100111000100"; -- -0.033267392670098844
	pesos_i(17223) := b"0000000000000000_0000000000000000_0001000100111110_0100011110100100"; -- 0.06735656497221947
	pesos_i(17224) := b"0000000000000000_0000000000000000_0001100111111011_1100001100010110"; -- 0.10149783402620229
	pesos_i(17225) := b"0000000000000000_0000000000000000_0000000100110111_1100101001111000"; -- 0.004757551396937791
	pesos_i(17226) := b"1111111111111111_1111111111111111_1101110000110010_0101101101001000"; -- -0.1398566198279723
	pesos_i(17227) := b"0000000000000000_0000000000000000_0001100000111101_1110010001111101"; -- 0.09469440502679843
	pesos_i(17228) := b"0000000000000000_0000000000000000_0010000111101110_0100001100001001"; -- 0.13254183734118968
	pesos_i(17229) := b"1111111111111111_1111111111111111_1110111100001000_1100001111011000"; -- -0.06627250645241027
	pesos_i(17230) := b"1111111111111111_1111111111111111_1110011110001111_1100011010110000"; -- -0.09546240043643983
	pesos_i(17231) := b"1111111111111111_1111111111111111_1111100101000101_1000110011110010"; -- -0.026282492599668594
	pesos_i(17232) := b"1111111111111111_1111111111111111_1111110011001110_1110011001100011"; -- -0.012467957444477904
	pesos_i(17233) := b"1111111111111111_1111111111111111_1111011001100011_1101111110001010"; -- -0.037538555977486836
	pesos_i(17234) := b"1111111111111111_1111111111111111_1110100011010110_1000011111100001"; -- -0.09047652010802806
	pesos_i(17235) := b"0000000000000000_0000000000000000_0010010100001000_1100001101111111"; -- 0.14466497285486038
	pesos_i(17236) := b"0000000000000000_0000000000000000_0000010110011101_1100010101110101"; -- 0.02193864931592275
	pesos_i(17237) := b"0000000000000000_0000000000000000_0000100010001001_1110110001101001"; -- 0.0333545453323498
	pesos_i(17238) := b"1111111111111111_1111111111111111_1111010001000011_1101010101000101"; -- -0.04583994937338093
	pesos_i(17239) := b"1111111111111111_1111111111111111_1101111101101110_1001100100110111"; -- -0.12721865086734965
	pesos_i(17240) := b"1111111111111111_1111111111111111_1111101110101110_1010101011110111"; -- -0.016866030293774942
	pesos_i(17241) := b"1111111111111111_1111111111111111_1111110011100000_0010010011101110"; -- -0.012204829999854285
	pesos_i(17242) := b"0000000000000000_0000000000000000_0001111100110001_0000000011101111"; -- 0.12184148642407612
	pesos_i(17243) := b"0000000000000000_0000000000000000_0000101001100101_1110100101000000"; -- 0.04061754047497202
	pesos_i(17244) := b"0000000000000000_0000000000000000_0001100111101010_1101101011011100"; -- 0.10123985157638465
	pesos_i(17245) := b"0000000000000000_0000000000000000_0010010101011101_1110001110011110"; -- 0.14596388442153316
	pesos_i(17246) := b"0000000000000000_0000000000000000_0001000001000111_0000011011001010"; -- 0.0635837786048085
	pesos_i(17247) := b"1111111111111111_1111111111111111_1111001000110011_0111110000000001"; -- -0.053901910462749524
	pesos_i(17248) := b"0000000000000000_0000000000000000_0001110111111100_0010100100100000"; -- 0.11712891611320736
	pesos_i(17249) := b"0000000000000000_0000000000000000_0000010010111001_1011100011101001"; -- 0.018458897581072997
	pesos_i(17250) := b"1111111111111111_1111111111111111_1111101011011000_0010011000100100"; -- -0.020139328214210644
	pesos_i(17251) := b"1111111111111111_1111111111111111_1110110001010100_0110011111000000"; -- -0.0768370778274992
	pesos_i(17252) := b"0000000000000000_0000000000000000_0000100001100110_1010111101011111"; -- 0.03281684931454516
	pesos_i(17253) := b"0000000000000000_0000000000000000_0001101111001010_0011000011101000"; -- 0.10855394042282476
	pesos_i(17254) := b"1111111111111111_1111111111111111_1110100100001100_1101100001100111"; -- -0.08964774599357177
	pesos_i(17255) := b"0000000000000000_0000000000000000_0000111000100001_1010010011001011"; -- 0.05520086256032106
	pesos_i(17256) := b"1111111111111111_1111111111111111_1111000000101111_0110010001101110"; -- -0.061776850901992156
	pesos_i(17257) := b"1111111111111111_1111111111111111_1110101010001010_0100100010010010"; -- -0.08382746154317532
	pesos_i(17258) := b"0000000000000000_0000000000000000_0000000000001011_1010011000110101"; -- 0.00017775347955149493
	pesos_i(17259) := b"1111111111111111_1111111111111111_1111001111011010_1011110010000011"; -- -0.04744359773166156
	pesos_i(17260) := b"0000000000000000_0000000000000000_0001000011111000_1101000100011100"; -- 0.0662966435563572
	pesos_i(17261) := b"0000000000000000_0000000000000000_0001010001110000_1111111000110100"; -- 0.07984913604904949
	pesos_i(17262) := b"1111111111111111_1111111111111111_1111100001010000_0100101100110010"; -- -0.030024814913514154
	pesos_i(17263) := b"1111111111111111_1111111111111111_1110000000010100_1110011011101101"; -- -0.1246810599803759
	pesos_i(17264) := b"0000000000000000_0000000000000000_0000111010100111_1100110100001000"; -- 0.05724793860624539
	pesos_i(17265) := b"0000000000000000_0000000000000000_0001011001100101_0011110110011010"; -- 0.08748230939949939
	pesos_i(17266) := b"1111111111111111_1111111111111111_1111011000000000_0011101100010011"; -- -0.0390589789129572
	pesos_i(17267) := b"1111111111111111_1111111111111111_1110000001111100_1100000010010010"; -- -0.12309643197128288
	pesos_i(17268) := b"0000000000000000_0000000000000000_0000010111111100_0010010101001101"; -- 0.023378688091296757
	pesos_i(17269) := b"1111111111111111_1111111111111111_1111001010010010_0001001000110000"; -- -0.052458632666862716
	pesos_i(17270) := b"1111111111111111_1111111111111111_1111010010000101_0101111101100010"; -- -0.044839895801420115
	pesos_i(17271) := b"0000000000000000_0000000000000000_0000110111111110_0011101011100000"; -- 0.05466049173793988
	pesos_i(17272) := b"0000000000000000_0000000000000000_0001010100010100_1101111001010111"; -- 0.08234967822719241
	pesos_i(17273) := b"1111111111111111_1111111111111111_1111011100100010_1100010101100001"; -- -0.03462568636329221
	pesos_i(17274) := b"0000000000000000_0000000000000000_0001110111100110_0101001000011111"; -- 0.11679566619794406
	pesos_i(17275) := b"1111111111111111_1111111111111111_1110110110001110_0000110000011011"; -- -0.07205128048590044
	pesos_i(17276) := b"0000000000000000_0000000000000000_0001010011110100_0100010101001010"; -- 0.08185227444086082
	pesos_i(17277) := b"0000000000000000_0000000000000000_0001011101000111_0111000000110100"; -- 0.09093381190630541
	pesos_i(17278) := b"1111111111111111_1111111111111111_1111111001111100_0101001101011010"; -- -0.005915442016982947
	pesos_i(17279) := b"1111111111111111_1111111111111111_1111011111110100_1011000100000011"; -- -0.03142255484414006
	pesos_i(17280) := b"0000000000000000_0000000000000000_0001011011100001_0001011101011000"; -- 0.0893721188569172
	pesos_i(17281) := b"1111111111111111_1111111111111111_1110110010101001_1101001111110111"; -- -0.07553363062633549
	pesos_i(17282) := b"1111111111111111_1111111111111111_1110010001000010_0001101000111100"; -- -0.10836635614433186
	pesos_i(17283) := b"1111111111111111_1111111111111111_1110001011001011_1011111110000010"; -- -0.11407855115215991
	pesos_i(17284) := b"0000000000000000_0000000000000000_0000101110011100_0011101110100101"; -- 0.04535267626633805
	pesos_i(17285) := b"1111111111111111_1111111111111111_1111011110101011_0110101110100101"; -- -0.03254058096608373
	pesos_i(17286) := b"1111111111111111_1111111111111111_1110011011010001_1101101100011101"; -- -0.09836035296433543
	pesos_i(17287) := b"0000000000000000_0000000000000000_0001110010001111_1111111101001000"; -- 0.11157222286899773
	pesos_i(17288) := b"0000000000000000_0000000000000000_0000101000101100_0001110101011111"; -- 0.03973563731514843
	pesos_i(17289) := b"0000000000000000_0000000000000000_0001000110010001_1110111011001000"; -- 0.06863300686323416
	pesos_i(17290) := b"0000000000000000_0000000000000000_0000001010001110_1110100101101111"; -- 0.009993161731255982
	pesos_i(17291) := b"0000000000000000_0000000000000000_0001101101001001_1010111101110110"; -- 0.10659310000401358
	pesos_i(17292) := b"1111111111111111_1111111111111111_1111011011101000_1010000110011000"; -- -0.035512829126665174
	pesos_i(17293) := b"0000000000000000_0000000000000000_0010001011000001_1101010100001010"; -- 0.13577014436071266
	pesos_i(17294) := b"0000000000000000_0000000000000000_0001010110000110_1100000110010100"; -- 0.08408746594979818
	pesos_i(17295) := b"0000000000000000_0000000000000000_0000001010001011_1101000000111011"; -- 0.00994588325560161
	pesos_i(17296) := b"1111111111111111_1111111111111111_1110101110100000_0100100100110110"; -- -0.07958548014665222
	pesos_i(17297) := b"1111111111111111_1111111111111111_1110000100001000_1011010111010010"; -- -0.12096084231828882
	pesos_i(17298) := b"0000000000000000_0000000000000000_0000011100100000_1111011000011100"; -- 0.027846700500703148
	pesos_i(17299) := b"0000000000000000_0000000000000000_0010011001100100_1110111101010000"; -- 0.149977642928354
	pesos_i(17300) := b"1111111111111111_1111111111111111_1110011100001000_1011100011100100"; -- -0.09752315939037329
	pesos_i(17301) := b"1111111111111111_1111111111111111_1111011111000111_0101010100101001"; -- -0.032114675112316395
	pesos_i(17302) := b"1111111111111111_1111111111111111_1111010101011000_0001101111111001"; -- -0.04162430933701398
	pesos_i(17303) := b"1111111111111111_1111111111111111_1111100001100000_0101101000011100"; -- -0.029779785202722814
	pesos_i(17304) := b"0000000000000000_0000000000000000_0001010011000011_1111111010100101"; -- 0.08111564196501912
	pesos_i(17305) := b"0000000000000000_0000000000000000_0000111101110010_0010011110111010"; -- 0.06033561987603112
	pesos_i(17306) := b"0000000000000000_0000000000000000_0010001111100101_1011110011100011"; -- 0.14022427127234244
	pesos_i(17307) := b"1111111111111111_1111111111111111_1110000011000010_0111110110111000"; -- -0.12203230143469164
	pesos_i(17308) := b"1111111111111111_1111111111111111_1111010111011101_0110111111010111"; -- -0.039589891506699594
	pesos_i(17309) := b"0000000000000000_0000000000000000_0000110111000110_1010111110000110"; -- 0.05381295222450405
	pesos_i(17310) := b"0000000000000000_0000000000000000_0001000101010011_1111011011100001"; -- 0.06768744453653355
	pesos_i(17311) := b"1111111111111111_1111111111111111_1111001101001000_0111000010000010"; -- -0.04967591129500181
	pesos_i(17312) := b"1111111111111111_1111111111111111_1101110010000000_1110100100111101"; -- -0.1386579729398581
	pesos_i(17313) := b"1111111111111111_1111111111111111_1110000110001001_0011010001111000"; -- -0.1190001684542584
	pesos_i(17314) := b"0000000000000000_0000000000000000_0001110011000001_0101100110011101"; -- 0.11232528761481651
	pesos_i(17315) := b"1111111111111111_1111111111111111_1110001110111100_0100010110010100"; -- -0.11040845057533849
	pesos_i(17316) := b"0000000000000000_0000000000000000_0000001111100111_1010110000100001"; -- 0.015253789888685285
	pesos_i(17317) := b"0000000000000000_0000000000000000_0010000011101001_1100011110100110"; -- 0.12856719785677645
	pesos_i(17318) := b"1111111111111111_1111111111111111_1110111100000001_1110000101111100"; -- -0.06637755138451985
	pesos_i(17319) := b"1111111111111111_1111111111111111_1110100010011011_0100101000101010"; -- -0.0913804671764796
	pesos_i(17320) := b"0000000000000000_0000000000000000_0001111110111111_1010110110101110"; -- 0.12401853080626357
	pesos_i(17321) := b"0000000000000000_0000000000000000_0000011001111101_1101110111111101"; -- 0.025358080262988258
	pesos_i(17322) := b"1111111111111111_1111111111111111_1110010110110101_0110001110100101"; -- -0.10270096983794363
	pesos_i(17323) := b"0000000000000000_0000000000000000_0001110011000001_0011101001000001"; -- 0.11232341841676345
	pesos_i(17324) := b"0000000000000000_0000000000000000_0001010100111100_0111100011000111"; -- 0.08295397623495042
	pesos_i(17325) := b"1111111111111111_1111111111111111_1101100110111000_0111000011000000"; -- -0.14952941236138925
	pesos_i(17326) := b"0000000000000000_0000000000000000_0000011010110101_1110101111001001"; -- 0.02621339465459627
	pesos_i(17327) := b"1111111111111111_1111111111111111_1111111100111001_1010011010010110"; -- -0.0030265697922698875
	pesos_i(17328) := b"0000000000000000_0000000000000000_0001110011101110_0101101101110100"; -- 0.1130120427296894
	pesos_i(17329) := b"0000000000000000_0000000000000000_0010010010111011_0000010001111011"; -- 0.14347866068800827
	pesos_i(17330) := b"1111111111111111_1111111111111111_1110000000000011_0011000011011000"; -- -0.12495131233458387
	pesos_i(17331) := b"0000000000000000_0000000000000000_0000110101010111_0010011001011110"; -- 0.052111051622386016
	pesos_i(17332) := b"1111111111111111_1111111111111111_1111000000101101_1000001110010110"; -- -0.06180551127155546
	pesos_i(17333) := b"0000000000000000_0000000000000000_0010000101011100_0101000010100010"; -- 0.13031486473706186
	pesos_i(17334) := b"1111111111111111_1111111111111111_1110111000110011_0110100011010000"; -- -0.06952805450235676
	pesos_i(17335) := b"0000000000000000_0000000000000000_0001000000011100_1010100111000011"; -- 0.06293736465346582
	pesos_i(17336) := b"0000000000000000_0000000000000000_0000110001101011_1111111100001010"; -- 0.04852289186308064
	pesos_i(17337) := b"0000000000000000_0000000000000000_0010001001111101_0010000000100011"; -- 0.1347217641506264
	pesos_i(17338) := b"0000000000000000_0000000000000000_0000000110010111_1110001110110010"; -- 0.006223898807940606
	pesos_i(17339) := b"1111111111111111_1111111111111111_1111010100000110_1011110110000010"; -- -0.04286590162644676
	pesos_i(17340) := b"1111111111111111_1111111111111111_1110100000111000_1010100101101100"; -- -0.09288540945500842
	pesos_i(17341) := b"1111111111111111_1111111111111111_1111010110011001_0010001010101001"; -- -0.04063208926575512
	pesos_i(17342) := b"1111111111111111_1111111111111111_1110010001100101_0010110110101100"; -- -0.10783114002423466
	pesos_i(17343) := b"0000000000000000_0000000000000000_0001001010100001_0111111111011010"; -- 0.07277678547694007
	pesos_i(17344) := b"0000000000000000_0000000000000000_0000011111100010_1100110101111000"; -- 0.030804483295958807
	pesos_i(17345) := b"1111111111111111_1111111111111111_1101110000000000_0001110110111000"; -- -0.14062322871340252
	pesos_i(17346) := b"0000000000000000_0000000000000000_0001100000111010_0110101110011001"; -- 0.09464142318800745
	pesos_i(17347) := b"0000000000000000_0000000000000000_0001111001011101_0010101100001100"; -- 0.11860913315254554
	pesos_i(17348) := b"1111111111111111_1111111111111111_1111110001000101_0101001101100100"; -- -0.014567173181809171
	pesos_i(17349) := b"1111111111111111_1111111111111111_1101111001100101_1110010110001110"; -- -0.131257679851276
	pesos_i(17350) := b"1111111111111111_1111111111111111_1110010000010110_1101100110010101"; -- -0.10902633776786753
	pesos_i(17351) := b"1111111111111111_1111111111111111_1111110010100000_1001011001110101"; -- -0.01317462585535942
	pesos_i(17352) := b"1111111111111111_1111111111111111_1111111010111001_0100100011100011"; -- -0.004985279687589614
	pesos_i(17353) := b"0000000000000000_0000000000000000_0000100000101011_0111010101111110"; -- 0.031913130998149304
	pesos_i(17354) := b"0000000000000000_0000000000000000_0000000010110011_1011101011111000"; -- 0.0027424674145326558
	pesos_i(17355) := b"1111111111111111_1111111111111111_1111101101000110_1101001110100010"; -- -0.01845052045589903
	pesos_i(17356) := b"0000000000000000_0000000000000000_0010001110111000_0011011011100011"; -- 0.1395296386956596
	pesos_i(17357) := b"0000000000000000_0000000000000000_0001100011010101_1001000100101011"; -- 0.09700877471733761
	pesos_i(17358) := b"1111111111111111_1111111111111111_1101110010101100_0101000001111100"; -- -0.13799569115015525
	pesos_i(17359) := b"1111111111111111_1111111111111111_1110010010110110_0010111001100010"; -- -0.10659513572082996
	pesos_i(17360) := b"0000000000000000_0000000000000000_0010000001110100_1000101111000111"; -- 0.1267783509063647
	pesos_i(17361) := b"0000000000000000_0000000000000000_0000010110011011_1011111000011101"; -- 0.021907693941972638
	pesos_i(17362) := b"0000000000000000_0000000000000000_0001010000000010_1111000011010101"; -- 0.07816987217457631
	pesos_i(17363) := b"0000000000000000_0000000000000000_0001110010101000_1001110111110001"; -- 0.11194789059303752
	pesos_i(17364) := b"1111111111111111_1111111111111111_1110001111010111_1000100011110100"; -- -0.1099924473920346
	pesos_i(17365) := b"1111111111111111_1111111111111111_1111010111100111_1101110101110001"; -- -0.03943077075234703
	pesos_i(17366) := b"1111111111111111_1111111111111111_1111010011010101_0010111101011110"; -- -0.043622054664882184
	pesos_i(17367) := b"1111111111111111_1111111111111111_1111010001000111_1100000101110100"; -- -0.04578009530361647
	pesos_i(17368) := b"0000000000000000_0000000000000000_0001111001000001_0101010001010010"; -- 0.11818434716300888
	pesos_i(17369) := b"1111111111111111_1111111111111111_1111000001011101_1110100000101000"; -- -0.06106709500317707
	pesos_i(17370) := b"0000000000000000_0000000000000000_0001111000001101_1110011011010100"; -- 0.11739962279698443
	pesos_i(17371) := b"1111111111111111_1111111111111111_1111100011100010_1101011000100000"; -- -0.027788750863569238
	pesos_i(17372) := b"1111111111111111_1111111111111111_1110001010010001_1101010111010100"; -- -0.11496223055120605
	pesos_i(17373) := b"1111111111111111_1111111111111111_1111011111101100_1011010110001001"; -- -0.03154435535168188
	pesos_i(17374) := b"0000000000000000_0000000000000000_0000111000010100_0100110000101001"; -- 0.05499721516956702
	pesos_i(17375) := b"1111111111111111_1111111111111111_1111011101011001_0010110111011001"; -- -0.033795485105734734
	pesos_i(17376) := b"0000000000000000_0000000000000000_0010011010100011_0000010100011100"; -- 0.1509249870772197
	pesos_i(17377) := b"1111111111111111_1111111111111111_1111010110110111_1010001101101101"; -- -0.04016665074540962
	pesos_i(17378) := b"0000000000000000_0000000000000000_0001111100000101_0001001001011110"; -- 0.12117113879546389
	pesos_i(17379) := b"1111111111111111_1111111111111111_1110100011110100_1110100111001001"; -- -0.0900129208062055
	pesos_i(17380) := b"0000000000000000_0000000000000000_0000100101011000_1110010011111000"; -- 0.036512671033701635
	pesos_i(17381) := b"1111111111111111_1111111111111111_1110100011100100_0100111000000110"; -- -0.09026634563840828
	pesos_i(17382) := b"1111111111111111_1111111111111111_1111001000100110_0000110100101011"; -- -0.05410688104524206
	pesos_i(17383) := b"1111111111111111_1111111111111111_1110000101010000_0100011010011100"; -- -0.11986883831829381
	pesos_i(17384) := b"0000000000000000_0000000000000000_0000010111101111_0111010011111001"; -- 0.023185072798360944
	pesos_i(17385) := b"1111111111111111_1111111111111111_1101110011001101_0000000000011111"; -- -0.1374969410313434
	pesos_i(17386) := b"0000000000000000_0000000000000000_0000100010001111_0111010010100101"; -- 0.033438959402631835
	pesos_i(17387) := b"1111111111111111_1111111111111111_1110110110101010_0111110100011000"; -- -0.07161729965531712
	pesos_i(17388) := b"1111111111111111_1111111111111111_1101110100111011_1110110011100010"; -- -0.13580436216335678
	pesos_i(17389) := b"1111111111111111_1111111111111111_1101110000110010_0010000001011101"; -- -0.1398601314885088
	pesos_i(17390) := b"1111111111111111_1111111111111111_1101111100100100_1000100101011011"; -- -0.12834874650717978
	pesos_i(17391) := b"1111111111111111_1111111111111111_1110000010010100_1101110010101000"; -- -0.12272854719567874
	pesos_i(17392) := b"0000000000000000_0000000000000000_0001011000010111_0101001111011111"; -- 0.08629345120169411
	pesos_i(17393) := b"1111111111111111_1111111111111111_1101110100011101_0000000011101000"; -- -0.13627619099172789
	pesos_i(17394) := b"1111111111111111_1111111111111111_1111100111100010_1100000001001011"; -- -0.023883802106310484
	pesos_i(17395) := b"1111111111111111_1111111111111111_1110111110010100_1000010000001101"; -- -0.06414007847733272
	pesos_i(17396) := b"1111111111111111_1111111111111111_1111100111100101_1100011101011000"; -- -0.023837605397665735
	pesos_i(17397) := b"0000000000000000_0000000000000000_0010010100011001_1010010100000101"; -- 0.1449225555699619
	pesos_i(17398) := b"1111111111111111_1111111111111111_1111010111111010_1001110011100101"; -- -0.03914470106045993
	pesos_i(17399) := b"1111111111111111_1111111111111111_1110100101100011_1000010001011010"; -- -0.08832524108930041
	pesos_i(17400) := b"0000000000000000_0000000000000000_0000101001100101_0000100001110101"; -- 0.04060414183065246
	pesos_i(17401) := b"0000000000000000_0000000000000000_0000111110001100_0101101010101010"; -- 0.06073538454362098
	pesos_i(17402) := b"1111111111111111_1111111111111111_1111101100010010_1100100010001010"; -- -0.019244638651316925
	pesos_i(17403) := b"1111111111111111_1111111111111111_1101110011111111_1011011010111001"; -- -0.1367231176327419
	pesos_i(17404) := b"0000000000000000_0000000000000000_0001110111110111_0001100100010101"; -- 0.11705166591170875
	pesos_i(17405) := b"0000000000000000_0000000000000000_0001001101100001_1111011011100001"; -- 0.07571356763773908
	pesos_i(17406) := b"0000000000000000_0000000000000000_0001001010010100_1110000110100001"; -- 0.07258424930991725
	pesos_i(17407) := b"0000000000000000_0000000000000000_0000110111001011_1111111011101000"; -- 0.05389397779534703
	pesos_i(17408) := b"0000000000000000_0000000000000000_0010000001000001_0110010101001011"; -- 0.12599785881041223
	pesos_i(17409) := b"0000000000000000_0000000000000000_0000010001011100_1000111101001010"; -- 0.017037349296805636
	pesos_i(17410) := b"1111111111111111_1111111111111111_1111010011100100_0011100101001010"; -- -0.04339258148337712
	pesos_i(17411) := b"1111111111111111_1111111111111111_1111111001001100_0011011000101010"; -- -0.006649603674977172
	pesos_i(17412) := b"0000000000000000_0000000000000000_0000001100001001_1110100001010111"; -- 0.011869927559300698
	pesos_i(17413) := b"0000000000000000_0000000000000000_0000001101101000_1011111011000100"; -- 0.013317034587469067
	pesos_i(17414) := b"1111111111111111_1111111111111111_1110101110010001_1111001011010001"; -- -0.0798042526945165
	pesos_i(17415) := b"1111111111111111_1111111111111111_1111001100001101_0100111101001000"; -- -0.05057816012074492
	pesos_i(17416) := b"1111111111111111_1111111111111111_1110001000010010_0011100100111011"; -- -0.11690943070071892
	pesos_i(17417) := b"0000000000000000_0000000000000000_0000011000000011_1110110001001110"; -- 0.02349736133272362
	pesos_i(17418) := b"1111111111111111_1111111111111111_1110110001100111_1110101000101000"; -- -0.07653938802944409
	pesos_i(17419) := b"1111111111111111_1111111111111111_1110010110111010_0100011001100111"; -- -0.10262641903886105
	pesos_i(17420) := b"1111111111111111_1111111111111111_1110011111100111_0011000100001111"; -- -0.09412854551404455
	pesos_i(17421) := b"0000000000000000_0000000000000000_0000001001100011_0110010100101101"; -- 0.009329150547290567
	pesos_i(17422) := b"0000000000000000_0000000000000000_0000000110110001_0011001100011010"; -- 0.006610101582855934
	pesos_i(17423) := b"0000000000000000_0000000000000000_0001011111101011_0110000101000011"; -- 0.0934353627364655
	pesos_i(17424) := b"1111111111111111_1111111111111111_1111010100001111_1011010111011100"; -- -0.04272902846899575
	pesos_i(17425) := b"0000000000000000_0000000000000000_0010100000111011_0111011101101011"; -- 0.15715738630818296
	pesos_i(17426) := b"0000000000000000_0000000000000000_0000011100111010_1000100101000001"; -- 0.028236940830202423
	pesos_i(17427) := b"0000000000000000_0000000000000000_0001000111100010_1010111001100100"; -- 0.06986513074587465
	pesos_i(17428) := b"0000000000000000_0000000000000000_0001010001111100_0100011000010111"; -- 0.08002126742859027
	pesos_i(17429) := b"0000000000000000_0000000000000000_0010001010110000_0001001010001001"; -- 0.1354991516821487
	pesos_i(17430) := b"1111111111111111_1111111111111111_1111001001111110_0001011000010110"; -- -0.0527635761144275
	pesos_i(17431) := b"1111111111111111_1111111111111111_1110111111010100_0100001100100000"; -- -0.06316738584110562
	pesos_i(17432) := b"0000000000000000_0000000000000000_0001101011110011_0111010010110000"; -- 0.10527734086928543
	pesos_i(17433) := b"1111111111111111_1111111111111111_1110011000111001_1010000111110100"; -- -0.10068309588646687
	pesos_i(17434) := b"0000000000000000_0000000000000000_0001110111011101_0011100111011001"; -- 0.11665689031935389
	pesos_i(17435) := b"1111111111111111_1111111111111111_1110111100000011_0000001010110001"; -- -0.0663603132848993
	pesos_i(17436) := b"1111111111111111_1111111111111111_1111101111100111_0110001111001000"; -- -0.016000522278357965
	pesos_i(17437) := b"0000000000000000_0000000000000000_0001100100010100_0100000001010110"; -- 0.09796526049673773
	pesos_i(17438) := b"1111111111111111_1111111111111111_1110110000011110_0100101010010111"; -- -0.07766279031404481
	pesos_i(17439) := b"1111111111111111_1111111111111111_1110101101110000_1101011101100101"; -- -0.08030942714004097
	pesos_i(17440) := b"0000000000000000_0000000000000000_0001111101000000_0101110100010000"; -- 0.12207585943978903
	pesos_i(17441) := b"1111111111111111_1111111111111111_1110100010010001_1110111101110101"; -- -0.0915232028055998
	pesos_i(17442) := b"1111111111111111_1111111111111111_1111110000111011_1000110000001100"; -- -0.014716384097483071
	pesos_i(17443) := b"1111111111111111_1111111111111111_1110001010010101_1010110011010000"; -- -0.11490363997384481
	pesos_i(17444) := b"1111111111111111_1111111111111111_1101111011110110_0001111101011100"; -- -0.12905696867612784
	pesos_i(17445) := b"1111111111111111_1111111111111111_1111101101110110_0111000101110101"; -- -0.01772395023116137
	pesos_i(17446) := b"1111111111111111_1111111111111111_1111010111100100_0010000100100110"; -- -0.039487770203557815
	pesos_i(17447) := b"0000000000000000_0000000000000000_0001011100000101_0011001100011000"; -- 0.08992308933280489
	pesos_i(17448) := b"0000000000000000_0000000000000000_0001010011011010_0101111100011000"; -- 0.0814570841463503
	pesos_i(17449) := b"0000000000000000_0000000000000000_0000001010100100_1110111100100011"; -- 0.01032919504107813
	pesos_i(17450) := b"1111111111111111_1111111111111111_1101101011001111_0101111001010111"; -- -0.14527330764875965
	pesos_i(17451) := b"0000000000000000_0000000000000000_0001010010001110_1000000011011110"; -- 0.08029942917212596
	pesos_i(17452) := b"0000000000000000_0000000000000000_0010000000101101_1101100010101000"; -- 0.12569955911101188
	pesos_i(17453) := b"0000000000000000_0000000000000000_0000011000011000_0001000100100100"; -- 0.023804732561742255
	pesos_i(17454) := b"1111111111111111_1111111111111111_1111110011111111_0010111110111010"; -- -0.011731164029230747
	pesos_i(17455) := b"0000000000000000_0000000000000000_0001011111100000_0010001111001110"; -- 0.09326385296912412
	pesos_i(17456) := b"1111111111111111_1111111111111111_1110101101100001_1001100110010100"; -- -0.0805419935165995
	pesos_i(17457) := b"0000000000000000_0000000000000000_0010010010001000_1100111000001110"; -- 0.142712477229458
	pesos_i(17458) := b"0000000000000000_0000000000000000_0001000110110001_0100110011110101"; -- 0.06911164269436777
	pesos_i(17459) := b"0000000000000000_0000000000000000_0010010010000110_0100010110000110"; -- 0.14267382157751768
	pesos_i(17460) := b"0000000000000000_0000000000000000_0000101001111100_0001011101101100"; -- 0.04095598587559661
	pesos_i(17461) := b"1111111111111111_1111111111111111_1111001101011000_1010101100110010"; -- -0.04942827263236264
	pesos_i(17462) := b"1111111111111111_1111111111111111_1110111010111011_0110101100011110"; -- -0.06745272166716014
	pesos_i(17463) := b"0000000000000000_0000000000000000_0010010100011110_1100010110000110"; -- 0.1450007869617132
	pesos_i(17464) := b"1111111111111111_1111111111111111_1110011001101001_0100110010101010"; -- -0.09995575759370934
	pesos_i(17465) := b"1111111111111111_1111111111111111_1111110001011110_1011000111101111"; -- -0.014180068054614907
	pesos_i(17466) := b"0000000000000000_0000000000000000_0000000001001100_0111100111111001"; -- 0.0011669381157720009
	pesos_i(17467) := b"0000000000000000_0000000000000000_0001100010000101_1011111110110001"; -- 0.09579084455612949
	pesos_i(17468) := b"0000000000000000_0000000000000000_0001110110111100_0110101100111111"; -- 0.11615629467510362
	pesos_i(17469) := b"1111111111111111_1111111111111111_1110100101011101_0011000011100111"; -- -0.08842176781635316
	pesos_i(17470) := b"0000000000000000_0000000000000000_0001111111101001_0111110100110000"; -- 0.12465650969508865
	pesos_i(17471) := b"0000000000000000_0000000000000000_0000110100010000_0101100110010011"; -- 0.05103072977892501
	pesos_i(17472) := b"1111111111111111_1111111111111111_1110111001100111_0001001000010111"; -- -0.06873976655859014
	pesos_i(17473) := b"1111111111111111_1111111111111111_1101110110101000_0100000001000101"; -- -0.13415144278086588
	pesos_i(17474) := b"1111111111111111_1111111111111111_1111010000110011_0011110101111100"; -- -0.04609313703528555
	pesos_i(17475) := b"0000000000000000_0000000000000000_0001101100111001_0011000100010101"; -- 0.10634142643485407
	pesos_i(17476) := b"0000000000000000_0000000000000000_0010000001110110_1101111101001001"; -- 0.12681384603396553
	pesos_i(17477) := b"0000000000000000_0000000000000000_0000011101100110_1101011100001001"; -- 0.028912963596326655
	pesos_i(17478) := b"1111111111111111_1111111111111111_1111110000111101_0110011001001001"; -- -0.014688117219973247
	pesos_i(17479) := b"0000000000000000_0000000000000000_0001000010111110_1101011100100011"; -- 0.0654119929727805
	pesos_i(17480) := b"0000000000000000_0000000000000000_0010000011110011_0111101000000011"; -- 0.12871515809231457
	pesos_i(17481) := b"1111111111111111_1111111111111111_1111110010000101_1010011101110110"; -- -0.013585599594603672
	pesos_i(17482) := b"1111111111111111_1111111111111111_1111111100101110_0001011001110011"; -- -0.0032030076053245642
	pesos_i(17483) := b"0000000000000000_0000000000000000_0001110110001101_0110001001101111"; -- 0.11543860644841929
	pesos_i(17484) := b"1111111111111111_1111111111111111_1110011101110011_1111100101011010"; -- -0.09588662663560749
	pesos_i(17485) := b"1111111111111111_1111111111111111_1111111000001000_0111100100011101"; -- -0.007683210880982236
	pesos_i(17486) := b"0000000000000000_0000000000000000_0001110110011110_0011101001010110"; -- 0.11569561583884119
	pesos_i(17487) := b"1111111111111111_1111111111111111_1110101110000111_0011111101000000"; -- -0.07996754342540237
	pesos_i(17488) := b"0000000000000000_0000000000000000_0001010110001101_1011110101001011"; -- 0.08419402200264678
	pesos_i(17489) := b"0000000000000000_0000000000000000_0000000100010100_1110001000111000"; -- 0.004224909477913598
	pesos_i(17490) := b"0000000000000000_0000000000000000_0010000111100110_1100110010100101"; -- 0.1324279692405129
	pesos_i(17491) := b"1111111111111111_1111111111111111_1110001111000000_1110001010101000"; -- -0.11033805281845038
	pesos_i(17492) := b"0000000000000000_0000000000000000_0000001001101011_0111100100011001"; -- 0.009452408385986577
	pesos_i(17493) := b"1111111111111111_1111111111111111_1111001001010110_1011000010110001"; -- -0.05336471251815542
	pesos_i(17494) := b"0000000000000000_0000000000000000_0010000011011101_1001101001101001"; -- 0.12838139592247616
	pesos_i(17495) := b"0000000000000000_0000000000000000_0000110110010111_0000001101101111"; -- 0.05308553171936846
	pesos_i(17496) := b"0000000000000000_0000000000000000_0001100110001001_0001011010000110"; -- 0.09974804655759616
	pesos_i(17497) := b"0000000000000000_0000000000000000_0000110101001010_1001011110101001"; -- 0.05191944004542677
	pesos_i(17498) := b"1111111111111111_1111111111111111_1110110001111100_1110001110110000"; -- -0.07621933891277814
	pesos_i(17499) := b"0000000000000000_0000000000000000_0010010010011011_0110111110000100"; -- 0.142996759130933
	pesos_i(17500) := b"0000000000000000_0000000000000000_0001001111110000_1001010011100010"; -- 0.07788973337307102
	pesos_i(17501) := b"1111111111111111_1111111111111111_1110111101000100_0001100000111100"; -- -0.06536720786674483
	pesos_i(17502) := b"0000000000000000_0000000000000000_0000011011010000_0100011110110100"; -- 0.026615602075801367
	pesos_i(17503) := b"1111111111111111_1111111111111111_1111000000000110_1111100000010001"; -- -0.062393661405527066
	pesos_i(17504) := b"0000000000000000_0000000000000000_0000010010111010_0011110110000011"; -- 0.018466801257321426
	pesos_i(17505) := b"1111111111111111_1111111111111111_1110101100011101_0101001111000110"; -- -0.08158375180351407
	pesos_i(17506) := b"1111111111111111_1111111111111111_1101111111010001_1111110011111111"; -- -0.12570208339381514
	pesos_i(17507) := b"1111111111111111_1111111111111111_1111000010000100_0010110010001110"; -- -0.0604831841076724
	pesos_i(17508) := b"0000000000000000_0000000000000000_0000110101111100_0111101010101001"; -- 0.05268065094328475
	pesos_i(17509) := b"0000000000000000_0000000000000000_0000101110110010_1110000111110101"; -- 0.045698282427332884
	pesos_i(17510) := b"1111111111111111_1111111111111111_1111001110100011_0001110010100101"; -- -0.048292359975649055
	pesos_i(17511) := b"1111111111111111_1111111111111111_1110100011110001_0001111010101000"; -- -0.09007080452947525
	pesos_i(17512) := b"0000000000000000_0000000000000000_0000000100101010_1101001110011001"; -- 0.004559731438710393
	pesos_i(17513) := b"1111111111111111_1111111111111111_1101111110001111_0001100111000010"; -- -0.12672270795760615
	pesos_i(17514) := b"0000000000000000_0000000000000000_0001011000000001_1110100001111111"; -- 0.08596661657355972
	pesos_i(17515) := b"1111111111111111_1111111111111111_1111101101001111_1010110110101001"; -- -0.018315454636715696
	pesos_i(17516) := b"0000000000000000_0000000000000000_0001100010101111_0110110100101010"; -- 0.0964267946938762
	pesos_i(17517) := b"0000000000000000_0000000000000000_0000101001000010_1101000000011100"; -- 0.040081984288467876
	pesos_i(17518) := b"1111111111111111_1111111111111111_1111001100110010_1010000000011000"; -- -0.050008768277994914
	pesos_i(17519) := b"1111111111111111_1111111111111111_1111000000010001_0000000101101101"; -- -0.06224051563851
	pesos_i(17520) := b"0000000000000000_0000000000000000_0000011001010000_0110000111111000"; -- 0.02466404259183307
	pesos_i(17521) := b"0000000000000000_0000000000000000_0001111101001010_0111010000001110"; -- 0.12222981775058424
	pesos_i(17522) := b"1111111111111111_1111111111111111_1111101110000111_1010001011100111"; -- -0.017461603634449162
	pesos_i(17523) := b"1111111111111111_1111111111111111_1111000010111110_1111011111011100"; -- -0.05958605655824282
	pesos_i(17524) := b"0000000000000000_0000000000000000_0001111000010101_0101110010001111"; -- 0.11751345149103236
	pesos_i(17525) := b"0000000000000000_0000000000000000_0000100010011001_0110001001100100"; -- 0.033590459366701325
	pesos_i(17526) := b"0000000000000000_0000000000000000_0010000101000001_0000001011001110"; -- 0.12989823844980036
	pesos_i(17527) := b"1111111111111111_1111111111111111_1110110111111001_0110111101011110"; -- -0.07041267344912441
	pesos_i(17528) := b"1111111111111111_1111111111111111_1110101110101000_1011000100100000"; -- -0.07945721605422587
	pesos_i(17529) := b"0000000000000000_0000000000000000_0001000011111110_1000010111000001"; -- 0.06638370469789749
	pesos_i(17530) := b"0000000000000000_0000000000000000_0000010010010100_0000100100101100"; -- 0.017883847403041
	pesos_i(17531) := b"0000000000000000_0000000000000000_0000010110001011_1011110001010000"; -- 0.02166344594836615
	pesos_i(17532) := b"0000000000000000_0000000000000000_0000011000000111_1001001000110110"; -- 0.023553026373765218
	pesos_i(17533) := b"0000000000000000_0000000000000000_0001001001101000_1111001010001001"; -- 0.07191387024735693
	pesos_i(17534) := b"1111111111111111_1111111111111111_1111000111110010_0000101010001010"; -- -0.054900494868476604
	pesos_i(17535) := b"0000000000000000_0000000000000000_0010011010111000_0011111110100000"; -- 0.1512489094636539
	pesos_i(17536) := b"1111111111111111_1111111111111111_1110101011100110_0001000010000110"; -- -0.0824269936005528
	pesos_i(17537) := b"1111111111111111_1111111111111111_1110110101010011_1001000111110111"; -- -0.07294357038725789
	pesos_i(17538) := b"0000000000000000_0000000000000000_0000111101111111_0001000110101011"; -- 0.06053266937700322
	pesos_i(17539) := b"0000000000000000_0000000000000000_0000110001110100_1101001111001110"; -- 0.048657644060887684
	pesos_i(17540) := b"1111111111111111_1111111111111111_1101111001111000_1000110111001011"; -- -0.1309729937293191
	pesos_i(17541) := b"0000000000000000_0000000000000000_0000110100111001_1100111010011011"; -- 0.0516633157154613
	pesos_i(17542) := b"0000000000000000_0000000000000000_0000110000000000_0010010011001011"; -- 0.0468771931086062
	pesos_i(17543) := b"0000000000000000_0000000000000000_0001101001111011_1000110101000011"; -- 0.1034477508499686
	pesos_i(17544) := b"0000000000000000_0000000000000000_0001000100110101_0100110011111000"; -- 0.06721955360761711
	pesos_i(17545) := b"1111111111111111_1111111111111111_1110000101010100_1111111010001011"; -- -0.11979683987949014
	pesos_i(17546) := b"1111111111111111_1111111111111111_1110000001110001_0101011100010110"; -- -0.12327056604898785
	pesos_i(17547) := b"0000000000000000_0000000000000000_0010010100001011_0100100001011001"; -- 0.14470340884257185
	pesos_i(17548) := b"0000000000000000_0000000000000000_0010010011101100_1010111111010001"; -- 0.14423655378775133
	pesos_i(17549) := b"0000000000000000_0000000000000000_0000010101010101_1101110111000010"; -- 0.02084146488984267
	pesos_i(17550) := b"1111111111111111_1111111111111111_1110000010100101_0111101000100111"; -- -0.12247501889252062
	pesos_i(17551) := b"0000000000000000_0000000000000000_0010010110101000_0001100101010100"; -- 0.14709623617043674
	pesos_i(17552) := b"0000000000000000_0000000000000000_0000111101111101_0000111110001001"; -- 0.06050202467179663
	pesos_i(17553) := b"1111111111111111_1111111111111111_1111110110000110_1101000101101011"; -- -0.009661590007644561
	pesos_i(17554) := b"0000000000000000_0000000000000000_0000100010100010_1001100111101101"; -- 0.03373109851259229
	pesos_i(17555) := b"0000000000000000_0000000000000000_0001011000110001_1111011000101101"; -- 0.08669985381385559
	pesos_i(17556) := b"1111111111111111_1111111111111111_1111111100100100_1011010100101110"; -- -0.0033461343902637776
	pesos_i(17557) := b"0000000000000000_0000000000000000_0001111110101100_1100000111001110"; -- 0.123729813293297
	pesos_i(17558) := b"0000000000000000_0000000000000000_0000000110011000_0100110101110011"; -- 0.006230202224485023
	pesos_i(17559) := b"1111111111111111_1111111111111111_1101100101000101_1100001110000101"; -- -0.1512792395893646
	pesos_i(17560) := b"1111111111111111_1111111111111111_1110011010000000_0110110011011001"; -- -0.09960288712236388
	pesos_i(17561) := b"0000000000000000_0000000000000000_0001100101011111_0111011110101101"; -- 0.099112968170867
	pesos_i(17562) := b"0000000000000000_0000000000000000_0001110100010110_1000110000011011"; -- 0.11362529423682559
	pesos_i(17563) := b"0000000000000000_0000000000000000_0000000001010100_0000111011110001"; -- 0.0012826288105762958
	pesos_i(17564) := b"1111111111111111_1111111111111111_1111001110111110_0000100100110111"; -- -0.04788153086729079
	pesos_i(17565) := b"0000000000000000_0000000000000000_0001100110010101_1111011101110010"; -- 0.099944558538668
	pesos_i(17566) := b"0000000000000000_0000000000000000_0000001011000101_1010110100111111"; -- 0.01082880774319984
	pesos_i(17567) := b"0000000000000000_0000000000000000_0001110111101111_0000101100100110"; -- 0.11692876500898321
	pesos_i(17568) := b"0000000000000000_0000000000000000_0010001010010111_1001100011011111"; -- 0.13512568897409555
	pesos_i(17569) := b"0000000000000000_0000000000000000_0001110010110000_0010011000001111"; -- 0.11206281527363543
	pesos_i(17570) := b"1111111111111111_1111111111111111_1111010010110011_0100110101000110"; -- -0.044139070824057554
	pesos_i(17571) := b"1111111111111111_1111111111111111_1111000011010111_0011101011111001"; -- -0.05921584527856845
	pesos_i(17572) := b"0000000000000000_0000000000000000_0001011101110000_1000010001101001"; -- 0.09156062655875227
	pesos_i(17573) := b"0000000000000000_0000000000000000_0001100111001110_0001000011100000"; -- 0.10080056648348237
	pesos_i(17574) := b"1111111111111111_1111111111111111_1111010110001111_1010000011101001"; -- -0.04077715217556028
	pesos_i(17575) := b"0000000000000000_0000000000000000_0000110101000011_1101111010010100"; -- 0.05181685544986227
	pesos_i(17576) := b"0000000000000000_0000000000000000_0000011111111010_0110000111110110"; -- 0.031164286255016754
	pesos_i(17577) := b"1111111111111111_1111111111111111_1111101011111111_0101100001010010"; -- -0.019541244506341225
	pesos_i(17578) := b"1111111111111111_1111111111111111_1110001011001100_1010001101000000"; -- -0.11406497659441768
	pesos_i(17579) := b"1111111111111111_1111111111111111_1110101101001001_0101110001100000"; -- -0.08091185244008105
	pesos_i(17580) := b"0000000000000000_0000000000000000_0010000011100001_1110100001111110"; -- 0.12844708506224695
	pesos_i(17581) := b"0000000000000000_0000000000000000_0010000111110001_0111100110000011"; -- 0.13259086081040267
	pesos_i(17582) := b"1111111111111111_1111111111111111_1111111111001001_0011110110101000"; -- -0.0008355583874728337
	pesos_i(17583) := b"0000000000000000_0000000000000000_0000111100110011_1110100110011100"; -- 0.05938587244921707
	pesos_i(17584) := b"0000000000000000_0000000000000000_0001110110100100_0111110101110001"; -- 0.11579116821243467
	pesos_i(17585) := b"1111111111111111_1111111111111111_1110001010010000_0100001110001000"; -- -0.11498620912001836
	pesos_i(17586) := b"0000000000000000_0000000000000000_0000100001110011_1000001001110010"; -- 0.03301253590762599
	pesos_i(17587) := b"0000000000000000_0000000000000000_0000010101100111_0000110100100100"; -- 0.02110368843137411
	pesos_i(17588) := b"0000000000000000_0000000000000000_0010001010001010_0011101011100101"; -- 0.13492172336366767
	pesos_i(17589) := b"0000000000000000_0000000000000000_0001100101001000_1100100101111010"; -- 0.09876689164616206
	pesos_i(17590) := b"0000000000000000_0000000000000000_0001100110010111_1110101001100001"; -- 0.09997429712936594
	pesos_i(17591) := b"0000000000000000_0000000000000000_0000110010110110_1101011110001000"; -- 0.049664946211576536
	pesos_i(17592) := b"0000000000000000_0000000000000000_0010010011001011_1000000101100001"; -- 0.14373024583686345
	pesos_i(17593) := b"1111111111111111_1111111111111111_1111101110101000_1100010100011100"; -- -0.01695602470442538
	pesos_i(17594) := b"0000000000000000_0000000000000000_0001100011001101_0110000001101110"; -- 0.09688379939814104
	pesos_i(17595) := b"0000000000000000_0000000000000000_0001001100011001_1000110011110001"; -- 0.07460862047347154
	pesos_i(17596) := b"1111111111111111_1111111111111111_1110001110010011_1100111000011100"; -- -0.1110259228952051
	pesos_i(17597) := b"1111111111111111_1111111111111111_1110011100101101_1110011100001100"; -- -0.09695583298249559
	pesos_i(17598) := b"1111111111111111_1111111111111111_1111010000110110_1001110100101010"; -- -0.046041657651460316
	pesos_i(17599) := b"0000000000000000_0000000000000000_0010011101110100_0101110110100010"; -- 0.15411935041364644
	pesos_i(17600) := b"1111111111111111_1111111111111111_1111101110011010_1010110010111100"; -- -0.017171100736463413
	pesos_i(17601) := b"1111111111111111_1111111111111111_1111100100110110_0000010000101011"; -- -0.02651952698280279
	pesos_i(17602) := b"0000000000000000_0000000000000000_0000101111001110_0101101010010100"; -- 0.04611745951498217
	pesos_i(17603) := b"1111111111111111_1111111111111111_1110101000101111_1100001110101101"; -- -0.08520867376875077
	pesos_i(17604) := b"0000000000000000_0000000000000000_0010010100001010_1100010110101101"; -- 0.1446956202526898
	pesos_i(17605) := b"0000000000000000_0000000000000000_0000000101100111_1010101101000000"; -- 0.00548811253890905
	pesos_i(17606) := b"1111111111111111_1111111111111111_1111011101010111_1011010100111101"; -- -0.033817932733865234
	pesos_i(17607) := b"1111111111111111_1111111111111111_1111111111000000_0110000010001011"; -- -0.0009708080126302399
	pesos_i(17608) := b"0000000000000000_0000000000000000_0001011011100111_0010110110010111"; -- 0.08946499755844493
	pesos_i(17609) := b"1111111111111111_1111111111111111_1110100001000101_0001011010001100"; -- -0.09269579967081581
	pesos_i(17610) := b"1111111111111111_1111111111111111_1110111100001101_1100110110011001"; -- -0.06619563116590896
	pesos_i(17611) := b"1111111111111111_1111111111111111_1111101110110010_1111111000000010"; -- -0.016800045394268888
	pesos_i(17612) := b"1111111111111111_1111111111111111_1110110010011101_1010011110111010"; -- -0.07571937290120845
	pesos_i(17613) := b"1111111111111111_1111111111111111_1101110000011111_0101010000000101"; -- -0.1401469696291789
	pesos_i(17614) := b"1111111111111111_1111111111111111_1111101100010000_1101111110010011"; -- -0.019273783281461107
	pesos_i(17615) := b"1111111111111111_1111111111111111_1111001000010101_0110000100001011"; -- -0.05436128126230909
	pesos_i(17616) := b"1111111111111111_1111111111111111_1101100111001101_1100110010000101"; -- -0.14920350786880635
	pesos_i(17617) := b"1111111111111111_1111111111111111_1110001111000011_1011111011110101"; -- -0.11029440424881413
	pesos_i(17618) := b"0000000000000000_0000000000000000_0001000011101110_1111001111101000"; -- 0.06614612984885504
	pesos_i(17619) := b"1111111111111111_1111111111111111_1110011101000001_0111001011001011"; -- -0.09665758647015708
	pesos_i(17620) := b"1111111111111111_1111111111111111_1101100111111111_1100001111011011"; -- -0.1484410848990893
	pesos_i(17621) := b"0000000000000000_0000000000000000_0001001100100111_1100011000111111"; -- 0.07482565909864858
	pesos_i(17622) := b"1111111111111111_1111111111111111_1110110101001010_1001000001010001"; -- -0.07308099773383896
	pesos_i(17623) := b"0000000000000000_0000000000000000_0000111101000011_1011110101110101"; -- 0.059627381281998744
	pesos_i(17624) := b"0000000000000000_0000000000000000_0000101011101111_1101011000011111"; -- 0.04272211319513259
	pesos_i(17625) := b"1111111111111111_1111111111111111_1111111011110110_1000100101010000"; -- -0.004050653423213574
	pesos_i(17626) := b"0000000000000000_0000000000000000_0001111111000110_0111000100110100"; -- 0.12412173762430646
	pesos_i(17627) := b"1111111111111111_1111111111111111_1101101110110000_1001111101110111"; -- -0.14183619822625493
	pesos_i(17628) := b"0000000000000000_0000000000000000_0001110010110110_0001011011000000"; -- 0.11215345571458485
	pesos_i(17629) := b"1111111111111111_1111111111111111_1101110000010100_0001011101100000"; -- -0.14031843095857216
	pesos_i(17630) := b"0000000000000000_0000000000000000_0001001001000010_1110000101110111"; -- 0.07133301881674342
	pesos_i(17631) := b"1111111111111111_1111111111111111_1111100110011011_0001111001010001"; -- -0.02497683063326364
	pesos_i(17632) := b"0000000000000000_0000000000000000_0001010111010111_0101010011111111"; -- 0.08531695590666871
	pesos_i(17633) := b"0000000000000000_0000000000000000_0000000101010101_1010111000100011"; -- 0.005213626427995418
	pesos_i(17634) := b"1111111111111111_1111111111111111_1111101101010101_0110000011100101"; -- -0.018228477497206925
	pesos_i(17635) := b"0000000000000000_0000000000000000_0000011111010010_1111010001000010"; -- 0.03056265452393781
	pesos_i(17636) := b"0000000000000000_0000000000000000_0010001010001111_1101000001100101"; -- 0.13500692811734483
	pesos_i(17637) := b"0000000000000000_0000000000000000_0000100010001100_0101010111101010"; -- 0.03339135126448249
	pesos_i(17638) := b"0000000000000000_0000000000000000_0001000001001010_0010111111101000"; -- 0.06363200573301785
	pesos_i(17639) := b"1111111111111111_1111111111111111_1110110111101100_1001111100100001"; -- -0.07060819090434087
	pesos_i(17640) := b"0000000000000000_0000000000000000_0000111100001001_0011111011000110"; -- 0.058734820646322204
	pesos_i(17641) := b"1111111111111111_1111111111111111_1110000110000101_0110100000110110"; -- -0.11905811970558276
	pesos_i(17642) := b"0000000000000000_0000000000000000_0001001101001100_1111000110110001"; -- 0.07539282385032685
	pesos_i(17643) := b"0000000000000000_0000000000000000_0010000011111111_1111010001110111"; -- 0.12890556236910902
	pesos_i(17644) := b"1111111111111111_1111111111111111_1111010010111010_0110101110110110"; -- -0.04403044520454606
	pesos_i(17645) := b"1111111111111111_1111111111111111_1111010110010000_0100110111101100"; -- -0.04076683994933711
	pesos_i(17646) := b"1111111111111111_1111111111111111_1111011001010111_1001000100110001"; -- -0.03772633117975565
	pesos_i(17647) := b"0000000000000000_0000000000000000_0010011001100100_1111100001001100"; -- 0.14997817848800107
	pesos_i(17648) := b"1111111111111111_1111111111111111_1111101101110011_1001101110011011"; -- -0.017767214436677968
	pesos_i(17649) := b"1111111111111111_1111111111111111_1101110000101101_1111100000011100"; -- -0.13992356610849907
	pesos_i(17650) := b"0000000000000000_0000000000000000_0000100110010111_0110110011110011"; -- 0.03746682105748901
	pesos_i(17651) := b"0000000000000000_0000000000000000_0000010001110011_1111111011011101"; -- 0.017394951673650856
	pesos_i(17652) := b"1111111111111111_1111111111111111_1111000101011100_0100011001000101"; -- -0.05718575300386697
	pesos_i(17653) := b"1111111111111111_1111111111111111_1111010000111010_0010010001011010"; -- -0.045987823473149995
	pesos_i(17654) := b"0000000000000000_0000000000000000_0000100111101101_0111111110010001"; -- 0.038780186594752186
	pesos_i(17655) := b"0000000000000000_0000000000000000_0001001000101100_1111011000001111"; -- 0.07099855306335402
	pesos_i(17656) := b"1111111111111111_1111111111111111_1110110101101011_1111101010010000"; -- -0.07257112482175133
	pesos_i(17657) := b"1111111111111111_1111111111111111_1101111000011001_1111111010011111"; -- -0.13241585358022792
	pesos_i(17658) := b"1111111111111111_1111111111111111_1110010111101101_1011011110111011"; -- -0.10184146589642636
	pesos_i(17659) := b"0000000000000000_0000000000000000_0001100010110111_1110110011110011"; -- 0.09655648178054188
	pesos_i(17660) := b"1111111111111111_1111111111111111_1110010100001100_0101101111101110"; -- -0.10528016513580545
	pesos_i(17661) := b"1111111111111111_1111111111111111_1111100000110101_1010010000111101"; -- -0.03043149483029126
	pesos_i(17662) := b"0000000000000000_0000000000000000_0000100011101110_1011001111001010"; -- 0.03489230798065553
	pesos_i(17663) := b"1111111111111111_1111111111111111_1101101100001000_0100110101010110"; -- -0.14440457015918132
	pesos_i(17664) := b"0000000000000000_0000000000000000_0000000011000110_1101110011011111"; -- 0.0030344052213444723
	pesos_i(17665) := b"1111111111111111_1111111111111111_1110101101011101_1000111111101010"; -- -0.080603604594893
	pesos_i(17666) := b"1111111111111111_1111111111111111_1110110000110000_1100110100111101"; -- -0.07738034494688023
	pesos_i(17667) := b"0000000000000000_0000000000000000_0000100011000011_1010001010000010"; -- 0.034235150195413545
	pesos_i(17668) := b"0000000000000000_0000000000000000_0000000110001010_1010010011001000"; -- 0.006021784577990407
	pesos_i(17669) := b"0000000000000000_0000000000000000_0000011111010111_1000001110011101"; -- 0.030632234432863663
	pesos_i(17670) := b"0000000000000000_0000000000000000_0001011001110110_0101000100010100"; -- 0.08774286982617956
	pesos_i(17671) := b"1111111111111111_1111111111111111_1110010111100010_1100110111101101"; -- -0.10200798955237009
	pesos_i(17672) := b"1111111111111111_1111111111111111_1111111110110010_0010000100100100"; -- -0.00118821026390189
	pesos_i(17673) := b"0000000000000000_0000000000000000_0000011111100101_0011100100101010"; -- 0.030841419891995365
	pesos_i(17674) := b"1111111111111111_1111111111111111_1110010000000010_1100011011000111"; -- -0.10933263446469867
	pesos_i(17675) := b"1111111111111111_1111111111111111_1110011110110011_1101001011010000"; -- -0.09491236125693023
	pesos_i(17676) := b"1111111111111111_1111111111111111_1101110110001010_1011111110111011"; -- -0.13460160910157956
	pesos_i(17677) := b"1111111111111111_1111111111111111_1110111001010011_0100111011010001"; -- -0.06904132266610088
	pesos_i(17678) := b"1111111111111111_1111111111111111_1111001101010100_1101101001001001"; -- -0.04948650087967925
	pesos_i(17679) := b"0000000000000000_0000000000000000_0000010100000110_0000101101001010"; -- 0.019623475609887114
	pesos_i(17680) := b"1111111111111111_1111111111111111_1111010111101001_0010010100000010"; -- -0.0394112463335512
	pesos_i(17681) := b"0000000000000000_0000000000000000_0000111100100011_1011010011111001"; -- 0.05913859443368878
	pesos_i(17682) := b"1111111111111111_1111111111111111_1110101110011100_0100011111011110"; -- -0.07964659517820977
	pesos_i(17683) := b"1111111111111111_1111111111111111_1111010011100011_1010111100010110"; -- -0.043400818977471375
	pesos_i(17684) := b"1111111111111111_1111111111111111_1110111110010111_0011011011011100"; -- -0.06409890296626738
	pesos_i(17685) := b"0000000000000000_0000000000000000_0000010001010000_0100011111110010"; -- 0.016849991510022286
	pesos_i(17686) := b"0000000000000000_0000000000000000_0010011011111001_1110001011110101"; -- 0.15225046628269426
	pesos_i(17687) := b"0000000000000000_0000000000000000_0001001000001110_0001100101101110"; -- 0.07052763887651826
	pesos_i(17688) := b"0000000000000000_0000000000000000_0000001100000101_0010100100011010"; -- 0.011797493813105972
	pesos_i(17689) := b"1111111111111111_1111111111111111_1111010010010101_0110010111110100"; -- -0.04459536366245752
	pesos_i(17690) := b"1111111111111111_1111111111111111_1110110100100100_0101010000011000"; -- -0.07366442127771118
	pesos_i(17691) := b"1111111111111111_1111111111111111_1110111111001010_0100100001101111"; -- -0.06331965723173597
	pesos_i(17692) := b"1111111111111111_1111111111111111_1111000101001011_1110000001001010"; -- -0.057435972051827225
	pesos_i(17693) := b"1111111111111111_1111111111111111_1111101010110110_1110000001111111"; -- -0.02064701940739398
	pesos_i(17694) := b"1111111111111111_1111111111111111_1101111001100110_1010001011000011"; -- -0.13124640215149963
	pesos_i(17695) := b"1111111111111111_1111111111111111_1110001000101101_0011011010011000"; -- -0.11649760040659904
	pesos_i(17696) := b"0000000000000000_0000000000000000_0010001100111000_0001100111000010"; -- 0.13757477747623167
	pesos_i(17697) := b"1111111111111111_1111111111111111_1101100010100011_1110011100011010"; -- -0.15374904276140883
	pesos_i(17698) := b"0000000000000000_0000000000000000_0001011010001011_0011100000000110"; -- 0.08806181084417787
	pesos_i(17699) := b"1111111111111111_1111111111111111_1101101101100100_1000111101011101"; -- -0.1429968259822875
	pesos_i(17700) := b"1111111111111111_1111111111111111_1111101010111100_1110100110101100"; -- -0.020554919760325457
	pesos_i(17701) := b"0000000000000000_0000000000000000_0001101011111101_1100010110111001"; -- 0.1054347589071187
	pesos_i(17702) := b"1111111111111111_1111111111111111_1110001101110101_0100111111001011"; -- -0.1114912157627965
	pesos_i(17703) := b"0000000000000000_0000000000000000_0010001000110000_1100101101100110"; -- 0.13355704527207116
	pesos_i(17704) := b"0000000000000000_0000000000000000_0001010111011111_0100101111100101"; -- 0.08543848373386459
	pesos_i(17705) := b"1111111111111111_1111111111111111_1111111000010111_1011111100110001"; -- -0.007450151852539827
	pesos_i(17706) := b"0000000000000000_0000000000000000_0001011001110011_1001101011010011"; -- 0.0877014889404214
	pesos_i(17707) := b"0000000000000000_0000000000000000_0000111100001101_0001110110101011"; -- 0.058793882722314526
	pesos_i(17708) := b"1111111111111111_1111111111111111_1110101001101101_1101001001101010"; -- -0.0842617502535938
	pesos_i(17709) := b"0000000000000000_0000000000000000_0001110101111110_1001111101000110"; -- 0.11521335085502857
	pesos_i(17710) := b"1111111111111111_1111111111111111_1111010010101000_0010111100000011"; -- -0.04430872134386599
	pesos_i(17711) := b"0000000000000000_0000000000000000_0010011101111001_1101000110101010"; -- 0.1542025605401058
	pesos_i(17712) := b"1111111111111111_1111111111111111_1101111111011101_1101000001010011"; -- -0.12552164043906214
	pesos_i(17713) := b"1111111111111111_1111111111111111_1110011101111110_0100111111010111"; -- -0.09572888372221053
	pesos_i(17714) := b"1111111111111111_1111111111111111_1111001011010010_1011001101110110"; -- -0.05147245763071411
	pesos_i(17715) := b"1111111111111111_1111111111111111_1110000100010010_1110011100011011"; -- -0.12080531682403209
	pesos_i(17716) := b"1111111111111111_1111111111111111_1111001001001000_0111101111100110"; -- -0.05358148228746308
	pesos_i(17717) := b"1111111111111111_1111111111111111_1111101001000010_0100101111011011"; -- -0.022425898610184822
	pesos_i(17718) := b"0000000000000000_0000000000000000_0010000110110111_1001101010111010"; -- 0.13170783089187205
	pesos_i(17719) := b"1111111111111111_1111111111111111_1111100111101010_0010011001111011"; -- -0.023770899726130522
	pesos_i(17720) := b"1111111111111111_1111111111111111_1111010111010101_1100110100111100"; -- -0.0397063951186075
	pesos_i(17721) := b"0000000000000000_0000000000000000_0000010111010010_1101010100011000"; -- 0.02274829699459798
	pesos_i(17722) := b"0000000000000000_0000000000000000_0000110001110110_1110110011010001"; -- 0.048689652388562994
	pesos_i(17723) := b"1111111111111111_1111111111111111_1101101011101111_1111111010101011"; -- -0.14477547009534822
	pesos_i(17724) := b"1111111111111111_1111111111111111_1110110101100101_1110101000110101"; -- -0.07266365247450239
	pesos_i(17725) := b"1111111111111111_1111111111111111_1111111000101000_0000010100100111"; -- -0.007201841320045428
	pesos_i(17726) := b"1111111111111111_1111111111111111_1101100101011101_0101000001101111"; -- -0.1509198884310904
	pesos_i(17727) := b"1111111111111111_1111111111111111_1111000100010100_1011001001010111"; -- -0.05827794436164392
	pesos_i(17728) := b"0000000000000000_0000000000000000_0001110111010010_1001000110001101"; -- 0.11649427127885305
	pesos_i(17729) := b"1111111111111111_1111111111111111_1101110110010000_0110101101110111"; -- -0.13451507888706118
	pesos_i(17730) := b"1111111111111111_1111111111111111_1110001001001100_0111110011001000"; -- -0.1160203945331602
	pesos_i(17731) := b"0000000000000000_0000000000000000_0000011000010100_0101000010011110"; -- 0.023747480912116183
	pesos_i(17732) := b"1111111111111111_1111111111111111_1110101010001010_0011000101001110"; -- -0.08382884830013572
	pesos_i(17733) := b"1111111111111111_1111111111111111_1111000011011011_1000010011100110"; -- -0.05915040388854934
	pesos_i(17734) := b"0000000000000000_0000000000000000_0000001101101100_0010110100001101"; -- 0.013369384562946528
	pesos_i(17735) := b"1111111111111111_1111111111111111_1111011101000100_1110111001110111"; -- -0.03410443869772821
	pesos_i(17736) := b"0000000000000000_0000000000000000_0001000101110101_1001000000110010"; -- 0.06820012311013239
	pesos_i(17737) := b"1111111111111111_1111111111111111_1110011000111011_0011100110111000"; -- -0.1006587911267504
	pesos_i(17738) := b"1111111111111111_1111111111111111_1111111101111101_1001011110011101"; -- -0.00198986456285312
	pesos_i(17739) := b"1111111111111111_1111111111111111_1110111001100100_1010111010011010"; -- -0.06877621404761106
	pesos_i(17740) := b"1111111111111111_1111111111111111_1111001011001001_0100010000011100"; -- -0.051616423705451275
	pesos_i(17741) := b"0000000000000000_0000000000000000_0000000000111001_1101101011011011"; -- 0.0008827958693474713
	pesos_i(17742) := b"1111111111111111_1111111111111111_1110001010110000_1100111110000001"; -- -0.11448958493578017
	pesos_i(17743) := b"1111111111111111_1111111111111111_1111111110101101_0110010011000100"; -- -0.001260473502578721
	pesos_i(17744) := b"1111111111111111_1111111111111111_1101111001100011_1101111001110111"; -- -0.13128862005214692
	pesos_i(17745) := b"0000000000000000_0000000000000000_0000010111100010_1010000001001001"; -- 0.02298929012438626
	pesos_i(17746) := b"0000000000000000_0000000000000000_0001111001010101_0110100010010010"; -- 0.1184907298366855
	pesos_i(17747) := b"1111111111111111_1111111111111111_1110111100000101_0101110100110100"; -- -0.06632440071346632
	pesos_i(17748) := b"1111111111111111_1111111111111111_1111001110110110_0111111000001000"; -- -0.047996638294304714
	pesos_i(17749) := b"1111111111111111_1111111111111111_1101101101110111_0000011010100101"; -- -0.14271505811412485
	pesos_i(17750) := b"0000000000000000_0000000000000000_0010010010101011_1110001010110111"; -- 0.1432477662681724
	pesos_i(17751) := b"1111111111111111_1111111111111111_1110010011100111_1011010000010000"; -- -0.10583948720749525
	pesos_i(17752) := b"1111111111111111_1111111111111111_1110010111010000_1000011001010110"; -- -0.10228691474493298
	pesos_i(17753) := b"1111111111111111_1111111111111111_1110110101100100_0100011100010110"; -- -0.07268863395568256
	pesos_i(17754) := b"0000000000000000_0000000000000000_0001111111011100_1100100101111011"; -- 0.12446269277040602
	pesos_i(17755) := b"1111111111111111_1111111111111111_1110011001011110_0100000001000001"; -- -0.1001243439640324
	pesos_i(17756) := b"0000000000000000_0000000000000000_0000110101100011_0111010000000110"; -- 0.05229878572795139
	pesos_i(17757) := b"0000000000000000_0000000000000000_0010000010010111_1010011100101011"; -- 0.1273140411640838
	pesos_i(17758) := b"1111111111111111_1111111111111111_1110111110010000_1100011100111100"; -- -0.06419710907466261
	pesos_i(17759) := b"0000000000000000_0000000000000000_0001000011000000_1010000100100100"; -- 0.06543929217633175
	pesos_i(17760) := b"0000000000000000_0000000000000000_0000100000110010_0110010000001101"; -- 0.03201890294974878
	pesos_i(17761) := b"1111111111111111_1111111111111111_1101111100100010_1001100001110111"; -- -0.1283783635962627
	pesos_i(17762) := b"0000000000000000_0000000000000000_0010000001110110_1101001001111110"; -- 0.1268130833223729
	pesos_i(17763) := b"0000000000000000_0000000000000000_0001001011011110_1011100010011100"; -- 0.0737109546787384
	pesos_i(17764) := b"0000000000000000_0000000000000000_0000100011011100_0111000110101000"; -- 0.03461370810920473
	pesos_i(17765) := b"0000000000000000_0000000000000000_0010000010011101_0100101111101100"; -- 0.12740015519187017
	pesos_i(17766) := b"1111111111111111_1111111111111111_1101101100011111_0010011110101110"; -- -0.1440558623350399
	pesos_i(17767) := b"1111111111111111_1111111111111111_1110100110010001_0110101010000101"; -- -0.08762487649228551
	pesos_i(17768) := b"1111111111111111_1111111111111111_1110110110000111_0110011011010000"; -- -0.07215268527285881
	pesos_i(17769) := b"1111111111111111_1111111111111111_1111001101010010_1000110101100101"; -- -0.0495216015639109
	pesos_i(17770) := b"1111111111111111_1111111111111111_1101110010110101_1011001111011110"; -- -0.13785243827365143
	pesos_i(17771) := b"1111111111111111_1111111111111111_1111101100100010_0011011000000010"; -- -0.019009232163460437
	pesos_i(17772) := b"1111111111111111_1111111111111111_1110011000100000_0011010111010100"; -- -0.10107101041432241
	pesos_i(17773) := b"0000000000000000_0000000000000000_0001100000101101_1000101100001100"; -- 0.09444493337837166
	pesos_i(17774) := b"1111111111111111_1111111111111111_1111000010101011_0000101001111011"; -- -0.05989012235741333
	pesos_i(17775) := b"0000000000000000_0000000000000000_0000111011101101_1010001101011001"; -- 0.058313569378552296
	pesos_i(17776) := b"0000000000000000_0000000000000000_0001111010010111_1010111100110101"; -- 0.11950202028561267
	pesos_i(17777) := b"1111111111111111_1111111111111111_1110101000110001_0011111110010001"; -- -0.085186030588593
	pesos_i(17778) := b"1111111111111111_1111111111111111_1111000011000001_1000101001110011"; -- -0.05954680139050747
	pesos_i(17779) := b"0000000000000000_0000000000000000_0001010000100000_0101011011001111"; -- 0.07861845538529305
	pesos_i(17780) := b"0000000000000000_0000000000000000_0001000000001001_1010110100010001"; -- 0.0626476447209363
	pesos_i(17781) := b"0000000000000000_0000000000000000_0000110001101110_1001001001110110"; -- 0.04856219665044088
	pesos_i(17782) := b"0000000000000000_0000000000000000_0000000001000010_0100000100100000"; -- 0.0010109618609553555
	pesos_i(17783) := b"1111111111111111_1111111111111111_1111011111010010_0100000011011011"; -- -0.031948038601938414
	pesos_i(17784) := b"0000000000000000_0000000000000000_0001101011100011_1101111111011100"; -- 0.10503958818899962
	pesos_i(17785) := b"0000000000000000_0000000000000000_0000110001110100_0101011011011010"; -- 0.04865019638517712
	pesos_i(17786) := b"1111111111111111_1111111111111111_1111110000111110_0111000010110101"; -- -0.0146722371978778
	pesos_i(17787) := b"0000000000000000_0000000000000000_0000110100110110_0101111111010001"; -- 0.05161093567451221
	pesos_i(17788) := b"0000000000000000_0000000000000000_0010001111111010_0111100111100100"; -- 0.14054071247978692
	pesos_i(17789) := b"1111111111111111_1111111111111111_1111011110101110_1010101010001001"; -- -0.03249105611296681
	pesos_i(17790) := b"1111111111111111_1111111111111111_1111011010111000_0010011011111100"; -- -0.03625255910366419
	pesos_i(17791) := b"0000000000000000_0000000000000000_0010010100111101_0111011001100111"; -- 0.14546909347077067
	pesos_i(17792) := b"0000000000000000_0000000000000000_0001100100010110_1110100000011010"; -- 0.09800577773475917
	pesos_i(17793) := b"0000000000000000_0000000000000000_0001011111111011_0101111111010100"; -- 0.09367941775211236
	pesos_i(17794) := b"1111111111111111_1111111111111111_1111110110100000_0110000110110110"; -- -0.009271519632724958
	pesos_i(17795) := b"0000000000000000_0000000000000000_0000011001110000_1010111001101101"; -- 0.02515688091162754
	pesos_i(17796) := b"0000000000000000_0000000000000000_0001010110000111_1111101110000001"; -- 0.08410617722513046
	pesos_i(17797) := b"1111111111111111_1111111111111111_1110111011111100_1100111101001011"; -- -0.0664549294740061
	pesos_i(17798) := b"0000000000000000_0000000000000000_0001010101110101_0011010110110111"; -- 0.08381972993646566
	pesos_i(17799) := b"0000000000000000_0000000000000000_0001010110011101_0000101010001100"; -- 0.0844275085110334
	pesos_i(17800) := b"1111111111111111_1111111111111111_1110111011011110_1011000101001101"; -- -0.0669144809811018
	pesos_i(17801) := b"0000000000000000_0000000000000000_0001100010000101_1010101101111000"; -- 0.09578963925480506
	pesos_i(17802) := b"1111111111111111_1111111111111111_1110110001111111_0001001101101011"; -- -0.07618597636264011
	pesos_i(17803) := b"1111111111111111_1111111111111111_1111000011111010_1111010101111000"; -- -0.0586706715816926
	pesos_i(17804) := b"0000000000000000_0000000000000000_0000000101101000_1001011100000101"; -- 0.005502165451078948
	pesos_i(17805) := b"0000000000000000_0000000000000000_0010001101110010_0111111100010010"; -- 0.1384658258288551
	pesos_i(17806) := b"0000000000000000_0000000000000000_0001010000100100_0101110010011101"; -- 0.07867983650125183
	pesos_i(17807) := b"0000000000000000_0000000000000000_0000110100000101_0100110110000001"; -- 0.05086216347896994
	pesos_i(17808) := b"1111111111111111_1111111111111111_1111010011110010_1110010000010111"; -- -0.043168777941501875
	pesos_i(17809) := b"1111111111111111_1111111111111111_1111100011110011_0001011100000001"; -- -0.027540743202400048
	pesos_i(17810) := b"1111111111111111_1111111111111111_1101001100010000_0001101001110010"; -- -0.17553553321670962
	pesos_i(17811) := b"0000000000000000_0000000000000000_0000110010011001_0110001110100101"; -- 0.0492155340767062
	pesos_i(17812) := b"1111111111111111_1111111111111111_1110010100010010_1010010001010110"; -- -0.10518429651746478
	pesos_i(17813) := b"0000000000000000_0000000000000000_0010000100110011_0111011001110101"; -- 0.12969150878997546
	pesos_i(17814) := b"0000000000000000_0000000000000000_0000110011010001_1101101110001011"; -- 0.05007717273896927
	pesos_i(17815) := b"1111111111111111_1111111111111111_1110100010101010_1111100111101000"; -- -0.09114111036768492
	pesos_i(17816) := b"0000000000000000_0000000000000000_0000100001100001_0000001110011011"; -- 0.03273031743857704
	pesos_i(17817) := b"1111111111111111_1111111111111111_1101011000111001_1010000000111100"; -- -0.16318319824735572
	pesos_i(17818) := b"1111111111111111_1111111111111111_1111100010110010_0110011101101111"; -- -0.028527770529561382
	pesos_i(17819) := b"0000000000000000_0000000000000000_0000011101011000_0010001000100100"; -- 0.028688558384103596
	pesos_i(17820) := b"1111111111111111_1111111111111111_1110101110000101_0110001111000111"; -- -0.07999588376293389
	pesos_i(17821) := b"0000000000000000_0000000000000000_0001101111101010_0001001100010000"; -- 0.10904044293121037
	pesos_i(17822) := b"1111111111111111_1111111111111111_1111010110001111_0100000101000110"; -- -0.04078285250144662
	pesos_i(17823) := b"0000000000000000_0000000000000000_0001010110100101_1101110001000110"; -- 0.08456207947843657
	pesos_i(17824) := b"1111111111111111_1111111111111111_1111010111111011_0101101001010001"; -- -0.03913341063048095
	pesos_i(17825) := b"0000000000000000_0000000000000000_0001101101100100_0010101010110001"; -- 0.10699717354363658
	pesos_i(17826) := b"0000000000000000_0000000000000000_0010011100010110_1110010001011110"; -- 0.15269305508760475
	pesos_i(17827) := b"1111111111111111_1111111111111111_1110110011001001_1101011111100111"; -- -0.07504511451478939
	pesos_i(17828) := b"0000000000000000_0000000000000000_0001101110110011_0010011111111111"; -- 0.10820245717038776
	pesos_i(17829) := b"0000000000000000_0000000000000000_0000011100111010_1100001011001011"; -- 0.028240370405667185
	pesos_i(17830) := b"1111111111111111_1111111111111111_1111111100001010_1111010100100000"; -- -0.003739051448910919
	pesos_i(17831) := b"0000000000000000_0000000000000000_0001100000111100_0000110111000100"; -- 0.09466634791885536
	pesos_i(17832) := b"1111111111111111_1111111111111111_1111111000001011_1000001101101011"; -- -0.007636820178386601
	pesos_i(17833) := b"1111111111111111_1111111111111111_1101110101000100_0111111000100011"; -- -0.13567363394820517
	pesos_i(17834) := b"0000000000000000_0000000000000000_0001100111101001_0101100101011000"; -- 0.10121687319299641
	pesos_i(17835) := b"1111111111111111_1111111111111111_1110011100110010_1000111010111100"; -- -0.09688480289960134
	pesos_i(17836) := b"1111111111111111_1111111111111111_1110000110000011_1001110010110001"; -- -0.1190855090110828
	pesos_i(17837) := b"1111111111111111_1111111111111111_1111001100101111_1011001110110011"; -- -0.050053375983534376
	pesos_i(17838) := b"1111111111111111_1111111111111111_1111010000101100_0000000101101100"; -- -0.04620352852076347
	pesos_i(17839) := b"0000000000000000_0000000000000000_0000001010011110_0010110100100110"; -- 0.010226079840888703
	pesos_i(17840) := b"0000000000000000_0000000000000000_0000010110101101_1101110101100111"; -- 0.022184217156571148
	pesos_i(17841) := b"0000000000000000_0000000000000000_0010000010101010_0001001100001000"; -- 0.12759512851200885
	pesos_i(17842) := b"1111111111111111_1111111111111111_1110110111001100_0000010001111010"; -- -0.07110569020266645
	pesos_i(17843) := b"1111111111111111_1111111111111111_1110100101001010_1011111000110010"; -- -0.08870326304189304
	pesos_i(17844) := b"0000000000000000_0000000000000000_0001001000010100_1101010110010000"; -- 0.07063040509168371
	pesos_i(17845) := b"1111111111111111_1111111111111111_1111000000010110_0010111001111011"; -- -0.06216153610580436
	pesos_i(17846) := b"0000000000000000_0000000000000000_0000111100100011_1000000001000111"; -- 0.05913545352387352
	pesos_i(17847) := b"0000000000000000_0000000000000000_0001000001001111_1110110011011000"; -- 0.06371956122289293
	pesos_i(17848) := b"1111111111111111_1111111111111111_1110100110000001_0000011101101111"; -- -0.0878749231670231
	pesos_i(17849) := b"0000000000000000_0000000000000000_0001010101101010_1001001100000000"; -- 0.0836574435787957
	pesos_i(17850) := b"0000000000000000_0000000000000000_0001101111111010_1010110100110101"; -- 0.10929377126104112
	pesos_i(17851) := b"1111111111111111_1111111111111111_1110110100011010_0000001011000011"; -- -0.07382185686601282
	pesos_i(17852) := b"1111111111111111_1111111111111111_1111010100100111_1001100010011001"; -- -0.04236456174487193
	pesos_i(17853) := b"0000000000000000_0000000000000000_0000110111011001_1100100001000000"; -- 0.05410434299100479
	pesos_i(17854) := b"1111111111111111_1111111111111111_1110110000111000_1110011110011011"; -- -0.07725670303584241
	pesos_i(17855) := b"1111111111111111_1111111111111111_1110100101101110_0011000000100100"; -- -0.08816241372182103
	pesos_i(17856) := b"0000000000000000_0000000000000000_0000010101001101_1110010110001000"; -- 0.02071985789583285
	pesos_i(17857) := b"0000000000000000_0000000000000000_0010000001001001_1010011010000010"; -- 0.12612381625528665
	pesos_i(17858) := b"0000000000000000_0000000000000000_0000011001011110_0101110011011011"; -- 0.024877360765634612
	pesos_i(17859) := b"1111111111111111_1111111111111111_1101001110101000_1010101010101110"; -- -0.17320760017025377
	pesos_i(17860) := b"0000000000000000_0000000000000000_0000101100100100_0001111001100011"; -- 0.043519877549198824
	pesos_i(17861) := b"0000000000000000_0000000000000000_0000101101111110_0000001010000011"; -- 0.04489150720378489
	pesos_i(17862) := b"0000000000000000_0000000000000000_0001000110010100_1000000110111111"; -- 0.06867228430837112
	pesos_i(17863) := b"1111111111111111_1111111111111111_1111011101010110_1010001100000011"; -- -0.03383427785035997
	pesos_i(17864) := b"0000000000000000_0000000000000000_0000111000010000_0010000110100001"; -- 0.054933645024850014
	pesos_i(17865) := b"1111111111111111_1111111111111111_1110101001000111_0110111010110011"; -- -0.08484752789355007
	pesos_i(17866) := b"0000000000000000_0000000000000000_0001001011010010_1101010110001110"; -- 0.07352957459398045
	pesos_i(17867) := b"1111111111111111_1111111111111111_1110111111100000_1100101101101001"; -- -0.0629761570928805
	pesos_i(17868) := b"0000000000000000_0000000000000000_0000100100110110_1100000110111001"; -- 0.03599177127213216
	pesos_i(17869) := b"0000000000000000_0000000000000000_0000100011010010_0000010001110110"; -- 0.034454611606941486
	pesos_i(17870) := b"0000000000000000_0000000000000000_0010001010010000_0101111001010011"; -- 0.13501538774646007
	pesos_i(17871) := b"1111111111111111_1111111111111111_1101011111011001_1111111101011110"; -- -0.15682987168957202
	pesos_i(17872) := b"1111111111111111_1111111111111111_1101111011110011_0101010100011000"; -- -0.1290995422279461
	pesos_i(17873) := b"0000000000000000_0000000000000000_0010010110101010_1100000010111001"; -- 0.1471367312422753
	pesos_i(17874) := b"1111111111111111_1111111111111111_1110110100100111_1101011100001100"; -- -0.07361083951658251
	pesos_i(17875) := b"0000000000000000_0000000000000000_0000000101101101_0000100101011001"; -- 0.0055700152093174134
	pesos_i(17876) := b"0000000000000000_0000000000000000_0001100110110101_0110011000100101"; -- 0.1004241792104625
	pesos_i(17877) := b"0000000000000000_0000000000000000_0000101011000001_1000100001010100"; -- 0.04201557215900325
	pesos_i(17878) := b"1111111111111111_1111111111111111_1111100100010011_0001001111011110"; -- -0.027052648902309996
	pesos_i(17879) := b"1111111111111111_1111111111111111_1101110011101111_1101111100110001"; -- -0.13696484609590345
	pesos_i(17880) := b"1111111111111111_1111111111111111_1101111011000111_0100011111011101"; -- -0.1297717175925239
	pesos_i(17881) := b"1111111111111111_1111111111111111_1111100011101001_0000000111100001"; -- -0.02769459015031236
	pesos_i(17882) := b"0000000000000000_0000000000000000_0001000100000011_0110111000001100"; -- 0.06645858555693206
	pesos_i(17883) := b"1111111111111111_1111111111111111_1111101001001101_0011101100010001"; -- -0.022259052590565525
	pesos_i(17884) := b"1111111111111111_1111111111111111_1110110101100011_0110011010001111"; -- -0.07270201699597299
	pesos_i(17885) := b"0000000000000000_0000000000000000_0001010001110011_0011100111011010"; -- 0.07988320899729942
	pesos_i(17886) := b"1111111111111111_1111111111111111_1110101011110100_1000100111110100"; -- -0.08220613276977014
	pesos_i(17887) := b"1111111111111111_1111111111111111_1110001101110010_1011101110101100"; -- -0.11153056187017707
	pesos_i(17888) := b"1111111111111111_1111111111111111_1110011100000110_0110110000000110"; -- -0.09755825851201798
	pesos_i(17889) := b"0000000000000000_0000000000000000_0001000110011010_1001101111001110"; -- 0.06876539009627956
	pesos_i(17890) := b"0000000000000000_0000000000000000_0001110010101001_0000110010010101"; -- 0.11195448532901511
	pesos_i(17891) := b"1111111111111111_1111111111111111_1111111101001001_0100010001000010"; -- -0.0027882898121181646
	pesos_i(17892) := b"0000000000000000_0000000000000000_0000110001011111_1111001001110110"; -- 0.04833903676012321
	pesos_i(17893) := b"1111111111111111_1111111111111111_1101110110110101_0101001010111000"; -- -0.13395197864696676
	pesos_i(17894) := b"0000000000000000_0000000000000000_0001001001101110_0001011011001000"; -- 0.07199232471100832
	pesos_i(17895) := b"0000000000000000_0000000000000000_0000111110001000_1001101000001010"; -- 0.060678126666806026
	pesos_i(17896) := b"0000000000000000_0000000000000000_0000001011011011_0100001111010010"; -- 0.01115821721035748
	pesos_i(17897) := b"1111111111111111_1111111111111111_1111110001101110_0001111000111000"; -- -0.013944731940116866
	pesos_i(17898) := b"1111111111111111_1111111111111111_1101111111111110_0101111011111000"; -- -0.1250248570593047
	pesos_i(17899) := b"1111111111111111_1111111111111111_1110010001001110_1001100111011001"; -- -0.10817564446430682
	pesos_i(17900) := b"0000000000000000_0000000000000000_0000011001111111_0111101001101010"; -- 0.025382662637946547
	pesos_i(17901) := b"0000000000000000_0000000000000000_0000101100110001_1001000110011010"; -- 0.043725109131419554
	pesos_i(17902) := b"1111111111111111_1111111111111111_1110101100111110_1011011101110011"; -- -0.08107427074837162
	pesos_i(17903) := b"1111111111111111_1111111111111111_1111011001011110_1101011100001000"; -- -0.037615356895731415
	pesos_i(17904) := b"1111111111111111_1111111111111111_1111000001001011_0111000000010010"; -- -0.06134891101154041
	pesos_i(17905) := b"0000000000000000_0000000000000000_0000010010001001_1111110001111000"; -- 0.017730502478226794
	pesos_i(17906) := b"0000000000000000_0000000000000000_0000001001011100_1010001010001101"; -- 0.009225997317372638
	pesos_i(17907) := b"0000000000000000_0000000000000000_0001011111100010_0101100001100110"; -- 0.09329750533162319
	pesos_i(17908) := b"1111111111111111_1111111111111111_1111010110110011_0100100101101000"; -- -0.040233051375608196
	pesos_i(17909) := b"1111111111111111_1111111111111111_1111001001111011_1111011011101010"; -- -0.05279595162374739
	pesos_i(17910) := b"1111111111111111_1111111111111111_1101100110010101_0010101111111110"; -- -0.15006756822020578
	pesos_i(17911) := b"0000000000000000_0000000000000000_0000111110101000_0100010011000010"; -- 0.06116132482896289
	pesos_i(17912) := b"0000000000000000_0000000000000000_0010011101011101_1010001101100110"; -- 0.15377255669543619
	pesos_i(17913) := b"0000000000000000_0000000000000000_0001010011000101_0100010101110101"; -- 0.08113512141605848
	pesos_i(17914) := b"0000000000000000_0000000000000000_0001110001101001_1111101001111010"; -- 0.11099210246577909
	pesos_i(17915) := b"1111111111111111_1111111111111111_1110011000000100_1000110100001000"; -- -0.10149305879948303
	pesos_i(17916) := b"1111111111111111_1111111111111111_1111010101111111_1110100010001111"; -- -0.0410170221173649
	pesos_i(17917) := b"1111111111111111_1111111111111111_1111010011100100_0010100101000100"; -- -0.043393536500625045
	pesos_i(17918) := b"0000000000000000_0000000000000000_0000011101011111_0011101001101001"; -- 0.028796816416252626
	pesos_i(17919) := b"1111111111111111_1111111111111111_1111100110010100_1001110010000111"; -- -0.025076119558415846
	pesos_i(17920) := b"0000000000000000_0000000000000000_0000111011010011_0100001011001110"; -- 0.05791108637697937
	pesos_i(17921) := b"0000000000000000_0000000000000000_0001010111010100_0001011101011011"; -- 0.08526750544267946
	pesos_i(17922) := b"0000000000000000_0000000000000000_0001110000001100_1110111011010011"; -- 0.10957234039219507
	pesos_i(17923) := b"0000000000000000_0000000000000000_0000101100100110_1000011100001010"; -- 0.04355663302881899
	pesos_i(17924) := b"0000000000000000_0000000000000000_0001000010111101_0100100110000111"; -- 0.06538829358812312
	pesos_i(17925) := b"0000000000000000_0000000000000000_0000001000000110_1001111001100110"; -- 0.007913493917534131
	pesos_i(17926) := b"1111111111111111_1111111111111111_1111010010010100_1001011101101101"; -- -0.04460767346186998
	pesos_i(17927) := b"1111111111111111_1111111111111111_1110001000100001_0101000101101001"; -- -0.11667910747907916
	pesos_i(17928) := b"1111111111111111_1111111111111111_1111000100110010_0011100001001000"; -- -0.05782745601831259
	pesos_i(17929) := b"0000000000000000_0000000000000000_0001001101010010_0001100100010101"; -- 0.07547146563349678
	pesos_i(17930) := b"0000000000000000_0000000000000000_0010000100100001_0000110001000001"; -- 0.12941052034030456
	pesos_i(17931) := b"0000000000000000_0000000000000000_0010000110110101_0001000011010111"; -- 0.13166909466432314
	pesos_i(17932) := b"1111111111111111_1111111111111111_1101111011001001_1101001001111111"; -- -0.12973293684056644
	pesos_i(17933) := b"1111111111111111_1111111111111111_1101110100001101_1011101010110010"; -- -0.13650925792848126
	pesos_i(17934) := b"1111111111111111_1111111111111111_1110000101101011_0101011111010001"; -- -0.11945582535738511
	pesos_i(17935) := b"0000000000000000_0000000000000000_0001011111011110_1010101010101001"; -- 0.09324137330464513
	pesos_i(17936) := b"0000000000000000_0000000000000000_0000011000100101_0010001101111000"; -- 0.024004189391874084
	pesos_i(17937) := b"0000000000000000_0000000000000000_0000010010011111_0101001110101101"; -- 0.01805613491656124
	pesos_i(17938) := b"0000000000000000_0000000000000000_0001101011011100_0011111111110100"; -- 0.10492324546479073
	pesos_i(17939) := b"1111111111111111_1111111111111111_1111100011110001_1110010010111001"; -- -0.02755899879238923
	pesos_i(17940) := b"0000000000000000_0000000000000000_0000001111010100_0100011010101111"; -- 0.014957826341179151
	pesos_i(17941) := b"0000000000000000_0000000000000000_0001010001100010_0000010110010110"; -- 0.07962069423908376
	pesos_i(17942) := b"1111111111111111_1111111111111111_1101100010100010_0101001100110110"; -- -0.15377311652570255
	pesos_i(17943) := b"0000000000000000_0000000000000000_0001100101110001_1000111100100111"; -- 0.09938902563639931
	pesos_i(17944) := b"1111111111111111_1111111111111111_1110111111111010_1101001001110000"; -- -0.06257900972828638
	pesos_i(17945) := b"1111111111111111_1111111111111111_1110011110100110_0001000011110011"; -- -0.09512228065271888
	pesos_i(17946) := b"1111111111111111_1111111111111111_1111110100011100_0000011101110000"; -- -0.011291060582950707
	pesos_i(17947) := b"0000000000000000_0000000000000000_0001111011001010_0001000011110001"; -- 0.12027078518513569
	pesos_i(17948) := b"1111111111111111_1111111111111111_1111001010000100_0010101011110100"; -- -0.05267077965056205
	pesos_i(17949) := b"0000000000000000_0000000000000000_0000010010111001_1101000001100101"; -- 0.018460297243741493
	pesos_i(17950) := b"0000000000000000_0000000000000000_0000010100010100_0101001010000001"; -- 0.019841343426847385
	pesos_i(17951) := b"1111111111111111_1111111111111111_1110001010101101_1100100100000110"; -- -0.11453574751406427
	pesos_i(17952) := b"1111111111111111_1111111111111111_1110111001001010_0111110110101110"; -- -0.0691758585172111
	pesos_i(17953) := b"0000000000000000_0000000000000000_0001100011000011_1001111010101011"; -- 0.09673492120380793
	pesos_i(17954) := b"0000000000000000_0000000000000000_0010011100010101_0010011111001101"; -- 0.15266655693910716
	pesos_i(17955) := b"1111111111111111_1111111111111111_1111011010010001_1110100100010011"; -- -0.03683608323542212
	pesos_i(17956) := b"1111111111111111_1111111111111111_1111001011000001_1010011110010110"; -- -0.05173256484879553
	pesos_i(17957) := b"1111111111111111_1111111111111111_1111100010010001_1011110010101110"; -- -0.029026229473934267
	pesos_i(17958) := b"0000000000000000_0000000000000000_0001010110000101_1001010111000011"; -- 0.08406959554006929
	pesos_i(17959) := b"1111111111111111_1111111111111111_1110100011000011_0111011001111000"; -- -0.09076747473824161
	pesos_i(17960) := b"0000000000000000_0000000000000000_0000110101101100_1010001101000100"; -- 0.052438930681071055
	pesos_i(17961) := b"1111111111111111_1111111111111111_1111011000111011_0111011111000011"; -- -0.03815509319955906
	pesos_i(17962) := b"1111111111111111_1111111111111111_1110011001101111_1100110010100111"; -- -0.09985657607505401
	pesos_i(17963) := b"0000000000000000_0000000000000000_0000000101111101_0110101000110100"; -- 0.005819928887083378
	pesos_i(17964) := b"0000000000000000_0000000000000000_0000110110100011_0011001001111111"; -- 0.05327144250154809
	pesos_i(17965) := b"1111111111111111_1111111111111111_1101101010001010_1001101111001010"; -- -0.1463225014503803
	pesos_i(17966) := b"0000000000000000_0000000000000000_0001000111011111_1010010110010000"; -- 0.0698188281971972
	pesos_i(17967) := b"0000000000000000_0000000000000000_0001110011101010_0110011100100110"; -- 0.11295170466447133
	pesos_i(17968) := b"1111111111111111_1111111111111111_1110100111100010_0110001111000111"; -- -0.08638931646310027
	pesos_i(17969) := b"0000000000000000_0000000000000000_0001111000110011_0111100110011100"; -- 0.11797294674672312
	pesos_i(17970) := b"0000000000000000_0000000000000000_0001000100001100_0010010101110110"; -- 0.06659158837769068
	pesos_i(17971) := b"1111111111111111_1111111111111111_1110111000010011_1101100110110000"; -- -0.07000960771494144
	pesos_i(17972) := b"1111111111111111_1111111111111111_1110100010011000_0111100010011100"; -- -0.09142347519250901
	pesos_i(17973) := b"0000000000000000_0000000000000000_0001101000000110_1010011100000011"; -- 0.10166400733628282
	pesos_i(17974) := b"0000000000000000_0000000000000000_0000110101110011_0111000110101000"; -- 0.05254278528452329
	pesos_i(17975) := b"0000000000000000_0000000000000000_0001111101101101_0000110001000111"; -- 0.12275768968816093
	pesos_i(17976) := b"0000000000000000_0000000000000000_0000001010111110_1111011001111101"; -- 0.010726361868181815
	pesos_i(17977) := b"1111111111111111_1111111111111111_1110100100010001_0000110010000101"; -- -0.08958360445854088
	pesos_i(17978) := b"1111111111111111_1111111111111111_1110010010000111_0111110101101001"; -- -0.10730758850138114
	pesos_i(17979) := b"0000000000000000_0000000000000000_0000001011001001_0100000101101111"; -- 0.010883416783440906
	pesos_i(17980) := b"0000000000000000_0000000000000000_0010100001001000_0110000100111011"; -- 0.15735442829270432
	pesos_i(17981) := b"1111111111111111_1111111111111111_1111010011101100_1001100100100011"; -- -0.043264798234724434
	pesos_i(17982) := b"0000000000000000_0000000000000000_0001000000100000_0011011000111101"; -- 0.06299151417949067
	pesos_i(17983) := b"0000000000000000_0000000000000000_0010010101001100_0110010000100000"; -- 0.1456968859208085
	pesos_i(17984) := b"0000000000000000_0000000000000000_0000110001001010_1001110001001101"; -- 0.0480134666810131
	pesos_i(17985) := b"1111111111111111_1111111111111111_1110100110010110_1110000111010110"; -- -0.08754147085397104
	pesos_i(17986) := b"0000000000000000_0000000000000000_0010011111010011_1010110011001110"; -- 0.15557365437156737
	pesos_i(17987) := b"1111111111111111_1111111111111111_1111111101100001_0001010000110110"; -- -0.0024249428969642353
	pesos_i(17988) := b"1111111111111111_1111111111111111_1111000010011100_1101001110110011"; -- -0.06010701061513625
	pesos_i(17989) := b"0000000000000000_0000000000000000_0001000010111010_1101010001010001"; -- 0.06535078987347134
	pesos_i(17990) := b"0000000000000000_0000000000000000_0001111110001010_1011110100010101"; -- 0.12321073297858022
	pesos_i(17991) := b"0000000000000000_0000000000000000_0001011111111111_1010011011010001"; -- 0.09374468423850513
	pesos_i(17992) := b"1111111111111111_1111111111111111_1111011111110001_0101100011101000"; -- -0.031473582713006015
	pesos_i(17993) := b"0000000000000000_0000000000000000_0000000100011010_0001110000110000"; -- 0.004304658732004818
	pesos_i(17994) := b"1111111111111111_1111111111111111_1101111110110101_0010101000010100"; -- -0.12614190108877343
	pesos_i(17995) := b"1111111111111111_1111111111111111_1110011010011011_1001101000011110"; -- -0.09918820166065513
	pesos_i(17996) := b"1111111111111111_1111111111111111_1110101100011011_0110110111111001"; -- -0.0816127078410478
	pesos_i(17997) := b"0000000000000000_0000000000000000_0001100001100111_0100100010011111"; -- 0.09532598379485943
	pesos_i(17998) := b"0000000000000000_0000000000000000_0000100101010011_0011110101101110"; -- 0.03642639099349819
	pesos_i(17999) := b"0000000000000000_0000000000000000_0001101100101000_1000011000010100"; -- 0.10608709324654522
	pesos_i(18000) := b"0000000000000000_0000000000000000_0001100011010111_1100111100110101"; -- 0.09704299022301718
	pesos_i(18001) := b"1111111111111111_1111111111111111_1111001010101111_1101100100010100"; -- -0.05200427308057483
	pesos_i(18002) := b"1111111111111111_1111111111111111_1111111101110000_1000111101000100"; -- -0.0021887263249850946
	pesos_i(18003) := b"0000000000000000_0000000000000000_0000111011011100_0010011010110110"; -- 0.05804674106165244
	pesos_i(18004) := b"1111111111111111_1111111111111111_1111011011111101_1011001011011111"; -- -0.035191364820860674
	pesos_i(18005) := b"0000000000000000_0000000000000000_0000110000111101_1101101010001010"; -- 0.04781881218505023
	pesos_i(18006) := b"0000000000000000_0000000000000000_0010001110001001_0110101010000001"; -- 0.1388155522901151
	pesos_i(18007) := b"1111111111111111_1111111111111111_1111100001111000_1101011111100110"; -- -0.029406076704251046
	pesos_i(18008) := b"1111111111111111_1111111111111111_1111111101101101_0111000111010011"; -- -0.0022362574370543165
	pesos_i(18009) := b"0000000000000000_0000000000000000_0000011000011000_1100001010101010"; -- 0.02381531388941663
	pesos_i(18010) := b"0000000000000000_0000000000000000_0010101001111111_0001101110101110"; -- 0.16600201608828025
	pesos_i(18011) := b"1111111111111111_1111111111111111_1101011001101000_1101111100000110"; -- -0.16246229270036378
	pesos_i(18012) := b"0000000000000000_0000000000000000_0000100001011011_0110101001011100"; -- 0.03264488937550258
	pesos_i(18013) := b"1111111111111111_1111111111111111_1110001100111100_0010100100000101"; -- -0.11236327758632618
	pesos_i(18014) := b"1111111111111111_1111111111111111_1111111000111111_1001111100101101"; -- -0.006841708642823159
	pesos_i(18015) := b"1111111111111111_1111111111111111_1111100101010111_0011111101011010"; -- -0.02601245934208227
	pesos_i(18016) := b"1111111111111111_1111111111111111_1111011010100110_1001111011011111"; -- -0.0365200716395704
	pesos_i(18017) := b"1111111111111111_1111111111111111_1101101111110100_1111010110010111"; -- -0.14079346725794956
	pesos_i(18018) := b"0000000000000000_0000000000000000_0001001100111110_0000110001101001"; -- 0.07516553455959019
	pesos_i(18019) := b"0000000000000000_0000000000000000_0001101110011011_1001001110010101"; -- 0.1078426589331389
	pesos_i(18020) := b"1111111111111111_1111111111111111_1101101010010101_0110001011110010"; -- -0.1461580429415646
	pesos_i(18021) := b"0000000000000000_0000000000000000_0001101010001011_0111111110100111"; -- 0.10369108027329962
	pesos_i(18022) := b"1111111111111111_1111111111111111_1110001100110010_0001010010010101"; -- -0.11251708370209684
	pesos_i(18023) := b"1111111111111111_1111111111111111_1101111000010110_0001100100011000"; -- -0.13247531102885127
	pesos_i(18024) := b"0000000000000000_0000000000000000_0001110110101100_1011100101011010"; -- 0.11591680955119343
	pesos_i(18025) := b"0000000000000000_0000000000000000_0001111000110110_0101110000110110"; -- 0.1180169708264445
	pesos_i(18026) := b"0000000000000000_0000000000000000_0001001110000010_1001101000000000"; -- 0.07621157169022084
	pesos_i(18027) := b"1111111111111111_1111111111111111_1111011110011101_0011000110010011"; -- -0.03275766520162678
	pesos_i(18028) := b"1111111111111111_1111111111111111_1110000010001110_0101100101010011"; -- -0.12282792771557961
	pesos_i(18029) := b"1111111111111111_1111111111111111_1111000111110001_1101000000001110"; -- -0.05490398085277344
	pesos_i(18030) := b"0000000000000000_0000000000000000_0001101001001010_1001110000110101"; -- 0.10270096093978678
	pesos_i(18031) := b"1111111111111111_1111111111111111_1110110000111000_0011001111001110"; -- -0.07726742000017156
	pesos_i(18032) := b"1111111111111111_1111111111111111_1111101100011010_1010000110101010"; -- -0.01912488545237156
	pesos_i(18033) := b"1111111111111111_1111111111111111_1101101011011000_1011010011110101"; -- -0.14513081556855825
	pesos_i(18034) := b"1111111111111111_1111111111111111_1111000100000111_0100101111101100"; -- -0.05848241316531641
	pesos_i(18035) := b"0000000000000000_0000000000000000_0001111001010001_1111100011011011"; -- 0.11843829479212263
	pesos_i(18036) := b"0000000000000000_0000000000000000_0010001011100111_0110101100111010"; -- 0.13634367141457007
	pesos_i(18037) := b"1111111111111111_1111111111111111_1110000001110100_0100111110000000"; -- -0.12322524179779921
	pesos_i(18038) := b"0000000000000000_0000000000000000_0001011101101100_1011111111011111"; -- 0.09150313571756892
	pesos_i(18039) := b"0000000000000000_0000000000000000_0010011000010000_0011001111001000"; -- 0.14868472693404142
	pesos_i(18040) := b"1111111111111111_1111111111111111_1111101101101100_0000000001010010"; -- -0.017883281692050317
	pesos_i(18041) := b"1111111111111111_1111111111111111_1111101110111000_0100000100100111"; -- -0.016719749315657405
	pesos_i(18042) := b"0000000000000000_0000000000000000_0001100000010001_1010000100111111"; -- 0.09401901040106496
	pesos_i(18043) := b"1111111111111111_1111111111111111_1101110110011001_0011010101100001"; -- -0.13438097366690663
	pesos_i(18044) := b"0000000000000000_0000000000000000_0000110011110011_0111000110010000"; -- 0.05058965470479969
	pesos_i(18045) := b"0000000000000000_0000000000000000_0000001100010101_1011101011101111"; -- 0.012050326582412806
	pesos_i(18046) := b"1111111111111111_1111111111111111_1111110100010100_0111101000000010"; -- -0.011406302083144169
	pesos_i(18047) := b"1111111111111111_1111111111111111_1101101011000101_1110100111011000"; -- -0.14541758042298342
	pesos_i(18048) := b"0000000000000000_0000000000000000_0000100011011101_1100101000111111"; -- 0.03463424721260635
	pesos_i(18049) := b"1111111111111111_1111111111111111_1110010010101101_0000101010100000"; -- -0.10673459614800422
	pesos_i(18050) := b"1111111111111111_1111111111111111_1101110001011011_0011011010101100"; -- -0.13923319142182675
	pesos_i(18051) := b"1111111111111111_1111111111111111_1111110001011001_1011111011111110"; -- -0.01425558370708698
	pesos_i(18052) := b"0000000000000000_0000000000000000_0001010010100010_0010100011000100"; -- 0.08059935363849778
	pesos_i(18053) := b"0000000000000000_0000000000000000_0001100011000110_1111110100010001"; -- 0.09678632405651559
	pesos_i(18054) := b"0000000000000000_0000000000000000_0001101001000001_0110111001101101"; -- 0.10256090314379451
	pesos_i(18055) := b"1111111111111111_1111111111111111_1111101000100010_0010101100101100"; -- -0.022916127817168563
	pesos_i(18056) := b"1111111111111111_1111111111111111_1110011110011111_0111111011111111"; -- -0.09522253291125403
	pesos_i(18057) := b"1111111111111111_1111111111111111_1111010100101011_0100011010101001"; -- -0.04230841050577719
	pesos_i(18058) := b"0000000000000000_0000000000000000_0000111111100001_1110111100011000"; -- 0.06204122859960524
	pesos_i(18059) := b"0000000000000000_0000000000000000_0010001111011100_0001101000011000"; -- 0.14007723894910637
	pesos_i(18060) := b"1111111111111111_1111111111111111_1111100100000111_1011101001011110"; -- -0.027225830193038147
	pesos_i(18061) := b"1111111111111111_1111111111111111_1110010000110101_1011001010010100"; -- -0.10855564012097849
	pesos_i(18062) := b"0000000000000000_0000000000000000_0010000001001010_1000100000101001"; -- 0.12613726619905202
	pesos_i(18063) := b"0000000000000000_0000000000000000_0010010000100110_1111011011000010"; -- 0.1412195418610019
	pesos_i(18064) := b"1111111111111111_1111111111111111_1101110001100111_0101100000101101"; -- -0.1390480890836499
	pesos_i(18065) := b"1111111111111111_1111111111111111_1110010111111101_0011111000010100"; -- -0.10160457633886594
	pesos_i(18066) := b"1111111111111111_1111111111111111_1111101110101111_0110111111111010"; -- -0.01685428750572973
	pesos_i(18067) := b"1111111111111111_1111111111111111_1110100011100101_1011010110100101"; -- -0.09024491045836097
	pesos_i(18068) := b"1111111111111111_1111111111111111_1110110111010000_0100010001111011"; -- -0.0710408401902363
	pesos_i(18069) := b"1111111111111111_1111111111111111_1110001101001111_1001001101101000"; -- -0.11206701966890587
	pesos_i(18070) := b"1111111111111111_1111111111111111_1111001111011000_1101011000001101"; -- -0.047472593049895574
	pesos_i(18071) := b"1111111111111111_1111111111111111_1101110100100101_1001010110001111"; -- -0.13614526033295105
	pesos_i(18072) := b"1111111111111111_1111111111111111_1110111000001101_1101011010110111"; -- -0.07010133784682228
	pesos_i(18073) := b"0000000000000000_0000000000000000_0001111110101011_1011111101010111"; -- 0.1237144076062496
	pesos_i(18074) := b"0000000000000000_0000000000000000_0010001111110000_1010110110101000"; -- 0.1403912100290616
	pesos_i(18075) := b"1111111111111111_1111111111111111_1110100111100001_0001110110110100"; -- -0.08640875212687239
	pesos_i(18076) := b"0000000000000000_0000000000000000_0001100001100101_0100100001000001"; -- 0.09529544444060083
	pesos_i(18077) := b"0000000000000000_0000000000000000_0001001000000100_1001000000111100"; -- 0.07038213211622209
	pesos_i(18078) := b"1111111111111111_1111111111111111_1111100010011110_1101111111010001"; -- -0.0288257708705716
	pesos_i(18079) := b"1111111111111111_1111111111111111_1110110010101010_1100110101010000"; -- -0.07551876819187152
	pesos_i(18080) := b"0000000000000000_0000000000000000_0010010010111001_0000000100100111"; -- 0.14344794465388158
	pesos_i(18081) := b"0000000000000000_0000000000000000_0010001001000100_0111011000100000"; -- 0.13385713846851666
	pesos_i(18082) := b"1111111111111111_1111111111111111_1101101011000110_0110011000001101"; -- -0.14541017718064736
	pesos_i(18083) := b"0000000000000000_0000000000000000_0000000101111010_1000101000011110"; -- 0.005776054763474346
	pesos_i(18084) := b"1111111111111111_1111111111111111_1110000001011001_1011100010111000"; -- -0.12363095764068646
	pesos_i(18085) := b"1111111111111111_1111111111111111_1110110110110100_1111101000101110"; -- -0.07145725616615801
	pesos_i(18086) := b"0000000000000000_0000000000000000_0001111111100101_0010110010001100"; -- 0.12459066784347295
	pesos_i(18087) := b"0000000000000000_0000000000000000_0001000110100011_0000101101010011"; -- 0.06889410758464086
	pesos_i(18088) := b"1111111111111111_1111111111111111_1110001001110001_1110010011010100"; -- -0.11544961762722412
	pesos_i(18089) := b"1111111111111111_1111111111111111_1111010101000001_0000000011010100"; -- -0.04197687935574046
	pesos_i(18090) := b"1111111111111111_1111111111111111_1110011000101011_1111000110101101"; -- -0.10089196696535387
	pesos_i(18091) := b"0000000000000000_0000000000000000_0010100101010000_1101011100111000"; -- 0.16138978105483692
	pesos_i(18092) := b"1111111111111111_1111111111111111_1111100111010100_1101100110100011"; -- -0.024095914495860352
	pesos_i(18093) := b"0000000000000000_0000000000000000_0001001111100110_0010011010010111"; -- 0.07773057168156265
	pesos_i(18094) := b"1111111111111111_1111111111111111_1111000101011110_1111001101000100"; -- -0.057144924113033804
	pesos_i(18095) := b"0000000000000000_0000000000000000_0000101110001000_0000011101000001"; -- 0.04504437757898207
	pesos_i(18096) := b"1111111111111111_1111111111111111_1111001111100110_1101010001110011"; -- -0.04725906566910501
	pesos_i(18097) := b"1111111111111111_1111111111111111_1111110101101111_1001100000000010"; -- -0.010015963926423253
	pesos_i(18098) := b"1111111111111111_1111111111111111_1111101010001010_0101000010111010"; -- -0.02132697547312295
	pesos_i(18099) := b"1111111111111111_1111111111111111_1110101001011000_0011111111011011"; -- -0.08459092040306022
	pesos_i(18100) := b"1111111111111111_1111111111111111_1101101001101010_1001001110100111"; -- -0.14681126758173882
	pesos_i(18101) := b"1111111111111111_1111111111111111_1111010110111110_1110000111100000"; -- -0.040056116976783095
	pesos_i(18102) := b"0000000000000000_0000000000000000_0001101111111110_1100110111001110"; -- 0.10935674931371164
	pesos_i(18103) := b"0000000000000000_0000000000000000_0001010100011111_0000111000111110"; -- 0.08250512124834741
	pesos_i(18104) := b"0000000000000000_0000000000000000_0001010011110000_0111110011110010"; -- 0.0817945567596036
	pesos_i(18105) := b"1111111111111111_1111111111111111_1111111001111011_0010011011111000"; -- -0.005933346227112792
	pesos_i(18106) := b"0000000000000000_0000000000000000_0010001001000110_1011111100010000"; -- 0.1338920034536765
	pesos_i(18107) := b"0000000000000000_0000000000000000_0000110110010101_1101100000001111"; -- 0.05306768774194115
	pesos_i(18108) := b"0000000000000000_0000000000000000_0000111001000111_1101110110110011"; -- 0.055784088430074735
	pesos_i(18109) := b"1111111111111111_1111111111111111_1111110100101000_0010111000000011"; -- -0.011105656009165833
	pesos_i(18110) := b"0000000000000000_0000000000000000_0000111111010010_0111111000000000"; -- 0.06180560581607011
	pesos_i(18111) := b"1111111111111111_1111111111111111_1101101110000000_0011000001101111"; -- -0.14257523822212503
	pesos_i(18112) := b"0000000000000000_0000000000000000_0000100100100111_0010101001101110"; -- 0.0357538718487
	pesos_i(18113) := b"0000000000000000_0000000000000000_0001110110110101_0011100010011111"; -- 0.11604646575469711
	pesos_i(18114) := b"0000000000000000_0000000000000000_0001000101100010_1010110000100100"; -- 0.06791187179982781
	pesos_i(18115) := b"0000000000000000_0000000000000000_0000111110011110_0101111010101010"; -- 0.06101028112922147
	pesos_i(18116) := b"1111111111111111_1111111111111111_1111001011100001_0001100101011111"; -- -0.05125276023982107
	pesos_i(18117) := b"0000000000000000_0000000000000000_0001111110011111_0010100010111011"; -- 0.12352232521693055
	pesos_i(18118) := b"0000000000000000_0000000000000000_0000000011010000_1101110001000101"; -- 0.0031869571060895116
	pesos_i(18119) := b"1111111111111111_1111111111111111_1110101111001111_1001111000110111"; -- -0.07886325030251319
	pesos_i(18120) := b"0000000000000000_0000000000000000_0001001111111111_1111010111001001"; -- 0.078124391150684
	pesos_i(18121) := b"0000000000000000_0000000000000000_0000101100001010_1100101111101100"; -- 0.043133492578806
	pesos_i(18122) := b"1111111111111111_1111111111111111_1110100011111001_1001001000101100"; -- -0.08994184894674752
	pesos_i(18123) := b"1111111111111111_1111111111111111_1101110100111000_1011000000101010"; -- -0.13585375768476776
	pesos_i(18124) := b"0000000000000000_0000000000000000_0000001010001001_1100010110000110"; -- 0.009914727528766007
	pesos_i(18125) := b"0000000000000000_0000000000000000_0001001110011000_0011101011110100"; -- 0.07654159972402153
	pesos_i(18126) := b"1111111111111111_1111111111111111_1111011110110001_0111101000101100"; -- -0.032448162418237975
	pesos_i(18127) := b"0000000000000000_0000000000000000_0010010001001010_1111010100110010"; -- 0.14176876510893396
	pesos_i(18128) := b"0000000000000000_0000000000000000_0000110010011010_1010100011100000"; -- 0.04923491918428444
	pesos_i(18129) := b"1111111111111111_1111111111111111_1111101010110010_0110111001010110"; -- -0.020714859003224558
	pesos_i(18130) := b"0000000000000000_0000000000000000_0010001011100110_0001000001111000"; -- 0.1363230031760628
	pesos_i(18131) := b"0000000000000000_0000000000000000_0010001100000011_1110110010110110"; -- 0.13677863545931462
	pesos_i(18132) := b"0000000000000000_0000000000000000_0000011000011111_0111000101000000"; -- 0.023917272700382596
	pesos_i(18133) := b"1111111111111111_1111111111111111_1101110111010011_0100101110000101"; -- -0.1334946442082578
	pesos_i(18134) := b"1111111111111111_1111111111111111_1111111111101111_0011100000001111"; -- -0.00025605809641659355
	pesos_i(18135) := b"1111111111111111_1111111111111111_1110101111110011_0010110010000101"; -- -0.07832071060276351
	pesos_i(18136) := b"1111111111111111_1111111111111111_1111010101110100_1011100100100110"; -- -0.04118769470813452
	pesos_i(18137) := b"0000000000000000_0000000000000000_0001111011010010_1010000001000000"; -- 0.12040139744894572
	pesos_i(18138) := b"1111111111111111_1111111111111111_1101110011000100_1001111001010001"; -- -0.13762484096381974
	pesos_i(18139) := b"0000000000000000_0000000000000000_0000011110000011_1001011110010110"; -- 0.029351686655232072
	pesos_i(18140) := b"1111111111111111_1111111111111111_1110111011110001_0101110001101111"; -- -0.0666296223900038
	pesos_i(18141) := b"1111111111111111_1111111111111111_1101100011011101_0111111000110101"; -- -0.15287028503642175
	pesos_i(18142) := b"1111111111111111_1111111111111111_1111110000010101_1001001010100000"; -- -0.01529582580184986
	pesos_i(18143) := b"1111111111111111_1111111111111111_1111000111011111_1011000001000110"; -- -0.05518053323045195
	pesos_i(18144) := b"0000000000000000_0000000000000000_0010001100100000_0101100100000101"; -- 0.1372123371355524
	pesos_i(18145) := b"0000000000000000_0000000000000000_0001010001001010_1110000001110100"; -- 0.0792675289431457
	pesos_i(18146) := b"0000000000000000_0000000000000000_0000000010110100_1000101101110101"; -- 0.002754894339781602
	pesos_i(18147) := b"1111111111111111_1111111111111111_1111110010111110_0001111010100111"; -- -0.01272400297454591
	pesos_i(18148) := b"0000000000000000_0000000000000000_0000101110111100_1100101001000000"; -- 0.045849457449952245
	pesos_i(18149) := b"0000000000000000_0000000000000000_0001011001000000_1111110000101110"; -- 0.0869290936522282
	pesos_i(18150) := b"1111111111111111_1111111111111111_1101101011111101_0111010011001110"; -- -0.14457006438169473
	pesos_i(18151) := b"1111111111111111_1111111111111111_1111000000011111_1100100101011000"; -- -0.06201497640883795
	pesos_i(18152) := b"1111111111111111_1111111111111111_1110101000001100_0111001000000111"; -- -0.08574759791578104
	pesos_i(18153) := b"0000000000000000_0000000000000000_0010011010010110_0100000011000010"; -- 0.15073017829569385
	pesos_i(18154) := b"0000000000000000_0000000000000000_0001100100001010_0001111111111101"; -- 0.09781074464820594
	pesos_i(18155) := b"1111111111111111_1111111111111111_1111011001110111_0101110110100101"; -- -0.037241122403947
	pesos_i(18156) := b"0000000000000000_0000000000000000_0000110001001011_1110011101110010"; -- 0.048033204462643524
	pesos_i(18157) := b"0000000000000000_0000000000000000_0001101001101101_1111011101111010"; -- 0.1032404588311373
	pesos_i(18158) := b"1111111111111111_1111111111111111_1111110101101000_0000101000000100"; -- -0.010131238963162426
	pesos_i(18159) := b"1111111111111111_1111111111111111_1101100011000100_1011001101001110"; -- -0.15324858986124423
	pesos_i(18160) := b"1111111111111111_1111111111111111_1111010011100000_1011110111000010"; -- -0.043445720902381316
	pesos_i(18161) := b"1111111111111111_1111111111111111_1110010111000101_1111110100111010"; -- -0.10244767518296671
	pesos_i(18162) := b"0000000000000000_0000000000000000_0000011101001100_1111000100001100"; -- 0.028517785450961397
	pesos_i(18163) := b"0000000000000000_0000000000000000_0000111111101110_1011001001100011"; -- 0.06223597439842164
	pesos_i(18164) := b"1111111111111111_1111111111111111_1111111000000000_1110000000001111"; -- -0.0077991451686938995
	pesos_i(18165) := b"1111111111111111_1111111111111111_1101100001110111_0101110111010000"; -- -0.15442861245977518
	pesos_i(18166) := b"1111111111111111_1111111111111111_1110110101101000_0111001011000101"; -- -0.07262499518330047
	pesos_i(18167) := b"1111111111111111_1111111111111111_1111110101001111_1011110110000111"; -- -0.010502008950965402
	pesos_i(18168) := b"1111111111111111_1111111111111111_1101101001101100_1101101001100100"; -- -0.1467765336966902
	pesos_i(18169) := b"1111111111111111_1111111111111111_1111111111000110_0100010100010110"; -- -0.0008808918893813028
	pesos_i(18170) := b"1111111111111111_1111111111111111_1101100110010101_1110110100111001"; -- -0.15005605082523407
	pesos_i(18171) := b"1111111111111111_1111111111111111_1110111001000001_1111010010000010"; -- -0.06930610499768591
	pesos_i(18172) := b"0000000000000000_0000000000000000_0001100011100100_0100001010111110"; -- 0.09723298211877429
	pesos_i(18173) := b"0000000000000000_0000000000000000_0010001000110111_0001001100011101"; -- 0.1336528725943222
	pesos_i(18174) := b"1111111111111111_1111111111111111_1110001110110000_0110111000000100"; -- -0.11058914563356083
	pesos_i(18175) := b"1111111111111111_1111111111111111_1110111110000010_0101010110110010"; -- -0.06441749965766021
	pesos_i(18176) := b"0000000000000000_0000000000000000_0010010111001001_1000010110111111"; -- 0.14760623859747354
	pesos_i(18177) := b"0000000000000000_0000000000000000_0000101011000011_0001100011001001"; -- 0.04203944120121291
	pesos_i(18178) := b"0000000000000000_0000000000000000_0000101101100000_0001100010111001"; -- 0.04443506726839291
	pesos_i(18179) := b"0000000000000000_0000000000000000_0001001011100111_0111001100010111"; -- 0.07384414025057229
	pesos_i(18180) := b"1111111111111111_1111111111111111_1110111011111001_1110100011010000"; -- -0.06649918480444567
	pesos_i(18181) := b"1111111111111111_1111111111111111_1110101011111001_0001101110111011"; -- -0.08213640867145432
	pesos_i(18182) := b"0000000000000000_0000000000000000_0001000000011001_0010010101001100"; -- 0.06288369276626514
	pesos_i(18183) := b"1111111111111111_1111111111111111_1111100001101100_1100101100101111"; -- -0.029589940104455644
	pesos_i(18184) := b"0000000000000000_0000000000000000_0010010101011011_0000010011000011"; -- 0.145920083735456
	pesos_i(18185) := b"1111111111111111_1111111111111111_1110010011111001_0100001110011010"; -- -0.10557153217828938
	pesos_i(18186) := b"1111111111111111_1111111111111111_1110000011111101_0000100101110010"; -- -0.12113896328234343
	pesos_i(18187) := b"1111111111111111_1111111111111111_1110111111111010_1100000100011001"; -- -0.06258004313623627
	pesos_i(18188) := b"0000000000000000_0000000000000000_0001000110110110_0011011110001010"; -- 0.06918666006888927
	pesos_i(18189) := b"0000000000000000_0000000000000000_0000100010011101_1001001100111111"; -- 0.0336544063855515
	pesos_i(18190) := b"1111111111111111_1111111111111111_1111111111110110_1011101000101110"; -- -0.00014149073407783894
	pesos_i(18191) := b"1111111111111111_1111111111111111_1111000001101111_0101001011111111"; -- -0.06080132755658558
	pesos_i(18192) := b"1111111111111111_1111111111111111_1110011000100001_1011011000100100"; -- -0.10104810355430328
	pesos_i(18193) := b"1111111111111111_1111111111111111_1110001101011110_1101000001110000"; -- -0.11183450006398814
	pesos_i(18194) := b"0000000000000000_0000000000000000_0001111110100110_1110010100101010"; -- 0.12364036824270183
	pesos_i(18195) := b"1111111111111111_1111111111111111_1101100001000000_1111100111010010"; -- -0.1552585469985085
	pesos_i(18196) := b"0000000000000000_0000000000000000_0000010101010110_0111110100101101"; -- 0.020850966981188167
	pesos_i(18197) := b"0000000000000000_0000000000000000_0001100011101111_1100010001101100"; -- 0.09740855829009316
	pesos_i(18198) := b"1111111111111111_1111111111111111_1110100110110001_0110010110010011"; -- -0.08713688996672894
	pesos_i(18199) := b"1111111111111111_1111111111111111_1101111111100010_0001111110110000"; -- -0.12545587487888665
	pesos_i(18200) := b"1111111111111111_1111111111111111_1110100001111110_1101101000101001"; -- -0.0918143892572802
	pesos_i(18201) := b"0000000000000000_0000000000000000_0001011111111000_0111110001101010"; -- 0.09363534540216235
	pesos_i(18202) := b"0000000000000000_0000000000000000_0010001000010111_1001110011011001"; -- 0.13317280103681678
	pesos_i(18203) := b"0000000000000000_0000000000000000_0000110000111011_1010010101110001"; -- 0.04778512960697948
	pesos_i(18204) := b"0000000000000000_0000000000000000_0000011011010110_0100111001010001"; -- 0.026707548982034434
	pesos_i(18205) := b"0000000000000000_0000000000000000_0010000011010010_0001110111000010"; -- 0.12820611931936587
	pesos_i(18206) := b"1111111111111111_1111111111111111_1110001011010111_1101111011001001"; -- -0.11389358134557846
	pesos_i(18207) := b"0000000000000000_0000000000000000_0000100100010110_0110111001000101"; -- 0.035498515842386925
	pesos_i(18208) := b"1111111111111111_1111111111111111_1111111010100100_0011111010111111"; -- -0.005306318598692488
	pesos_i(18209) := b"0000000000000000_0000000000000000_0000111010101100_0100011000111111"; -- 0.05731619866352455
	pesos_i(18210) := b"0000000000000000_0000000000000000_0010100001110011_1010110110001010"; -- 0.1580151044209669
	pesos_i(18211) := b"1111111111111111_1111111111111111_1110001110110101_1111101001011101"; -- -0.11050448635269854
	pesos_i(18212) := b"1111111111111111_1111111111111111_1101111000000111_1000000010111100"; -- -0.13269801536355597
	pesos_i(18213) := b"0000000000000000_0000000000000000_0000110111001101_1100100001100001"; -- 0.05392124533315015
	pesos_i(18214) := b"1111111111111111_1111111111111111_1111101011000101_1111110111010111"; -- -0.020416388573204915
	pesos_i(18215) := b"1111111111111111_1111111111111111_1101100000101011_0011101110001101"; -- -0.1555903224639912
	pesos_i(18216) := b"0000000000000000_0000000000000000_0010010000101000_0011100100110001"; -- 0.14123876047400186
	pesos_i(18217) := b"1111111111111111_1111111111111111_1101110010101001_1111011011101111"; -- -0.13803154619665894
	pesos_i(18218) := b"1111111111111111_1111111111111111_1101011110001010_1111111000001001"; -- -0.15803539546666565
	pesos_i(18219) := b"0000000000000000_0000000000000000_0000100000000110_0010111100100010"; -- 0.031344362182159996
	pesos_i(18220) := b"1111111111111111_1111111111111111_1111010100010000_1110010010101000"; -- -0.042710980437417216
	pesos_i(18221) := b"0000000000000000_0000000000000000_0001101110100100_0001111110010111"; -- 0.10797307434975255
	pesos_i(18222) := b"0000000000000000_0000000000000000_0010000001101100_1100001100000111"; -- 0.12665957373094677
	pesos_i(18223) := b"0000000000000000_0000000000000000_0010001000001001_0101011101100101"; -- 0.1329550381416415
	pesos_i(18224) := b"0000000000000000_0000000000000000_0000111100101101_1101001000000100"; -- 0.05929291344291534
	pesos_i(18225) := b"0000000000000000_0000000000000000_0000111101011110_0001110001100011"; -- 0.06002976805002514
	pesos_i(18226) := b"1111111111111111_1111111111111111_1110000101000111_1011010100010110"; -- -0.11999958238974118
	pesos_i(18227) := b"0000000000000000_0000000000000000_0010001101101111_1101101111110110"; -- 0.13842558618697592
	pesos_i(18228) := b"1111111111111111_1111111111111111_1110100010000001_1010001011101111"; -- -0.0917719046394181
	pesos_i(18229) := b"0000000000000000_0000000000000000_0001000011000110_0100000111111010"; -- 0.06552517263642717
	pesos_i(18230) := b"0000000000000000_0000000000000000_0000010000001000_0111001110010000"; -- 0.015753958260440595
	pesos_i(18231) := b"1111111111111111_1111111111111111_1111011000101000_1100000000001101"; -- -0.03844070143097705
	pesos_i(18232) := b"1111111111111111_1111111111111111_1111010010101010_0111110101011001"; -- -0.04427353444797283
	pesos_i(18233) := b"1111111111111111_1111111111111111_1110101100010001_0001001110111100"; -- -0.08177067422307292
	pesos_i(18234) := b"1111111111111111_1111111111111111_1111010000010111_1000111011011001"; -- -0.046515533564303206
	pesos_i(18235) := b"0000000000000000_0000000000000000_0000010111111000_1001110011110101"; -- 0.023324784978771076
	pesos_i(18236) := b"1111111111111111_1111111111111111_1101101101100001_0000010110100000"; -- -0.14305081207134357
	pesos_i(18237) := b"1111111111111111_1111111111111111_1101110011011100_1111011000000100"; -- -0.13725340273666226
	pesos_i(18238) := b"1111111111111111_1111111111111111_1110010110001001_0011000001101100"; -- -0.10337540974376505
	pesos_i(18239) := b"1111111111111111_1111111111111111_1111100100101011_0010011100001011"; -- -0.026685295042151978
	pesos_i(18240) := b"1111111111111111_1111111111111111_1111001011111111_0000101110000001"; -- -0.050795823117853744
	pesos_i(18241) := b"1111111111111111_1111111111111111_1110111010010100_1100010100100010"; -- -0.06804244917351075
	pesos_i(18242) := b"1111111111111111_1111111111111111_1110011111000110_1111110111000111"; -- -0.0946198835473755
	pesos_i(18243) := b"0000000000000000_0000000000000000_0000111111111111_1001001110101100"; -- 0.06249354321052993
	pesos_i(18244) := b"0000000000000000_0000000000000000_0010000101001111_0010100100011010"; -- 0.13011414413538777
	pesos_i(18245) := b"1111111111111111_1111111111111111_1101111010110111_1111110110011001"; -- -0.13000502606451814
	pesos_i(18246) := b"0000000000000000_0000000000000000_0000101001111011_0010111111101011"; -- 0.04094218715475227
	pesos_i(18247) := b"1111111111111111_1111111111111111_1101110000100100_0000011011111001"; -- -0.14007526808736
	pesos_i(18248) := b"1111111111111111_1111111111111111_1101110000000110_1111000001011000"; -- -0.14051912176983927
	pesos_i(18249) := b"1111111111111111_1111111111111111_1111100100001111_0110010010010110"; -- -0.0271088727413804
	pesos_i(18250) := b"0000000000000000_0000000000000000_0000110111011001_0000101101101101"; -- 0.05409308821330565
	pesos_i(18251) := b"0000000000000000_0000000000000000_0000101100101101_0101010000000001"; -- 0.04366040242593532
	pesos_i(18252) := b"0000000000000000_0000000000000000_0000001100000100_0010100101111101"; -- 0.011782258131835954
	pesos_i(18253) := b"0000000000000000_0000000000000000_0001010001011110_0110010000101101"; -- 0.07956529710605743
	pesos_i(18254) := b"0000000000000000_0000000000000000_0001001011010101_0001011111000010"; -- 0.07356403823377643
	pesos_i(18255) := b"0000000000000000_0000000000000000_0000100100010000_0101000110101111"; -- 0.03540525939481123
	pesos_i(18256) := b"0000000000000000_0000000000000000_0000101111101000_1100010011101000"; -- 0.046520525608106024
	pesos_i(18257) := b"0000000000000000_0000000000000000_0001110111111100_1001100111011011"; -- 0.11713563536922758
	pesos_i(18258) := b"1111111111111111_1111111111111111_1110101101100000_1011010000100110"; -- -0.0805556686347302
	pesos_i(18259) := b"0000000000000000_0000000000000000_0000010111101001_1101110100000010"; -- 0.023099721043351215
	pesos_i(18260) := b"0000000000000000_0000000000000000_0000010110111011_1100001101101000"; -- 0.02239629070727741
	pesos_i(18261) := b"0000000000000000_0000000000000000_0000100011000111_0011110101011001"; -- 0.03429015559497483
	pesos_i(18262) := b"0000000000000000_0000000000000000_0001101010111110_0110110110001011"; -- 0.10446819920378526
	pesos_i(18263) := b"1111111111111111_1111111111111111_1110001100111001_0101000111000010"; -- -0.11240662583794425
	pesos_i(18264) := b"1111111111111111_1111111111111111_1110000110100101_0101001001000000"; -- -0.1185711473216663
	pesos_i(18265) := b"1111111111111111_1111111111111111_1110110010001101_0010101001110001"; -- -0.07597098105902687
	pesos_i(18266) := b"0000000000000000_0000000000000000_0000111101011001_0101010000101010"; -- 0.059956798724618225
	pesos_i(18267) := b"0000000000000000_0000000000000000_0001001001000001_1110110011010011"; -- 0.07131843712924833
	pesos_i(18268) := b"0000000000000000_0000000000000000_0001011000100010_1001111011100100"; -- 0.08646576941773504
	pesos_i(18269) := b"0000000000000000_0000000000000000_0010011010100101_1111011011001000"; -- 0.1509699094305101
	pesos_i(18270) := b"0000000000000000_0000000000000000_0001001011001001_1010010011011101"; -- 0.07338934312386684
	pesos_i(18271) := b"1111111111111111_1111111111111111_1111011010000011_0011100101111011"; -- -0.037060172614949184
	pesos_i(18272) := b"0000000000000000_0000000000000000_0001000110110000_0011001101111000"; -- 0.06909486473155768
	pesos_i(18273) := b"1111111111111111_1111111111111111_1111011100001110_0001001001111110"; -- -0.0349415247973331
	pesos_i(18274) := b"1111111111111111_1111111111111111_1111110011011000_1110111111001000"; -- -0.012314809533888471
	pesos_i(18275) := b"1111111111111111_1111111111111111_1111001100011000_0010000000100000"; -- -0.050413124169218185
	pesos_i(18276) := b"1111111111111111_1111111111111111_1111100010101111_1001101011011111"; -- -0.028570480761793252
	pesos_i(18277) := b"0000000000000000_0000000000000000_0010001101111110_1110100111100110"; -- 0.13865529876154337
	pesos_i(18278) := b"1111111111111111_1111111111111111_1111100000101100_0101000101001010"; -- -0.03057376816653111
	pesos_i(18279) := b"0000000000000000_0000000000000000_0000101111011101_1000100011100110"; -- 0.04634910211093119
	pesos_i(18280) := b"0000000000000000_0000000000000000_0000010001000101_1100110110011000"; -- 0.01669011080463517
	pesos_i(18281) := b"1111111111111111_1111111111111111_1110100001010110_1001011011000111"; -- -0.09242875707252705
	pesos_i(18282) := b"1111111111111111_1111111111111111_1111011110011110_1001011001110011"; -- -0.032736393903628355
	pesos_i(18283) := b"0000000000000000_0000000000000000_0000010010001101_0001110001101101"; -- 0.017778183520716907
	pesos_i(18284) := b"1111111111111111_1111111111111111_1110001100001011_0001111001100111"; -- -0.11311159129330882
	pesos_i(18285) := b"0000000000000000_0000000000000000_0000000111100011_0110000000111110"; -- 0.007375731596945751
	pesos_i(18286) := b"1111111111111111_1111111111111111_1111100011111110_0010001101101100"; -- -0.02737215638204402
	pesos_i(18287) := b"1111111111111111_1111111111111111_1111000100100011_0100101011011110"; -- -0.05805522987464827
	pesos_i(18288) := b"0000000000000000_0000000000000000_0001000110100001_1111110101010011"; -- 0.06887801442375
	pesos_i(18289) := b"1111111111111111_1111111111111111_1110010011010111_1001011111101111"; -- -0.1060853043302241
	pesos_i(18290) := b"0000000000000000_0000000000000000_0001010101101001_0011110001111101"; -- 0.08363702813674086
	pesos_i(18291) := b"0000000000000000_0000000000000000_0001000011111101_0111000000101000"; -- 0.06636715873942971
	pesos_i(18292) := b"1111111111111111_1111111111111111_1111011011001001_0011100101100101"; -- -0.03599206249059067
	pesos_i(18293) := b"0000000000000000_0000000000000000_0010101101111110_0000101111010010"; -- 0.1698920620110062
	pesos_i(18294) := b"0000000000000000_0000000000000000_0000000000001001_0110111011111101"; -- 0.00014394442703801456
	pesos_i(18295) := b"0000000000000000_0000000000000000_0010000100000001_1110101001110101"; -- 0.12893548352592638
	pesos_i(18296) := b"0000000000000000_0000000000000000_0000111001101011_1110011000000101"; -- 0.056333900570589804
	pesos_i(18297) := b"1111111111111111_1111111111111111_1110000111101100_1010100000011100"; -- -0.11748265572301649
	pesos_i(18298) := b"0000000000000000_0000000000000000_0000100101000010_0001100000100101"; -- 0.03616476921148134
	pesos_i(18299) := b"1111111111111111_1111111111111111_1101110100101101_0111111111000010"; -- -0.13602448949032242
	pesos_i(18300) := b"0000000000000000_0000000000000000_0000110000001000_0010000001100100"; -- 0.046999000910878226
	pesos_i(18301) := b"0000000000000000_0000000000000000_0000011111111111_0101110101011111"; -- 0.03124030646926699
	pesos_i(18302) := b"0000000000000000_0000000000000000_0001010010111011_0011101001011100"; -- 0.08098187202851505
	pesos_i(18303) := b"0000000000000000_0000000000000000_0001110001011101_1011100010000111"; -- 0.1108050660713207
	pesos_i(18304) := b"1111111111111111_1111111111111111_1110001000010010_1101110010010110"; -- -0.11689969374689341
	pesos_i(18305) := b"1111111111111111_1111111111111111_1111001010100110_1001111011011001"; -- -0.05214507298328112
	pesos_i(18306) := b"1111111111111111_1111111111111111_1111110111010010_0011101101100110"; -- -0.008510863958493957
	pesos_i(18307) := b"1111111111111111_1111111111111111_1110111000110000_0110100010011110"; -- -0.06957384255379341
	pesos_i(18308) := b"0000000000000000_0000000000000000_0000110010110001_0110001001001100"; -- 0.04958166451122973
	pesos_i(18309) := b"0000000000000000_0000000000000000_0000011111010110_1100010010110011"; -- 0.030620854936601976
	pesos_i(18310) := b"0000000000000000_0000000000000000_0000001110100000_1001000011100111"; -- 0.01416879304833929
	pesos_i(18311) := b"0000000000000000_0000000000000000_0000000011111101_0111110011011110"; -- 0.0038679161906017712
	pesos_i(18312) := b"0000000000000000_0000000000000000_0001001111110100_1110100011111001"; -- 0.07795578068751235
	pesos_i(18313) := b"0000000000000000_0000000000000000_0001000001110101_1001100001000101"; -- 0.06429435423630485
	pesos_i(18314) := b"1111111111111111_1111111111111111_1110010010101011_0010010110000000"; -- -0.10676351194407825
	pesos_i(18315) := b"1111111111111111_1111111111111111_1110011101100001_1000101100001100"; -- -0.09616785953567349
	pesos_i(18316) := b"0000000000000000_0000000000000000_0000011100000101_1010100000110010"; -- 0.027430069149138148
	pesos_i(18317) := b"1111111111111111_1111111111111111_1111011110011001_0100000111100110"; -- -0.03281772737054304
	pesos_i(18318) := b"1111111111111111_1111111111111111_1101110110100110_1101010111110100"; -- -0.13417303844336148
	pesos_i(18319) := b"0000000000000000_0000000000000000_0001100000011000_1111111010110010"; -- 0.09413139187733872
	pesos_i(18320) := b"1111111111111111_1111111111111111_1111100111111100_0101110010000111"; -- -0.023493020130474
	pesos_i(18321) := b"0000000000000000_0000000000000000_0010001110000001_1100101010000001"; -- 0.1386992039749548
	pesos_i(18322) := b"0000000000000000_0000000000000000_0001100011111110_1111101100001100"; -- 0.09764069598925736
	pesos_i(18323) := b"0000000000000000_0000000000000000_0010001110111001_0000011111000000"; -- 0.13954208786685007
	pesos_i(18324) := b"0000000000000000_0000000000000000_0000011001010001_1110010100000010"; -- 0.024687111912234615
	pesos_i(18325) := b"0000000000000000_0000000000000000_0000111111011101_0101101110111001"; -- 0.06197140954707293
	pesos_i(18326) := b"0000000000000000_0000000000000000_0000101001110000_0010000111111110"; -- 0.040773510524993166
	pesos_i(18327) := b"0000000000000000_0000000000000000_0010010111101111_1001010001001100"; -- 0.14818693976391367
	pesos_i(18328) := b"1111111111111111_1111111111111111_1111010110100001_0110100011111100"; -- -0.0405058273944226
	pesos_i(18329) := b"0000000000000000_0000000000000000_0001000100001001_0001110001100000"; -- 0.06654527028812406
	pesos_i(18330) := b"1111111111111111_1111111111111111_1101101000100101_1001101100000100"; -- -0.147863685183037
	pesos_i(18331) := b"1111111111111111_1111111111111111_1111111101001001_0110101011011100"; -- -0.002785989012148037
	pesos_i(18332) := b"1111111111111111_1111111111111111_1101111101011110_1110011000111010"; -- -0.1274582013141852
	pesos_i(18333) := b"1111111111111111_1111111111111111_1110011100101011_1110011001111101"; -- -0.09698638394118321
	pesos_i(18334) := b"0000000000000000_0000000000000000_0000111100000110_0000100011111011"; -- 0.058685837938477876
	pesos_i(18335) := b"1111111111111111_1111111111111111_1111011000111110_0001101101010000"; -- -0.038114827139819896
	pesos_i(18336) := b"0000000000000000_0000000000000000_0001110111001101_1001001011111111"; -- 0.11641806340595313
	pesos_i(18337) := b"1111111111111111_1111111111111111_1110111110001111_1010101111000010"; -- -0.06421400551135523
	pesos_i(18338) := b"0000000000000000_0000000000000000_0001010110110011_0011000000000111"; -- 0.08476543585937119
	pesos_i(18339) := b"0000000000000000_0000000000000000_0001011110000101_1011010111100111"; -- 0.09188401113392045
	pesos_i(18340) := b"1111111111111111_1111111111111111_1111100011111111_0101101010100110"; -- -0.0273536056376753
	pesos_i(18341) := b"1111111111111111_1111111111111111_1111011010101110_0010001000011100"; -- -0.036405437570248826
	pesos_i(18342) := b"1111111111111111_1111111111111111_1101100000000000_0000000101110001"; -- -0.1562499141607071
	pesos_i(18343) := b"1111111111111111_1111111111111111_1110111111100001_1010110011011011"; -- -0.06296271939431196
	pesos_i(18344) := b"0000000000000000_0000000000000000_0000001101111110_1100011101001001"; -- 0.01365323563724744
	pesos_i(18345) := b"0000000000000000_0000000000000000_0001000101100000_0100110010101110"; -- 0.06787566422550909
	pesos_i(18346) := b"0000000000000000_0000000000000000_0010000100100110_1001100010001011"; -- 0.12949517625336798
	pesos_i(18347) := b"0000000000000000_0000000000000000_0001010000001100_0010111111101111"; -- 0.07831096250142337
	pesos_i(18348) := b"1111111111111111_1111111111111111_1110110100000100_1111010010101111"; -- -0.07414313052020444
	pesos_i(18349) := b"0000000000000000_0000000000000000_0000001110011001_1001111110110000"; -- 0.01406286276822963
	pesos_i(18350) := b"1111111111111111_1111111111111111_1110101100111011_1011001101100101"; -- -0.08112028878467323
	pesos_i(18351) := b"1111111111111111_1111111111111111_1111000000111111_0010111001110111"; -- -0.0615359267962272
	pesos_i(18352) := b"1111111111111111_1111111111111111_1110100010010101_0101010011001001"; -- -0.09147138693244915
	pesos_i(18353) := b"0000000000000000_0000000000000000_0010010010001010_1011001001011111"; -- 0.14274134468266714
	pesos_i(18354) := b"0000000000000000_0000000000000000_0001001110010111_0001000110011000"; -- 0.07652387592323744
	pesos_i(18355) := b"0000000000000000_0000000000000000_0010011000100110_0100011000000001"; -- 0.14902150656455845
	pesos_i(18356) := b"0000000000000000_0000000000000000_0001001010111100_1110110111010110"; -- 0.07319532841293547
	pesos_i(18357) := b"1111111111111111_1111111111111111_1111111111011101_1101001000111000"; -- -0.0005215275517735135
	pesos_i(18358) := b"0000000000000000_0000000000000000_0001111111000101_1101010001100011"; -- 0.12411239069051534
	pesos_i(18359) := b"0000000000000000_0000000000000000_0000111000010110_1111110011100000"; -- 0.055038265875161245
	pesos_i(18360) := b"0000000000000000_0000000000000000_0000101001001000_0111010011110111"; -- 0.04016810448358907
	pesos_i(18361) := b"0000000000000000_0000000000000000_0001000101011010_0111000000001110"; -- 0.06778621997095943
	pesos_i(18362) := b"0000000000000000_0000000000000000_0010000001010101_0111111111010110"; -- 0.12630461661083137
	pesos_i(18363) := b"1111111111111111_1111111111111111_1110110100011110_0000100101010010"; -- -0.07376043086222278
	pesos_i(18364) := b"0000000000000000_0000000000000000_0001111100010111_1010000111000100"; -- 0.12145434413956117
	pesos_i(18365) := b"0000000000000000_0000000000000000_0001000001011111_1110000001000100"; -- 0.06396295233125406
	pesos_i(18366) := b"0000000000000000_0000000000000000_0001110111110011_0010110110110011"; -- 0.11699185962965153
	pesos_i(18367) := b"1111111111111111_1111111111111111_1111110011001111_0001011110010011"; -- -0.012465025423522753
	pesos_i(18368) := b"0000000000000000_0000000000000000_0000101101100111_0100011000111110"; -- 0.04454459196621891
	pesos_i(18369) := b"0000000000000000_0000000000000000_0010011110110000_1101100111010000"; -- 0.15504227939571547
	pesos_i(18370) := b"1111111111111111_1111111111111111_1110010110011011_0010011101011110"; -- -0.10310129127216107
	pesos_i(18371) := b"1111111111111111_1111111111111111_1101010101101100_0000011001011000"; -- -0.1663204226808688
	pesos_i(18372) := b"0000000000000000_0000000000000000_0000000101111101_1010100010011001"; -- 0.005823647723299726
	pesos_i(18373) := b"1111111111111111_1111111111111111_1111010010001010_0000010010001101"; -- -0.044769015927557644
	pesos_i(18374) := b"0000000000000000_0000000000000000_0000100010000000_1010111011001011"; -- 0.033213543585700354
	pesos_i(18375) := b"1111111111111111_1111111111111111_1111000001000110_0001111100000111"; -- -0.06143003548585724
	pesos_i(18376) := b"0000000000000000_0000000000000000_0000000000111100_1000101100011101"; -- 0.0009238191885113322
	pesos_i(18377) := b"0000000000000000_0000000000000000_0000111110110101_1101000010111010"; -- 0.06136803183547332
	pesos_i(18378) := b"0000000000000000_0000000000000000_0000001110100100_1011111110000000"; -- 0.014232605777746273
	pesos_i(18379) := b"1111111111111111_1111111111111111_1111111111010110_1110100110111101"; -- -0.0006269372292615222
	pesos_i(18380) := b"1111111111111111_1111111111111111_1101110111101101_1001010001000000"; -- -0.13309358056219592
	pesos_i(18381) := b"1111111111111111_1111111111111111_1110111001011001_0111100110000110"; -- -0.06894722434040103
	pesos_i(18382) := b"1111111111111111_1111111111111111_1101100101101000_1011001111000010"; -- -0.1507461215106802
	pesos_i(18383) := b"1111111111111111_1111111111111111_1111100010010100_0001010101000011"; -- -0.02899043203541305
	pesos_i(18384) := b"1111111111111111_1111111111111111_1110010001000000_1000001111110100"; -- -0.10839057242412635
	pesos_i(18385) := b"1111111111111111_1111111111111111_1111001000111001_1011010000011111"; -- -0.053807012903424614
	pesos_i(18386) := b"0000000000000000_0000000000000000_0000000101100110_0010000101101101"; -- 0.005464638848788495
	pesos_i(18387) := b"1111111111111111_1111111111111111_1110111111001000_1000011110000011"; -- -0.06334641495985263
	pesos_i(18388) := b"1111111111111111_1111111111111111_1111010011011110_1011001001000110"; -- -0.043476922970860025
	pesos_i(18389) := b"0000000000000000_0000000000000000_0001111110100001_1110111011101101"; -- 0.1235646560253243
	pesos_i(18390) := b"0000000000000000_0000000000000000_0000110110011100_0100001110010000"; -- 0.05316564812858459
	pesos_i(18391) := b"1111111111111111_1111111111111111_1111011100001101_0000011001101110"; -- -0.0349575025079323
	pesos_i(18392) := b"1111111111111111_1111111111111111_1101110100101001_0011001110001100"; -- -0.13609006729647433
	pesos_i(18393) := b"0000000000000000_0000000000000000_0001100101100101_1101010001001100"; -- 0.0992100414654155
	pesos_i(18394) := b"1111111111111111_1111111111111111_1111011101000011_0100000010001011"; -- -0.03413006405762892
	pesos_i(18395) := b"1111111111111111_1111111111111111_1111101001111111_0110101110111110"; -- -0.021493211875646335
	pesos_i(18396) := b"1111111111111111_1111111111111111_1111111110010110_1110111010100101"; -- -0.0016032072169293772
	pesos_i(18397) := b"1111111111111111_1111111111111111_1110111111111100_1100011001110011"; -- -0.06254920677518296
	pesos_i(18398) := b"1111111111111111_1111111111111111_1111101000110000_0101101100010101"; -- -0.022699649219498325
	pesos_i(18399) := b"1111111111111111_1111111111111111_1111000111100101_1100110110011101"; -- -0.05508723174411865
	pesos_i(18400) := b"0000000000000000_0000000000000000_0001110111010000_1110011001101101"; -- 0.11646881251258413
	pesos_i(18401) := b"0000000000000000_0000000000000000_0010000100110011_1100100101001110"; -- 0.12969644685551102
	pesos_i(18402) := b"1111111111111111_1111111111111111_1110000000111110_1011001001001111"; -- -0.12404332708138022
	pesos_i(18403) := b"1111111111111111_1111111111111111_1110111001101010_0100100011101001"; -- -0.06869072262354393
	pesos_i(18404) := b"0000000000000000_0000000000000000_0010011011101110_0000010000000101"; -- 0.15206933142693715
	pesos_i(18405) := b"0000000000000000_0000000000000000_0001000101001101_0101000010111001"; -- 0.06758598818294288
	pesos_i(18406) := b"0000000000000000_0000000000000000_0000100111010011_0110011011000100"; -- 0.03838197973432653
	pesos_i(18407) := b"0000000000000000_0000000000000000_0000000100110011_0000111011111010"; -- 0.004685340839785233
	pesos_i(18408) := b"1111111111111111_1111111111111111_1101100110111110_0000110111111001"; -- -0.14944374726969167
	pesos_i(18409) := b"0000000000000000_0000000000000000_0001111001110011_1111011111010100"; -- 0.1189570324101547
	pesos_i(18410) := b"0000000000000000_0000000000000000_0000010011010101_1010010111100111"; -- 0.018885010555010327
	pesos_i(18411) := b"1111111111111111_1111111111111111_1111000110011010_0101010101101001"; -- -0.056238805659882735
	pesos_i(18412) := b"1111111111111111_1111111111111111_1111101010010110_0010010010110110"; -- -0.021146493612114247
	pesos_i(18413) := b"1111111111111111_1111111111111111_1101110101110000_0110100000010001"; -- -0.13500356277855155
	pesos_i(18414) := b"0000000000000000_0000000000000000_0001111001111100_0100100011001111"; -- 0.11908392954277591
	pesos_i(18415) := b"0000000000000000_0000000000000000_0010001010011111_0010010100111111"; -- 0.13524086739973676
	pesos_i(18416) := b"1111111111111111_1111111111111111_1111101101011111_0011000001001111"; -- -0.01807878567679704
	pesos_i(18417) := b"1111111111111111_1111111111111111_1110100111000111_0111111000100000"; -- -0.08679973334879526
	pesos_i(18418) := b"1111111111111111_1111111111111111_1111110101101011_0000110010010111"; -- -0.010085309243599351
	pesos_i(18419) := b"0000000000000000_0000000000000000_0001001000100010_1101110000010101"; -- 0.07084441679280579
	pesos_i(18420) := b"0000000000000000_0000000000000000_0010001001010000_0010111000111100"; -- 0.13403595883065628
	pesos_i(18421) := b"1111111111111111_1111111111111111_1111010110111101_0110100100000110"; -- -0.04007857891329046
	pesos_i(18422) := b"0000000000000000_0000000000000000_0010011001011100_0111111010010110"; -- 0.14984885375887916
	pesos_i(18423) := b"0000000000000000_0000000000000000_0000101111011111_0110111010010100"; -- 0.04637805103148161
	pesos_i(18424) := b"0000000000000000_0000000000000000_0000101110001111_0110000100101111"; -- 0.04515654953133462
	pesos_i(18425) := b"0000000000000000_0000000000000000_0000010011010101_0111000101011101"; -- 0.018881878966589553
	pesos_i(18426) := b"0000000000000000_0000000000000000_0001001111010101_0101000010110011"; -- 0.07747368203148004
	pesos_i(18427) := b"1111111111111111_1111111111111111_1111110010110111_0011010001000110"; -- -0.012829525902218726
	pesos_i(18428) := b"1111111111111111_1111111111111111_1110011010011111_1100101110011101"; -- -0.09912421626066463
	pesos_i(18429) := b"1111111111111111_1111111111111111_1111010011110111_0010000001110111"; -- -0.0431041439768102
	pesos_i(18430) := b"0000000000000000_0000000000000000_0000100011010110_0011010001110011"; -- 0.03451850701513193
	pesos_i(18431) := b"0000000000000000_0000000000000000_0001100001111100_1010000011000010"; -- 0.0956516718455851
	pesos_i(18432) := b"1111111111111111_1111111111111111_1101011010011010_1111000100110101"; -- -0.16169826933459408
	pesos_i(18433) := b"1111111111111111_1111111111111111_1111000100001100_0110100101001001"; -- -0.05840436902923686
	pesos_i(18434) := b"0000000000000000_0000000000000000_0001000100101111_0100011011111111"; -- 0.06712764477994297
	pesos_i(18435) := b"1111111111111111_1111111111111111_1101111110101100_1001001100001011"; -- -0.12627297385441866
	pesos_i(18436) := b"0000000000000000_0000000000000000_0001000011101101_1111100100110100"; -- 0.0661311866350213
	pesos_i(18437) := b"0000000000000000_0000000000000000_0000001110011010_1110010110111101"; -- 0.014082296936417743
	pesos_i(18438) := b"1111111111111111_1111111111111111_1110000101001011_0011010111001000"; -- -0.11994613532436638
	pesos_i(18439) := b"1111111111111111_1111111111111111_1110001010011100_0001011001111011"; -- -0.11480578901424571
	pesos_i(18440) := b"0000000000000000_0000000000000000_0001000010010101_0101011010010011"; -- 0.06477871972572755
	pesos_i(18441) := b"1111111111111111_1111111111111111_1110000011001001_0000111001101011"; -- -0.12193212404498512
	pesos_i(18442) := b"1111111111111111_1111111111111111_1110100101011110_0100100101111011"; -- -0.08840504411297304
	pesos_i(18443) := b"0000000000000000_0000000000000000_0001000001100010_1100101110111111"; -- 0.0640075055170206
	pesos_i(18444) := b"0000000000000000_0000000000000000_0010000101001000_1100100001000001"; -- 0.13001681881071547
	pesos_i(18445) := b"1111111111111111_1111111111111111_1101110000100100_1001011100110110"; -- -0.14006667081081184
	pesos_i(18446) := b"0000000000000000_0000000000000000_0000000110011001_0111110100110111"; -- 0.006248308138912824
	pesos_i(18447) := b"0000000000000000_0000000000000000_0000010101010111_1101100000100000"; -- 0.02087164681023069
	pesos_i(18448) := b"0000000000000000_0000000000000000_0010011111110010_1000010111101011"; -- 0.15604435898939276
	pesos_i(18449) := b"1111111111111111_1111111111111111_1111010110100110_0110011101011001"; -- -0.04042963096900651
	pesos_i(18450) := b"0000000000000000_0000000000000000_0001110110111001_0100000010100100"; -- 0.11610797874399677
	pesos_i(18451) := b"1111111111111111_1111111111111111_1101111010100001_1101001010101111"; -- -0.13034327724643088
	pesos_i(18452) := b"1111111111111111_1111111111111111_1111010011010010_0001011011001010"; -- -0.04366929602385666
	pesos_i(18453) := b"0000000000000000_0000000000000000_0001100010111100_1010001111110111"; -- 0.09662842547065591
	pesos_i(18454) := b"1111111111111111_1111111111111111_1110001111011001_1010101100010010"; -- -0.10995989622978485
	pesos_i(18455) := b"1111111111111111_1111111111111111_1111011000111000_0001100101101000"; -- -0.0382064935370009
	pesos_i(18456) := b"1111111111111111_1111111111111111_1111011110101111_0010111011100101"; -- -0.03248316682139545
	pesos_i(18457) := b"0000000000000000_0000000000000000_0000111100101011_0111000100101001"; -- 0.05925662288858573
	pesos_i(18458) := b"1111111111111111_1111111111111111_1110110100111101_1001000111110100"; -- -0.07327926446219654
	pesos_i(18459) := b"0000000000000000_0000000000000000_0001111101101101_0100001010010110"; -- 0.12276092691140124
	pesos_i(18460) := b"0000000000000000_0000000000000000_0000100011101110_1111010000010100"; -- 0.034896140092429015
	pesos_i(18461) := b"0000000000000000_0000000000000000_0010001010101100_0101011111000000"; -- 0.13544224208218827
	pesos_i(18462) := b"1111111111111111_1111111111111111_1111100101011111_0001011010000011"; -- -0.02589282321496745
	pesos_i(18463) := b"1111111111111111_1111111111111111_1110001100100011_0111110101011001"; -- -0.11273972098894562
	pesos_i(18464) := b"0000000000000000_0000000000000000_0000010011000100_1011011101100110"; -- 0.01862665405883988
	pesos_i(18465) := b"1111111111111111_1111111111111111_1111011100111000_1011100111011011"; -- -0.034290679901939077
	pesos_i(18466) := b"1111111111111111_1111111111111111_1111111101111101_0101000100101111"; -- -0.001994062340202191
	pesos_i(18467) := b"1111111111111111_1111111111111111_1110001111101100_0101110110110101"; -- -0.10967459047614757
	pesos_i(18468) := b"1111111111111111_1111111111111111_1101110111000011_0011011001010001"; -- -0.13374004865365677
	pesos_i(18469) := b"1111111111111111_1111111111111111_1111000010001100_1011011000100110"; -- -0.06035291265121518
	pesos_i(18470) := b"1111111111111111_1111111111111111_1111111111011100_1011110011111011"; -- -0.0005380523345092267
	pesos_i(18471) := b"0000000000000000_0000000000000000_0001000101101110_0100111010101010"; -- 0.06808940558232743
	pesos_i(18472) := b"0000000000000000_0000000000000000_0000000100100101_0100100110000100"; -- 0.0044752070179712375
	pesos_i(18473) := b"1111111111111111_1111111111111111_1111101101111010_1010110010001001"; -- -0.017659393761038773
	pesos_i(18474) := b"1111111111111111_1111111111111111_1111111101100001_0101011001011100"; -- -0.002420999960232902
	pesos_i(18475) := b"1111111111111111_1111111111111111_1110111011000110_0111101100111001"; -- -0.0672839150672987
	pesos_i(18476) := b"0000000000000000_0000000000000000_0001101011010000_0001110000100101"; -- 0.10473800571768993
	pesos_i(18477) := b"1111111111111111_1111111111111111_1111100010100111_1101110111111101"; -- -0.028688550740048
	pesos_i(18478) := b"1111111111111111_1111111111111111_1101110001110110_1100001000001110"; -- -0.13881289633879898
	pesos_i(18479) := b"1111111111111111_1111111111111111_1111101001000000_0011010010110010"; -- -0.022457796689076635
	pesos_i(18480) := b"0000000000000000_0000000000000000_0001111010000011_1000100001110010"; -- 0.11919453425732161
	pesos_i(18481) := b"1111111111111111_1111111111111111_1111111011001000_1111001100110100"; -- -0.004746246235926547
	pesos_i(18482) := b"1111111111111111_1111111111111111_1101110001010001_1011010011000101"; -- -0.13937826344738571
	pesos_i(18483) := b"1111111111111111_1111111111111111_1101110100011000_0011110001001101"; -- -0.13634894490272553
	pesos_i(18484) := b"1111111111111111_1111111111111111_1101101010000111_1011100000110001"; -- -0.14636658484674814
	pesos_i(18485) := b"1111111111111111_1111111111111111_1110100100000010_1110011110111010"; -- -0.08979942033567098
	pesos_i(18486) := b"0000000000000000_0000000000000000_0000100100100010_1011001101010100"; -- 0.03568573765983039
	pesos_i(18487) := b"0000000000000000_0000000000000000_0010000010111101_1010010001100000"; -- 0.1278937085675676
	pesos_i(18488) := b"0000000000000000_0000000000000000_0010000011011100_0001101111000110"; -- 0.12835858891163432
	pesos_i(18489) := b"0000000000000000_0000000000000000_0000001001101101_0100101101100001"; -- 0.009480200927798528
	pesos_i(18490) := b"0000000000000000_0000000000000000_0001110111010001_0010011010101011"; -- 0.1164726418208684
	pesos_i(18491) := b"0000000000000000_0000000000000000_0000100011011111_1110110101110101"; -- 0.0346668635632585
	pesos_i(18492) := b"0000000000000000_0000000000000000_0000000110010110_1011011011001011"; -- 0.006205963612238759
	pesos_i(18493) := b"1111111111111111_1111111111111111_1110010111111111_1101111011100001"; -- -0.10156447427226735
	pesos_i(18494) := b"0000000000000000_0000000000000000_0000010101101100_1000010100010101"; -- 0.02118713142039958
	pesos_i(18495) := b"1111111111111111_1111111111111111_1110111000101001_0000110000100011"; -- -0.06968616632560734
	pesos_i(18496) := b"0000000000000000_0000000000000000_0000011001001110_1111000011010001"; -- 0.024642039277267314
	pesos_i(18497) := b"1111111111111111_1111111111111111_1111100100001011_0101000000000011"; -- -0.02717113431393039
	pesos_i(18498) := b"1111111111111111_1111111111111111_1101111000010000_0011110011010011"; -- -0.1325647340180042
	pesos_i(18499) := b"1111111111111111_1111111111111111_1111001110100011_1110011001001110"; -- -0.04828034011298936
	pesos_i(18500) := b"1111111111111111_1111111111111111_1111110000000110_1100101010101101"; -- -0.015521366951252422
	pesos_i(18501) := b"1111111111111111_1111111111111111_1101110100111100_1101101101000111"; -- -0.13579015266481798
	pesos_i(18502) := b"0000000000000000_0000000000000000_0000000011111010_1000010100011000"; -- 0.003822630374894476
	pesos_i(18503) := b"0000000000000000_0000000000000000_0001100101010011_1000000100001010"; -- 0.0989304207388043
	pesos_i(18504) := b"0000000000000000_0000000000000000_0000100001011001_1011010101100101"; -- 0.032618844120014916
	pesos_i(18505) := b"1111111111111111_1111111111111111_1110111111001000_0010010001100000"; -- -0.06335232418362349
	pesos_i(18506) := b"0000000000000000_0000000000000000_0010010001001001_0101000110100110"; -- 0.1417437581727964
	pesos_i(18507) := b"0000000000000000_0000000000000000_0001011011101010_1001101111100110"; -- 0.08951734881657909
	pesos_i(18508) := b"1111111111111111_1111111111111111_1110000001010110_0001111000001011"; -- -0.12368595335119924
	pesos_i(18509) := b"1111111111111111_1111111111111111_1111110101111101_0011011011111010"; -- -0.00980812443895292
	pesos_i(18510) := b"0000000000000000_0000000000000000_0000100000110000_1010000010011000"; -- 0.0319919939790142
	pesos_i(18511) := b"1111111111111111_1111111111111111_1110101010101010_0110110101101001"; -- -0.08333698449870186
	pesos_i(18512) := b"1111111111111111_1111111111111111_1111010110000000_0000001111010101"; -- -0.04101539647848442
	pesos_i(18513) := b"0000000000000000_0000000000000000_0000011000001101_1011111101010111"; -- 0.023647269090403097
	pesos_i(18514) := b"1111111111111111_1111111111111111_1110001010111110_1100000011001001"; -- -0.11427683922940543
	pesos_i(18515) := b"1111111111111111_1111111111111111_1110111100100100_0010100111111110"; -- -0.06585443073648227
	pesos_i(18516) := b"0000000000000000_0000000000000000_0000000001100001_1011110001101011"; -- 0.0014913331896465865
	pesos_i(18517) := b"1111111111111111_1111111111111111_1110000110000011_1011100001110000"; -- -0.11908385541287887
	pesos_i(18518) := b"0000000000000000_0000000000000000_0000101001111010_1001101111101100"; -- 0.04093336586689728
	pesos_i(18519) := b"1111111111111111_1111111111111111_1110000100010110_0100001010000010"; -- -0.12075409256447582
	pesos_i(18520) := b"1111111111111111_1111111111111111_1111110000101100_0111010011011001"; -- -0.014946648590032575
	pesos_i(18521) := b"1111111111111111_1111111111111111_1111111110100111_0101011001111000"; -- -0.001352878203349517
	pesos_i(18522) := b"0000000000000000_0000000000000000_0010010010000100_0110010111001101"; -- 0.14264522796299517
	pesos_i(18523) := b"1111111111111111_1111111111111111_1110110111010110_1111001011001100"; -- -0.0709388972614971
	pesos_i(18524) := b"1111111111111111_1111111111111111_1111001110000101_0110011100101000"; -- -0.048745682362097434
	pesos_i(18525) := b"0000000000000000_0000000000000000_0000000011010010_1010100100011011"; -- 0.0032144251786831468
	pesos_i(18526) := b"1111111111111111_1111111111111111_1101101110111111_1101110011010001"; -- -0.14160365960568522
	pesos_i(18527) := b"1111111111111111_1111111111111111_1110101110111110_1010000101010010"; -- -0.07912246469658227
	pesos_i(18528) := b"1111111111111111_1111111111111111_1111101110011010_0111001001001011"; -- -0.017174584035227074
	pesos_i(18529) := b"1111111111111111_1111111111111111_1101011101100111_0111011000011100"; -- -0.15857755497212447
	pesos_i(18530) := b"0000000000000000_0000000000000000_0010001100000010_1010001101011100"; -- 0.1367590044733976
	pesos_i(18531) := b"1111111111111111_1111111111111111_1110101010101011_0010101000001101"; -- -0.08332574073750978
	pesos_i(18532) := b"0000000000000000_0000000000000000_0010010000111100_1100010111111010"; -- 0.141552327582647
	pesos_i(18533) := b"0000000000000000_0000000000000000_0001111001010010_1001001101110111"; -- 0.1184475101854294
	pesos_i(18534) := b"1111111111111111_1111111111111111_1111000110110100_0101011010101000"; -- -0.055842002738011084
	pesos_i(18535) := b"1111111111111111_1111111111111111_1110001010100011_1110011010100001"; -- -0.11468657079422195
	pesos_i(18536) := b"0000000000000000_0000000000000000_0001110111000101_0011100011001111"; -- 0.11629061761424404
	pesos_i(18537) := b"1111111111111111_1111111111111111_1101111110101110_1010001111101001"; -- -0.12624145091888658
	pesos_i(18538) := b"0000000000000000_0000000000000000_0001100110011000_0001001000111101"; -- 0.09997667309630624
	pesos_i(18539) := b"1111111111111111_1111111111111111_1111100010001001_0010110111001110"; -- -0.029156815678312634
	pesos_i(18540) := b"0000000000000000_0000000000000000_0000001100101100_0010110111101001"; -- 0.012392873175461214
	pesos_i(18541) := b"0000000000000000_0000000000000000_0001110111010111_0011001011000100"; -- 0.11656491548296963
	pesos_i(18542) := b"0000000000000000_0000000000000000_0001000011110011_1101010001010010"; -- 0.06622054111073208
	pesos_i(18543) := b"0000000000000000_0000000000000000_0000101001010000_0001000111001000"; -- 0.040284262948940455
	pesos_i(18544) := b"0000000000000000_0000000000000000_0010000111101101_0111111111011100"; -- 0.13253020390799147
	pesos_i(18545) := b"1111111111111111_1111111111111111_1111000101111000_0110011110010011"; -- -0.056756521840224956
	pesos_i(18546) := b"0000000000000000_0000000000000000_0000000011111010_1000010111100100"; -- 0.003822677876467451
	pesos_i(18547) := b"1111111111111111_1111111111111111_1110100001000101_0111100010001011"; -- -0.09268995866307055
	pesos_i(18548) := b"1111111111111111_1111111111111111_1111100000001101_0111000001011111"; -- -0.031044937989575073
	pesos_i(18549) := b"0000000000000000_0000000000000000_0001000101111000_0011111000000110"; -- 0.06824100161496229
	pesos_i(18550) := b"0000000000000000_0000000000000000_0000000111001011_0111000011000111"; -- 0.007010506186391269
	pesos_i(18551) := b"0000000000000000_0000000000000000_0001000101110110_1010011010010101"; -- 0.06821671621392121
	pesos_i(18552) := b"1111111111111111_1111111111111111_1111010011010111_1110110111110110"; -- -0.043580176851582685
	pesos_i(18553) := b"0000000000000000_0000000000000000_0000101101010111_0101001011000000"; -- 0.044301196882061196
	pesos_i(18554) := b"1111111111111111_1111111111111111_1110110001001111_1100001110100100"; -- -0.07690789463335898
	pesos_i(18555) := b"1111111111111111_1111111111111111_1110110101100110_0100111001011100"; -- -0.07265768286712913
	pesos_i(18556) := b"0000000000000000_0000000000000000_0001100010000110_1010011000101101"; -- 0.09580458261406756
	pesos_i(18557) := b"1111111111111111_1111111111111111_1101100101010001_0011100011101110"; -- -0.15110439483077362
	pesos_i(18558) := b"1111111111111111_1111111111111111_1110010000001011_0111000111000001"; -- -0.10920037305788302
	pesos_i(18559) := b"0000000000000000_0000000000000000_0001101010110101_1010011110110001"; -- 0.10433433605597396
	pesos_i(18560) := b"0000000000000000_0000000000000000_0000011000100111_1011011011001100"; -- 0.024043488401447214
	pesos_i(18561) := b"0000000000000000_0000000000000000_0001111001001010_1111111100000010"; -- 0.11833185005149184
	pesos_i(18562) := b"1111111111111111_1111111111111111_1110010100000100_1010100010010011"; -- -0.10539766706675342
	pesos_i(18563) := b"1111111111111111_1111111111111111_1110100010101010_0101000111100100"; -- -0.09115112472933141
	pesos_i(18564) := b"0000000000000000_0000000000000000_0000101100011001_0111010010000110"; -- 0.04335716497573153
	pesos_i(18565) := b"0000000000000000_0000000000000000_0010001010011111_0101110110100101"; -- 0.13524422900148972
	pesos_i(18566) := b"0000000000000000_0000000000000000_0000001100001110_1101011000110010"; -- 0.011945140142822117
	pesos_i(18567) := b"1111111111111111_1111111111111111_1111101000111010_1001001110000010"; -- -0.022543698163413187
	pesos_i(18568) := b"1111111111111111_1111111111111111_1101101111111111_1000101000111101"; -- -0.14063201918959653
	pesos_i(18569) := b"1111111111111111_1111111111111111_1110101100100001_1000000100001000"; -- -0.0815200190998463
	pesos_i(18570) := b"0000000000000000_0000000000000000_0000001101100010_0011000000000100"; -- 0.01321697332425362
	pesos_i(18571) := b"0000000000000000_0000000000000000_0001101110100100_0010011010101001"; -- 0.1079734957520155
	pesos_i(18572) := b"0000000000000000_0000000000000000_0001101110001100_0110011111101001"; -- 0.10761117388917836
	pesos_i(18573) := b"0000000000000000_0000000000000000_0001011001111111_0011011011110110"; -- 0.08787864212256553
	pesos_i(18574) := b"0000000000000000_0000000000000000_0000001010010010_0100000110101100"; -- 0.010044197479749828
	pesos_i(18575) := b"0000000000000000_0000000000000000_0001000011101111_0110001101001001"; -- 0.06615276854314248
	pesos_i(18576) := b"0000000000000000_0000000000000000_0010010100001001_0011111011001111"; -- 0.14467232276153003
	pesos_i(18577) := b"1111111111111111_1111111111111111_1111010111001000_0010110100011011"; -- -0.039914303669425014
	pesos_i(18578) := b"0000000000000000_0000000000000000_0010000000110000_0101110000010000"; -- 0.12573790913417401
	pesos_i(18579) := b"0000000000000000_0000000000000000_0000111101110100_0011101011000100"; -- 0.06036727224083085
	pesos_i(18580) := b"0000000000000000_0000000000000000_0000101010011011_0110100110110101"; -- 0.04143391283016748
	pesos_i(18581) := b"0000000000000000_0000000000000000_0001001000011101_1111110000000000"; -- 0.07077002532697678
	pesos_i(18582) := b"1111111111111111_1111111111111111_1101111110100100_1001000011111101"; -- -0.12639516665371112
	pesos_i(18583) := b"0000000000000000_0000000000000000_0000011001110100_0001001010110100"; -- 0.02520863434998182
	pesos_i(18584) := b"0000000000000000_0000000000000000_0000100101101001_0011111110111010"; -- 0.036762221172873345
	pesos_i(18585) := b"0000000000000000_0000000000000000_0000110000001000_1111110101010011"; -- 0.04701216958369354
	pesos_i(18586) := b"1111111111111111_1111111111111111_1111111010101100_1001100100100011"; -- -0.005178860652659967
	pesos_i(18587) := b"1111111111111111_1111111111111111_1101110001101000_0111110011101110"; -- -0.13903063958360976
	pesos_i(18588) := b"0000000000000000_0000000000000000_0000111010000110_0011011110101010"; -- 0.0567354956516701
	pesos_i(18589) := b"1111111111111111_1111111111111111_1111000001111111_0101001110111000"; -- -0.06055714375077458
	pesos_i(18590) := b"0000000000000000_0000000000000000_0001001010000010_0101110100110001"; -- 0.07230169732853338
	pesos_i(18591) := b"1111111111111111_1111111111111111_1110101001111101_1100011000001110"; -- -0.08401834636473374
	pesos_i(18592) := b"0000000000000000_0000000000000000_0000110000111100_0100101010100000"; -- 0.04779497529746826
	pesos_i(18593) := b"0000000000000000_0000000000000000_0010100100110001_0001111100110010"; -- 0.16090579001426403
	pesos_i(18594) := b"1111111111111111_1111111111111111_1111011011101111_1101001011000110"; -- -0.0354030863784362
	pesos_i(18595) := b"1111111111111111_1111111111111111_1111000111000110_0101111010001010"; -- -0.05556687479297038
	pesos_i(18596) := b"1111111111111111_1111111111111111_1110110100111011_1001111111110110"; -- -0.07330894698060797
	pesos_i(18597) := b"1111111111111111_1111111111111111_1110000001101010_0111100001001011"; -- -0.12337539826522506
	pesos_i(18598) := b"0000000000000000_0000000000000000_0000010011101010_1010000110110110"; -- 0.019205195288128054
	pesos_i(18599) := b"1111111111111111_1111111111111111_1111010010000000_0111010001110101"; -- -0.04491493371907691
	pesos_i(18600) := b"1111111111111111_1111111111111111_1111101000011010_1000111111100110"; -- -0.02303219450155957
	pesos_i(18601) := b"0000000000000000_0000000000000000_0001101010000001_1101000111011101"; -- 0.1035433926046432
	pesos_i(18602) := b"0000000000000000_0000000000000000_0000000010000010_0001100001100001"; -- 0.001985095685341801
	pesos_i(18603) := b"1111111111111111_1111111111111111_1111101100011000_0101011111100101"; -- -0.019159800223860383
	pesos_i(18604) := b"1111111111111111_1111111111111111_1111010001000101_1010100110000101"; -- -0.04581203951863932
	pesos_i(18605) := b"0000000000000000_0000000000000000_0000111000111000_1011101011010001"; -- 0.055553127366327074
	pesos_i(18606) := b"0000000000000000_0000000000000000_0000000100100100_0011100001111001"; -- 0.0044589325209517215
	pesos_i(18607) := b"1111111111111111_1111111111111111_1101100011011111_1011101000111010"; -- -0.15283619002129942
	pesos_i(18608) := b"1111111111111111_1111111111111111_1101111010001010_1110001101000010"; -- -0.13069324154112882
	pesos_i(18609) := b"0000000000000000_0000000000000000_0001011101001111_0011111110001101"; -- 0.09105298236075572
	pesos_i(18610) := b"1111111111111111_1111111111111111_1110011111100111_0000110000011110"; -- -0.09413074754413642
	pesos_i(18611) := b"1111111111111111_1111111111111111_1101110100101010_1110100010100111"; -- -0.13606401360429543
	pesos_i(18612) := b"0000000000000000_0000000000000000_0001110101100001_1110010111100111"; -- 0.11477505570347295
	pesos_i(18613) := b"0000000000000000_0000000000000000_0001000110111000_0111000011001010"; -- 0.06922058999417743
	pesos_i(18614) := b"1111111111111111_1111111111111111_1111000110100001_0101001010001110"; -- -0.05613216423034888
	pesos_i(18615) := b"0000000000000000_0000000000000000_0010010010000111_1111011100011010"; -- 0.14269966497076514
	pesos_i(18616) := b"0000000000000000_0000000000000000_0001011100001001_1011111110101010"; -- 0.0899925032740418
	pesos_i(18617) := b"1111111111111111_1111111111111111_1110111101100010_1010011101011001"; -- -0.06490091387109362
	pesos_i(18618) := b"1111111111111111_1111111111111111_1110001101011110_1111100101010101"; -- -0.11183206249680568
	pesos_i(18619) := b"1111111111111111_1111111111111111_1110001010110001_0110110000010000"; -- -0.11448025321117146
	pesos_i(18620) := b"0000000000000000_0000000000000000_0000110000000010_0101001000111100"; -- 0.0469104191701934
	pesos_i(18621) := b"1111111111111111_1111111111111111_1110101010110111_0011111001101111"; -- -0.08314142038347434
	pesos_i(18622) := b"0000000000000000_0000000000000000_0010000100111000_0110001000011001"; -- 0.1297665892552909
	pesos_i(18623) := b"0000000000000000_0000000000000000_0000000110110101_0011110100011010"; -- 0.0066717327876560685
	pesos_i(18624) := b"0000000000000000_0000000000000000_0000011101000000_0000100100110100"; -- 0.028320861038210885
	pesos_i(18625) := b"0000000000000000_0000000000000000_0000010101111100_1111111110010100"; -- 0.02143857344113781
	pesos_i(18626) := b"1111111111111111_1111111111111111_1110101000001100_1001100101000111"; -- -0.08574525843136345
	pesos_i(18627) := b"0000000000000000_0000000000000000_0001010001111110_1110111011001011"; -- 0.08006184070483387
	pesos_i(18628) := b"0000000000000000_0000000000000000_0001001010100011_0101110100101100"; -- 0.07280523598187051
	pesos_i(18629) := b"1111111111111111_1111111111111111_1111110110001001_1000001110010111"; -- -0.009620452621071994
	pesos_i(18630) := b"1111111111111111_1111111111111111_1110101000011111_1110010101011010"; -- -0.08545080709581522
	pesos_i(18631) := b"1111111111111111_1111111111111111_1110001011010100_0110101000011000"; -- -0.11394631314377739
	pesos_i(18632) := b"1111111111111111_1111111111111111_1111101101001111_1011111110100010"; -- -0.018314383356450564
	pesos_i(18633) := b"1111111111111111_1111111111111111_1110110101001110_0010111000001011"; -- -0.07302581998366997
	pesos_i(18634) := b"1111111111111111_1111111111111111_1111110010100001_1000000100001101"; -- -0.013160642863885266
	pesos_i(18635) := b"1111111111111111_1111111111111111_1110000111010101_1000011111011001"; -- -0.11783553078333782
	pesos_i(18636) := b"0000000000000000_0000000000000000_0000000100010010_0001110100101111"; -- 0.004182647666589442
	pesos_i(18637) := b"0000000000000000_0000000000000000_0001110101010001_1010011000110001"; -- 0.11452711778309824
	pesos_i(18638) := b"1111111111111111_1111111111111111_1110010111110110_1001010101011001"; -- -0.10170618597564564
	pesos_i(18639) := b"1111111111111111_1111111111111111_1101101011110010_1010110001000000"; -- -0.14473460607591873
	pesos_i(18640) := b"1111111111111111_1111111111111111_1111111111001011_1111001010001110"; -- -0.0007942583259567971
	pesos_i(18641) := b"1111111111111111_1111111111111111_1111000001100011_0001110100001011"; -- -0.06098764876415752
	pesos_i(18642) := b"0000000000000000_0000000000000000_0001000000011001_1101000001010010"; -- 0.06289388646935483
	pesos_i(18643) := b"1111111111111111_1111111111111111_1111101100100110_1100010101001111"; -- -0.018939655550953314
	pesos_i(18644) := b"0000000000000000_0000000000000000_0000101110111101_0110001010011100"; -- 0.04585853863533134
	pesos_i(18645) := b"1111111111111111_1111111111111111_1111000011011111_1101110100101100"; -- -0.05908410718473014
	pesos_i(18646) := b"0000000000000000_0000000000000000_0010001110000011_0110100111010011"; -- 0.13872395909422283
	pesos_i(18647) := b"1111111111111111_1111111111111111_1101100101000011_1000111011010100"; -- -0.15131289783515153
	pesos_i(18648) := b"1111111111111111_1111111111111111_1111000100101001_1010000101101110"; -- -0.057958517615960777
	pesos_i(18649) := b"1111111111111111_1111111111111111_1101101010010101_1101010011011100"; -- -0.14615125302824133
	pesos_i(18650) := b"1111111111111111_1111111111111111_1110100011110010_0100111110011010"; -- -0.09005262851363337
	pesos_i(18651) := b"0000000000000000_0000000000000000_0001101001111110_0110110100110100"; -- 0.10349161633125216
	pesos_i(18652) := b"0000000000000000_0000000000000000_0010001100101100_1011000000101010"; -- 0.13740063694449006
	pesos_i(18653) := b"1111111111111111_1111111111111111_1111101100000100_0000000001100001"; -- -0.019470192264375363
	pesos_i(18654) := b"1111111111111111_1111111111111111_1101111110111011_1101010001010110"; -- -0.12604020030679355
	pesos_i(18655) := b"0000000000000000_0000000000000000_0010010100101100_0000101101101111"; -- 0.14520331828771665
	pesos_i(18656) := b"0000000000000000_0000000000000000_0010010000001011_0111111111001001"; -- 0.1408004633614573
	pesos_i(18657) := b"0000000000000000_0000000000000000_0001011000010010_1110000000100000"; -- 0.08622551714698057
	pesos_i(18658) := b"0000000000000000_0000000000000000_0000010001000100_0010100011110110"; -- 0.016665039003192286
	pesos_i(18659) := b"1111111111111111_1111111111111111_1111111000011111_0011101101010100"; -- -0.007335941386452526
	pesos_i(18660) := b"0000000000000000_0000000000000000_0000000010101100_0110011100011110"; -- 0.002630658021217371
	pesos_i(18661) := b"1111111111111111_1111111111111111_1110001000011001_1101100110011001"; -- -0.11679306041517032
	pesos_i(18662) := b"0000000000000000_0000000000000000_0000001011010010_0011011111111010"; -- 0.011020182156132288
	pesos_i(18663) := b"0000000000000000_0000000000000000_0010001101001011_0010101010111011"; -- 0.1378657061007508
	pesos_i(18664) := b"0000000000000000_0000000000000000_0001001110000010_0011010011010011"; -- 0.07620554118091094
	pesos_i(18665) := b"1111111111111111_1111111111111111_1111010011001110_1100001010100100"; -- -0.043720088054096586
	pesos_i(18666) := b"1111111111111111_1111111111111111_1111010011101110_0110001011110101"; -- -0.04323750986967929
	pesos_i(18667) := b"0000000000000000_0000000000000000_0000110010010011_1011101000100010"; -- 0.049129136294950596
	pesos_i(18668) := b"0000000000000000_0000000000000000_0000010010000011_0110010111100101"; -- 0.01762997476223438
	pesos_i(18669) := b"0000000000000000_0000000000000000_0010011001011100_1101111010001000"; -- 0.14985457237916788
	pesos_i(18670) := b"1111111111111111_1111111111111111_1101010100111011_1000001101101000"; -- -0.167060648982371
	pesos_i(18671) := b"0000000000000000_0000000000000000_0010000100100000_1110000010011010"; -- 0.12940791855898873
	pesos_i(18672) := b"1111111111111111_1111111111111111_1101101101110010_1000100001101111"; -- -0.14278361593992653
	pesos_i(18673) := b"1111111111111111_1111111111111111_1110110101110110_1111111000110110"; -- -0.07240306081039143
	pesos_i(18674) := b"0000000000000000_0000000000000000_0001000110110101_1101101110000101"; -- 0.06918117522556624
	pesos_i(18675) := b"1111111111111111_1111111111111111_1101110110010011_1001010010000001"; -- -0.13446685651819246
	pesos_i(18676) := b"1111111111111111_1111111111111111_1101010111001111_0101001110100111"; -- -0.1648051946439838
	pesos_i(18677) := b"1111111111111111_1111111111111111_1110101000011000_0111110100001001"; -- -0.08556383630199575
	pesos_i(18678) := b"0000000000000000_0000000000000000_0000111111000000_0111111001011000"; -- 0.06153096812293327
	pesos_i(18679) := b"1111111111111111_1111111111111111_1111110110111001_0101001000011010"; -- -0.008890980312454257
	pesos_i(18680) := b"1111111111111111_1111111111111111_1111111011111011_0010110100000111"; -- -0.003979860054626265
	pesos_i(18681) := b"1111111111111111_1111111111111111_1111000011110101_0100101110111100"; -- -0.05875708257711604
	pesos_i(18682) := b"1111111111111111_1111111111111111_1110001111000001_1100110101000111"; -- -0.11032406823305489
	pesos_i(18683) := b"0000000000000000_0000000000000000_0000010001011100_1101010110100101"; -- 0.017041542846420055
	pesos_i(18684) := b"1111111111111111_1111111111111111_1101101000011100_1101011010010100"; -- -0.14799746395921423
	pesos_i(18685) := b"1111111111111111_1111111111111111_1110100000110100_1111110101001111"; -- -0.09294144451278478
	pesos_i(18686) := b"1111111111111111_1111111111111111_1110010011111110_1101001100111010"; -- -0.10548667739156753
	pesos_i(18687) := b"0000000000000000_0000000000000000_0000111010100011_1000010010111010"; -- 0.05718259369946181
	pesos_i(18688) := b"1111111111111111_1111111111111111_1110000011010100_1000000111110110"; -- -0.12175739033244569
	pesos_i(18689) := b"0000000000000000_0000000000000000_0001001100011000_0010110110111111"; -- 0.07458768763723668
	pesos_i(18690) := b"1111111111111111_1111111111111111_1110001111110010_0001001001101000"; -- -0.10958752592647165
	pesos_i(18691) := b"1111111111111111_1111111111111111_1110001101000111_0011100100101111"; -- -0.11219446767680007
	pesos_i(18692) := b"0000000000000000_0000000000000000_0010010111100101_1111101000010111"; -- 0.14804041925694378
	pesos_i(18693) := b"1111111111111111_1111111111111111_1111000111100001_0000011111100101"; -- -0.0551600518138729
	pesos_i(18694) := b"1111111111111111_1111111111111111_1101111111000010_1111000100111011"; -- -0.12593166648743154
	pesos_i(18695) := b"1111111111111111_1111111111111111_1110111011101100_1110011100111100"; -- -0.06669764312026255
	pesos_i(18696) := b"1111111111111111_1111111111111111_1111110101101010_0001101001110001"; -- -0.010099742347976757
	pesos_i(18697) := b"0000000000000000_0000000000000000_0000101001111101_1000011000101101"; -- 0.040977846226960664
	pesos_i(18698) := b"0000000000000000_0000000000000000_0001000101001000_1111000111110111"; -- 0.0675193051119273
	pesos_i(18699) := b"1111111111111111_1111111111111111_1111000010101100_1010110011100100"; -- -0.05986518329132479
	pesos_i(18700) := b"0000000000000000_0000000000000000_0000111000111010_0010001101100100"; -- 0.055574619290103815
	pesos_i(18701) := b"1111111111111111_1111111111111111_1110001010001001_0111101011111110"; -- -0.11508971501574994
	pesos_i(18702) := b"0000000000000000_0000000000000000_0000001100000111_0111110100101001"; -- 0.011833021635147975
	pesos_i(18703) := b"1111111111111111_1111111111111111_1110110011111011_0100000000010001"; -- -0.0742912252845664
	pesos_i(18704) := b"0000000000000000_0000000000000000_0000110100001000_0011111101100000"; -- 0.0509070977325957
	pesos_i(18705) := b"0000000000000000_0000000000000000_0001101100101111_0000101011000011"; -- 0.10618655460210792
	pesos_i(18706) := b"0000000000000000_0000000000000000_0010001111010101_0101000100110100"; -- 0.13997371212534795
	pesos_i(18707) := b"0000000000000000_0000000000000000_0000100101010011_1010100110110100"; -- 0.03643284453740907
	pesos_i(18708) := b"1111111111111111_1111111111111111_1110010100000111_0001111011000001"; -- -0.10536010533565558
	pesos_i(18709) := b"1111111111111111_1111111111111111_1110011100011101_0000110111110110"; -- -0.0972129128684579
	pesos_i(18710) := b"1111111111111111_1111111111111111_1111001110000101_0110111011000110"; -- -0.048745228418871016
	pesos_i(18711) := b"0000000000000000_0000000000000000_0000101001100010_1110011001100001"; -- 0.040571592960678464
	pesos_i(18712) := b"1111111111111111_1111111111111111_1110100011001110_1010001010100111"; -- -0.09059699470308756
	pesos_i(18713) := b"0000000000000000_0000000000000000_0001110001101100_1001101110111100"; -- 0.111032231702692
	pesos_i(18714) := b"0000000000000000_0000000000000000_0000101010001111_1001101010011000"; -- 0.04125372142959966
	pesos_i(18715) := b"0000000000000000_0000000000000000_0001110010111111_1110100101110000"; -- 0.11230334262095203
	pesos_i(18716) := b"0000000000000000_0000000000000000_0010001101010101_0100001101101101"; -- 0.13801976593451054
	pesos_i(18717) := b"0000000000000000_0000000000000000_0001111101110010_1010111111110100"; -- 0.12284373966234041
	pesos_i(18718) := b"1111111111111111_1111111111111111_1101110111010110_0011001101100011"; -- -0.1334503062675391
	pesos_i(18719) := b"0000000000000000_0000000000000000_0000011111011111_0111110110101011"; -- 0.030753950358173583
	pesos_i(18720) := b"1111111111111111_1111111111111111_1101101111101110_1100100100100000"; -- -0.1408876701309022
	pesos_i(18721) := b"0000000000000000_0000000000000000_0001001110111100_1001011000001101"; -- 0.0770963461071128
	pesos_i(18722) := b"0000000000000000_0000000000000000_0001010101000110_1011000101010100"; -- 0.08310993490512085
	pesos_i(18723) := b"1111111111111111_1111111111111111_1110101000011001_0111001001000011"; -- -0.08554921973465336
	pesos_i(18724) := b"0000000000000000_0000000000000000_0010001110101001_1100100011000100"; -- 0.139309451828943
	pesos_i(18725) := b"1111111111111111_1111111111111111_1110001111000100_1010110111110100"; -- -0.11028015902028881
	pesos_i(18726) := b"0000000000000000_0000000000000000_0001101011100110_0111010100110111"; -- 0.1050790080749166
	pesos_i(18727) := b"1111111111111111_1111111111111111_1110110111110110_1011010011100000"; -- -0.07045430687694378
	pesos_i(18728) := b"1111111111111111_1111111111111111_1111111011011100_1111000111000000"; -- -0.004441156947971604
	pesos_i(18729) := b"0000000000000000_0000000000000000_0000000100101010_0001001110001110"; -- 0.004548284666480122
	pesos_i(18730) := b"1111111111111111_1111111111111111_1110100100001010_1010011110000000"; -- -0.08968117834782106
	pesos_i(18731) := b"0000000000000000_0000000000000000_0001100010010101_1010111101000000"; -- 0.09603400539651778
	pesos_i(18732) := b"0000000000000000_0000000000000000_0010011010011000_0110101111010000"; -- 0.15076326196917786
	pesos_i(18733) := b"0000000000000000_0000000000000000_0000001111101010_0101010000010101"; -- 0.01529431832222831
	pesos_i(18734) := b"0000000000000000_0000000000000000_0001110110101011_0111101010101100"; -- 0.1158978146442145
	pesos_i(18735) := b"1111111111111111_1111111111111111_1111001010010001_1001101101101010"; -- -0.052465712097771476
	pesos_i(18736) := b"1111111111111111_1111111111111111_1110011101110010_0100111011010010"; -- -0.0959120500422205
	pesos_i(18737) := b"1111111111111111_1111111111111111_1111110011110011_1011010110110011"; -- -0.011906284228731608
	pesos_i(18738) := b"0000000000000000_0000000000000000_0000010100100100_0100011111011101"; -- 0.020084849678310757
	pesos_i(18739) := b"1111111111111111_1111111111111111_1110111011101011_1110011001101001"; -- -0.06671295108437961
	pesos_i(18740) := b"0000000000000000_0000000000000000_0000010011011110_0011010000100110"; -- 0.019015559482884022
	pesos_i(18741) := b"0000000000000000_0000000000000000_0001011111110101_1011101001100111"; -- 0.09359326369201491
	pesos_i(18742) := b"1111111111111111_1111111111111111_1110000011100010_0101011001010100"; -- -0.12154636815822654
	pesos_i(18743) := b"0000000000000000_0000000000000000_0001101000110110_0000000010001010"; -- 0.10238650674966404
	pesos_i(18744) := b"1111111111111111_1111111111111111_1111000011110101_1010010000100111"; -- -0.058751812351055775
	pesos_i(18745) := b"1111111111111111_1111111111111111_1111110001001010_1000110011110100"; -- -0.014487448081784636
	pesos_i(18746) := b"1111111111111111_1111111111111111_1111010101001001_0001011011101011"; -- -0.04185349243494914
	pesos_i(18747) := b"1111111111111111_1111111111111111_1111111110110100_1100011010111011"; -- -0.0011478226652818647
	pesos_i(18748) := b"1111111111111111_1111111111111111_1111100111011011_0111111100000111"; -- -0.023994503721378294
	pesos_i(18749) := b"0000000000000000_0000000000000000_0000011101001110_0101100011011010"; -- 0.028539231501719553
	pesos_i(18750) := b"1111111111111111_1111111111111111_1110110100010010_1110010001100010"; -- -0.07393047911748238
	pesos_i(18751) := b"0000000000000000_0000000000000000_0000010100000010_1011010110000110"; -- 0.019572587271859135
	pesos_i(18752) := b"0000000000000000_0000000000000000_0010001100010001_1111101001100000"; -- 0.13699307292034588
	pesos_i(18753) := b"0000000000000000_0000000000000000_0001111001000000_1101000100111000"; -- 0.11817653280067308
	pesos_i(18754) := b"0000000000000000_0000000000000000_0000001001011011_1000111111101110"; -- 0.009209628710630724
	pesos_i(18755) := b"0000000000000000_0000000000000000_0010001001101111_1001100111010001"; -- 0.13451539371849866
	pesos_i(18756) := b"1111111111111111_1111111111111111_1111101011101100_0000101101001111"; -- -0.01983575166357714
	pesos_i(18757) := b"0000000000000000_0000000000000000_0010011000001000_1101110111100001"; -- 0.14857279532924447
	pesos_i(18758) := b"1111111111111111_1111111111111111_1110101111000111_1100101001010100"; -- -0.0789826911890403
	pesos_i(18759) := b"1111111111111111_1111111111111111_1111010001010011_0100001011110001"; -- -0.045604530516536596
	pesos_i(18760) := b"0000000000000000_0000000000000000_0001100000011010_0001111101011011"; -- 0.09414859739663448
	pesos_i(18761) := b"1111111111111111_1111111111111111_1111110010011100_0001000001100010"; -- -0.013243652339641039
	pesos_i(18762) := b"1111111111111111_1111111111111111_1111000111010001_1011111010011010"; -- -0.05539330228789527
	pesos_i(18763) := b"1111111111111111_1111111111111111_1110001110110110_1010000010111111"; -- -0.11049456907793702
	pesos_i(18764) := b"0000000000000000_0000000000000000_0000100101110010_1011011010000000"; -- 0.03690662973912206
	pesos_i(18765) := b"1111111111111111_1111111111111111_1110001011000000_1111111100010110"; -- -0.11424260816490645
	pesos_i(18766) := b"1111111111111111_1111111111111111_1101100011000011_1111101010110010"; -- -0.15325959354220828
	pesos_i(18767) := b"1111111111111111_1111111111111111_1110110010010100_1001111100011111"; -- -0.07585721476142851
	pesos_i(18768) := b"0000000000000000_0000000000000000_0001010000011111_0011000011111101"; -- 0.07860094234903987
	pesos_i(18769) := b"1111111111111111_1111111111111111_1111000101010000_0000110111000010"; -- -0.05737222673408685
	pesos_i(18770) := b"1111111111111111_1111111111111111_1110010011111000_1010100110111001"; -- -0.10558070411840365
	pesos_i(18771) := b"1111111111111111_1111111111111111_1111011110011000_0100011000001010"; -- -0.03283273951909032
	pesos_i(18772) := b"1111111111111111_1111111111111111_1110001100101010_0100110001001111"; -- -0.11263583248646354
	pesos_i(18773) := b"0000000000000000_0000000000000000_0010000100111111_0010111111000000"; -- 0.1298703997411407
	pesos_i(18774) := b"0000000000000000_0000000000000000_0001000011101010_0100010010000111"; -- 0.06607464121073214
	pesos_i(18775) := b"1111111111111111_1111111111111111_1110000101011001_1010110010100101"; -- -0.11972542736319747
	pesos_i(18776) := b"1111111111111111_1111111111111111_1111100101011000_0101100100011001"; -- -0.02599566589626449
	pesos_i(18777) := b"0000000000000000_0000000000000000_0001000011111101_0011101000111010"; -- 0.0663639441456882
	pesos_i(18778) := b"1111111111111111_1111111111111111_1110010000000110_1110100101010110"; -- -0.10926953938314544
	pesos_i(18779) := b"0000000000000000_0000000000000000_0010001001100101_0111011010101110"; -- 0.1343607114634737
	pesos_i(18780) := b"0000000000000000_0000000000000000_0000011101111000_0000011110100011"; -- 0.029175259924582767
	pesos_i(18781) := b"0000000000000000_0000000000000000_0001101100111100_0111000010101101"; -- 0.10639099333285305
	pesos_i(18782) := b"1111111111111111_1111111111111111_1111011010001111_1101110001110110"; -- -0.03686735255391565
	pesos_i(18783) := b"0000000000000000_0000000000000000_0001010000001111_1011010100101001"; -- 0.07836467990480923
	pesos_i(18784) := b"1111111111111111_1111111111111111_1110110001001010_1101011010110000"; -- -0.07698305326599802
	pesos_i(18785) := b"0000000000000000_0000000000000000_0010101011111000_1000111110111001"; -- 0.16785524630097062
	pesos_i(18786) := b"0000000000000000_0000000000000000_0000011101011100_0101110001101000"; -- 0.028753066442672247
	pesos_i(18787) := b"1111111111111111_1111111111111111_1111111101100111_0010110111000011"; -- -0.002331867229597103
	pesos_i(18788) := b"0000000000000000_0000000000000000_0000011101000111_1110101110111010"; -- 0.028441174318643073
	pesos_i(18789) := b"1111111111111111_1111111111111111_1101111011000110_0001100011010001"; -- -0.12978978051929452
	pesos_i(18790) := b"1111111111111111_1111111111111111_1111011110100100_1101111100101100"; -- -0.03264050661965218
	pesos_i(18791) := b"1111111111111111_1111111111111111_1110100001101100_0001100000110111"; -- -0.0921006075535168
	pesos_i(18792) := b"0000000000000000_0000000000000000_0000100001010111_1010100010111001"; -- 0.03258757139105299
	pesos_i(18793) := b"0000000000000000_0000000000000000_0001001100111001_1000111011000110"; -- 0.07509701092664224
	pesos_i(18794) := b"0000000000000000_0000000000000000_0001111110001100_0101111101011010"; -- 0.12323566391441647
	pesos_i(18795) := b"0000000000000000_0000000000000000_0000101101110101_1011101001110010"; -- 0.04476514131804277
	pesos_i(18796) := b"0000000000000000_0000000000000000_0000101001100110_0001110110000101"; -- 0.040620656067891545
	pesos_i(18797) := b"0000000000000000_0000000000000000_0000101011111000_1010100101101001"; -- 0.042856777235731655
	pesos_i(18798) := b"1111111111111111_1111111111111111_1111101001011101_0111111111000011"; -- -0.02201081747050131
	pesos_i(18799) := b"1111111111111111_1111111111111111_1110101101000001_1010000101101111"; -- -0.08102980650751261
	pesos_i(18800) := b"0000000000000000_0000000000000000_0000000011000001_1010100011000000"; -- 0.0029550045245781203
	pesos_i(18801) := b"0000000000000000_0000000000000000_0001101011000110_1001101100001101"; -- 0.10459298197332327
	pesos_i(18802) := b"0000000000000000_0000000000000000_0010100100000010_1011001011011010"; -- 0.16019742795061326
	pesos_i(18803) := b"0000000000000000_0000000000000000_0000001000001011_1011110111011001"; -- 0.007991662365680701
	pesos_i(18804) := b"1111111111111111_1111111111111111_1110111001010100_1111100101000111"; -- -0.0690159037209033
	pesos_i(18805) := b"1111111111111111_1111111111111111_1110010010000100_1111101101001100"; -- -0.10734586144637989
	pesos_i(18806) := b"0000000000000000_0000000000000000_0010010111101000_1100010001100000"; -- 0.14808299384888754
	pesos_i(18807) := b"1111111111111111_1111111111111111_1111111111011101_0100011000111100"; -- -0.0005298712443750961
	pesos_i(18808) := b"1111111111111111_1111111111111111_1101111101011010_0111100110000010"; -- -0.12752571662720652
	pesos_i(18809) := b"1111111111111111_1111111111111111_1111001000010110_1011000011110011"; -- -0.05434125967962772
	pesos_i(18810) := b"1111111111111111_1111111111111111_1101101000101001_0100000111001110"; -- -0.1478079674647458
	pesos_i(18811) := b"0000000000000000_0000000000000000_0010000111111001_1001001011110000"; -- 0.1327144467227223
	pesos_i(18812) := b"1111111111111111_1111111111111111_1101011110111011_0101111001010110"; -- -0.1572972336962843
	pesos_i(18813) := b"1111111111111111_1111111111111111_1111000101101010_1111110100001011"; -- -0.056961235831285664
	pesos_i(18814) := b"0000000000000000_0000000000000000_0000110010000001_0010000000001100"; -- 0.04884529403108572
	pesos_i(18815) := b"0000000000000000_0000000000000000_0010010010110110_1010100001010001"; -- 0.1434121320530365
	pesos_i(18816) := b"0000000000000000_0000000000000000_0000100011110010_1011010111111000"; -- 0.03495347317502851
	pesos_i(18817) := b"0000000000000000_0000000000000000_0000100011100111_1011011001000000"; -- 0.03478564314372375
	pesos_i(18818) := b"0000000000000000_0000000000000000_0000101111100110_1100100111011010"; -- 0.04649030276690075
	pesos_i(18819) := b"1111111111111111_1111111111111111_1110000111111010_0100001010110000"; -- -0.1172750778942945
	pesos_i(18820) := b"0000000000000000_0000000000000000_0000100010100100_0110010111111011"; -- 0.033758519974602524
	pesos_i(18821) := b"0000000000000000_0000000000000000_0000111001110001_0111001000000110"; -- 0.056418539520244504
	pesos_i(18822) := b"0000000000000000_0000000000000000_0000111101100110_0100011000010100"; -- 0.06015432357031417
	pesos_i(18823) := b"1111111111111111_1111111111111111_1111010100000001_1101111000100011"; -- -0.042940250795633884
	pesos_i(18824) := b"1111111111111111_1111111111111111_1111001000100001_1110000110101101"; -- -0.05417050873767823
	pesos_i(18825) := b"1111111111111111_1111111111111111_1111101100101010_0010100011011010"; -- -0.01888794590870235
	pesos_i(18826) := b"1111111111111111_1111111111111111_1110111011100011_0110011100001011"; -- -0.06684261305897257
	pesos_i(18827) := b"1111111111111111_1111111111111111_1110000010110101_1011011111110110"; -- -0.12222719427238811
	pesos_i(18828) := b"0000000000000000_0000000000000000_0000000110000001_0110010010100001"; -- 0.005880631773180021
	pesos_i(18829) := b"0000000000000000_0000000000000000_0010000011011111_0111101110111001"; -- 0.1284100843363569
	pesos_i(18830) := b"0000000000000000_0000000000000000_0010010110101110_1000001111111011"; -- 0.14719414588674917
	pesos_i(18831) := b"0000000000000000_0000000000000000_0000011101001010_1101010111001110"; -- 0.0284856442159321
	pesos_i(18832) := b"1111111111111111_1111111111111111_1110101100001000_0001001111100001"; -- -0.08190799487044353
	pesos_i(18833) := b"1111111111111111_1111111111111111_1101010101111001_1001011110100010"; -- -0.16611339851332407
	pesos_i(18834) := b"1111111111111111_1111111111111111_1110100001010101_0010110100100100"; -- -0.0924503122586402
	pesos_i(18835) := b"0000000000000000_0000000000000000_0000110010101001_1010010111001110"; -- 0.04946361808647633
	pesos_i(18836) := b"1111111111111111_1111111111111111_1111111110001010_1111111000111101"; -- -0.0017853833535559493
	pesos_i(18837) := b"1111111111111111_1111111111111111_1111011010110110_1100100110110000"; -- -0.03627337883174614
	pesos_i(18838) := b"0000000000000000_0000000000000000_0000111001101010_1011001011110011"; -- 0.05631559786645931
	pesos_i(18839) := b"0000000000000000_0000000000000000_0000110100000100_1010010100110101"; -- 0.050852132272185775
	pesos_i(18840) := b"0000000000000000_0000000000000000_0010000111100101_0111111101010010"; -- 0.13240810163630282
	pesos_i(18841) := b"1111111111111111_1111111111111111_1110010110101100_1111010110001010"; -- -0.10282960309804814
	pesos_i(18842) := b"1111111111111111_1111111111111111_1101110011000100_0100100001000101"; -- -0.1376299697707722
	pesos_i(18843) := b"1111111111111111_1111111111111111_1111110110100101_0000001110011111"; -- -0.009200834043371334
	pesos_i(18844) := b"0000000000000000_0000000000000000_0001110001001100_0110001010100100"; -- 0.11054054729345779
	pesos_i(18845) := b"1111111111111111_1111111111111111_1110001000110001_1101101010101000"; -- -0.11642678637682462
	pesos_i(18846) := b"1111111111111111_1111111111111111_1111101100100111_1001001100111001"; -- -0.01892738204160568
	pesos_i(18847) := b"1111111111111111_1111111111111111_1101111100011001_1101001111110110"; -- -0.12851214646872933
	pesos_i(18848) := b"1111111111111111_1111111111111111_1110100111101011_1001000001101001"; -- -0.08624932700456135
	pesos_i(18849) := b"1111111111111111_1111111111111111_1101011111100010_1001011011100100"; -- -0.15669876994612625
	pesos_i(18850) := b"1111111111111111_1111111111111111_1111111000001101_0011001101110011"; -- -0.007611069017695454
	pesos_i(18851) := b"0000000000000000_0000000000000000_0000010100000000_1101101011110101"; -- 0.019544300931249856
	pesos_i(18852) := b"0000000000000000_0000000000000000_0000001000010001_0101010000001011"; -- 0.008076908781140394
	pesos_i(18853) := b"0000000000000000_0000000000000000_0000110001111000_0111000000110001"; -- 0.04871274170410467
	pesos_i(18854) := b"0000000000000000_0000000000000000_0001011000001001_0001000110101101"; -- 0.08607588257628321
	pesos_i(18855) := b"1111111111111111_1111111111111111_1110110100101010_1101100110111110"; -- -0.07356490231867956
	pesos_i(18856) := b"1111111111111111_1111111111111111_1111111001111101_0010001010000001"; -- -0.005903094799476105
	pesos_i(18857) := b"0000000000000000_0000000000000000_0000011010010100_0011111001110100"; -- 0.025699523191496224
	pesos_i(18858) := b"1111111111111111_1111111111111111_1111010001001001_0100000101001000"; -- -0.045757217343767684
	pesos_i(18859) := b"0000000000000000_0000000000000000_0000110101000011_1101110011110111"; -- 0.0518167593243287
	pesos_i(18860) := b"0000000000000000_0000000000000000_0001110011110011_0111000001010000"; -- 0.11308958004397836
	pesos_i(18861) := b"0000000000000000_0000000000000000_0010010010001011_0110000011111101"; -- 0.14275175264155496
	pesos_i(18862) := b"1111111111111111_1111111111111111_1101110000110000_1111000000011001"; -- -0.1398782672810553
	pesos_i(18863) := b"0000000000000000_0000000000000000_0000010100110010_1011001011001100"; -- 0.020304846575455344
	pesos_i(18864) := b"0000000000000000_0000000000000000_0010010101010000_0011111100010011"; -- 0.14575571256280365
	pesos_i(18865) := b"1111111111111111_1111111111111111_1111011110000100_0111110000001101"; -- -0.03313469575359446
	pesos_i(18866) := b"1111111111111111_1111111111111111_1110101000101110_1111110111100111"; -- -0.08522046200795609
	pesos_i(18867) := b"0000000000000000_0000000000000000_0001101011011110_0110100011000110"; -- 0.10495619618606633
	pesos_i(18868) := b"0000000000000000_0000000000000000_0001010011110011_0000000000110001"; -- 0.08183289716983971
	pesos_i(18869) := b"0000000000000000_0000000000000000_0010101000110011_1111100101110010"; -- 0.16485556632552312
	pesos_i(18870) := b"0000000000000000_0000000000000000_0001000110111000_1000010111110111"; -- 0.06922185222731038
	pesos_i(18871) := b"0000000000000000_0000000000000000_0001110000010100_1100100111100100"; -- 0.10969220941325718
	pesos_i(18872) := b"1111111111111111_1111111111111111_1110101011111000_0110010001011100"; -- -0.08214733831325503
	pesos_i(18873) := b"0000000000000000_0000000000000000_0000001000110011_1001110100000100"; -- 0.008600057076934816
	pesos_i(18874) := b"0000000000000000_0000000000000000_0001110000101110_1101001011010101"; -- 0.11008947083399125
	pesos_i(18875) := b"1111111111111111_1111111111111111_1111001101001000_1011111101011111"; -- -0.049671210676952
	pesos_i(18876) := b"1111111111111111_1111111111111111_1110010000001101_0001010111011111"; -- -0.109175332209364
	pesos_i(18877) := b"1111111111111111_1111111111111111_1110101000100100_1110100101010100"; -- -0.08537427607614138
	pesos_i(18878) := b"1111111111111111_1111111111111111_1110111000010001_1100011101011110"; -- -0.07004121728373412
	pesos_i(18879) := b"0000000000000000_0000000000000000_0000001111001011_1111111001010111"; -- 0.014831443965420571
	pesos_i(18880) := b"0000000000000000_0000000000000000_0000011000101001_1101010100110101"; -- 0.024075818480160233
	pesos_i(18881) := b"0000000000000000_0000000000000000_0000100100001110_1001111000100110"; -- 0.03537929952499426
	pesos_i(18882) := b"1111111111111111_1111111111111111_1110100111010011_0111100110011000"; -- -0.08661689794109668
	pesos_i(18883) := b"1111111111111111_1111111111111111_1110000011000111_1000100000100001"; -- -0.12195538699942193
	pesos_i(18884) := b"1111111111111111_1111111111111111_1111010100000011_1111010101001000"; -- -0.042908353758812676
	pesos_i(18885) := b"0000000000000000_0000000000000000_0000000111000011_0110100101010001"; -- 0.006887991218040125
	pesos_i(18886) := b"1111111111111111_1111111111111111_1111101101100000_1000010101100001"; -- -0.018058456227623504
	pesos_i(18887) := b"1111111111111111_1111111111111111_1111111111110100_0010110100000000"; -- -0.00018042334906107467
	pesos_i(18888) := b"0000000000000000_0000000000000000_0001001011000110_1101101010100011"; -- 0.07334677195696349
	pesos_i(18889) := b"1111111111111111_1111111111111111_1110100001001100_1010000110100000"; -- -0.09258069833646256
	pesos_i(18890) := b"1111111111111111_1111111111111111_1110100010000001_0111011000111101"; -- -0.09177456861683703
	pesos_i(18891) := b"1111111111111111_1111111111111111_1101111000001100_0010010011001101"; -- -0.13262720101651035
	pesos_i(18892) := b"1111111111111111_1111111111111111_1110101110110110_0001100001111110"; -- -0.07925269057613774
	pesos_i(18893) := b"0000000000000000_0000000000000000_0010000100000001_1000101001011111"; -- 0.128929756454206
	pesos_i(18894) := b"0000000000000000_0000000000000000_0000110111101011_0101010111000100"; -- 0.054372177347093424
	pesos_i(18895) := b"1111111111111111_1111111111111111_1110011101100110_0000010001100001"; -- -0.09609959255001678
	pesos_i(18896) := b"1111111111111111_1111111111111111_1101011010101011_0100001101001010"; -- -0.16144923644007853
	pesos_i(18897) := b"1111111111111111_1111111111111111_1110110110011101_1010001011111000"; -- -0.07181340644160514
	pesos_i(18898) := b"1111111111111111_1111111111111111_1111110000011000_0110011101111101"; -- -0.015252620619153237
	pesos_i(18899) := b"0000000000000000_0000000000000000_0000101010011011_0000010110100110"; -- 0.041427949010540935
	pesos_i(18900) := b"0000000000000000_0000000000000000_0000100000001110_0111011100100001"; -- 0.03147072365190217
	pesos_i(18901) := b"1111111111111111_1111111111111111_1111000100000110_1100111010001001"; -- -0.05848988680279829
	pesos_i(18902) := b"0000000000000000_0000000000000000_0010000011111101_0101110000011000"; -- 0.12886596290881525
	pesos_i(18903) := b"1111111111111111_1111111111111111_1101111110101110_1010101011100110"; -- -0.126241034401027
	pesos_i(18904) := b"1111111111111111_1111111111111111_1110110011101100_0101001001111000"; -- -0.07451901026432643
	pesos_i(18905) := b"1111111111111111_1111111111111111_1110011000100100_1101001000100001"; -- -0.10100065899310866
	pesos_i(18906) := b"1111111111111111_1111111111111111_1101010011101000_1010011001001010"; -- -0.16832504933091497
	pesos_i(18907) := b"0000000000000000_0000000000000000_0001100000011001_0111010111011110"; -- 0.09413849524969951
	pesos_i(18908) := b"1111111111111111_1111111111111111_1111011110111001_1110101010110011"; -- -0.03231938477920443
	pesos_i(18909) := b"0000000000000000_0000000000000000_0010000110001100_0100101011011010"; -- 0.13104694192188213
	pesos_i(18910) := b"1111111111111111_1111111111111111_1111000011000110_1110000101110110"; -- -0.05946532120725988
	pesos_i(18911) := b"0000000000000000_0000000000000000_0000110010010000_0011000001100010"; -- 0.04907514947610872
	pesos_i(18912) := b"0000000000000000_0000000000000000_0000010101011010_0110010100111010"; -- 0.020910574633125775
	pesos_i(18913) := b"1111111111111111_1111111111111111_1111011110111111_0001001101110101"; -- -0.032240661465030025
	pesos_i(18914) := b"1111111111111111_1111111111111111_1110010001101001_1101111111110110"; -- -0.10775947793401743
	pesos_i(18915) := b"0000000000000000_0000000000000000_0000101101010000_0000001101010111"; -- 0.04418965223716902
	pesos_i(18916) := b"0000000000000000_0000000000000000_0001100011110011_1110101100110001"; -- 0.09747190431671278
	pesos_i(18917) := b"0000000000000000_0000000000000000_0010001011011100_0101010001011100"; -- 0.1361744618400428
	pesos_i(18918) := b"0000000000000000_0000000000000000_0000000101001010_0000010100111010"; -- 0.005035711978232039
	pesos_i(18919) := b"1111111111111111_1111111111111111_1110011010100101_1001101001111101"; -- -0.09903559153407682
	pesos_i(18920) := b"0000000000000000_0000000000000000_0001011000001110_0100100110101100"; -- 0.08615551412066369
	pesos_i(18921) := b"1111111111111111_1111111111111111_1111001110001111_0000010100101101"; -- -0.04859893457470923
	pesos_i(18922) := b"1111111111111111_1111111111111111_1110101101110010_1010111001111101"; -- -0.08028134769472371
	pesos_i(18923) := b"0000000000000000_0000000000000000_0010010001011100_1001111011001111"; -- 0.14203827423393384
	pesos_i(18924) := b"1111111111111111_1111111111111111_1111001000010111_1111100111100000"; -- -0.054321654199769545
	pesos_i(18925) := b"0000000000000000_0000000000000000_0000000111100011_0010001101000001"; -- 0.007372096355986154
	pesos_i(18926) := b"0000000000000000_0000000000000000_0001101111101001_1101110111101010"; -- 0.10903727503533191
	pesos_i(18927) := b"0000000000000000_0000000000000000_0000110001010000_1010000111000010"; -- 0.04810534471606429
	pesos_i(18928) := b"0000000000000000_0000000000000000_0000100111101111_1000001001010111"; -- 0.03881086956048975
	pesos_i(18929) := b"1111111111111111_1111111111111111_1111100000010110_1010101111101001"; -- -0.03090406010171315
	pesos_i(18930) := b"0000000000000000_0000000000000000_0010100000100011_1110010001101001"; -- 0.1567976718170889
	pesos_i(18931) := b"1111111111111111_1111111111111111_1110011101110110_0110000110101001"; -- -0.0958498919959239
	pesos_i(18932) := b"0000000000000000_0000000000000000_0001001011001000_1010001100000001"; -- 0.07337397364620098
	pesos_i(18933) := b"0000000000000000_0000000000000000_0001001001011011_0010010111010110"; -- 0.0717033049034711
	pesos_i(18934) := b"0000000000000000_0000000000000000_0001110001011001_0101111101011000"; -- 0.11073871514978995
	pesos_i(18935) := b"0000000000000000_0000000000000000_0001110110100001_1111110110100100"; -- 0.11575303310217387
	pesos_i(18936) := b"1111111111111111_1111111111111111_1111010011100111_0100111000000101"; -- -0.04334556941507549
	pesos_i(18937) := b"1111111111111111_1111111111111111_1111000011110101_0101101011000101"; -- -0.05875618632099325
	pesos_i(18938) := b"1111111111111111_1111111111111111_1110100110010110_1011011011001101"; -- -0.08754403585167177
	pesos_i(18939) := b"0000000000000000_0000000000000000_0000101101001010_1010001110110011"; -- 0.04410765755679168
	pesos_i(18940) := b"1111111111111111_1111111111111111_1110001000111111_0001100000001000"; -- -0.116224763824842
	pesos_i(18941) := b"1111111111111111_1111111111111111_1111011000001011_1001000111001010"; -- -0.03888596368405848
	pesos_i(18942) := b"1111111111111111_1111111111111111_1110010111111011_1100011010111000"; -- -0.10162694949127209
	pesos_i(18943) := b"1111111111111111_1111111111111111_1110010010111010_0101010100011010"; -- -0.10653179275929807
	pesos_i(18944) := b"1111111111111111_1111111111111111_1110001101100101_0100010001010011"; -- -0.1117360399640837
	pesos_i(18945) := b"1111111111111111_1111111111111111_1111010011100011_1110100000000101"; -- -0.04339742540086265
	pesos_i(18946) := b"1111111111111111_1111111111111111_1110010001110011_0000101011010001"; -- -0.10761959457755622
	pesos_i(18947) := b"0000000000000000_0000000000000000_0000111010100100_1000010100010001"; -- 0.057197872772373946
	pesos_i(18948) := b"1111111111111111_1111111111111111_1101111011101110_1010111000100111"; -- -0.12917052802328116
	pesos_i(18949) := b"0000000000000000_0000000000000000_0001101001001000_0010110000001001"; -- 0.10266375759885706
	pesos_i(18950) := b"0000000000000000_0000000000000000_0010000011111101_1100001100101010"; -- 0.12887210643175206
	pesos_i(18951) := b"0000000000000000_0000000000000000_0000011001101111_1100011010010110"; -- 0.02514306212433918
	pesos_i(18952) := b"1111111111111111_1111111111111111_1101111111010000_0010001100000011"; -- -0.1257303349058013
	pesos_i(18953) := b"1111111111111111_1111111111111111_1101101011001101_0001011111101011"; -- -0.14530802255130956
	pesos_i(18954) := b"1111111111111111_1111111111111111_1111000011110011_1101011111111001"; -- -0.05877924123212805
	pesos_i(18955) := b"1111111111111111_1111111111111111_1111001001000110_1011011011011100"; -- -0.05360848545961571
	pesos_i(18956) := b"0000000000000000_0000000000000000_0000111001101001_0101100011010110"; -- 0.05629496796910307
	pesos_i(18957) := b"0000000000000000_0000000000000000_0000001001110100_0100010100010100"; -- 0.009586636801781658
	pesos_i(18958) := b"0000000000000000_0000000000000000_0001110001011101_0000110111101011"; -- 0.1107948969129259
	pesos_i(18959) := b"1111111111111111_1111111111111111_1101100000101011_0110000010011010"; -- -0.1555881142242738
	pesos_i(18960) := b"1111111111111111_1111111111111111_1110001010100111_0110011100110000"; -- -0.1146331317537112
	pesos_i(18961) := b"1111111111111111_1111111111111111_1111111101001111_0100000000111101"; -- -0.002696976715242974
	pesos_i(18962) := b"1111111111111111_1111111111111111_1111000001000001_1001101100110110"; -- -0.06149892738029989
	pesos_i(18963) := b"0000000000000000_0000000000000000_0001001100101001_0010011010101111"; -- 0.07484666602210191
	pesos_i(18964) := b"0000000000000000_0000000000000000_0000101111001110_0000101010000100"; -- 0.04611268723580918
	pesos_i(18965) := b"1111111111111111_1111111111111111_1101111100100001_0101010111101100"; -- -0.12839758870840884
	pesos_i(18966) := b"0000000000000000_0000000000000000_0000011010011101_1101000010110011"; -- 0.02584556927591715
	pesos_i(18967) := b"0000000000000000_0000000000000000_0001111010101111_1000110010110010"; -- 0.11986617427784368
	pesos_i(18968) := b"1111111111111111_1111111111111111_1111110100010100_1001000000100110"; -- -0.011404982267089704
	pesos_i(18969) := b"1111111111111111_1111111111111111_1101110110101000_1001110000010010"; -- -0.13414597086957175
	pesos_i(18970) := b"1111111111111111_1111111111111111_1101100100000101_1001110100001100"; -- -0.15225809535934026
	pesos_i(18971) := b"1111111111111111_1111111111111111_1111100010010011_1000101100101010"; -- -0.028998663130457084
	pesos_i(18972) := b"0000000000000000_0000000000000000_0001100000110101_0010101011111111"; -- 0.09456127854061144
	pesos_i(18973) := b"0000000000000000_0000000000000000_0010001110110101_1001000111100000"; -- 0.13948928567892172
	pesos_i(18974) := b"0000000000000000_0000000000000000_0001111110001110_0001010111111101"; -- 0.1232618086532659
	pesos_i(18975) := b"1111111111111111_1111111111111111_1111111110000100_0101010111000001"; -- -0.0018869785293519497
	pesos_i(18976) := b"0000000000000000_0000000000000000_0010100110101110_0101100101101111"; -- 0.16281660989963215
	pesos_i(18977) := b"0000000000000000_0000000000000000_0001011101111010_0111111111001101"; -- 0.09171293982603697
	pesos_i(18978) := b"1111111111111111_1111111111111111_1111000010011100_0011101101100110"; -- -0.06011608842620901
	pesos_i(18979) := b"0000000000000000_0000000000000000_0000100011100010_0000011110111010"; -- 0.03469894682938607
	pesos_i(18980) := b"0000000000000000_0000000000000000_0010000100100000_1101010100101011"; -- 0.1294072370989033
	pesos_i(18981) := b"0000000000000000_0000000000000000_0000100100001011_1100011101011000"; -- 0.03533597847127364
	pesos_i(18982) := b"0000000000000000_0000000000000000_0000010100101010_0100101101011100"; -- 0.02017661090974372
	pesos_i(18983) := b"0000000000000000_0000000000000000_0001011011000001_1101101010000010"; -- 0.0888954702780862
	pesos_i(18984) := b"0000000000000000_0000000000000000_0001101100001100_0010010001000000"; -- 0.10565401619297249
	pesos_i(18985) := b"0000000000000000_0000000000000000_0001011111010110_0101101100111011"; -- 0.09311456866743677
	pesos_i(18986) := b"1111111111111111_1111111111111111_1111011001110100_1010010101101011"; -- -0.03728262083475757
	pesos_i(18987) := b"1111111111111111_1111111111111111_1111101010011001_1101110011011111"; -- -0.02108974040620202
	pesos_i(18988) := b"0000000000000000_0000000000000000_0001110000110100_1100010110101000"; -- 0.11018023827724664
	pesos_i(18989) := b"0000000000000000_0000000000000000_0000100101000000_1001010001001100"; -- 0.036141651611920914
	pesos_i(18990) := b"1111111111111111_1111111111111111_1110101010100001_1001111101101001"; -- -0.08347133342877741
	pesos_i(18991) := b"0000000000000000_0000000000000000_0001101010000001_1000110001001110"; -- 0.10353924671027412
	pesos_i(18992) := b"0000000000000000_0000000000000000_0010010010001100_1011100101001100"; -- 0.14277227504218976
	pesos_i(18993) := b"1111111111111111_1111111111111111_1111100010100111_0010011110011100"; -- -0.028699421369034726
	pesos_i(18994) := b"1111111111111111_1111111111111111_1111011111001111_0100111100110010"; -- -0.031992960215603695
	pesos_i(18995) := b"1111111111111111_1111111111111111_1110000010011000_1111101010100110"; -- -0.12266572420601309
	pesos_i(18996) := b"1111111111111111_1111111111111111_1101111000100000_0001101000001000"; -- -0.13232266713208413
	pesos_i(18997) := b"0000000000000000_0000000000000000_0010001110100110_1011000010011001"; -- 0.1392622351325532
	pesos_i(18998) := b"1111111111111111_1111111111111111_1111000001010111_1110010110111011"; -- -0.06115879240761014
	pesos_i(18999) := b"1111111111111111_1111111111111111_1110100100010011_0110001111101101"; -- -0.08954787704244167
	pesos_i(19000) := b"1111111111111111_1111111111111111_1111010001111110_1011101110011110"; -- -0.04494120968896157
	pesos_i(19001) := b"0000000000000000_0000000000000000_0001101001001010_0000001010101000"; -- 0.10269180875623388
	pesos_i(19002) := b"1111111111111111_1111111111111111_1110010111011111_0010100100110000"; -- -0.10206358499387902
	pesos_i(19003) := b"0000000000000000_0000000000000000_0000101010110000_0000011101010011"; -- 0.04174848344883743
	pesos_i(19004) := b"1111111111111111_1111111111111111_1110101101011111_1010110000111100"; -- -0.08057139896789592
	pesos_i(19005) := b"1111111111111111_1111111111111111_1101111010010101_1000100100101011"; -- -0.13053076450588325
	pesos_i(19006) := b"1111111111111111_1111111111111111_1101011111000101_1010100001101100"; -- -0.15714022983508846
	pesos_i(19007) := b"0000000000000000_0000000000000000_0010010010001101_1000100100100001"; -- 0.14278466275791116
	pesos_i(19008) := b"1111111111111111_1111111111111111_1110110111011110_0111011101111101"; -- -0.07082417685947263
	pesos_i(19009) := b"0000000000000000_0000000000000000_0001110011010001_1011111110011000"; -- 0.1125755068365617
	pesos_i(19010) := b"1111111111111111_1111111111111111_1101101100111101_0010001111111010"; -- -0.14359831958672417
	pesos_i(19011) := b"0000000000000000_0000000000000000_0001111010101010_0110111011110010"; -- 0.11978810701992414
	pesos_i(19012) := b"0000000000000000_0000000000000000_0000000001011001_1011111001110100"; -- 0.0013693841662793256
	pesos_i(19013) := b"1111111111111111_1111111111111111_1110001110100101_1011011111010010"; -- -0.1107525931640867
	pesos_i(19014) := b"0000000000000000_0000000000000000_0010000100100111_1100010010000101"; -- 0.1295130561667293
	pesos_i(19015) := b"0000000000000000_0000000000000000_0000110000101101_0000011011111111"; -- 0.04756206247381663
	pesos_i(19016) := b"0000000000000000_0000000000000000_0001100111000100_1101011011111111"; -- 0.10065978749062336
	pesos_i(19017) := b"0000000000000000_0000000000000000_0001001101001101_0100010011010110"; -- 0.07539777966611638
	pesos_i(19018) := b"0000000000000000_0000000000000000_0000101011101011_1000011010100111"; -- 0.04265634144408293
	pesos_i(19019) := b"1111111111111111_1111111111111111_1101111100000111_1101011101000111"; -- -0.12878660688084465
	pesos_i(19020) := b"0000000000000000_0000000000000000_0000110100011001_0110110001011110"; -- 0.05116917902536401
	pesos_i(19021) := b"1111111111111111_1111111111111111_1101111011100011_1101100001101010"; -- -0.12933585569981879
	pesos_i(19022) := b"1111111111111111_1111111111111111_1111010111100100_0100001110001101"; -- -0.03948571973282612
	pesos_i(19023) := b"1111111111111111_1111111111111111_1111001111011101_0011101010100101"; -- -0.04740556210566649
	pesos_i(19024) := b"0000000000000000_0000000000000000_0000101100000101_0110100000000100"; -- 0.0430512436849204
	pesos_i(19025) := b"1111111111111111_1111111111111111_1110100110110100_1000011001101100"; -- -0.08708915578207517
	pesos_i(19026) := b"1111111111111111_1111111111111111_1110010011000111_1001010001100011"; -- -0.10632965637000412
	pesos_i(19027) := b"0000000000000000_0000000000000000_0001100000111111_1110010101011100"; -- 0.09472497448001667
	pesos_i(19028) := b"1111111111111111_1111111111111111_1110011110100101_1000100111100110"; -- -0.09513033030593214
	pesos_i(19029) := b"0000000000000000_0000000000000000_0000010010110101_0100010010110001"; -- 0.018390935222327674
	pesos_i(19030) := b"0000000000000000_0000000000000000_0001101011111111_1011110110111110"; -- 0.10546480066818537
	pesos_i(19031) := b"1111111111111111_1111111111111111_1110110001001101_0000100111010000"; -- -0.07694948843256122
	pesos_i(19032) := b"0000000000000000_0000000000000000_0001100001110001_0111100010001010"; -- 0.09548142790540394
	pesos_i(19033) := b"0000000000000000_0000000000000000_0001110010110101_1010100101100110"; -- 0.11214693784518809
	pesos_i(19034) := b"0000000000000000_0000000000000000_0000011101010100_0110010000110000"; -- 0.028631460013552757
	pesos_i(19035) := b"1111111111111111_1111111111111111_1110110101010001_0110100000111110"; -- -0.07297657469916988
	pesos_i(19036) := b"0000000000000000_0000000000000000_0001000100100000_0000010100001001"; -- 0.06689483125929341
	pesos_i(19037) := b"0000000000000000_0000000000000000_0001011110001011_1100011100000000"; -- 0.09197658308093051
	pesos_i(19038) := b"0000000000000000_0000000000000000_0010001110001010_1000011111010100"; -- 0.13883255898326616
	pesos_i(19039) := b"0000000000000000_0000000000000000_0001110010101111_0001101000010001"; -- 0.11204684176661864
	pesos_i(19040) := b"1111111111111111_1111111111111111_1111111010011111_0011101110111100"; -- -0.0053827921038231055
	pesos_i(19041) := b"1111111111111111_1111111111111111_1111010000000001_0010011011100000"; -- -0.04685742410133881
	pesos_i(19042) := b"0000000000000000_0000000000000000_0001100001110001_0011001111011000"; -- 0.0954773333390738
	pesos_i(19043) := b"0000000000000000_0000000000000000_0001101000101101_1001010100001110"; -- 0.10225802980840239
	pesos_i(19044) := b"0000000000000000_0000000000000000_0010001110011100_0000010111101001"; -- 0.1390994733620495
	pesos_i(19045) := b"0000000000000000_0000000000000000_0001011100010000_1001000011001010"; -- 0.09009652067839345
	pesos_i(19046) := b"0000000000000000_0000000000000000_0001111011010111_1110010010001001"; -- 0.12048176140856526
	pesos_i(19047) := b"0000000000000000_0000000000000000_0010000011100100_1100111011011010"; -- 0.12849133315912542
	pesos_i(19048) := b"0000000000000000_0000000000000000_0001000001110101_1001111111110010"; -- 0.06429481185906563
	pesos_i(19049) := b"1111111111111111_1111111111111111_1111010101001100_0011011101011001"; -- -0.04180578310297692
	pesos_i(19050) := b"0000000000000000_0000000000000000_0000100100010111_0001100101111110"; -- 0.03550872154732395
	pesos_i(19051) := b"0000000000000000_0000000000000000_0001010011011111_1011111111010100"; -- 0.0815391437981729
	pesos_i(19052) := b"0000000000000000_0000000000000000_0001101011111001_0110100101010101"; -- 0.10536821666109279
	pesos_i(19053) := b"1111111111111111_1111111111111111_1110101101001001_1011000001100110"; -- -0.08090684418476772
	pesos_i(19054) := b"1111111111111111_1111111111111111_1110110111101111_0110000000011110"; -- -0.07056617029541624
	pesos_i(19055) := b"0000000000000000_0000000000000000_0001100001001111_1110011001001001"; -- 0.09496917039026642
	pesos_i(19056) := b"0000000000000000_0000000000000000_0001111010111101_1001000100101100"; -- 0.12008006408954684
	pesos_i(19057) := b"0000000000000000_0000000000000000_0010100101100011_1011101111111110"; -- 0.16167807530488335
	pesos_i(19058) := b"1111111111111111_1111111111111111_1111011111111110_1001001101000001"; -- -0.03127174066442976
	pesos_i(19059) := b"1111111111111111_1111111111111111_1101101111110000_0001010001111110"; -- -0.14086791911084645
	pesos_i(19060) := b"0000000000000000_0000000000000000_0000001110001001_1100000001001100"; -- 0.013820665884613767
	pesos_i(19061) := b"0000000000000000_0000000000000000_0000111011101000_0111100111000010"; -- 0.05823479631153501
	pesos_i(19062) := b"0000000000000000_0000000000000000_0010001110111011_1110110101010111"; -- 0.13958629004217857
	pesos_i(19063) := b"1111111111111111_1111111111111111_1111111011110110_0001111010110000"; -- -0.004057008761838308
	pesos_i(19064) := b"1111111111111111_1111111111111111_1110000100000100_0110110010100111"; -- -0.12102623858692485
	pesos_i(19065) := b"1111111111111111_1111111111111111_1110001111111001_1111101110010011"; -- -0.10946681657029687
	pesos_i(19066) := b"1111111111111111_1111111111111111_1110101000101110_0101101000000000"; -- -0.08523023137753301
	pesos_i(19067) := b"0000000000000000_0000000000000000_0001000011110100_0100111011110110"; -- 0.06622785103046928
	pesos_i(19068) := b"0000000000000000_0000000000000000_0001101110001011_0000100111111111"; -- 0.10759031758820287
	pesos_i(19069) := b"0000000000000000_0000000000000000_0000001000010111_1001100000100011"; -- 0.008172520165306042
	pesos_i(19070) := b"1111111111111111_1111111111111111_1111010010010001_1110111100111100"; -- -0.04464821607679171
	pesos_i(19071) := b"0000000000000000_0000000000000000_0010001100101011_0010000100100100"; -- 0.1373768533692579
	pesos_i(19072) := b"0000000000000000_0000000000000000_0000011100111000_1100010001010111"; -- 0.028209945063663568
	pesos_i(19073) := b"0000000000000000_0000000000000000_0001011011000111_0001001111100000"; -- 0.08897518372548781
	pesos_i(19074) := b"1111111111111111_1111111111111111_1111001001110101_0010010000000001"; -- -0.052900075580816996
	pesos_i(19075) := b"0000000000000000_0000000000000000_0001000010001000_0011000111011000"; -- 0.06457816617514778
	pesos_i(19076) := b"1111111111111111_1111111111111111_1111111101000010_1101001011110011"; -- -0.002886596363340627
	pesos_i(19077) := b"1111111111111111_1111111111111111_1110010111000111_0111100101101001"; -- -0.10242501448003352
	pesos_i(19078) := b"1111111111111111_1111111111111111_1101111010011010_1101001010000000"; -- -0.13045009968637278
	pesos_i(19079) := b"0000000000000000_0000000000000000_0001010100001000_1110000001001011"; -- 0.08216668926558035
	pesos_i(19080) := b"1111111111111111_1111111111111111_1111010111100100_1011101010110011"; -- -0.039478618035208836
	pesos_i(19081) := b"0000000000000000_0000000000000000_0000001001101110_1010101111100001"; -- 0.009501211664058585
	pesos_i(19082) := b"0000000000000000_0000000000000000_0000101100011100_1000111110101101"; -- 0.04340455990455489
	pesos_i(19083) := b"0000000000000000_0000000000000000_0010011010000110_1011101011001000"; -- 0.15049331071326333
	pesos_i(19084) := b"0000000000000000_0000000000000000_0010000101010011_1110010111111011"; -- 0.1301864373759242
	pesos_i(19085) := b"1111111111111111_1111111111111111_1110101010011001_0001101111110010"; -- -0.08360123963069635
	pesos_i(19086) := b"0000000000000000_0000000000000000_0001110001111101_1111001010100110"; -- 0.11129681150239346
	pesos_i(19087) := b"0000000000000000_0000000000000000_0000111111000010_0100111111111100"; -- 0.061558722538226716
	pesos_i(19088) := b"0000000000000000_0000000000000000_0010000011000101_1011100001000111"; -- 0.1280169651969639
	pesos_i(19089) := b"1111111111111111_1111111111111111_1110111100011101_1110100010010101"; -- -0.06594988215094198
	pesos_i(19090) := b"0000000000000000_0000000000000000_0000011010101100_1101000000111110"; -- 0.02607442390938673
	pesos_i(19091) := b"1111111111111111_1111111111111111_1101100111011001_1011010001001001"; -- -0.1490218468634272
	pesos_i(19092) := b"0000000000000000_0000000000000000_0000001001010101_0011001000000110"; -- 0.009112478769998775
	pesos_i(19093) := b"0000000000000000_0000000000000000_0001111010110000_0000110011101000"; -- 0.11987381611411305
	pesos_i(19094) := b"1111111111111111_1111111111111111_1111001010111001_1001110111111001"; -- -0.05185520809839902
	pesos_i(19095) := b"0000000000000000_0000000000000000_0010011111010001_1111100011001111"; -- 0.15554766713749002
	pesos_i(19096) := b"1111111111111111_1111111111111111_1110110000010100_1011111001110100"; -- -0.07780847224473322
	pesos_i(19097) := b"0000000000000000_0000000000000000_0000000100000001_0001101000010001"; -- 0.003923062556797178
	pesos_i(19098) := b"0000000000000000_0000000000000000_0001001010010111_0010110001111111"; -- 0.07261922926878119
	pesos_i(19099) := b"1111111111111111_1111111111111111_1101101110111000_0011101011101111"; -- -0.14172012014619673
	pesos_i(19100) := b"1111111111111111_1111111111111111_1110010110010010_0110101000011111"; -- -0.10323464159091301
	pesos_i(19101) := b"0000000000000000_0000000000000000_0001100001010001_1101101011010000"; -- 0.09499900411581287
	pesos_i(19102) := b"1111111111111111_1111111111111111_1110010010001001_0001011110011100"; -- -0.10728313867390296
	pesos_i(19103) := b"0000000000000000_0000000000000000_0000011001000101_1011101001010011"; -- 0.024501462275991995
	pesos_i(19104) := b"0000000000000000_0000000000000000_0001001000101101_0101100111110010"; -- 0.07100450661326074
	pesos_i(19105) := b"1111111111111111_1111111111111111_1111010011001111_1110010011011101"; -- -0.043702789242783785
	pesos_i(19106) := b"1111111111111111_1111111111111111_1110011000101011_1001111000001100"; -- -0.10089695166323243
	pesos_i(19107) := b"1111111111111111_1111111111111111_1111001110111110_0110011010100000"; -- -0.04787596325128281
	pesos_i(19108) := b"1111111111111111_1111111111111111_1110011100110000_0011000110110010"; -- -0.0969208660645631
	pesos_i(19109) := b"0000000000000000_0000000000000000_0000100011101000_1101111001011001"; -- 0.03480329190859209
	pesos_i(19110) := b"0000000000000000_0000000000000000_0001101000101101_0010000010110000"; -- 0.10225109385132682
	pesos_i(19111) := b"0000000000000000_0000000000000000_0001100101000101_0111000101111000"; -- 0.09871586981111577
	pesos_i(19112) := b"1111111111111111_1111111111111111_1111011010000001_1001100101000101"; -- -0.037084980647492154
	pesos_i(19113) := b"1111111111111111_1111111111111111_1111110100101000_0011000000000110"; -- -0.01110553609953818
	pesos_i(19114) := b"1111111111111111_1111111111111111_1111011111110111_0101000000001011"; -- -0.031382558216590535
	pesos_i(19115) := b"0000000000000000_0000000000000000_0001111111111110_1100100000001110"; -- 0.12498140662348003
	pesos_i(19116) := b"1111111111111111_1111111111111111_1111111010010100_0001000110101001"; -- -0.005553146692771674
	pesos_i(19117) := b"0000000000000000_0000000000000000_0000001011101011_1101101001001000"; -- 0.011411325994440889
	pesos_i(19118) := b"1111111111111111_1111111111111111_1101110011101000_1000000110001000"; -- -0.13707724029273324
	pesos_i(19119) := b"1111111111111111_1111111111111111_1110001010101011_1111001100100100"; -- -0.11456375486876579
	pesos_i(19120) := b"1111111111111111_1111111111111111_1111110001101100_1011111101101000"; -- -0.013965642168460144
	pesos_i(19121) := b"0000000000000000_0000000000000000_0000001001111110_1001110100111101"; -- 0.009744479523034769
	pesos_i(19122) := b"1111111111111111_1111111111111111_1101111000010111_0110011010111001"; -- -0.13245542514832637
	pesos_i(19123) := b"1111111111111111_1111111111111111_1111100101010110_0101111101111001"; -- -0.02602580358521734
	pesos_i(19124) := b"0000000000000000_0000000000000000_0010011001001001_0101110111100110"; -- 0.149556988368492
	pesos_i(19125) := b"0000000000000000_0000000000000000_0001000011100000_1110001110111110"; -- 0.06593154318792632
	pesos_i(19126) := b"0000000000000000_0000000000000000_0000000100001110_0100101001111001"; -- 0.004124312004427952
	pesos_i(19127) := b"1111111111111111_1111111111111111_1101110100111111_0100010001110100"; -- -0.1357533661948056
	pesos_i(19128) := b"1111111111111111_1111111111111111_1111101000110111_0011111011100101"; -- -0.02259451774618633
	pesos_i(19129) := b"1111111111111111_1111111111111111_1111110011100011_1001011101011011"; -- -0.012152233397282563
	pesos_i(19130) := b"0000000000000000_0000000000000000_0001101001000011_0101100101100000"; -- 0.10259016606439016
	pesos_i(19131) := b"0000000000000000_0000000000000000_0000011101101001_1000111000000000"; -- 0.028954386632706993
	pesos_i(19132) := b"0000000000000000_0000000000000000_0001100100100010_1011010011010101"; -- 0.09818582724604523
	pesos_i(19133) := b"0000000000000000_0000000000000000_0001000110000001_0110110010100100"; -- 0.06838110925124441
	pesos_i(19134) := b"0000000000000000_0000000000000000_0001111110110101_1010000001110000"; -- 0.12386515373386496
	pesos_i(19135) := b"1111111111111111_1111111111111111_1111011101101101_1110011011101110"; -- -0.03347927761473703
	pesos_i(19136) := b"0000000000000000_0000000000000000_0010011000110011_0110100111011101"; -- 0.14922200811206687
	pesos_i(19137) := b"1111111111111111_1111111111111111_1101101100010001_1001001011100010"; -- -0.14426309560751222
	pesos_i(19138) := b"1111111111111111_1111111111111111_1111101111101011_0110101010011001"; -- -0.015939080935001643
	pesos_i(19139) := b"1111111111111111_1111111111111111_1111011001111001_1110000001110010"; -- -0.03720280848434469
	pesos_i(19140) := b"1111111111111111_1111111111111111_1110010110001011_1011010000010111"; -- -0.10333704422738961
	pesos_i(19141) := b"0000000000000000_0000000000000000_0001000011001010_1100111000111111"; -- 0.0655945686543387
	pesos_i(19142) := b"1111111111111111_1111111111111111_1110011011000101_1001011000111100"; -- -0.09854756382092233
	pesos_i(19143) := b"0000000000000000_0000000000000000_0001000100101000_0110110011000110"; -- 0.06702308492523544
	pesos_i(19144) := b"0000000000000000_0000000000000000_0001000010100000_0011100111000110"; -- 0.06494484973523745
	pesos_i(19145) := b"0000000000000000_0000000000000000_0010000000000101_1100001101111000"; -- 0.12508794475809148
	pesos_i(19146) := b"1111111111111111_1111111111111111_1101110111101011_1100101100010001"; -- -0.13312083084406182
	pesos_i(19147) := b"1111111111111111_1111111111111111_1110001111010010_0000101010111101"; -- -0.11007626432008434
	pesos_i(19148) := b"0000000000000000_0000000000000000_0001110101110010_1111101101101000"; -- 0.11503573692563974
	pesos_i(19149) := b"0000000000000000_0000000000000000_0010010011100110_0010110111111000"; -- 0.1441372613957569
	pesos_i(19150) := b"1111111111111111_1111111111111111_1110110100110110_0001111010010111"; -- -0.0733929522010748
	pesos_i(19151) := b"0000000000000000_0000000000000000_0010010011011011_1100000001101011"; -- 0.143978143693045
	pesos_i(19152) := b"0000000000000000_0000000000000000_0010100001001101_1011111111110101"; -- 0.15743636831599772
	pesos_i(19153) := b"1111111111111111_1111111111111111_1111001010011000_1001100110001011"; -- -0.05235901214882646
	pesos_i(19154) := b"0000000000000000_0000000000000000_0010000111111111_0010000111011011"; -- 0.13279925905183823
	pesos_i(19155) := b"1111111111111111_1111111111111111_1101111101111001_1101010011111111"; -- -0.12704724103202328
	pesos_i(19156) := b"0000000000000000_0000000000000000_0001001000111110_0000101001011110"; -- 0.07125916284743608
	pesos_i(19157) := b"0000000000000000_0000000000000000_0001001001001011_1001000001001110"; -- 0.07146551041069688
	pesos_i(19158) := b"1111111111111111_1111111111111111_1111101000001111_1011100011101110"; -- -0.023197595470778095
	pesos_i(19159) := b"1111111111111111_1111111111111111_1111110011011010_0111010111100001"; -- -0.012291557790182445
	pesos_i(19160) := b"0000000000000000_0000000000000000_0000101011010100_0101101010110000"; -- 0.04230276858717712
	pesos_i(19161) := b"0000000000000000_0000000000000000_0000110110110100_1000101101100010"; -- 0.053536139870688504
	pesos_i(19162) := b"1111111111111111_1111111111111111_1110000010110110_0100010000110111"; -- -0.1222188345737565
	pesos_i(19163) := b"1111111111111111_1111111111111111_1111100100101000_0010111110011001"; -- -0.0267305614540589
	pesos_i(19164) := b"0000000000000000_0000000000000000_0001101010110000_0001000110110110"; -- 0.10424910242292498
	pesos_i(19165) := b"0000000000000000_0000000000000000_0000001011000011_0000110001100110"; -- 0.010788702959396067
	pesos_i(19166) := b"0000000000000000_0000000000000000_0001101110000110_1101010111101011"; -- 0.10752617814626626
	pesos_i(19167) := b"0000000000000000_0000000000000000_0010100000101010_1000111111000010"; -- 0.15689943778523635
	pesos_i(19168) := b"0000000000000000_0000000000000000_0010010100110000_1011010101010101"; -- 0.14527448013223876
	pesos_i(19169) := b"1111111111111111_1111111111111111_1110100101001001_1111000011011101"; -- -0.08871550190369046
	pesos_i(19170) := b"1111111111111111_1111111111111111_1111100100000010_0110111001011100"; -- -0.027306654486658317
	pesos_i(19171) := b"0000000000000000_0000000000000000_0000000001111001_1110011001010001"; -- 0.0018600413155028975
	pesos_i(19172) := b"0000000000000000_0000000000000000_0001111001001111_1000001000100100"; -- 0.11840070131701118
	pesos_i(19173) := b"1111111111111111_1111111111111111_1110110010111001_0000000011100100"; -- -0.07530207083233693
	pesos_i(19174) := b"1111111111111111_1111111111111111_1111110100110001_0010111010111000"; -- -0.010968284745432887
	pesos_i(19175) := b"1111111111111111_1111111111111111_1110011011011110_1101001111101101"; -- -0.0981624170572653
	pesos_i(19176) := b"0000000000000000_0000000000000000_0000101111000001_1111110000010011"; -- 0.045928721181239994
	pesos_i(19177) := b"0000000000000000_0000000000000000_0000010100100100_0000100101100001"; -- 0.020081125415651508
	pesos_i(19178) := b"1111111111111111_1111111111111111_1111010001111110_0010101001011001"; -- -0.044949868541966316
	pesos_i(19179) := b"1111111111111111_1111111111111111_1110011010101110_1101010101110010"; -- -0.09889474825690833
	pesos_i(19180) := b"1111111111111111_1111111111111111_1110001110010111_1111000011110011"; -- -0.11096281116423216
	pesos_i(19181) := b"0000000000000000_0000000000000000_0001101111101000_0111001101100101"; -- 0.10901566703867586
	pesos_i(19182) := b"1111111111111111_1111111111111111_1111010100001001_1001000110001111"; -- -0.04282274489588677
	pesos_i(19183) := b"1111111111111111_1111111111111111_1110000100011111_0100100001011011"; -- -0.12061641491699057
	pesos_i(19184) := b"0000000000000000_0000000000000000_0001100100101011_0101011010000101"; -- 0.09831753491836734
	pesos_i(19185) := b"1111111111111111_1111111111111111_1111001111001001_0100010001110100"; -- -0.04771015331189088
	pesos_i(19186) := b"1111111111111111_1111111111111111_1111010011111110_0001101010100010"; -- -0.04299768021155646
	pesos_i(19187) := b"1111111111111111_1111111111111111_1101101000110001_1001010010001011"; -- -0.14768096546875406
	pesos_i(19188) := b"0000000000000000_0000000000000000_0001100011111010_0111111011010000"; -- 0.09757225598952664
	pesos_i(19189) := b"1111111111111111_1111111111111111_1110100111011011_0001010111111000"; -- -0.08650076584751523
	pesos_i(19190) := b"0000000000000000_0000000000000000_0010001011001001_1101111100000000"; -- 0.13589280833342765
	pesos_i(19191) := b"0000000000000000_0000000000000000_0001000101100101_1000111111011011"; -- 0.06795596213953842
	pesos_i(19192) := b"0000000000000000_0000000000000000_0000010011001010_1011101110011101"; -- 0.018718457940226696
	pesos_i(19193) := b"1111111111111111_1111111111111111_1110001101010000_0101010110000000"; -- -0.11205545070132308
	pesos_i(19194) := b"0000000000000000_0000000000000000_0001101001011111_1101110101001100"; -- 0.10302527520155051
	pesos_i(19195) := b"1111111111111111_1111111111111111_1111110000001110_0011011010100110"; -- -0.015408119704747581
	pesos_i(19196) := b"1111111111111111_1111111111111111_1110100010111110_1110100101011001"; -- -0.0908369213577844
	pesos_i(19197) := b"1111111111111111_1111111111111111_1110010000101010_1010000010100001"; -- -0.10872455665731848
	pesos_i(19198) := b"0000000000000000_0000000000000000_0010100100110101_1101011101010111"; -- 0.1609778010432159
	pesos_i(19199) := b"0000000000000000_0000000000000000_0000100001100111_1011100010100010"; -- 0.032832660293427095
	pesos_i(19200) := b"0000000000000000_0000000000000000_0000110001001000_0011100101011101"; -- 0.04797705190487069
	pesos_i(19201) := b"1111111111111111_1111111111111111_1111100100111011_1110010011011000"; -- -0.026429841271870962
	pesos_i(19202) := b"0000000000000000_0000000000000000_0001110001101110_0001100001100101"; -- 0.11105492079329936
	pesos_i(19203) := b"0000000000000000_0000000000000000_0010001001100001_1010001010011110"; -- 0.1343022952040894
	pesos_i(19204) := b"0000000000000000_0000000000000000_0001010001011100_1010001000100110"; -- 0.07953847332865321
	pesos_i(19205) := b"1111111111111111_1111111111111111_1111000011111001_0101010001110001"; -- -0.058695528503463254
	pesos_i(19206) := b"0000000000000000_0000000000000000_0001010111101000_1011100010110000"; -- 0.08558229737733167
	pesos_i(19207) := b"1111111111111111_1111111111111111_1111111111000000_0111011110101110"; -- -0.0009694291051839792
	pesos_i(19208) := b"0000000000000000_0000000000000000_0000010011011011_0001101011000110"; -- 0.01896827066714994
	pesos_i(19209) := b"0000000000000000_0000000000000000_0001000011100101_0101111001111111"; -- 0.0659998950790018
	pesos_i(19210) := b"0000000000000000_0000000000000000_0001000000011001_0000001011100111"; -- 0.06288164268385459
	pesos_i(19211) := b"0000000000000000_0000000000000000_0010001010011000_1101000100100100"; -- 0.13514430162621427
	pesos_i(19212) := b"0000000000000000_0000000000000000_0000100100100011_1001111100000101"; -- 0.0356997860110847
	pesos_i(19213) := b"0000000000000000_0000000000000000_0001111010011100_1010011110100111"; -- 0.11957786404835416
	pesos_i(19214) := b"0000000000000000_0000000000000000_0001100010101010_0101101010111111"; -- 0.09634940307385294
	pesos_i(19215) := b"1111111111111111_1111111111111111_1101101111101011_1010010111010000"; -- -0.14093555139219
	pesos_i(19216) := b"1111111111111111_1111111111111111_1110010011101110_0010111001111111"; -- -0.10574063688101833
	pesos_i(19217) := b"0000000000000000_0000000000000000_0000111110011000_1111001110000100"; -- 0.060927600588867994
	pesos_i(19218) := b"0000000000000000_0000000000000000_0000011111101110_0000111100000111"; -- 0.03097623754024572
	pesos_i(19219) := b"0000000000000000_0000000000000000_0010001000000000_1010010100000111"; -- 0.13282233641706923
	pesos_i(19220) := b"1111111111111111_1111111111111111_1101110110011110_1101011000100011"; -- -0.13429509781599272
	pesos_i(19221) := b"0000000000000000_0000000000000000_0000001000100011_0101111001111100"; -- 0.008352189260360817
	pesos_i(19222) := b"0000000000000000_0000000000000000_0001111111010011_0010101100110011"; -- 0.12431592939554262
	pesos_i(19223) := b"1111111111111111_1111111111111111_1111011111100101_0100010110010011"; -- -0.031657840420750614
	pesos_i(19224) := b"0000000000000000_0000000000000000_0001001110111110_1101101100110110"; -- 0.07713098588027169
	pesos_i(19225) := b"0000000000000000_0000000000000000_0010100011110000_0010001110100101"; -- 0.15991423402712365
	pesos_i(19226) := b"1111111111111111_1111111111111111_1110111101110101_1100000001101101"; -- -0.06460950214745571
	pesos_i(19227) := b"0000000000000000_0000000000000000_0010001010110011_1001001000100100"; -- 0.13555253398880257
	pesos_i(19228) := b"0000000000000000_0000000000000000_0010000001000001_0010101100111110"; -- 0.12599439883895175
	pesos_i(19229) := b"1111111111111111_1111111111111111_1110100010000111_1000111111100000"; -- -0.09168148778599997
	pesos_i(19230) := b"0000000000000000_0000000000000000_0010000001101110_0000001000001010"; -- 0.1266785883703954
	pesos_i(19231) := b"1111111111111111_1111111111111111_1101101101100111_0010101110011010"; -- -0.14295699588145716
	pesos_i(19232) := b"1111111111111111_1111111111111111_1111101110101110_0010000001010101"; -- -0.01687429364328009
	pesos_i(19233) := b"0000000000000000_0000000000000000_0010011110011100_0011001111000011"; -- 0.154727206218094
	pesos_i(19234) := b"1111111111111111_1111111111111111_1110010001110101_1000000111001010"; -- -0.1075819857151368
	pesos_i(19235) := b"0000000000000000_0000000000000000_0000100000110101_0010110110011000"; -- 0.032061433488215385
	pesos_i(19236) := b"1111111111111111_1111111111111111_1111001111110010_0101001010100010"; -- -0.04708369770371063
	pesos_i(19237) := b"0000000000000000_0000000000000000_0001111011001100_1010100011000010"; -- 0.12031035181445318
	pesos_i(19238) := b"1111111111111111_1111111111111111_1110010100100001_1000001001010010"; -- -0.10495744221200742
	pesos_i(19239) := b"0000000000000000_0000000000000000_0001010001001111_0100000101000011"; -- 0.07933433431199097
	pesos_i(19240) := b"1111111111111111_1111111111111111_1101111111100100_0111000001011100"; -- -0.12542054899414665
	pesos_i(19241) := b"0000000000000000_0000000000000000_0001011111001001_1100100010101010"; -- 0.09292272715304167
	pesos_i(19242) := b"1111111111111111_1111111111111111_1110000110110011_0000011010110001"; -- -0.1183620278128555
	pesos_i(19243) := b"0000000000000000_0000000000000000_0001011001010110_0101101111100101"; -- 0.08725523320330844
	pesos_i(19244) := b"0000000000000000_0000000000000000_0010011001000110_0010111000101110"; -- 0.14950836780457388
	pesos_i(19245) := b"1111111111111111_1111111111111111_1101111010001100_0111001010110101"; -- -0.1306694325050016
	pesos_i(19246) := b"0000000000000000_0000000000000000_0001000000010000_0011101010101000"; -- 0.06274763683442064
	pesos_i(19247) := b"0000000000000000_0000000000000000_0000000110001011_0000110111100111"; -- 0.006028050267491384
	pesos_i(19248) := b"1111111111111111_1111111111111111_1111010010110100_0001100000110110"; -- -0.04412697480968298
	pesos_i(19249) := b"0000000000000000_0000000000000000_0001001011101011_1101001110010110"; -- 0.07391092703237825
	pesos_i(19250) := b"0000000000000000_0000000000000000_0001010111101010_0110100110111111"; -- 0.0856081095120176
	pesos_i(19251) := b"1111111111111111_1111111111111111_1110101111010100_0110001100011011"; -- -0.07879047952802613
	pesos_i(19252) := b"0000000000000000_0000000000000000_0000000000111101_0101010111000000"; -- 0.0009358972479577242
	pesos_i(19253) := b"0000000000000000_0000000000000000_0000001000110011_0001101100100110"; -- 0.008592316348897603
	pesos_i(19254) := b"1111111111111111_1111111111111111_1110101011101101_1101000110110101"; -- -0.08230866741384645
	pesos_i(19255) := b"0000000000000000_0000000000000000_0010011000010010_1001000110101110"; -- 0.14872084138189184
	pesos_i(19256) := b"0000000000000000_0000000000000000_0001000110000011_0010000100111101"; -- 0.06840713262192091
	pesos_i(19257) := b"0000000000000000_0000000000000000_0000100101101001_1100100011100111"; -- 0.036770397654248534
	pesos_i(19258) := b"0000000000000000_0000000000000000_0000001110001011_0010100110111101"; -- 0.013842209383071796
	pesos_i(19259) := b"0000000000000000_0000000000000000_0001101010101110_0010111100010110"; -- 0.10422033573407766
	pesos_i(19260) := b"1111111111111111_1111111111111111_1110011001111000_1010000100000110"; -- -0.09972184746917592
	pesos_i(19261) := b"0000000000000000_0000000000000000_0000111001110100_1110011110001101"; -- 0.056471320982931505
	pesos_i(19262) := b"0000000000000000_0000000000000000_0000011001110001_1111011111001010"; -- 0.02517651245262835
	pesos_i(19263) := b"0000000000000000_0000000000000000_0001111110000101_0011110011111010"; -- 0.12312680353880183
	pesos_i(19264) := b"0000000000000000_0000000000000000_0010000100111110_0100011100001100"; -- 0.12985652975824816
	pesos_i(19265) := b"1111111111111111_1111111111111111_1110110010011100_1100110010001111"; -- -0.07573243620383498
	pesos_i(19266) := b"1111111111111111_1111111111111111_1110011010000100_0111011000001110"; -- -0.09954130324587505
	pesos_i(19267) := b"1111111111111111_1111111111111111_1111110110100010_1011010100100010"; -- -0.00923602984125374
	pesos_i(19268) := b"1111111111111111_1111111111111111_1110111010110000_1101110010001001"; -- -0.06761380819987613
	pesos_i(19269) := b"1111111111111111_1111111111111111_1111100110101001_0101011000001001"; -- -0.02475988661375801
	pesos_i(19270) := b"0000000000000000_0000000000000000_0001110011010100_0101001110011100"; -- 0.11261484682188981
	pesos_i(19271) := b"0000000000000000_0000000000000000_0001100110101101_0000111100001100"; -- 0.10029691742506461
	pesos_i(19272) := b"1111111111111111_1111111111111111_1111010010000010_1101000001000011"; -- -0.04487894397895173
	pesos_i(19273) := b"0000000000000000_0000000000000000_0000100001011101_0011111100101100"; -- 0.03267283275545167
	pesos_i(19274) := b"1111111111111111_1111111111111111_1110011000010100_1000001100110101"; -- -0.10124950375450326
	pesos_i(19275) := b"1111111111111111_1111111111111111_1101101001110001_0000101001111001"; -- -0.14671263262027223
	pesos_i(19276) := b"1111111111111111_1111111111111111_1111110110010010_0001010000001111"; -- -0.009489771218118942
	pesos_i(19277) := b"1111111111111111_1111111111111111_1101101010000110_0000001111110000"; -- -0.14639258758342788
	pesos_i(19278) := b"0000000000000000_0000000000000000_0000000011110101_1111001111100101"; -- 0.003752940476386687
	pesos_i(19279) := b"1111111111111111_1111111111111111_1111101011000010_0100111011100011"; -- -0.020472592864030876
	pesos_i(19280) := b"1111111111111111_1111111111111111_1111001101010110_0011100010100101"; -- -0.04946561786071159
	pesos_i(19281) := b"0000000000000000_0000000000000000_0000101100010111_0111010111010011"; -- 0.04332672490928441
	pesos_i(19282) := b"1111111111111111_1111111111111111_1101100101110111_1101111111101010"; -- -0.15051460772627634
	pesos_i(19283) := b"0000000000000000_0000000000000000_0000110101011110_0101010110011111"; -- 0.05222067956642081
	pesos_i(19284) := b"0000000000000000_0000000000000000_0001000001111011_1000011010100101"; -- 0.06438485660257771
	pesos_i(19285) := b"1111111111111111_1111111111111111_1111101110010110_0000001111000100"; -- -0.01724220714368252
	pesos_i(19286) := b"0000000000000000_0000000000000000_0001001110100100_1011011010101010"; -- 0.07673207895033902
	pesos_i(19287) := b"1111111111111111_1111111111111111_1110101001101100_0100101101101001"; -- -0.08428505608614172
	pesos_i(19288) := b"1111111111111111_1111111111111111_1110101100111110_0111100011011100"; -- -0.08107800135511972
	pesos_i(19289) := b"1111111111111111_1111111111111111_1101101110000010_1001001000011011"; -- -0.14253889888411378
	pesos_i(19290) := b"1111111111111111_1111111111111111_1110110011111110_1001011111110100"; -- -0.07424021046319161
	pesos_i(19291) := b"1111111111111111_1111111111111111_1111011001111111_0111111111001001"; -- -0.037117017313711205
	pesos_i(19292) := b"0000000000000000_0000000000000000_0001110101100001_1110000110010001"; -- 0.11477479737906802
	pesos_i(19293) := b"0000000000000000_0000000000000000_0001010100100001_1000001001100000"; -- 0.08254256103511624
	pesos_i(19294) := b"0000000000000000_0000000000000000_0001010111110110_0100011101110111"; -- 0.08578917173435555
	pesos_i(19295) := b"0000000000000000_0000000000000000_0001111010111001_1111101100001111"; -- 0.12002534031182616
	pesos_i(19296) := b"0000000000000000_0000000000000000_0001100000100101_0101100011010010"; -- 0.09431986926960642
	pesos_i(19297) := b"1111111111111111_1111111111111111_1110010011111101_0001100110111010"; -- -0.10551299287213269
	pesos_i(19298) := b"1111111111111111_1111111111111111_1110110001100110_1011100111111101"; -- -0.07655751782360548
	pesos_i(19299) := b"1111111111111111_1111111111111111_1101111010110001_0101101010011110"; -- -0.13010629306766788
	pesos_i(19300) := b"1111111111111111_1111111111111111_1111110100001101_0110011101000011"; -- -0.011514230797432736
	pesos_i(19301) := b"1111111111111111_1111111111111111_1111101100011101_1110011111001001"; -- -0.019074929726227097
	pesos_i(19302) := b"1111111111111111_1111111111111111_1111011010010000_1101101101001100"; -- -0.03685216335706533
	pesos_i(19303) := b"1111111111111111_1111111111111111_1111000010110101_0011100100011100"; -- -0.05973475520193944
	pesos_i(19304) := b"1111111111111111_1111111111111111_1111111100110110_0011110101100111"; -- -0.0030786155366765086
	pesos_i(19305) := b"1111111111111111_1111111111111111_1110011110011001_1101100101101001"; -- -0.09530869654813347
	pesos_i(19306) := b"1111111111111111_1111111111111111_1111001010101011_1001111110010110"; -- -0.05206873502737782
	pesos_i(19307) := b"0000000000000000_0000000000000000_0001101111000101_0100110100110100"; -- 0.10847933304207824
	pesos_i(19308) := b"0000000000000000_0000000000000000_0001010110001101_0110101101000000"; -- 0.08418913182078092
	pesos_i(19309) := b"0000000000000000_0000000000000000_0010001000111000_1011111100010010"; -- 0.1336783809601225
	pesos_i(19310) := b"0000000000000000_0000000000000000_0001000111011100_1111000111100011"; -- 0.06977760120698515
	pesos_i(19311) := b"0000000000000000_0000000000000000_0001011100101101_1001110101000100"; -- 0.09053976934269328
	pesos_i(19312) := b"0000000000000000_0000000000000000_0001110101100001_0110111011001010"; -- 0.11476795607501002
	pesos_i(19313) := b"1111111111111111_1111111111111111_1101110010101010_0101110000100001"; -- -0.13802551452652995
	pesos_i(19314) := b"0000000000000000_0000000000000000_0000101110001111_1011000101000100"; -- 0.045161322738708626
	pesos_i(19315) := b"1111111111111111_1111111111111111_1110000110110110_0111101001111110"; -- -0.1183093493731475
	pesos_i(19316) := b"0000000000000000_0000000000000000_0001001011111010_0011110000101001"; -- 0.07413078308033876
	pesos_i(19317) := b"1111111111111111_1111111111111111_1110011100000101_0101110001010000"; -- -0.09757445376055554
	pesos_i(19318) := b"1111111111111111_1111111111111111_1101100101001001_1001000111101010"; -- -0.15122116120333773
	pesos_i(19319) := b"1111111111111111_1111111111111111_1110110111101001_0001111111100111"; -- -0.07066155060641088
	pesos_i(19320) := b"0000000000000000_0000000000000000_0001110111110001_0010000100100000"; -- 0.11696059249226641
	pesos_i(19321) := b"0000000000000000_0000000000000000_0010000001101000_0011100011011010"; -- 0.12659030257607395
	pesos_i(19322) := b"0000000000000000_0000000000000000_0001001001010001_0011101010001101"; -- 0.07155195188351662
	pesos_i(19323) := b"0000000000000000_0000000000000000_0000001100111001_1011010111011000"; -- 0.012599339731614317
	pesos_i(19324) := b"0000000000000000_0000000000000000_0000100011100100_1000101110010000"; -- 0.03473732249992829
	pesos_i(19325) := b"0000000000000000_0000000000000000_0001011011010001_1110000101011101"; -- 0.08914001951625097
	pesos_i(19326) := b"0000000000000000_0000000000000000_0001010101111111_0100100010100110"; -- 0.08397344642063474
	pesos_i(19327) := b"0000000000000000_0000000000000000_0001110001101111_1001100000101111"; -- 0.11107779633389353
	pesos_i(19328) := b"1111111111111111_1111111111111111_1101110111000010_1100011001100100"; -- -0.13374671986222844
	pesos_i(19329) := b"0000000000000000_0000000000000000_0001011010000100_0101111111101100"; -- 0.0879573775048625
	pesos_i(19330) := b"0000000000000000_0000000000000000_0001110011101000_1011001100111100"; -- 0.11292572229778132
	pesos_i(19331) := b"1111111111111111_1111111111111111_1111000101110101_0110000001011110"; -- -0.056802727644560284
	pesos_i(19332) := b"0000000000000000_0000000000000000_0000111101100011_0010001110100011"; -- 0.06010649419913299
	pesos_i(19333) := b"1111111111111111_1111111111111111_1111100011010101_0100000010010001"; -- -0.027996029412541236
	pesos_i(19334) := b"1111111111111111_1111111111111111_1110000000011100_1110000111110000"; -- -0.12455928703594674
	pesos_i(19335) := b"1111111111111111_1111111111111111_1111000001011110_0000110110101111"; -- -0.06106485820111494
	pesos_i(19336) := b"1111111111111111_1111111111111111_1101110000000111_1110110110010011"; -- -0.14050402792857772
	pesos_i(19337) := b"0000000000000000_0000000000000000_0001111100100101_0101000111100101"; -- 0.12166320647415371
	pesos_i(19338) := b"0000000000000000_0000000000000000_0000000111111100_0000010100111001"; -- 0.007751776095424405
	pesos_i(19339) := b"1111111111111111_1111111111111111_1111011111010011_1110001011011011"; -- -0.031923123783396574
	pesos_i(19340) := b"1111111111111111_1111111111111111_1110010010111100_1110000100001111"; -- -0.10649293303931637
	pesos_i(19341) := b"1111111111111111_1111111111111111_1111111011000111_1000110100111011"; -- -0.004767582882728918
	pesos_i(19342) := b"0000000000000000_0000000000000000_0000000101001101_1100100111000011"; -- 0.0050932027936441615
	pesos_i(19343) := b"0000000000000000_0000000000000000_0000000000100100_0101101001010000"; -- 0.0005546994158137712
	pesos_i(19344) := b"0000000000000000_0000000000000000_0000101000110000_0100110110110000"; -- 0.039799552466120824
	pesos_i(19345) := b"0000000000000000_0000000000000000_0010000110011101_0010100110110000"; -- 0.13130436475050283
	pesos_i(19346) := b"1111111111111111_1111111111111111_1111000001011001_0010100001101111"; -- -0.061139557732789236
	pesos_i(19347) := b"1111111111111111_1111111111111111_1110010101000111_1101010000010110"; -- -0.10437273466142141
	pesos_i(19348) := b"0000000000000000_0000000000000000_0000011010010110_1000110111111100"; -- 0.02573478123243211
	pesos_i(19349) := b"1111111111111111_1111111111111111_1110101001011111_0111000111101101"; -- -0.0844811245595109
	pesos_i(19350) := b"1111111111111111_1111111111111111_1110010111101001_0000100110000110"; -- -0.10191288456791153
	pesos_i(19351) := b"0000000000000000_0000000000000000_0000101101001101_0110011011001010"; -- 0.0441498034784122
	pesos_i(19352) := b"0000000000000000_0000000000000000_0001011011110110_1101100111101001"; -- 0.08970415059294227
	pesos_i(19353) := b"0000000000000000_0000000000000000_0001001010111111_1100100100010111"; -- 0.07323891455285571
	pesos_i(19354) := b"0000000000000000_0000000000000000_0000000100110001_1110000100011110"; -- 0.00466734869187239
	pesos_i(19355) := b"1111111111111111_1111111111111111_1110010100100011_1011010001001001"; -- -0.10492394666349356
	pesos_i(19356) := b"1111111111111111_1111111111111111_1101111100000110_0101000110010101"; -- -0.12880983454953004
	pesos_i(19357) := b"1111111111111111_1111111111111111_1111101010010100_1111111011111010"; -- -0.021164001337048426
	pesos_i(19358) := b"1111111111111111_1111111111111111_1101110000101000_1011100111000001"; -- -0.1400035765850514
	pesos_i(19359) := b"0000000000000000_0000000000000000_0001001010011000_0011111111111010"; -- 0.0726356492432005
	pesos_i(19360) := b"1111111111111111_1111111111111111_1110010110000111_1011011111100100"; -- -0.10339785283843127
	pesos_i(19361) := b"0000000000000000_0000000000000000_0010001001101000_1000110010110110"; -- 0.13440780097319685
	pesos_i(19362) := b"0000000000000000_0000000000000000_0001111001001011_1110111110111011"; -- 0.11834619818069174
	pesos_i(19363) := b"1111111111111111_1111111111111111_1111100100010000_1011100111010000"; -- -0.02708853403654106
	pesos_i(19364) := b"1111111111111111_1111111111111111_1111000001110111_0111110100011100"; -- -0.06067674695606523
	pesos_i(19365) := b"0000000000000000_0000000000000000_0001110010100011_0100011110100011"; -- 0.11186645255333882
	pesos_i(19366) := b"0000000000000000_0000000000000000_0001110110011110_1011110000100110"; -- 0.11570335325254626
	pesos_i(19367) := b"0000000000000000_0000000000000000_0001101011101101_1011100110111011"; -- 0.10518990332456096
	pesos_i(19368) := b"0000000000000000_0000000000000000_0010000101100100_1100111101010101"; -- 0.1304444869666308
	pesos_i(19369) := b"1111111111111111_1111111111111111_1111110100100000_0100000101010110"; -- -0.011226574366047671
	pesos_i(19370) := b"1111111111111111_1111111111111111_1111101011001101_0110010110011001"; -- -0.02030339255765881
	pesos_i(19371) := b"0000000000000000_0000000000000000_0000011110100111_1110011000100010"; -- 0.029905684727949765
	pesos_i(19372) := b"1111111111111111_1111111111111111_1111000111111111_0011010100011001"; -- -0.054699594036659506
	pesos_i(19373) := b"1111111111111111_1111111111111111_1101111111111101_1111001100011110"; -- -0.12503128556549742
	pesos_i(19374) := b"0000000000000000_0000000000000000_0000011100101000_1001111001000000"; -- 0.027963534000885228
	pesos_i(19375) := b"1111111111111111_1111111111111111_1110011110010101_0100111000111101"; -- -0.09537802717925468
	pesos_i(19376) := b"0000000000000000_0000000000000000_0000111001101001_1100100101011010"; -- 0.05630167429643885
	pesos_i(19377) := b"0000000000000000_0000000000000000_0001110100001111_1100110001101100"; -- 0.11352231622370183
	pesos_i(19378) := b"0000000000000000_0000000000000000_0000001011001100_0000101010001111"; -- 0.010925922335022936
	pesos_i(19379) := b"0000000000000000_0000000000000000_0010000010001001_0000001110101111"; -- 0.12709067359848225
	pesos_i(19380) := b"0000000000000000_0000000000000000_0000100110001001_0110111111011111"; -- 0.037253372071492354
	pesos_i(19381) := b"0000000000000000_0000000000000000_0001001001010000_1011011101011000"; -- 0.07154413132193824
	pesos_i(19382) := b"0000000000000000_0000000000000000_0001110000001001_0110101001110011"; -- 0.10951867401766488
	pesos_i(19383) := b"1111111111111111_1111111111111111_1111111110101111_1100110010011110"; -- -0.0012237657231737203
	pesos_i(19384) := b"0000000000000000_0000000000000000_0001010010000001_0011111001100001"; -- 0.08009710187895593
	pesos_i(19385) := b"1111111111111111_1111111111111111_1111010010000101_1001100100001101"; -- -0.04483645846408021
	pesos_i(19386) := b"1111111111111111_1111111111111111_1111010000001100_0110000011100111"; -- -0.04668611878781251
	pesos_i(19387) := b"1111111111111111_1111111111111111_1111100010001110_1101011101101001"; -- -0.029070412542479086
	pesos_i(19388) := b"0000000000000000_0000000000000000_0000100011011001_0010010011001110"; -- 0.03456335096100035
	pesos_i(19389) := b"0000000000000000_0000000000000000_0001000110010000_0111000001010000"; -- 0.06861020994425655
	pesos_i(19390) := b"0000000000000000_0000000000000000_0000101010010110_0010001001000001"; -- 0.04135336001635001
	pesos_i(19391) := b"0000000000000000_0000000000000000_0000001111010011_0111110110101101"; -- 0.014945845277816523
	pesos_i(19392) := b"0000000000000000_0000000000000000_0000011101100010_1000100011011001"; -- 0.028847268109486193
	pesos_i(19393) := b"1111111111111111_1111111111111111_1111101110100000_0000101100011101"; -- -0.017089181328184728
	pesos_i(19394) := b"1111111111111111_1111111111111111_1110011000100101_1100111100110100"; -- -0.10098557456264115
	pesos_i(19395) := b"1111111111111111_1111111111111111_1110100011110110_0010010111111101"; -- -0.08999407354588664
	pesos_i(19396) := b"1111111111111111_1111111111111111_1110001101011101_0101000100000000"; -- -0.1118573546343854
	pesos_i(19397) := b"1111111111111111_1111111111111111_1111111100001110_1000010101100010"; -- -0.0036846766685802255
	pesos_i(19398) := b"1111111111111111_1111111111111111_1110101011101010_0111101101101110"; -- -0.08235958643148951
	pesos_i(19399) := b"1111111111111111_1111111111111111_1110110000011110_1000000101110011"; -- -0.07765952051282171
	pesos_i(19400) := b"1111111111111111_1111111111111111_1110010111101100_1011111101101100"; -- -0.1018562662562976
	pesos_i(19401) := b"1111111111111111_1111111111111111_1111110101010110_1011101111000111"; -- -0.010395301645305513
	pesos_i(19402) := b"1111111111111111_1111111111111111_1111111100100111_1110010111111011"; -- -0.0032974494030252074
	pesos_i(19403) := b"0000000000000000_0000000000000000_0001100010011101_1110011000000100"; -- 0.09615933979735626
	pesos_i(19404) := b"1111111111111111_1111111111111111_1101111000111010_1101000011011110"; -- -0.1319150407243056
	pesos_i(19405) := b"1111111111111111_1111111111111111_1110011010100100_1000110011001000"; -- -0.09905166740614438
	pesos_i(19406) := b"1111111111111111_1111111111111111_1110001111001000_0011010000010011"; -- -0.11022638838515268
	pesos_i(19407) := b"0000000000000000_0000000000000000_0000000111110111_0000110011101011"; -- 0.0076759409633809575
	pesos_i(19408) := b"0000000000000000_0000000000000000_0000101100001100_1011011101000110"; -- 0.04316277952526145
	pesos_i(19409) := b"0000000000000000_0000000000000000_0000100000010001_1111010100010001"; -- 0.03152400646297704
	pesos_i(19410) := b"0000000000000000_0000000000000000_0001101101010000_0100010100111100"; -- 0.10669357984115456
	pesos_i(19411) := b"0000000000000000_0000000000000000_0000111000110001_0110110000010011"; -- 0.05544162249521404
	pesos_i(19412) := b"0000000000000000_0000000000000000_0000010110010110_1000001101101101"; -- 0.021827901903946966
	pesos_i(19413) := b"0000000000000000_0000000000000000_0000000111111111_1111011000100110"; -- 0.007811912721081469
	pesos_i(19414) := b"1111111111111111_1111111111111111_1110111101001001_1011011010100010"; -- -0.06528147273419792
	pesos_i(19415) := b"1111111111111111_1111111111111111_1111111101000110_1111010111101011"; -- -0.0028234768718031185
	pesos_i(19416) := b"1111111111111111_1111111111111111_1111000011100110_1101010011010011"; -- -0.058977793091104375
	pesos_i(19417) := b"1111111111111111_1111111111111111_1111001010101001_0000011111000110"; -- -0.052108301372056846
	pesos_i(19418) := b"0000000000000000_0000000000000000_0000001101100100_0000001111100011"; -- 0.013244860543687988
	pesos_i(19419) := b"0000000000000000_0000000000000000_0000110100000001_0100010110000011"; -- 0.050800652072550176
	pesos_i(19420) := b"1111111111111111_1111111111111111_1101110110101011_0010100001001101"; -- -0.13410709489388703
	pesos_i(19421) := b"1111111111111111_1111111111111111_1101110001111101_0001101001100011"; -- -0.13871607855294443
	pesos_i(19422) := b"1111111111111111_1111111111111111_1111011111101000_0110010001110110"; -- -0.03161022311118778
	pesos_i(19423) := b"0000000000000000_0000000000000000_0001001111111011_1111101100110001"; -- 0.07806367825063275
	pesos_i(19424) := b"1111111111111111_1111111111111111_1101011100111111_0110110101000100"; -- -0.1591884336331145
	pesos_i(19425) := b"1111111111111111_1111111111111111_1110111000010110_0100110010011100"; -- -0.06997224025126536
	pesos_i(19426) := b"0000000000000000_0000000000000000_0010001101110111_0001101111011110"; -- 0.1385362068524007
	pesos_i(19427) := b"0000000000000000_0000000000000000_0010000111001011_1001110010100110"; -- 0.13201312106043342
	pesos_i(19428) := b"1111111111111111_1111111111111111_1111011100010110_1111001011100001"; -- -0.034806080006899436
	pesos_i(19429) := b"1111111111111111_1111111111111111_1101101111100010_1011100000000011"; -- -0.14107179575465523
	pesos_i(19430) := b"1111111111111111_1111111111111111_1111101001101111_0110100101101000"; -- -0.021737491740950337
	pesos_i(19431) := b"1111111111111111_1111111111111111_1101011111010001_1001001000011111"; -- -0.15695845356812146
	pesos_i(19432) := b"1111111111111111_1111111111111111_1110100001111010_1001110111101100"; -- -0.0918790148195158
	pesos_i(19433) := b"1111111111111111_1111111111111111_1101101001000101_0000011110100111"; -- -0.14738418742414425
	pesos_i(19434) := b"1111111111111111_1111111111111111_1101110011011110_0100000101011000"; -- -0.13723365395970105
	pesos_i(19435) := b"0000000000000000_0000000000000000_0000111111010100_0100011001110011"; -- 0.06183281233898333
	pesos_i(19436) := b"0000000000000000_0000000000000000_0000001101101110_1000101100000101"; -- 0.01340550297931709
	pesos_i(19437) := b"0000000000000000_0000000000000000_0000101001101010_0001011011111110"; -- 0.04068130201713187
	pesos_i(19438) := b"1111111111111111_1111111111111111_1111010101111100_0101010110101100"; -- -0.04107155370003765
	pesos_i(19439) := b"1111111111111111_1111111111111111_1110010001011010_1001000101110100"; -- -0.10799303921765299
	pesos_i(19440) := b"0000000000000000_0000000000000000_0010011010110001_0000100010011110"; -- 0.15113881919986596
	pesos_i(19441) := b"0000000000000000_0000000000000000_0001100101100011_0000010100110101"; -- 0.09916718056851043
	pesos_i(19442) := b"0000000000000000_0000000000000000_0000100110110000_0101010000010101"; -- 0.037846808482554846
	pesos_i(19443) := b"0000000000000000_0000000000000000_0000100000111001_1111000101111011"; -- 0.032134144433788085
	pesos_i(19444) := b"1111111111111111_1111111111111111_1111000011000001_1110100000011001"; -- -0.05954121963620491
	pesos_i(19445) := b"1111111111111111_1111111111111111_1110001010111110_0000100110100010"; -- -0.11428775584377994
	pesos_i(19446) := b"0000000000000000_0000000000000000_0001100011001110_1101101100000111"; -- 0.09690636553201609
	pesos_i(19447) := b"0000000000000000_0000000000000000_0001101001100011_1101011111011011"; -- 0.10308598619191506
	pesos_i(19448) := b"0000000000000000_0000000000000000_0010011000110011_0100000010110010"; -- 0.14921955432575246
	pesos_i(19449) := b"0000000000000000_0000000000000000_0000001011110111_1001110001001101"; -- 0.01159073716714224
	pesos_i(19450) := b"0000000000000000_0000000000000000_0000101101110010_0001100111100001"; -- 0.04470979454406487
	pesos_i(19451) := b"0000000000000000_0000000000000000_0000001010100111_0110000011011000"; -- 0.010366490094991928
	pesos_i(19452) := b"0000000000000000_0000000000000000_0000010001100011_1110000000000111"; -- 0.01714897309197274
	pesos_i(19453) := b"1111111111111111_1111111111111111_1110101001100010_0001001010011100"; -- -0.08444102946041575
	pesos_i(19454) := b"0000000000000000_0000000000000000_0010000101110100_1100000110110111"; -- 0.13068781579940814
	pesos_i(19455) := b"0000000000000000_0000000000000000_0000000100101010_1011001111001111"; -- 0.004557836588619244
	pesos_i(19456) := b"1111111111111111_1111111111111111_1110000101101111_0100010110100101"; -- -0.11939587328928218
	pesos_i(19457) := b"0000000000000000_0000000000000000_0000000111010000_0010000101101110"; -- 0.007082070624554103
	pesos_i(19458) := b"1111111111111111_1111111111111111_1110111111101101_0100000100001111"; -- -0.06278603919871792
	pesos_i(19459) := b"0000000000000000_0000000000000000_0001010111001111_0001000000001010"; -- 0.08519077524741232
	pesos_i(19460) := b"0000000000000000_0000000000000000_0000001000000011_0101101010010110"; -- 0.007863675741856466
	pesos_i(19461) := b"1111111111111111_1111111111111111_1110000111011011_1110110011001101"; -- -0.11773796079259988
	pesos_i(19462) := b"0000000000000000_0000000000000000_0001100000111001_1011111011010001"; -- 0.09463112456560975
	pesos_i(19463) := b"1111111111111111_1111111111111111_1110101010001010_1110000101001110"; -- -0.08381835801647526
	pesos_i(19464) := b"1111111111111111_1111111111111111_1110100000100000_1100011100001010"; -- -0.09324985506024254
	pesos_i(19465) := b"1111111111111111_1111111111111111_1110001011111100_0001000111000011"; -- -0.1133412265314049
	pesos_i(19466) := b"0000000000000000_0000000000000000_0000011001100000_0100000110000001"; -- 0.024906248013705844
	pesos_i(19467) := b"1111111111111111_1111111111111111_1111100110101101_0101111110000111"; -- -0.024698285537640915
	pesos_i(19468) := b"0000000000000000_0000000000000000_0001101011110001_0010000101111000"; -- 0.10524186302593293
	pesos_i(19469) := b"0000000000000000_0000000000000000_0000011110011000_0101100001100001"; -- 0.029668353778822595
	pesos_i(19470) := b"0000000000000000_0000000000000000_0001100000001000_0111000001001011"; -- 0.09387876338588938
	pesos_i(19471) := b"1111111111111111_1111111111111111_1111111100110111_0001010100101010"; -- -0.0030657550102221073
	pesos_i(19472) := b"0000000000000000_0000000000000000_0010000110111001_1010110001010110"; -- 0.1317393979156381
	pesos_i(19473) := b"1111111111111111_1111111111111111_1110111011001011_1011011000111000"; -- -0.0672041046636495
	pesos_i(19474) := b"0000000000000000_0000000000000000_0010101101010100_0110010110011000"; -- 0.16925654383695377
	pesos_i(19475) := b"1111111111111111_1111111111111111_1111000100101110_0011001110101000"; -- -0.05788876671733134
	pesos_i(19476) := b"1111111111111111_1111111111111111_1110100010010010_1011000101110000"; -- -0.09151164068442856
	pesos_i(19477) := b"0000000000000000_0000000000000000_0001010110100010_0110111010011100"; -- 0.08450976671542856
	pesos_i(19478) := b"0000000000000000_0000000000000000_0010000010101001_0110000011000110"; -- 0.12758450360305892
	pesos_i(19479) := b"0000000000000000_0000000000000000_0001010101011001_1000101000101001"; -- 0.08339751729736497
	pesos_i(19480) := b"1111111111111111_1111111111111111_1110010110011100_1001000001001001"; -- -0.1030797788452342
	pesos_i(19481) := b"1111111111111111_1111111111111111_1111111010101110_1111010100110011"; -- -0.005142855719494839
	pesos_i(19482) := b"1111111111111111_1111111111111111_1110000100010111_1110010100011001"; -- -0.120729142626489
	pesos_i(19483) := b"1111111111111111_1111111111111111_1111000010111111_0010110110101100"; -- -0.0595828491173624
	pesos_i(19484) := b"0000000000000000_0000000000000000_0000110000010010_0100010110100011"; -- 0.04715380890152758
	pesos_i(19485) := b"1111111111111111_1111111111111111_1101101001101101_1110101101101110"; -- -0.1467602592405372
	pesos_i(19486) := b"0000000000000000_0000000000000000_0010001000101110_0011010101000110"; -- 0.13351757965435587
	pesos_i(19487) := b"0000000000000000_0000000000000000_0001101010011000_0001000011110000"; -- 0.10388284555226628
	pesos_i(19488) := b"0000000000000000_0000000000000000_0001011110100110_0100110111010100"; -- 0.09238134785978064
	pesos_i(19489) := b"0000000000000000_0000000000000000_0010001111000000_0011000101010010"; -- 0.1396513771486138
	pesos_i(19490) := b"1111111111111111_1111111111111111_1110000000111001_0011010010010011"; -- -0.1241271154306859
	pesos_i(19491) := b"0000000000000000_0000000000000000_0010001110001101_1111000000110101"; -- 0.13888455670327543
	pesos_i(19492) := b"1111111111111111_1111111111111111_1101111100110011_1001100101111000"; -- -0.128118904214447
	pesos_i(19493) := b"0000000000000000_0000000000000000_0001010101011111_0000001111010111"; -- 0.08348106387053633
	pesos_i(19494) := b"0000000000000000_0000000000000000_0001011010010111_1010111110111000"; -- 0.08825205070903681
	pesos_i(19495) := b"0000000000000000_0000000000000000_0010100101110011_0111011001000111"; -- 0.16191806068956846
	pesos_i(19496) := b"1111111111111111_1111111111111111_1101101101110101_1100000101001000"; -- -0.14273445123270298
	pesos_i(19497) := b"1111111111111111_1111111111111111_1111111010111000_0010001000111101"; -- -0.005002841988904691
	pesos_i(19498) := b"1111111111111111_1111111111111111_1110010010111111_0011110011100000"; -- -0.10645694274548284
	pesos_i(19499) := b"0000000000000000_0000000000000000_0000101001010101_0110000010111011"; -- 0.04036526260425506
	pesos_i(19500) := b"1111111111111111_1111111111111111_1111101000111110_1011001010100110"; -- -0.02248080687198473
	pesos_i(19501) := b"0000000000000000_0000000000000000_0001110010001100_1100010100101101"; -- 0.11152298295789972
	pesos_i(19502) := b"0000000000000000_0000000000000000_0010001010111101_1110011110010000"; -- 0.1357102133493465
	pesos_i(19503) := b"0000000000000000_0000000000000000_0000000101100100_0001001000011111"; -- 0.005433208919969634
	pesos_i(19504) := b"0000000000000000_0000000000000000_0000101011000011_1010110001110110"; -- 0.04204824345064213
	pesos_i(19505) := b"1111111111111111_1111111111111111_1101110101111111_0101111010100010"; -- -0.13477524317212605
	pesos_i(19506) := b"1111111111111111_1111111111111111_1110000101111111_1001000011111001"; -- -0.11914724265172609
	pesos_i(19507) := b"0000000000000000_0000000000000000_0000011001011110_1011001011100001"; -- 0.024882488291618852
	pesos_i(19508) := b"1111111111111111_1111111111111111_1111001101100011_0010000010010101"; -- -0.04926868778119451
	pesos_i(19509) := b"0000000000000000_0000000000000000_0000101010011101_1010100000010010"; -- 0.041468147644760645
	pesos_i(19510) := b"1111111111111111_1111111111111111_1110001001110101_0010000000001100"; -- -0.11540031150218899
	pesos_i(19511) := b"1111111111111111_1111111111111111_1111101111110111_0101110001000001"; -- -0.01575683036231379
	pesos_i(19512) := b"1111111111111111_1111111111111111_1110010000100100_1000101010000000"; -- -0.10881742823708607
	pesos_i(19513) := b"1111111111111111_1111111111111111_1111011101001010_1011010010011100"; -- -0.03401633455323274
	pesos_i(19514) := b"0000000000000000_0000000000000000_0001110001010110_0111100111000011"; -- 0.110694513520021
	pesos_i(19515) := b"1111111111111111_1111111111111111_1110010101100000_0011101000001110"; -- -0.10400044599257399
	pesos_i(19516) := b"1111111111111111_1111111111111111_1110100001110100_1110000000110110"; -- -0.0919666165661957
	pesos_i(19517) := b"1111111111111111_1111111111111111_1110010001100011_0010010000001111"; -- -0.10786223065639848
	pesos_i(19518) := b"0000000000000000_0000000000000000_0000111110100101_0100010111000110"; -- 0.06111560903709295
	pesos_i(19519) := b"1111111111111111_1111111111111111_1101110010101101_0110010110010111"; -- -0.1379791742569878
	pesos_i(19520) := b"0000000000000000_0000000000000000_0000001010100110_1110010111101100"; -- 0.01035916336087927
	pesos_i(19521) := b"1111111111111111_1111111111111111_1110101111110000_1100111101101011"; -- -0.07835677745373522
	pesos_i(19522) := b"1111111111111111_1111111111111111_1110000111001010_1001101000011000"; -- -0.11800228997349035
	pesos_i(19523) := b"0000000000000000_0000000000000000_0010101110100100_0000000011110011"; -- 0.17047124788511475
	pesos_i(19524) := b"0000000000000000_0000000000000000_0001001000011001_1000101011100000"; -- 0.07070224741027217
	pesos_i(19525) := b"1111111111111111_1111111111111111_1110001010110111_1011111101011111"; -- -0.11438373490324741
	pesos_i(19526) := b"1111111111111111_1111111111111111_1111011100001111_1111100001001110"; -- -0.03491256798067499
	pesos_i(19527) := b"0000000000000000_0000000000000000_0001101000100010_0010111001110110"; -- 0.10208406807014206
	pesos_i(19528) := b"0000000000000000_0000000000000000_0001001111110001_1100100111110111"; -- 0.07790815618065475
	pesos_i(19529) := b"0000000000000000_0000000000000000_0000110101000100_1111110110001111"; -- 0.05183396083227513
	pesos_i(19530) := b"1111111111111111_1111111111111111_1111100010000010_1110100111010101"; -- -0.029252420032271024
	pesos_i(19531) := b"1111111111111111_1111111111111111_1101110100100110_0011100001101011"; -- -0.13613555320647128
	pesos_i(19532) := b"1111111111111111_1111111111111111_1110001110110101_1011101111001100"; -- -0.11050821571715573
	pesos_i(19533) := b"1111111111111111_1111111111111111_1111011100000001_1010000110001000"; -- -0.03513136312167222
	pesos_i(19534) := b"1111111111111111_1111111111111111_1101111011000000_1000001010110000"; -- -0.12987502302032874
	pesos_i(19535) := b"1111111111111111_1111111111111111_1110000010101010_0101001000000000"; -- -0.12240111832272407
	pesos_i(19536) := b"1111111111111111_1111111111111111_1101100100111101_1001111011110010"; -- -0.15140348997537187
	pesos_i(19537) := b"1111111111111111_1111111111111111_1111000111010000_0011100111001101"; -- -0.055416476630092054
	pesos_i(19538) := b"1111111111111111_1111111111111111_1101111100001001_0100000010011010"; -- -0.12876507024400358
	pesos_i(19539) := b"0000000000000000_0000000000000000_0000101001010100_1001110000001100"; -- 0.04035353942411834
	pesos_i(19540) := b"1111111111111111_1111111111111111_1110011010100101_1100111111000000"; -- -0.09903241699921358
	pesos_i(19541) := b"0000000000000000_0000000000000000_0000100001001001_0001011100010010"; -- 0.03236526663584555
	pesos_i(19542) := b"1111111111111111_1111111111111111_1110111000000011_1111100011001000"; -- -0.07025189513648057
	pesos_i(19543) := b"0000000000000000_0000000000000000_0000001010100001_0110101100010001"; -- 0.010275546636061325
	pesos_i(19544) := b"0000000000000000_0000000000000000_0001010100010011_0111010111110010"; -- 0.08232819701658178
	pesos_i(19545) := b"0000000000000000_0000000000000000_0001000110100001_0101110001101110"; -- 0.0688684242034115
	pesos_i(19546) := b"1111111111111111_1111111111111111_1110011000101111_1101110110111010"; -- -0.10083212094772943
	pesos_i(19547) := b"0000000000000000_0000000000000000_0001101111001101_0001000010010010"; -- 0.10859778953838556
	pesos_i(19548) := b"1111111111111111_1111111111111111_1111101001110011_0111111000101010"; -- -0.02167521933529663
	pesos_i(19549) := b"1111111111111111_1111111111111111_1111000111110111_0011001110011011"; -- -0.05482175324911715
	pesos_i(19550) := b"1111111111111111_1111111111111111_1101011001100111_0111111100101111"; -- -0.16248326399520716
	pesos_i(19551) := b"0000000000000000_0000000000000000_0000101101011010_1110111110000010"; -- 0.04435631680939551
	pesos_i(19552) := b"1111111111111111_1111111111111111_1111000111100101_0100000000011001"; -- -0.05509566675994011
	pesos_i(19553) := b"1111111111111111_1111111111111111_1110000101100010_0100000000111010"; -- -0.11959456037615256
	pesos_i(19554) := b"1111111111111111_1111111111111111_1111001110011101_1001101100110110"; -- -0.04837636882809664
	pesos_i(19555) := b"1111111111111111_1111111111111111_1101100100110010_1101000010110011"; -- -0.15156837107471666
	pesos_i(19556) := b"0000000000000000_0000000000000000_0010000001100100_0100111111000101"; -- 0.1265306336233879
	pesos_i(19557) := b"1111111111111111_1111111111111111_1111100011101111_1010111110001101"; -- -0.02759268575124306
	pesos_i(19558) := b"0000000000000000_0000000000000000_0001000011011000_0110001001110001"; -- 0.0658017660490454
	pesos_i(19559) := b"1111111111111111_1111111111111111_1111111110000010_1011001000010110"; -- -0.0019119925848599267
	pesos_i(19560) := b"0000000000000000_0000000000000000_0001111001001000_1110001100000011"; -- 0.11829966387477117
	pesos_i(19561) := b"0000000000000000_0000000000000000_0010001010111100_0000100011000000"; -- 0.13568167386473676
	pesos_i(19562) := b"0000000000000000_0000000000000000_0001001101010101_1010100011011001"; -- 0.0755258111511911
	pesos_i(19563) := b"1111111111111111_1111111111111111_1111111111110011_0101110010111001"; -- -0.00019283744676629584
	pesos_i(19564) := b"0000000000000000_0000000000000000_0001100111011100_1000110100000001"; -- 0.10102158809763519
	pesos_i(19565) := b"1111111111111111_1111111111111111_1111011001011000_0100001011101101"; -- -0.037715737565393294
	pesos_i(19566) := b"1111111111111111_1111111111111111_1110000000110010_1001101111011000"; -- -0.12422777157419851
	pesos_i(19567) := b"1111111111111111_1111111111111111_1111100000001111_0011001001001010"; -- -0.031018120815342512
	pesos_i(19568) := b"0000000000000000_0000000000000000_0010000101100000_1110000101111101"; -- 0.13038453389949886
	pesos_i(19569) := b"0000000000000000_0000000000000000_0000001011001111_1100001111001101"; -- 0.010982739900700558
	pesos_i(19570) := b"1111111111111111_1111111111111111_1101110100100101_0111100101101010"; -- -0.13614693802839842
	pesos_i(19571) := b"0000000000000000_0000000000000000_0010011111111001_1001111010110000"; -- 0.1561526469961057
	pesos_i(19572) := b"0000000000000000_0000000000000000_0001110101010100_0000011000000001"; -- 0.11456334608937682
	pesos_i(19573) := b"1111111111111111_1111111111111111_1101010000100000_1011011110110111"; -- -0.17137576853570172
	pesos_i(19574) := b"1111111111111111_1111111111111111_1111110100001001_1110101101010100"; -- -0.0115673942364337
	pesos_i(19575) := b"1111111111111111_1111111111111111_1101110011100111_0111000111110011"; -- -0.1370934277396005
	pesos_i(19576) := b"0000000000000000_0000000000000000_0010000110111000_1010010000010110"; -- 0.13172364742580436
	pesos_i(19577) := b"0000000000000000_0000000000000000_0000011010010010_0011000001011100"; -- 0.02566816559527588
	pesos_i(19578) := b"1111111111111111_1111111111111111_1111100110001111_0111100000000101"; -- -0.025154589420812033
	pesos_i(19579) := b"1111111111111111_1111111111111111_1111001101010001_1110111010010011"; -- -0.049531067933969844
	pesos_i(19580) := b"1111111111111111_1111111111111111_1110110110101100_1010110110011011"; -- -0.07158389051014093
	pesos_i(19581) := b"0000000000000000_0000000000000000_0000101011010111_0010101100100011"; -- 0.042345710712499054
	pesos_i(19582) := b"1111111111111111_1111111111111111_1111110110010110_1001101001001001"; -- -0.009420735591876029
	pesos_i(19583) := b"1111111111111111_1111111111111111_1111101111100001_1110000010110111"; -- -0.016084628398578903
	pesos_i(19584) := b"0000000000000000_0000000000000000_0001011000110110_1001000110101010"; -- 0.08677015697394268
	pesos_i(19585) := b"1111111111111111_1111111111111111_1101110101101111_1110000101110100"; -- -0.13501158624446838
	pesos_i(19586) := b"0000000000000000_0000000000000000_0001011000000110_1110001101100101"; -- 0.08604260642403634
	pesos_i(19587) := b"1111111111111111_1111111111111111_1110011100100101_0111100111110101"; -- -0.0970844055221458
	pesos_i(19588) := b"1111111111111111_1111111111111111_1111101110101101_0011000001001011"; -- -0.01688860106550457
	pesos_i(19589) := b"0000000000000000_0000000000000000_0010100101011100_0001011100111110"; -- 0.16156144394291505
	pesos_i(19590) := b"0000000000000000_0000000000000000_0000000110010010_1101001000001110"; -- 0.0061465533783269955
	pesos_i(19591) := b"0000000000000000_0000000000000000_0001010001110000_1111011000010000"; -- 0.07984865080621921
	pesos_i(19592) := b"1111111111111111_1111111111111111_1111000010011011_0110111010010110"; -- -0.06012829633755674
	pesos_i(19593) := b"0000000000000000_0000000000000000_0001000010000111_0010000010001000"; -- 0.06456187547407656
	pesos_i(19594) := b"0000000000000000_0000000000000000_0001001001000110_0101110100111100"; -- 0.07138617243951796
	pesos_i(19595) := b"1111111111111111_1111111111111111_1110111011110011_0101110100110101"; -- -0.06659905857388915
	pesos_i(19596) := b"0000000000000000_0000000000000000_0001010110101100_1100110000111000"; -- 0.08466793410042994
	pesos_i(19597) := b"1111111111111111_1111111111111111_1110101111101110_1010111110100101"; -- -0.07838918903397869
	pesos_i(19598) := b"1111111111111111_1111111111111111_1111000010100000_1111000110101101"; -- -0.06004418885891854
	pesos_i(19599) := b"0000000000000000_0000000000000000_0001110100011101_1101011110011010"; -- 0.11373660566440902
	pesos_i(19600) := b"1111111111111111_1111111111111111_1110001110000101_0001000000010100"; -- -0.11125087262219674
	pesos_i(19601) := b"0000000000000000_0000000000000000_0000011011001001_0110111110010100"; -- 0.026511167262061184
	pesos_i(19602) := b"0000000000000000_0000000000000000_0000101011001001_1101100011110001"; -- 0.04214244741479471
	pesos_i(19603) := b"0000000000000000_0000000000000000_0000111010010011_0101010010011110"; -- 0.05693558567369741
	pesos_i(19604) := b"0000000000000000_0000000000000000_0001010110110100_1100111011010011"; -- 0.08479015972303636
	pesos_i(19605) := b"0000000000000000_0000000000000000_0001110110010011_1011101011000111"; -- 0.1155354248889943
	pesos_i(19606) := b"1111111111111111_1111111111111111_1110000011111001_0110010100111000"; -- -0.12119452834929462
	pesos_i(19607) := b"1111111111111111_1111111111111111_1101110000011000_1100101011101111"; -- -0.14024669330912884
	pesos_i(19608) := b"1111111111111111_1111111111111111_1110010100011000_0001111000111110"; -- -0.10510073648712948
	pesos_i(19609) := b"0000000000000000_0000000000000000_0001010000010010_1000111010001101"; -- 0.0784081549426906
	pesos_i(19610) := b"1111111111111111_1111111111111111_1110001000001001_0111100011101000"; -- -0.11704296440366956
	pesos_i(19611) := b"1111111111111111_1111111111111111_1111100001100011_0001101011010100"; -- -0.029737780865585203
	pesos_i(19612) := b"1111111111111111_1111111111111111_1110000011111100_1101000011010100"; -- -0.12114233800545073
	pesos_i(19613) := b"1111111111111111_1111111111111111_1110001000001011_0111001100010001"; -- -0.11701279475747935
	pesos_i(19614) := b"1111111111111111_1111111111111111_1101101101011101_0001010001010100"; -- -0.1431109709144698
	pesos_i(19615) := b"1111111111111111_1111111111111111_1111010011000011_0000111101000010"; -- -0.04389862679893559
	pesos_i(19616) := b"0000000000000000_0000000000000000_0000010100010001_0110011000100111"; -- 0.019796738187292485
	pesos_i(19617) := b"0000000000000000_0000000000000000_0001111011110010_0011011011000100"; -- 0.1208833912776539
	pesos_i(19618) := b"0000000000000000_0000000000000000_0001001000101100_1001011111100100"; -- 0.07099294019789111
	pesos_i(19619) := b"1111111111111111_1111111111111111_1101111111011101_1000100100111000"; -- -0.12552587882627522
	pesos_i(19620) := b"0000000000000000_0000000000000000_0001011100011111_1100011000111110"; -- 0.09032858870683826
	pesos_i(19621) := b"1111111111111111_1111111111111111_1101101101000101_0100100010001011"; -- -0.1434740695479463
	pesos_i(19622) := b"0000000000000000_0000000000000000_0001000100001011_1011001100010100"; -- 0.06658477049979876
	pesos_i(19623) := b"1111111111111111_1111111111111111_1111110101100100_1011111100101100"; -- -0.010181476327207516
	pesos_i(19624) := b"1111111111111111_1111111111111111_1111111001001001_1000110100001101"; -- -0.006690201142628109
	pesos_i(19625) := b"1111111111111111_1111111111111111_1111100000111101_0011111011010001"; -- -0.030315469613923732
	pesos_i(19626) := b"0000000000000000_0000000000000000_0000100010110110_1100111101000101"; -- 0.03403945391565788
	pesos_i(19627) := b"1111111111111111_1111111111111111_1110101000111101_0000001001100011"; -- -0.08500657151284251
	pesos_i(19628) := b"1111111111111111_1111111111111111_1111101100101011_1110100111100100"; -- -0.01886118110292871
	pesos_i(19629) := b"1111111111111111_1111111111111111_1110110101110010_0100011110011011"; -- -0.07247498008614904
	pesos_i(19630) := b"1111111111111111_1111111111111111_1101110011011101_0000101010000111"; -- -0.13725218004310444
	pesos_i(19631) := b"0000000000000000_0000000000000000_0001100011010011_1100110010001001"; -- 0.09698179564181061
	pesos_i(19632) := b"1111111111111111_1111111111111111_1111101100100110_1101011100111001"; -- -0.018938587749821663
	pesos_i(19633) := b"1111111111111111_1111111111111111_1110100110011101_1011010100011010"; -- -0.0874373256911332
	pesos_i(19634) := b"1111111111111111_1111111111111111_1110010011011110_0100010011101100"; -- -0.10598344072741059
	pesos_i(19635) := b"1111111111111111_1111111111111111_1111101010110001_0011110000001110"; -- -0.020733114784778024
	pesos_i(19636) := b"0000000000000000_0000000000000000_0001000001000100_1010101100101000"; -- 0.06354779930101341
	pesos_i(19637) := b"0000000000000000_0000000000000000_0001001001000111_0001100101101001"; -- 0.07139738862553846
	pesos_i(19638) := b"1111111111111111_1111111111111111_1110001000100001_1011000011100111"; -- -0.11667341578457067
	pesos_i(19639) := b"0000000000000000_0000000000000000_0010011011001100_0000100010100010"; -- 0.15155080746403785
	pesos_i(19640) := b"0000000000000000_0000000000000000_0000101111011100_1011100011101000"; -- 0.04633670487137338
	pesos_i(19641) := b"0000000000000000_0000000000000000_0000110010000000_0101101011010000"; -- 0.04883353791132612
	pesos_i(19642) := b"1111111111111111_1111111111111111_1110011101000100_1110100001110010"; -- -0.09660479751359305
	pesos_i(19643) := b"1111111111111111_1111111111111111_1111010000101010_0110011111100110"; -- -0.04622793812585266
	pesos_i(19644) := b"0000000000000000_0000000000000000_0001101100001011_1100000011010110"; -- 0.10564809060195046
	pesos_i(19645) := b"1111111111111111_1111111111111111_1110010100010110_0010010001111100"; -- -0.1051308819430082
	pesos_i(19646) := b"0000000000000000_0000000000000000_0010000001001101_1000110101101110"; -- 0.12618335662273775
	pesos_i(19647) := b"1111111111111111_1111111111111111_1101101001101101_1010001101100110"; -- -0.14676455263509805
	pesos_i(19648) := b"1111111111111111_1111111111111111_1110010100001101_1101100010000110"; -- -0.10525747989358601
	pesos_i(19649) := b"1111111111111111_1111111111111111_1110000101100111_1101001001000000"; -- -0.11950956285911322
	pesos_i(19650) := b"0000000000000000_0000000000000000_0000011000100101_0101100000110001"; -- 0.024007331771903395
	pesos_i(19651) := b"1111111111111111_1111111111111111_1111000101111100_1111001001110100"; -- -0.056687208827517474
	pesos_i(19652) := b"1111111111111111_1111111111111111_1111000010111010_0000001010000100"; -- -0.05966171529113729
	pesos_i(19653) := b"1111111111111111_1111111111111111_1111110111010101_0101001010000100"; -- -0.008463709649986542
	pesos_i(19654) := b"0000000000000000_0000000000000000_0001100100100001_0101101000100010"; -- 0.09816516246859609
	pesos_i(19655) := b"1111111111111111_1111111111111111_1110010101000101_0101000000100101"; -- -0.1044111164711198
	pesos_i(19656) := b"1111111111111111_1111111111111111_1111001100100001_1010101011100101"; -- -0.05026752378056549
	pesos_i(19657) := b"1111111111111111_1111111111111111_1101111110010011_0011110000101000"; -- -0.1266596223968886
	pesos_i(19658) := b"1111111111111111_1111111111111111_1111000001111000_1000111100100101"; -- -0.06066041315169821
	pesos_i(19659) := b"1111111111111111_1111111111111111_1110110110000010_1101000101010011"; -- -0.07222263073659464
	pesos_i(19660) := b"0000000000000000_0000000000000000_0010001011000101_0110100100101110"; -- 0.1358247506860469
	pesos_i(19661) := b"1111111111111111_1111111111111111_1110100010101100_1011000001111101"; -- -0.09111496865092909
	pesos_i(19662) := b"0000000000000000_0000000000000000_0000111001111111_0110110101000000"; -- 0.05663187792836309
	pesos_i(19663) := b"0000000000000000_0000000000000000_0000101110000011_1110000111110110"; -- 0.044981119651479974
	pesos_i(19664) := b"0000000000000000_0000000000000000_0010000000000000_1000010111011100"; -- 0.1250079785944467
	pesos_i(19665) := b"1111111111111111_1111111111111111_1110110101000101_1110001010010010"; -- -0.07315238883536553
	pesos_i(19666) := b"1111111111111111_1111111111111111_1110011110110110_1101000100111111"; -- -0.09486667841258994
	pesos_i(19667) := b"0000000000000000_0000000000000000_0001011111011110_0000101111011100"; -- 0.09323190793139835
	pesos_i(19668) := b"0000000000000000_0000000000000000_0000110001100101_1101011111110000"; -- 0.048429008550889746
	pesos_i(19669) := b"1111111111111111_1111111111111111_1110011111001111_1011111100101110"; -- -0.09448628538116696
	pesos_i(19670) := b"0000000000000000_0000000000000000_0000100001001101_1000011101010111"; -- 0.032432993744958775
	pesos_i(19671) := b"0000000000000000_0000000000000000_0000000010101011_1010001000011010"; -- 0.0026189148964495517
	pesos_i(19672) := b"0000000000000000_0000000000000000_0001010011011111_0010100001110110"; -- 0.08153012167070293
	pesos_i(19673) := b"0000000000000000_0000000000000000_0000101001111000_0101101110100111"; -- 0.04089901763906044
	pesos_i(19674) := b"1111111111111111_1111111111111111_1111000001001110_1010011111110010"; -- -0.061299804019686405
	pesos_i(19675) := b"1111111111111111_1111111111111111_1101110000001100_1100100001110101"; -- -0.14042994631996783
	pesos_i(19676) := b"0000000000000000_0000000000000000_0010010100110111_1001110010011110"; -- 0.14537981857748578
	pesos_i(19677) := b"1111111111111111_1111111111111111_1111011100011110_0111001100110111"; -- -0.0346916190305915
	pesos_i(19678) := b"0000000000000000_0000000000000000_0010010000000000_0111000000001111"; -- 0.14063167916818506
	pesos_i(19679) := b"0000000000000000_0000000000000000_0001001100000110_1001011100001010"; -- 0.07431930530076492
	pesos_i(19680) := b"0000000000000000_0000000000000000_0001111010010010_0111101101100011"; -- 0.11942263756146505
	pesos_i(19681) := b"1111111111111111_1111111111111111_1111100101100100_1011001111101100"; -- -0.025807146917632563
	pesos_i(19682) := b"1111111111111111_1111111111111111_1110101011001010_0001000001111011"; -- -0.08285424224236289
	pesos_i(19683) := b"0000000000000000_0000000000000000_0001100001111111_1001000001111011"; -- 0.095696477970399
	pesos_i(19684) := b"1111111111111111_1111111111111111_1110110101010101_1000010101011101"; -- -0.07291380376238804
	pesos_i(19685) := b"1111111111111111_1111111111111111_1101101100000010_0110011100010011"; -- -0.1444945887965005
	pesos_i(19686) := b"1111111111111111_1111111111111111_1101111001000110_0000011001111111"; -- -0.13174399754511706
	pesos_i(19687) := b"1111111111111111_1111111111111111_1111110011000011_0100000001111011"; -- -0.012645692859219269
	pesos_i(19688) := b"1111111111111111_1111111111111111_1110010001111011_0011111001001010"; -- -0.1074944561844888
	pesos_i(19689) := b"0000000000000000_0000000000000000_0000100001101000_0010001110111101"; -- 0.0328390442238059
	pesos_i(19690) := b"1111111111111111_1111111111111111_1110010011100110_0111011101001110"; -- -0.10585836747210638
	pesos_i(19691) := b"1111111111111111_1111111111111111_1110001011001100_1101111000001011"; -- -0.1140614721437697
	pesos_i(19692) := b"0000000000000000_0000000000000000_0000101100000001_1010010101011110"; -- 0.04299386546337727
	pesos_i(19693) := b"0000000000000000_0000000000000000_0001001101111001_1001110111110010"; -- 0.07607447764105567
	pesos_i(19694) := b"0000000000000000_0000000000000000_0010001000110011_0111100000111000"; -- 0.13359786376798266
	pesos_i(19695) := b"0000000000000000_0000000000000000_0001100110110000_0110101010010001"; -- 0.10034814875327842
	pesos_i(19696) := b"0000000000000000_0000000000000000_0000000111000000_1000001010000001"; -- 0.0068437161569123136
	pesos_i(19697) := b"1111111111111111_1111111111111111_1101111011110111_1111000111110111"; -- -0.1290291569561372
	pesos_i(19698) := b"0000000000000000_0000000000000000_0001000100000110_0111000001100101"; -- 0.06650450191438587
	pesos_i(19699) := b"0000000000000000_0000000000000000_0001001111110110_1100001010110101"; -- 0.07798401761732487
	pesos_i(19700) := b"1111111111111111_1111111111111111_1111110011111111_0101110000101100"; -- -0.011728514884932073
	pesos_i(19701) := b"0000000000000000_0000000000000000_0010010000011100_1001010011001110"; -- 0.14106111554019765
	pesos_i(19702) := b"1111111111111111_1111111111111111_1110011010111101_1111100001111100"; -- -0.09866377794241406
	pesos_i(19703) := b"0000000000000000_0000000000000000_0001001011000111_1001001100111100"; -- 0.07335777492193248
	pesos_i(19704) := b"1111111111111111_1111111111111111_1101111110000100_1100011110011111"; -- -0.12688019143390536
	pesos_i(19705) := b"1111111111111111_1111111111111111_1101101011010100_1011000010010011"; -- -0.14519211199510557
	pesos_i(19706) := b"1111111111111111_1111111111111111_1101110110111011_1100100100101001"; -- -0.13385336644301654
	pesos_i(19707) := b"0000000000000000_0000000000000000_0000010010010100_0110011100000101"; -- 0.017889441231241525
	pesos_i(19708) := b"1111111111111111_1111111111111111_1101100101110101_1010110001001010"; -- -0.15054820239858774
	pesos_i(19709) := b"0000000000000000_0000000000000000_0001011000000111_1101011011110111"; -- 0.08605712436963363
	pesos_i(19710) := b"1111111111111111_1111111111111111_1110101100110000_0010001110101100"; -- -0.08129670191578581
	pesos_i(19711) := b"0000000000000000_0000000000000000_0001011010110110_0101000100110110"; -- 0.0887194400538712
	pesos_i(19712) := b"1111111111111111_1111111111111111_1111011010000011_0011011001111000"; -- -0.03706035208924502
	pesos_i(19713) := b"1111111111111111_1111111111111111_1110010110011001_1100100001011101"; -- -0.10312221276868543
	pesos_i(19714) := b"1111111111111111_1111111111111111_1110101101111110_0000001101000100"; -- -0.08010844784063963
	pesos_i(19715) := b"1111111111111111_1111111111111111_1111000100010110_1101000101010111"; -- -0.058245578966695195
	pesos_i(19716) := b"0000000000000000_0000000000000000_0000000010001011_0111101010011000"; -- 0.0021282787424598735
	pesos_i(19717) := b"1111111111111111_1111111111111111_1111100100110110_1010110111111010"; -- -0.026509405593720958
	pesos_i(19718) := b"0000000000000000_0000000000000000_0000101111000100_0001100001001001"; -- 0.04596092015806477
	pesos_i(19719) := b"1111111111111111_1111111111111111_1110010011100111_0111110100111110"; -- -0.1058427546806174
	pesos_i(19720) := b"0000000000000000_0000000000000000_0001011110111110_0110100011000101"; -- 0.09274916461959276
	pesos_i(19721) := b"1111111111111111_1111111111111111_1111001101000000_0110100101100010"; -- -0.04979840623585591
	pesos_i(19722) := b"1111111111111111_1111111111111111_1111011101010101_0001011010001010"; -- -0.03385790953851184
	pesos_i(19723) := b"0000000000000000_0000000000000000_0010001110000010_1000011010001110"; -- 0.13871041262593392
	pesos_i(19724) := b"1111111111111111_1111111111111111_1101101110000011_1100011011011010"; -- -0.1425204962524636
	pesos_i(19725) := b"1111111111111111_1111111111111111_1111010110101100_0010110100000010"; -- -0.04034155553653289
	pesos_i(19726) := b"1111111111111111_1111111111111111_1110010010000110_0111001110000001"; -- -0.10732343765258462
	pesos_i(19727) := b"1111111111111111_1111111111111111_1110001111010110_1101100110100010"; -- -0.11000289720665658
	pesos_i(19728) := b"1111111111111111_1111111111111111_1111100110111101_0110100101011011"; -- -0.024453559219034922
	pesos_i(19729) := b"0000000000000000_0000000000000000_0000101001001001_1010001111011111"; -- 0.040186159117559635
	pesos_i(19730) := b"1111111111111111_1111111111111111_1101100000100110_1011011101000011"; -- -0.1556592428364903
	pesos_i(19731) := b"0000000000000000_0000000000000000_0001010110111000_0100110001111011"; -- 0.08484342578149859
	pesos_i(19732) := b"0000000000000000_0000000000000000_0001110111110010_1100110101111110"; -- 0.11698612518293681
	pesos_i(19733) := b"1111111111111111_1111111111111111_1111011010010001_1101001010010000"; -- -0.03683742513992154
	pesos_i(19734) := b"1111111111111111_1111111111111111_1110001000101001_0101101010010100"; -- -0.11655649085821262
	pesos_i(19735) := b"1111111111111111_1111111111111111_1110100101000011_1000101110000011"; -- -0.08881309549308831
	pesos_i(19736) := b"1111111111111111_1111111111111111_1110010001000101_1011001010011000"; -- -0.10831149854298543
	pesos_i(19737) := b"0000000000000000_0000000000000000_0001001100001011_0001101100101110"; -- 0.07438821679081785
	pesos_i(19738) := b"1111111111111111_1111111111111111_1111110101111100_0111001001000110"; -- -0.009819849032483513
	pesos_i(19739) := b"1111111111111111_1111111111111111_1110001100000101_1011110100001101"; -- -0.11319368786038682
	pesos_i(19740) := b"0000000000000000_0000000000000000_0001001001000100_0110001000100111"; -- 0.0713559479467842
	pesos_i(19741) := b"1111111111111111_1111111111111111_1111011101100010_1111101111010100"; -- -0.03364587857978416
	pesos_i(19742) := b"1111111111111111_1111111111111111_1110011101000011_0011110111001000"; -- -0.09663022866943241
	pesos_i(19743) := b"1111111111111111_1111111111111111_1110010110000001_1001110110111000"; -- -0.10349096534005638
	pesos_i(19744) := b"0000000000000000_0000000000000000_0010010010100011_1110101101001001"; -- 0.14312620675015225
	pesos_i(19745) := b"1111111111111111_1111111111111111_1110110111011101_1011000011110010"; -- -0.07083601085249738
	pesos_i(19746) := b"1111111111111111_1111111111111111_1110110101010011_1110001010011111"; -- -0.07293876273317423
	pesos_i(19747) := b"0000000000000000_0000000000000000_0000110001010101_0101100000000110"; -- 0.04817724364983503
	pesos_i(19748) := b"1111111111111111_1111111111111111_1111010101111101_0110111111111011"; -- -0.04105472670590248
	pesos_i(19749) := b"1111111111111111_1111111111111111_1101111110011111_1100011100101000"; -- -0.12646823197945484
	pesos_i(19750) := b"0000000000000000_0000000000000000_0001111101010100_0011011011010000"; -- 0.12237875542778215
	pesos_i(19751) := b"0000000000000000_0000000000000000_0010011010100010_1000101001011110"; -- 0.15091767106684612
	pesos_i(19752) := b"0000000000000000_0000000000000000_0001111110101111_1011001100010010"; -- 0.12377471147152841
	pesos_i(19753) := b"1111111111111111_1111111111111111_1110001011110011_1000011100001001"; -- -0.1134715654912206
	pesos_i(19754) := b"0000000000000000_0000000000000000_0000000011110001_0001100100111111"; -- 0.003678873054924719
	pesos_i(19755) := b"1111111111111111_1111111111111111_1101110110000011_1000101110101111"; -- -0.13471152277560294
	pesos_i(19756) := b"0000000000000000_0000000000000000_0010001001110000_0101110000001000"; -- 0.1345269699504076
	pesos_i(19757) := b"1111111111111111_1111111111111111_1111010010100011_1000101110000000"; -- -0.04437950252116685
	pesos_i(19758) := b"0000000000000000_0000000000000000_0001101100000101_1100101110010110"; -- 0.10555717868950971
	pesos_i(19759) := b"1111111111111111_1111111111111111_1111111110000011_0001011101000101"; -- -0.0019059616215805339
	pesos_i(19760) := b"0000000000000000_0000000000000000_0000110011001110_0001110100111000"; -- 0.05002005209094092
	pesos_i(19761) := b"1111111111111111_1111111111111111_1111110011100111_1111001010000011"; -- -0.01208576500023192
	pesos_i(19762) := b"1111111111111111_1111111111111111_1111000001000101_1111011011010001"; -- -0.06143243204861865
	pesos_i(19763) := b"1111111111111111_1111111111111111_1111100000000100_0111100101001100"; -- -0.03118173509202223
	pesos_i(19764) := b"1111111111111111_1111111111111111_1110011111001110_0011101010010100"; -- -0.09450944798329163
	pesos_i(19765) := b"1111111111111111_1111111111111111_1101111001010011_1011000011011110"; -- -0.1315354783773985
	pesos_i(19766) := b"0000000000000000_0000000000000000_0001000110100011_1101001011001110"; -- 0.06890599751403893
	pesos_i(19767) := b"0000000000000000_0000000000000000_0010001010100001_1110001001101101"; -- 0.13528266105496825
	pesos_i(19768) := b"1111111111111111_1111111111111111_1111001000010111_1101110101110001"; -- -0.054323348928928754
	pesos_i(19769) := b"0000000000000000_0000000000000000_0010010110000001_1111001100111111"; -- 0.14651413227642454
	pesos_i(19770) := b"0000000000000000_0000000000000000_0001100111111010_1101111010110110"; -- 0.10148422188754029
	pesos_i(19771) := b"0000000000000000_0000000000000000_0001000011100111_1001010000101101"; -- 0.06603361212573584
	pesos_i(19772) := b"0000000000000000_0000000000000000_0000000111110101_0101011001000111"; -- 0.007649795963418362
	pesos_i(19773) := b"1111111111111111_1111111111111111_1111011100101010_0011110111010111"; -- -0.034511694823670426
	pesos_i(19774) := b"1111111111111111_1111111111111111_1110011101001110_0001000111011000"; -- -0.09646500088642587
	pesos_i(19775) := b"0000000000000000_0000000000000000_0001000011010010_0001011000100011"; -- 0.06570566522575119
	pesos_i(19776) := b"1111111111111111_1111111111111111_1110010011011100_0010000010010100"; -- -0.10601612471051618
	pesos_i(19777) := b"0000000000000000_0000000000000000_0001101001011011_1100100011010100"; -- 0.10296302018185503
	pesos_i(19778) := b"1111111111111111_1111111111111111_1111101110001111_1101001101100110"; -- -0.01733664290021472
	pesos_i(19779) := b"0000000000000000_0000000000000000_0000100110111100_1111111001011011"; -- 0.038040063199023394
	pesos_i(19780) := b"1111111111111111_1111111111111111_1110010101001011_1110111001011111"; -- -0.10431013273922607
	pesos_i(19781) := b"1111111111111111_1111111111111111_1110110010011011_0110001001010010"; -- -0.0757540273446125
	pesos_i(19782) := b"1111111111111111_1111111111111111_1110101110100111_1001100011110101"; -- -0.07947391535967159
	pesos_i(19783) := b"1111111111111111_1111111111111111_1110101110111101_1010001000100001"; -- -0.07913767523849449
	pesos_i(19784) := b"0000000000000000_0000000000000000_0000000000001110_0100110110001010"; -- 0.0002182446799417032
	pesos_i(19785) := b"1111111111111111_1111111111111111_1111111110110001_1000011101001100"; -- -0.001197380105215468
	pesos_i(19786) := b"0000000000000000_0000000000000000_0001110000001110_1001111001101001"; -- 0.10959806514158504
	pesos_i(19787) := b"0000000000000000_0000000000000000_0000011110000100_0111000110101101"; -- 0.0293646857975206
	pesos_i(19788) := b"0000000000000000_0000000000000000_0000000100100111_1100001000001000"; -- 0.004512907854768011
	pesos_i(19789) := b"0000000000000000_0000000000000000_0010001001000000_0011101111111011"; -- 0.13379263765331895
	pesos_i(19790) := b"0000000000000000_0000000000000000_0001100111111010_0101010001110111"; -- 0.1014759817717246
	pesos_i(19791) := b"0000000000000000_0000000000000000_0001001100000001_1101101111101000"; -- 0.07424711613139734
	pesos_i(19792) := b"0000000000000000_0000000000000000_0000011111000111_1010000111010101"; -- 0.030389894938969098
	pesos_i(19793) := b"1111111111111111_1111111111111111_1110111110011010_0001011100000001"; -- -0.06405502536200898
	pesos_i(19794) := b"0000000000000000_0000000000000000_0000111100001001_0100011100010111"; -- 0.05873531643963836
	pesos_i(19795) := b"0000000000000000_0000000000000000_0000110100010010_0111011111010111"; -- 0.051063051293887794
	pesos_i(19796) := b"1111111111111111_1111111111111111_1111110010101011_0101000010000100"; -- -0.013010947898484657
	pesos_i(19797) := b"1111111111111111_1111111111111111_1111011110111001_0101101100100110"; -- -0.03232794106245163
	pesos_i(19798) := b"1111111111111111_1111111111111111_1110100100110010_0110110010001001"; -- -0.08907434144000519
	pesos_i(19799) := b"0000000000000000_0000000000000000_0001111010111111_1110100001010111"; -- 0.12011577717153725
	pesos_i(19800) := b"1111111111111111_1111111111111111_1111001011111100_1111011001111010"; -- -0.050827593973900125
	pesos_i(19801) := b"1111111111111111_1111111111111111_1101101001101011_1111110101011001"; -- -0.14678970883609532
	pesos_i(19802) := b"0000000000000000_0000000000000000_0010000000101101_1011110100111001"; -- 0.12569792405118307
	pesos_i(19803) := b"1111111111111111_1111111111111111_1110000010100100_1110100010000111"; -- -0.12248369881250434
	pesos_i(19804) := b"0000000000000000_0000000000000000_0000001111010111_0111100001100001"; -- 0.015006564838551924
	pesos_i(19805) := b"1111111111111111_1111111111111111_1110000010111001_1001011011001110"; -- -0.12216813541658042
	pesos_i(19806) := b"1111111111111111_1111111111111111_1111000011101100_0010011111000101"; -- -0.058896555234233955
	pesos_i(19807) := b"0000000000000000_0000000000000000_0001011000010111_1001111111111100"; -- 0.08629798792206478
	pesos_i(19808) := b"0000000000000000_0000000000000000_0010001011101000_0110001111001110"; -- 0.13635848782460464
	pesos_i(19809) := b"0000000000000000_0000000000000000_0001000011111110_0100101000001000"; -- 0.06638014494464944
	pesos_i(19810) := b"0000000000000000_0000000000000000_0000010011101000_0010001011110100"; -- 0.01916712252473495
	pesos_i(19811) := b"0000000000000000_0000000000000000_0010001011010110_1000100000011001"; -- 0.13608599298631385
	pesos_i(19812) := b"1111111111111111_1111111111111111_1110100001010000_1001011110101011"; -- -0.09252025676819632
	pesos_i(19813) := b"1111111111111111_1111111111111111_1101111001000011_1000011111110100"; -- -0.13178205771129814
	pesos_i(19814) := b"1111111111111111_1111111111111111_1111100010011010_1111100001010001"; -- -0.028885345696806966
	pesos_i(19815) := b"1111111111111111_1111111111111111_1111111110010111_0110110000001011"; -- -0.0015957328919002675
	pesos_i(19816) := b"1111111111111111_1111111111111111_1110100011110111_1010111111011010"; -- -0.08997059755843503
	pesos_i(19817) := b"0000000000000000_0000000000000000_0000100000111111_1111111101101011"; -- 0.03222652781914199
	pesos_i(19818) := b"1111111111111111_1111111111111111_1110001101101110_0001000001111001"; -- -0.11160180141338627
	pesos_i(19819) := b"1111111111111111_1111111111111111_1111100000001111_0110011101001100"; -- -0.031014961180232257
	pesos_i(19820) := b"0000000000000000_0000000000000000_0000101111000111_1010010000111011"; -- 0.04601503781256992
	pesos_i(19821) := b"0000000000000000_0000000000000000_0001101100000000_1100110001101111"; -- 0.1054809352165294
	pesos_i(19822) := b"1111111111111111_1111111111111111_1110000111110110_0101001100010010"; -- -0.11733513643191115
	pesos_i(19823) := b"0000000000000000_0000000000000000_0000100011111010_1011001111110101"; -- 0.035075423548638254
	pesos_i(19824) := b"1111111111111111_1111111111111111_1110100011101110_1000010110101010"; -- -0.09011044125820034
	pesos_i(19825) := b"1111111111111111_1111111111111111_1111000110100001_0100100100001011"; -- -0.056132731170193864
	pesos_i(19826) := b"0000000000000000_0000000000000000_0000100010100001_1010000111010111"; -- 0.03371631148857848
	pesos_i(19827) := b"1111111111111111_1111111111111111_1110000101010011_0010111101011101"; -- -0.11982444744366294
	pesos_i(19828) := b"1111111111111111_1111111111111111_1101100000111010_0010110100100011"; -- -0.1553622998032522
	pesos_i(19829) := b"0000000000000000_0000000000000000_0001010101101111_0010010010011100"; -- 0.08372715767277797
	pesos_i(19830) := b"1111111111111111_1111111111111111_1101111001100000_1010001001001000"; -- -0.13133798348852238
	pesos_i(19831) := b"0000000000000000_0000000000000000_0000100101111010_0110111101100101"; -- 0.03702446192683654
	pesos_i(19832) := b"0000000000000000_0000000000000000_0001001111100101_1111101110011010"; -- 0.07772800928880186
	pesos_i(19833) := b"0000000000000000_0000000000000000_0000101011111011_1011101001011010"; -- 0.042903563380042
	pesos_i(19834) := b"0000000000000000_0000000000000000_0000011101101011_1001101100000100"; -- 0.028985679965395195
	pesos_i(19835) := b"0000000000000000_0000000000000000_0010001011011100_0000001000111110"; -- 0.1361695673065099
	pesos_i(19836) := b"0000000000000000_0000000000000000_0000110000100000_1100011101111101"; -- 0.047375171695283144
	pesos_i(19837) := b"0000000000000000_0000000000000000_0001111111100011_1101011111011001"; -- 0.1245703607168472
	pesos_i(19838) := b"1111111111111111_1111111111111111_1111001010011011_1001010010110100"; -- -0.052313524209093513
	pesos_i(19839) := b"0000000000000000_0000000000000000_0000011000111001_0010000110010110"; -- 0.024309252867162727
	pesos_i(19840) := b"1111111111111111_1111111111111111_1110100011110100_0101101110110100"; -- -0.09002138942246056
	pesos_i(19841) := b"1111111111111111_1111111111111111_1111011000001110_0110110000101101"; -- -0.0388424291885149
	pesos_i(19842) := b"1111111111111111_1111111111111111_1110000101011100_0111011010100110"; -- -0.11968286951077205
	pesos_i(19843) := b"1111111111111111_1111111111111111_1111001011010001_0010101100001110"; -- -0.05149584690404889
	pesos_i(19844) := b"0000000000000000_0000000000000000_0010010110100101_1001110011000010"; -- 0.14705829378321075
	pesos_i(19845) := b"1111111111111111_1111111111111111_1111001011011001_1110001110001010"; -- -0.05136278031046295
	pesos_i(19846) := b"0000000000000000_0000000000000000_0000111010000001_0101111100101001"; -- 0.0566615557940164
	pesos_i(19847) := b"0000000000000000_0000000000000000_0001101110110101_1011100101001110"; -- 0.1082416358444861
	pesos_i(19848) := b"0000000000000000_0000000000000000_0001100001011110_1011101010000111"; -- 0.09519544396056015
	pesos_i(19849) := b"0000000000000000_0000000000000000_0000110110100101_1110010101011110"; -- 0.053312621634143686
	pesos_i(19850) := b"0000000000000000_0000000000000000_0001101001111110_1111010010000110"; -- 0.1034996820645012
	pesos_i(19851) := b"0000000000000000_0000000000000000_0000100010110010_0100101010011001"; -- 0.033970510927741525
	pesos_i(19852) := b"0000000000000000_0000000000000000_0010000010000001_0110101001010011"; -- 0.12697472128312462
	pesos_i(19853) := b"1111111111111111_1111111111111111_1101110010100001_0011011000000000"; -- -0.13816511635195908
	pesos_i(19854) := b"1111111111111111_1111111111111111_1110010010110001_1100101000111111"; -- -0.10666213941766073
	pesos_i(19855) := b"0000000000000000_0000000000000000_0001011010100111_0000111110010101"; -- 0.08848664645766544
	pesos_i(19856) := b"1111111111111111_1111111111111111_1111111000011000_0010100111000010"; -- -0.0074438002079169775
	pesos_i(19857) := b"1111111111111111_1111111111111111_1101101111010110_0000000011010100"; -- -0.14126581978328162
	pesos_i(19858) := b"1111111111111111_1111111111111111_1101100100101001_0010011010001110"; -- -0.15171584161389165
	pesos_i(19859) := b"0000000000000000_0000000000000000_0001111110110010_0011101101000100"; -- 0.12381334702100301
	pesos_i(19860) := b"0000000000000000_0000000000000000_0000010010001101_1100110000101000"; -- 0.017788657894803907
	pesos_i(19861) := b"1111111111111111_1111111111111111_1110111011010101_1001101111001111"; -- -0.06705309094237186
	pesos_i(19862) := b"1111111111111111_1111111111111111_1111111111001100_0011100101100011"; -- -0.0007900365710109145
	pesos_i(19863) := b"0000000000000000_0000000000000000_0010010000001111_0011110100100001"; -- 0.14085752551849004
	pesos_i(19864) := b"1111111111111111_1111111111111111_1111101101110011_0110110111110000"; -- -0.01776993647767509
	pesos_i(19865) := b"0000000000000000_0000000000000000_0001010011010011_1000111110111111"; -- 0.08135317232842951
	pesos_i(19866) := b"0000000000000000_0000000000000000_0000111101111110_1110110101000111"; -- 0.06053050016960181
	pesos_i(19867) := b"0000000000000000_0000000000000000_0000100001011000_0110100101000000"; -- 0.03259904675882667
	pesos_i(19868) := b"1111111111111111_1111111111111111_1111100001011101_0110001001000100"; -- -0.029825075430437324
	pesos_i(19869) := b"1111111111111111_1111111111111111_1111010011101000_0111111001100001"; -- -0.04332742827620958
	pesos_i(19870) := b"1111111111111111_1111111111111111_1101101110010111_1111011010111011"; -- -0.1422124666714996
	pesos_i(19871) := b"0000000000000000_0000000000000000_0001110111100000_1011100101100010"; -- 0.11671026837127328
	pesos_i(19872) := b"1111111111111111_1111111111111111_1111001010010010_0001111000001000"; -- -0.052457926904240774
	pesos_i(19873) := b"1111111111111111_1111111111111111_1111100110110010_1001010011111110"; -- -0.02461880500727615
	pesos_i(19874) := b"0000000000000000_0000000000000000_0010001000111111_1110111110111000"; -- 0.13378809199654734
	pesos_i(19875) := b"0000000000000000_0000000000000000_0000010111001100_0110110010010001"; -- 0.022650514047046055
	pesos_i(19876) := b"0000000000000000_0000000000000000_0000011001011010_1010100101000101"; -- 0.024820880240406993
	pesos_i(19877) := b"0000000000000000_0000000000000000_0001101111110010_0010100000101010"; -- 0.10916377081809628
	pesos_i(19878) := b"1111111111111111_1111111111111111_1111011011110100_1010101000101000"; -- -0.03532921332601842
	pesos_i(19879) := b"0000000000000000_0000000000000000_0001001010001010_1001001111100101"; -- 0.0724270281160487
	pesos_i(19880) := b"0000000000000000_0000000000000000_0001101101110000_1100111101001101"; -- 0.1071900904757616
	pesos_i(19881) := b"1111111111111111_1111111111111111_1111111001011010_1000111010010111"; -- -0.006430710002035024
	pesos_i(19882) := b"0000000000000000_0000000000000000_0001110100010000_1100000000000101"; -- 0.11353683576838582
	pesos_i(19883) := b"0000000000000000_0000000000000000_0000110001011110_0010100100010010"; -- 0.04831177414063391
	pesos_i(19884) := b"0000000000000000_0000000000000000_0000000010000100_0101111110101111"; -- 0.002019863386354599
	pesos_i(19885) := b"0000000000000000_0000000000000000_0001011011010110_0011001010101110"; -- 0.0892059016861187
	pesos_i(19886) := b"0000000000000000_0000000000000000_0001100011100011_1110111011000001"; -- 0.09722797601628877
	pesos_i(19887) := b"0000000000000000_0000000000000000_0001100010010110_1101100101101010"; -- 0.09605177723824668
	pesos_i(19888) := b"0000000000000000_0000000000000000_0001101000001100_0000100110010000"; -- 0.10174617546826606
	pesos_i(19889) := b"0000000000000000_0000000000000000_0001100100011100_1100100111011000"; -- 0.0980955270078449
	pesos_i(19890) := b"0000000000000000_0000000000000000_0001010110001111_0100010101001110"; -- 0.08421738772631664
	pesos_i(19891) := b"0000000000000000_0000000000000000_0000010110110110_0100000101011001"; -- 0.022312244620410326
	pesos_i(19892) := b"0000000000000000_0000000000000000_0001101001100011_1010001100110001"; -- 0.1030828470493096
	pesos_i(19893) := b"0000000000000000_0000000000000000_0001111111010111_1001100110011111"; -- 0.12438354610139674
	pesos_i(19894) := b"1111111111111111_1111111111111111_1111011110101111_1000100010011111"; -- -0.03247781864962376
	pesos_i(19895) := b"0000000000000000_0000000000000000_0000101001000010_0100010111011111"; -- 0.04007374469199289
	pesos_i(19896) := b"1111111111111111_1111111111111111_1110111101010011_1010011001000000"; -- -0.06512986114853789
	pesos_i(19897) := b"0000000000000000_0000000000000000_0001100110011101_1101001111100110"; -- 0.10006451000865575
	pesos_i(19898) := b"1111111111111111_1111111111111111_1111011001001110_1010010000010001"; -- -0.03786253530807794
	pesos_i(19899) := b"1111111111111111_1111111111111111_1110101111101101_1011001111110010"; -- -0.07840419135117233
	pesos_i(19900) := b"0000000000000000_0000000000000000_0001111111001010_1011011011001100"; -- 0.12418692097196393
	pesos_i(19901) := b"0000000000000000_0000000000000000_0010001101011101_1110011111001110"; -- 0.13815163392540034
	pesos_i(19902) := b"1111111111111111_1111111111111111_1110100000101001_1101011101111010"; -- -0.09311154627927822
	pesos_i(19903) := b"0000000000000000_0000000000000000_0000001111000110_0010100011001110"; -- 0.0147424223847767
	pesos_i(19904) := b"0000000000000000_0000000000000000_0000000111000011_1011000000100011"; -- 0.00689221245442572
	pesos_i(19905) := b"0000000000000000_0000000000000000_0001111011101000_1110111101100110"; -- 0.12074180836122479
	pesos_i(19906) := b"0000000000000000_0000000000000000_0010000101010111_1001111100001101"; -- 0.1302432448447539
	pesos_i(19907) := b"0000000000000000_0000000000000000_0010011001110001_1100111111000011"; -- 0.15017412678848113
	pesos_i(19908) := b"0000000000000000_0000000000000000_0010011001100010_0100110000010110"; -- 0.14993739647196205
	pesos_i(19909) := b"1111111111111111_1111111111111111_1111010111000100_0000001001010000"; -- -0.03997788950418939
	pesos_i(19910) := b"1111111111111111_1111111111111111_1101101100001101_0000001001001000"; -- -0.1443327498396678
	pesos_i(19911) := b"1111111111111111_1111111111111111_1110100101101000_1010001101011010"; -- -0.08824709937241262
	pesos_i(19912) := b"1111111111111111_1111111111111111_1111100100110110_0110001110111001"; -- -0.026513831481212786
	pesos_i(19913) := b"1111111111111111_1111111111111111_1110101111111111_0110111011101101"; -- -0.07813364699213371
	pesos_i(19914) := b"1111111111111111_1111111111111111_1110111100000110_0110110011111101"; -- -0.06630820097947196
	pesos_i(19915) := b"1111111111111111_1111111111111111_1111000011111011_0000101110001100"; -- -0.05866935573500086
	pesos_i(19916) := b"0000000000000000_0000000000000000_0001000111010101_1010001000110011"; -- 0.06966603978859724
	pesos_i(19917) := b"0000000000000000_0000000000000000_0001110000011101_1000000000001000"; -- 0.10982513615316429
	pesos_i(19918) := b"1111111111111111_1111111111111111_1101101110000001_0110111001101011"; -- -0.14255628477508372
	pesos_i(19919) := b"0000000000000000_0000000000000000_0010010011000001_1011110100000100"; -- 0.14358121251760597
	pesos_i(19920) := b"0000000000000000_0000000000000000_0010011000101110_1111010001001100"; -- 0.14915396556666066
	pesos_i(19921) := b"1111111111111111_1111111111111111_1111001010000000_0000100101000100"; -- -0.05273382273489137
	pesos_i(19922) := b"1111111111111111_1111111111111111_1110010100111010_0111101110110011"; -- -0.1045763671951948
	pesos_i(19923) := b"0000000000000000_0000000000000000_0000001010000101_0111111000011010"; -- 0.009849435257573869
	pesos_i(19924) := b"0000000000000000_0000000000000000_0001111011010001_1100110011000101"; -- 0.1203887921401788
	pesos_i(19925) := b"1111111111111111_1111111111111111_1110100110000110_1110010101001011"; -- -0.08778540532099033
	pesos_i(19926) := b"1111111111111111_1111111111111111_1110010110110000_0100111010001010"; -- -0.10277852193250883
	pesos_i(19927) := b"1111111111111111_1111111111111111_1111011110100000_0000111100000011"; -- -0.03271394886957225
	pesos_i(19928) := b"0000000000000000_0000000000000000_0001100011111111_0110001111100111"; -- 0.0976469458396979
	pesos_i(19929) := b"0000000000000000_0000000000000000_0001010011101100_1000110001011110"; -- 0.0817344407447217
	pesos_i(19930) := b"0000000000000000_0000000000000000_0000010100100101_0100101110100000"; -- 0.020100332830493135
	pesos_i(19931) := b"1111111111111111_1111111111111111_1110100101000101_1110101100110110"; -- -0.08877687396083106
	pesos_i(19932) := b"0000000000000000_0000000000000000_0000001101010000_1011111111110101"; -- 0.012950894744915812
	pesos_i(19933) := b"0000000000000000_0000000000000000_0001011000001011_0000111010101001"; -- 0.086106220401063
	pesos_i(19934) := b"1111111111111111_1111111111111111_1111000110010101_0110100000001011"; -- -0.056313988931755724
	pesos_i(19935) := b"0000000000000000_0000000000000000_0001100101110001_1001011101000011"; -- 0.09938950899136241
	pesos_i(19936) := b"1111111111111111_1111111111111111_1110000111111001_1000100101001101"; -- -0.11728612785760241
	pesos_i(19937) := b"0000000000000000_0000000000000000_0010001100111001_0010000111011001"; -- 0.13759051846896803
	pesos_i(19938) := b"1111111111111111_1111111111111111_1110111010101111_0101010011000001"; -- -0.06763716009086855
	pesos_i(19939) := b"0000000000000000_0000000000000000_0001001110011100_0010110100010110"; -- 0.0766018084675865
	pesos_i(19940) := b"0000000000000000_0000000000000000_0001101100110111_0011100101011111"; -- 0.10631140290888229
	pesos_i(19941) := b"0000000000000000_0000000000000000_0001100010010001_1001110000100100"; -- 0.09597183111754738
	pesos_i(19942) := b"1111111111111111_1111111111111111_1111001001001010_0101110100001100"; -- -0.05355280357083393
	pesos_i(19943) := b"1111111111111111_1111111111111111_1110110011010110_1001111100000010"; -- -0.07485014155639573
	pesos_i(19944) := b"0000000000000000_0000000000000000_0000101001111101_1101011011100000"; -- 0.04098265619576479
	pesos_i(19945) := b"0000000000000000_0000000000000000_0001101011011111_1100010001001110"; -- 0.10497691059590497
	pesos_i(19946) := b"0000000000000000_0000000000000000_0010011110110010_1111111101001101"; -- 0.1550750314719135
	pesos_i(19947) := b"0000000000000000_0000000000000000_0000100110001000_1111101001000110"; -- 0.03724636271456455
	pesos_i(19948) := b"0000000000000000_0000000000000000_0001111101010000_1110101000101001"; -- 0.12232841025423674
	pesos_i(19949) := b"1111111111111111_1111111111111111_1110111100011001_0010111011100101"; -- -0.06602198511893645
	pesos_i(19950) := b"0000000000000000_0000000000000000_0010010110100101_0111101100110100"; -- 0.1470562937839362
	pesos_i(19951) := b"0000000000000000_0000000000000000_0000010100011111_1010100010110000"; -- 0.02001432699216988
	pesos_i(19952) := b"0000000000000000_0000000000000000_0000110101100011_0001110110101010"; -- 0.05229363824168173
	pesos_i(19953) := b"1111111111111111_1111111111111111_1111111101011101_0110010110111010"; -- -0.002481119275230335
	pesos_i(19954) := b"1111111111111111_1111111111111111_1110101011111101_0111110111110111"; -- -0.08206951821351792
	pesos_i(19955) := b"1111111111111111_1111111111111111_1110011011010010_0001110111011001"; -- -0.09835637533779491
	pesos_i(19956) := b"1111111111111111_1111111111111111_1110110110011011_0011101001000001"; -- -0.07185016540150164
	pesos_i(19957) := b"1111111111111111_1111111111111111_1101111100110101_0001000111001100"; -- -0.12809647337619176
	pesos_i(19958) := b"1111111111111111_1111111111111111_1110101001010110_0010000111010110"; -- -0.08462322742038524
	pesos_i(19959) := b"0000000000000000_0000000000000000_0000010001001000_1011010110100110"; -- 0.016734459888057766
	pesos_i(19960) := b"0000000000000000_0000000000000000_0000111010111100_1000001001101101"; -- 0.05756392643823162
	pesos_i(19961) := b"0000000000000000_0000000000000000_0001110111100101_1111000010011110"; -- 0.11678985469194239
	pesos_i(19962) := b"1111111111111111_1111111111111111_1101110100011001_0001100110010001"; -- -0.1363357564803869
	pesos_i(19963) := b"0000000000000000_0000000000000000_0001101000000010_1010011111011000"; -- 0.1016030217454543
	pesos_i(19964) := b"0000000000000000_0000000000000000_0000000101001010_0111000000100000"; -- 0.005042083623542979
	pesos_i(19965) := b"1111111111111111_1111111111111111_1111101011001100_1001001001110101"; -- -0.0203159774746459
	pesos_i(19966) := b"0000000000000000_0000000000000000_0000100011100111_1110111100100100"; -- 0.03478903419121265
	pesos_i(19967) := b"0000000000000000_0000000000000000_0000011011100110_0000010111100111"; -- 0.026947373283562986
	pesos_i(19968) := b"1111111111111111_1111111111111111_1111101110001011_1010001110010010"; -- -0.0174005288023267
	pesos_i(19969) := b"0000000000000000_0000000000000000_0000000101110111_0110110010000100"; -- 0.005728513991830031
	pesos_i(19970) := b"0000000000000000_0000000000000000_0001010111101011_1011011001000010"; -- 0.08562792884716115
	pesos_i(19971) := b"0000000000000000_0000000000000000_0000001110111110_1001000110011111"; -- 0.014626599590955337
	pesos_i(19972) := b"0000000000000000_0000000000000000_0001111010110111_0101010011001111"; -- 0.11998491346902006
	pesos_i(19973) := b"1111111111111111_1111111111111111_1110101010010010_1111000001010000"; -- -0.08369539313842564
	pesos_i(19974) := b"1111111111111111_1111111111111111_1111111000010010_1011001011100101"; -- -0.007527178799901114
	pesos_i(19975) := b"1111111111111111_1111111111111111_1110010001111101_0100101000101110"; -- -0.10746323002828319
	pesos_i(19976) := b"1111111111111111_1111111111111111_1111001111000101_0110111000110100"; -- -0.04776869997126765
	pesos_i(19977) := b"1111111111111111_1111111111111111_1110101110101001_0001001011011010"; -- -0.07945139103695702
	pesos_i(19978) := b"0000000000000000_0000000000000000_0001110110001101_1010110000101100"; -- 0.11544300145382388
	pesos_i(19979) := b"1111111111111111_1111111111111111_1111011000110100_1100111111010011"; -- -0.03825665573597711
	pesos_i(19980) := b"0000000000000000_0000000000000000_0000001001001011_1010100110011001"; -- 0.008967017944056363
	pesos_i(19981) := b"0000000000000000_0000000000000000_0000001000100001_0010001001110010"; -- 0.00831809310822272
	pesos_i(19982) := b"0000000000000000_0000000000000000_0000110100010111_1110100101111001"; -- 0.05114611819297961
	pesos_i(19983) := b"0000000000000000_0000000000000000_0000000001001001_1000001100111000"; -- 0.0011217128225489196
	pesos_i(19984) := b"0000000000000000_0000000000000000_0000110110001011_0001001101001011"; -- 0.05290337160868775
	pesos_i(19985) := b"1111111111111111_1111111111111111_1110111010111111_1110101010000100"; -- -0.06738409295412114
	pesos_i(19986) := b"0000000000000000_0000000000000000_0001011101010101_1111110101101111"; -- 0.09115585278443432
	pesos_i(19987) := b"1111111111111111_1111111111111111_1110000000000111_0011010100001101"; -- -0.12489002642123945
	pesos_i(19988) := b"1111111111111111_1111111111111111_1110110101111100_1011110011010010"; -- -0.07231540559612643
	pesos_i(19989) := b"1111111111111111_1111111111111111_1111001110010111_0110011000000001"; -- -0.04847109284239153
	pesos_i(19990) := b"1111111111111111_1111111111111111_1110010001001111_0000111001101011"; -- -0.10816869619866025
	pesos_i(19991) := b"0000000000000000_0000000000000000_0000000011111111_0100111101011101"; -- 0.003895721669341989
	pesos_i(19992) := b"0000000000000000_0000000000000000_0001011010111101_0101101110101001"; -- 0.08882687457726299
	pesos_i(19993) := b"0000000000000000_0000000000000000_0001101000110010_1010111010100101"; -- 0.1023358491737942
	pesos_i(19994) := b"0000000000000000_0000000000000000_0010001111011111_0011101100101100"; -- 0.1401249869077219
	pesos_i(19995) := b"0000000000000000_0000000000000000_0000000000111110_0000001110100011"; -- 0.0009462615710233489
	pesos_i(19996) := b"1111111111111111_1111111111111111_1111110011101100_0011000000001110"; -- -0.012021061526719553
	pesos_i(19997) := b"1111111111111111_1111111111111111_1111000100110010_0110110101111111"; -- -0.05782428405077303
	pesos_i(19998) := b"0000000000000000_0000000000000000_0000011100111100_1010101100011101"; -- 0.028269476478986803
	pesos_i(19999) := b"1111111111111111_1111111111111111_1101110110111011_0010110110100001"; -- -0.13386263674823634
	pesos_i(20000) := b"0000000000000000_0000000000000000_0000001101011110_0011111011100101"; -- 0.013156825030402263
	pesos_i(20001) := b"0000000000000000_0000000000000000_0010001000011001_0100001001011001"; -- 0.13319792435481578
	pesos_i(20002) := b"0000000000000000_0000000000000000_0001001011100111_0011001110110010"; -- 0.07384036156774282
	pesos_i(20003) := b"0000000000000000_0000000000000000_0000010000000111_1110100110101101"; -- 0.015745739598692316
	pesos_i(20004) := b"1111111111111111_1111111111111111_1101100001011110_1000111111000000"; -- -0.15480710576228826
	pesos_i(20005) := b"1111111111111111_1111111111111111_1111010100100111_1110010001000100"; -- -0.04236005146047179
	pesos_i(20006) := b"0000000000000000_0000000000000000_0000011001111101_0111100110011111"; -- 0.025352097720029568
	pesos_i(20007) := b"1111111111111111_1111111111111111_1110001011001111_1011000010010000"; -- -0.11401840672022487
	pesos_i(20008) := b"1111111111111111_1111111111111111_1101111010110100_0101001000000010"; -- -0.1300610299574111
	pesos_i(20009) := b"0000000000000000_0000000000000000_0000111101001010_1011111110001001"; -- 0.0597343166856575
	pesos_i(20010) := b"0000000000000000_0000000000000000_0001110011010110_1110100000010000"; -- 0.11265421286935882
	pesos_i(20011) := b"1111111111111111_1111111111111111_1111100010001010_1100111011010000"; -- -0.029131960071433913
	pesos_i(20012) := b"0000000000000000_0000000000000000_0010010000101010_1111101000000110"; -- 0.14128077166055766
	pesos_i(20013) := b"1111111111111111_1111111111111111_1110010101001100_1111010001110100"; -- -0.10429451150317566
	pesos_i(20014) := b"0000000000000000_0000000000000000_0000001010000101_0011011110011100"; -- 0.009845233473010626
	pesos_i(20015) := b"0000000000000000_0000000000000000_0000010000101001_0100000111111100"; -- 0.016254543303294157
	pesos_i(20016) := b"1111111111111111_1111111111111111_1110001000010111_0011101101100110"; -- -0.11683300748885936
	pesos_i(20017) := b"1111111111111111_1111111111111111_1111101000101100_0010001110111111"; -- -0.022763982573172237
	pesos_i(20018) := b"1111111111111111_1111111111111111_1110110101100111_0110000011111001"; -- -0.07264131470031539
	pesos_i(20019) := b"1111111111111111_1111111111111111_1101100110110110_1000001011011000"; -- -0.14955885144994055
	pesos_i(20020) := b"0000000000000000_0000000000000000_0001001101100001_0101011000001000"; -- 0.07570398034284628
	pesos_i(20021) := b"1111111111111111_1111111111111111_1110010110101101_1000001001101111"; -- -0.10282120503759996
	pesos_i(20022) := b"0000000000000000_0000000000000000_0001100100100110_0010101100100000"; -- 0.09823865446267808
	pesos_i(20023) := b"1111111111111111_1111111111111111_1110001100011101_1000001101010110"; -- -0.11283091693850901
	pesos_i(20024) := b"0000000000000000_0000000000000000_0000001010111110_1010001101100111"; -- 0.010721409458324829
	pesos_i(20025) := b"0000000000000000_0000000000000000_0000110000010110_0010110100100001"; -- 0.04721338334244112
	pesos_i(20026) := b"1111111111111111_1111111111111111_1101101000101100_1101111100011001"; -- -0.14775281560141115
	pesos_i(20027) := b"0000000000000000_0000000000000000_0001000010110110_1101011001111010"; -- 0.06528988342393191
	pesos_i(20028) := b"1111111111111111_1111111111111111_1111000011110101_1000100001111110"; -- -0.058753461151709645
	pesos_i(20029) := b"1111111111111111_1111111111111111_1111111011000011_1110000010001010"; -- -0.004823652581244754
	pesos_i(20030) := b"1111111111111111_1111111111111111_1111000000000111_0001100100001100"; -- -0.06239169556395102
	pesos_i(20031) := b"1111111111111111_1111111111111111_1110100100010101_1110110010000101"; -- -0.08950921776659586
	pesos_i(20032) := b"1111111111111111_1111111111111111_1110001000011101_0101100111001000"; -- -0.11673964379498428
	pesos_i(20033) := b"0000000000000000_0000000000000000_0000110110010010_1100100110111110"; -- 0.05302105803364877
	pesos_i(20034) := b"1111111111111111_1111111111111111_1101101111000010_0111010000101100"; -- -0.14156412042492697
	pesos_i(20035) := b"0000000000000000_0000000000000000_0000011010011011_1101100111101100"; -- 0.02581560154076341
	pesos_i(20036) := b"0000000000000000_0000000000000000_0001010010001110_0110100011000000"; -- 0.08029799174098252
	pesos_i(20037) := b"1111111111111111_1111111111111111_1110001110101010_1001001010011000"; -- -0.11067851817831156
	pesos_i(20038) := b"1111111111111111_1111111111111111_1101100111111101_0000000011000111"; -- -0.14848323007768296
	pesos_i(20039) := b"0000000000000000_0000000000000000_0000000110111010_1110000010000011"; -- 0.006757766607337817
	pesos_i(20040) := b"0000000000000000_0000000000000000_0000001000010001_0001011010111101"; -- 0.008073254645793773
	pesos_i(20041) := b"1111111111111111_1111111111111111_1101110101010100_0110111111100001"; -- -0.1354303431944627
	pesos_i(20042) := b"1111111111111111_1111111111111111_1110100101110000_0110110110101000"; -- -0.0881282297179889
	pesos_i(20043) := b"1111111111111111_1111111111111111_1110011101101101_0101111100011011"; -- -0.09598737328892153
	pesos_i(20044) := b"1111111111111111_1111111111111111_1111001001010000_0001001010010100"; -- -0.05346568959175914
	pesos_i(20045) := b"1111111111111111_1111111111111111_1110100100110000_0111000011111011"; -- -0.08910459389430066
	pesos_i(20046) := b"0000000000000000_0000000000000000_0000011100001000_1101010100110110"; -- 0.027478528571642444
	pesos_i(20047) := b"0000000000000000_0000000000000000_0001101011010000_0000101011111000"; -- 0.10473698186526083
	pesos_i(20048) := b"1111111111111111_1111111111111111_1101011000111000_1101110010000001"; -- -0.16319486483532705
	pesos_i(20049) := b"1111111111111111_1111111111111111_1111011111000011_0011101010001110"; -- -0.03217729597622754
	pesos_i(20050) := b"0000000000000000_0000000000000000_0000011000010111_0010000010100101"; -- 0.023790397999050302
	pesos_i(20051) := b"0000000000000000_0000000000000000_0000010110001001_1011101110101110"; -- 0.021632890761989276
	pesos_i(20052) := b"0000000000000000_0000000000000000_0001110111001101_0100110111000011"; -- 0.11641393680607746
	pesos_i(20053) := b"1111111111111111_1111111111111111_1110111000101000_0001000011111110"; -- -0.06970113554171431
	pesos_i(20054) := b"0000000000000000_0000000000000000_0000110011011101_0001011101000010"; -- 0.05024857875391946
	pesos_i(20055) := b"1111111111111111_1111111111111111_1111111100011111_1101010111110011"; -- -0.003420475181624699
	pesos_i(20056) := b"0000000000000000_0000000000000000_0001111110100000_1011011101000100"; -- 0.1235460796991803
	pesos_i(20057) := b"0000000000000000_0000000000000000_0010001000011010_0110110101001011"; -- 0.1332157428212356
	pesos_i(20058) := b"0000000000000000_0000000000000000_0000001000111011_0011011001110001"; -- 0.00871601354148663
	pesos_i(20059) := b"1111111111111111_1111111111111111_1111001110111110_1101111100111100"; -- -0.04786877435916079
	pesos_i(20060) := b"1111111111111111_1111111111111111_1101110010110011_1011111010110100"; -- -0.1378823099320004
	pesos_i(20061) := b"1111111111111111_1111111111111111_1110101100001111_0001000110101000"; -- -0.08180131586745142
	pesos_i(20062) := b"1111111111111111_1111111111111111_1101110011100110_1000111011001001"; -- -0.1371069677670767
	pesos_i(20063) := b"1111111111111111_1111111111111111_1110011100010101_1011101101001100"; -- -0.09732465165026115
	pesos_i(20064) := b"1111111111111111_1111111111111111_1111011011011000_0111000111001110"; -- -0.035759818364979844
	pesos_i(20065) := b"0000000000000000_0000000000000000_0000000110000000_1111101000000000"; -- 0.005874276141906777
	pesos_i(20066) := b"1111111111111111_1111111111111111_1110011110101000_1000001100001111"; -- -0.0950849618087036
	pesos_i(20067) := b"0000000000000000_0000000000000000_0010000111011111_0000101001001000"; -- 0.13230957285275113
	pesos_i(20068) := b"1111111111111111_1111111111111111_1101101010001111_0001100001110101"; -- -0.14625403537528542
	pesos_i(20069) := b"0000000000000000_0000000000000000_0001000101101111_1100000110000110"; -- 0.0681115104302077
	pesos_i(20070) := b"1111111111111111_1111111111111111_1111001111001101_1111101000010010"; -- -0.04763829285402462
	pesos_i(20071) := b"0000000000000000_0000000000000000_0000111100100001_1111011101001011"; -- 0.059112029796787466
	pesos_i(20072) := b"1111111111111111_1111111111111111_1111010010001110_0011110010111101"; -- -0.04470463161585031
	pesos_i(20073) := b"1111111111111111_1111111111111111_1101111110110101_1101011001011011"; -- -0.12613163255133164
	pesos_i(20074) := b"1111111111111111_1111111111111111_1110000001011011_1010011011011011"; -- -0.12360150480752753
	pesos_i(20075) := b"1111111111111111_1111111111111111_1110100101100110_1100001100110100"; -- -0.08827571842265526
	pesos_i(20076) := b"1111111111111111_1111111111111111_1101111010000010_0111010011100000"; -- -0.13082189107319409
	pesos_i(20077) := b"0000000000000000_0000000000000000_0000000011001000_1000111011101011"; -- 0.003060276424858098
	pesos_i(20078) := b"0000000000000000_0000000000000000_0000110001000111_1011110001000011"; -- 0.04796959524546876
	pesos_i(20079) := b"0000000000000000_0000000000000000_0001111110100111_1110010011111000"; -- 0.12365561534215393
	pesos_i(20080) := b"0000000000000000_0000000000000000_0001000000101011_1000111011110000"; -- 0.06316464768910765
	pesos_i(20081) := b"1111111111111111_1111111111111111_1111001010001110_1101101101110000"; -- -0.05250767250408424
	pesos_i(20082) := b"1111111111111111_1111111111111111_1111101000110011_0001001010001010"; -- -0.022658196717245345
	pesos_i(20083) := b"1111111111111111_1111111111111111_1111101101101001_0001011111010001"; -- -0.017927657536093173
	pesos_i(20084) := b"0000000000000000_0000000000000000_0001111110000000_0001010001000001"; -- 0.12304808219432495
	pesos_i(20085) := b"0000000000000000_0000000000000000_0000010000110100_1110101010110010"; -- 0.01643244604218034
	pesos_i(20086) := b"1111111111111111_1111111111111111_1111001111011111_0101001100100011"; -- -0.047373584713594645
	pesos_i(20087) := b"1111111111111111_1111111111111111_1101111001001000_0000100000110100"; -- -0.13171337816250028
	pesos_i(20088) := b"0000000000000000_0000000000000000_0001100010101010_0111001011111001"; -- 0.09635084694775531
	pesos_i(20089) := b"1111111111111111_1111111111111111_1111000100101001_0000000011100000"; -- -0.057968087434151036
	pesos_i(20090) := b"1111111111111111_1111111111111111_1110011111111011_1010000101100001"; -- -0.09381667491058734
	pesos_i(20091) := b"0000000000000000_0000000000000000_0001000101111010_1011110100111011"; -- 0.0682791012775516
	pesos_i(20092) := b"1111111111111111_1111111111111111_1110100101110100_1111010110000101"; -- -0.08805909639476049
	pesos_i(20093) := b"0000000000000000_0000000000000000_0001000011000000_1111111001001111"; -- 0.06544484553568067
	pesos_i(20094) := b"1111111111111111_1111111111111111_1111111000111111_1011011111110010"; -- -0.006840232369064005
	pesos_i(20095) := b"1111111111111111_1111111111111111_1111001100110111_1101101011001100"; -- -0.049928975334695765
	pesos_i(20096) := b"0000000000000000_0000000000000000_0001000110100001_0110110011100100"; -- 0.06886940534192261
	pesos_i(20097) := b"0000000000000000_0000000000000000_0000001111111100_1010010101100001"; -- 0.015573822263584669
	pesos_i(20098) := b"0000000000000000_0000000000000000_0000010001111000_1101011011010101"; -- 0.017468859568737137
	pesos_i(20099) := b"0000000000000000_0000000000000000_0000100011110000_1111011011111000"; -- 0.034926829750096165
	pesos_i(20100) := b"1111111111111111_1111111111111111_1110001101011000_1101011101110000"; -- -0.11192563556852356
	pesos_i(20101) := b"1111111111111111_1111111111111111_1110000110110010_1100001011110111"; -- -0.11836606480179059
	pesos_i(20102) := b"1111111111111111_1111111111111111_1111001000111101_0000100110001100"; -- -0.05375614484843285
	pesos_i(20103) := b"0000000000000000_0000000000000000_0010001111110001_0111100000111111"; -- 0.1404032854172572
	pesos_i(20104) := b"1111111111111111_1111111111111111_1110110100110101_1111011010010101"; -- -0.07339533675436045
	pesos_i(20105) := b"1111111111111111_1111111111111111_1110110110111000_0110111100101011"; -- -0.07140450657828597
	pesos_i(20106) := b"0000000000000000_0000000000000000_0001001000111000_0110011110001001"; -- 0.07117316344013726
	pesos_i(20107) := b"1111111111111111_1111111111111111_1110000111011011_1011011000011111"; -- -0.11774121998180108
	pesos_i(20108) := b"1111111111111111_1111111111111111_1101110011011011_1010000001111011"; -- -0.13727375984969975
	pesos_i(20109) := b"1111111111111111_1111111111111111_1111101110110100_0110010001111111"; -- -0.01677867792938936
	pesos_i(20110) := b"1111111111111111_1111111111111111_1110010110000111_1110001110000001"; -- -0.10339525313147685
	pesos_i(20111) := b"1111111111111111_1111111111111111_1111110100100100_0101101110101110"; -- -0.011163969166527624
	pesos_i(20112) := b"0000000000000000_0000000000000000_0001011110111010_0101010111111110"; -- 0.09268701026811962
	pesos_i(20113) := b"0000000000000000_0000000000000000_0001011011011111_1010111000110001"; -- 0.08935059256534814
	pesos_i(20114) := b"1111111111111111_1111111111111111_1111001100101101_1101010110011100"; -- -0.05008187241345333
	pesos_i(20115) := b"1111111111111111_1111111111111111_1111001101111100_1110101110110010"; -- -0.04887511153110056
	pesos_i(20116) := b"1111111111111111_1111111111111111_1110101111001100_0100000110010001"; -- -0.07891454890133118
	pesos_i(20117) := b"0000000000000000_0000000000000000_0001010010110111_1000111101111000"; -- 0.08092590974796907
	pesos_i(20118) := b"0000000000000000_0000000000000000_0000010111011110_0000000000111010"; -- 0.022918714698200678
	pesos_i(20119) := b"0000000000000000_0000000000000000_0000000010001100_0110111011001111"; -- 0.002142835161597093
	pesos_i(20120) := b"0000000000000000_0000000000000000_0000101100100001_0010010101111111"; -- 0.043474524887946155
	pesos_i(20121) := b"1111111111111111_1111111111111111_1110111111000110_0011110111010001"; -- -0.06338132519356547
	pesos_i(20122) := b"1111111111111111_1111111111111111_1111111001011010_1000110011000010"; -- -0.006430819178178409
	pesos_i(20123) := b"0000000000000000_0000000000000000_0010000111110011_1000000110011101"; -- 0.13262186118594024
	pesos_i(20124) := b"0000000000000000_0000000000000000_0000001100001011_0110100001100100"; -- 0.011892818891088975
	pesos_i(20125) := b"1111111111111111_1111111111111111_1110000111110111_1011101101101101"; -- -0.11731365766483513
	pesos_i(20126) := b"1111111111111111_1111111111111111_1110101000011100_1000110101000011"; -- -0.08550183397977147
	pesos_i(20127) := b"1111111111111111_1111111111111111_1111101000000110_0001010011100011"; -- -0.023344702415945513
	pesos_i(20128) := b"0000000000000000_0000000000000000_0000000000111110_1110111110000000"; -- 0.0009603202573450769
	pesos_i(20129) := b"1111111111111111_1111111111111111_1110111111100011_1001110011100101"; -- -0.06293315319670642
	pesos_i(20130) := b"1111111111111111_1111111111111111_1110111110111111_0000100011101110"; -- -0.06349128900196722
	pesos_i(20131) := b"0000000000000000_0000000000000000_0001001100111100_0011011111111011"; -- 0.07513761415207618
	pesos_i(20132) := b"1111111111111111_1111111111111111_1111001001010110_0001100001011010"; -- -0.05337379271773901
	pesos_i(20133) := b"1111111111111111_1111111111111111_1111110101100011_1110011111010011"; -- -0.010194311984229308
	pesos_i(20134) := b"0000000000000000_0000000000000000_0001110100100011_0111000001101100"; -- 0.11382200852819344
	pesos_i(20135) := b"1111111111111111_1111111111111111_1111010101011000_0010100010000101"; -- -0.04162356144725114
	pesos_i(20136) := b"0000000000000000_0000000000000000_0001110100110101_0000101100010101"; -- 0.1140906262461795
	pesos_i(20137) := b"0000000000000000_0000000000000000_0000011000001011_0000111110101010"; -- 0.02360628043206355
	pesos_i(20138) := b"1111111111111111_1111111111111111_1101110011010000_0110101001101111"; -- -0.13744482803343086
	pesos_i(20139) := b"0000000000000000_0000000000000000_0001010111111001_0110111011000100"; -- 0.08583729070804848
	pesos_i(20140) := b"1111111111111111_1111111111111111_1110111110011101_0000101000111100"; -- -0.06401001009858802
	pesos_i(20141) := b"1111111111111111_1111111111111111_1110111001111110_0100111011000010"; -- -0.06838519825727862
	pesos_i(20142) := b"1111111111111111_1111111111111111_1101111101100000_0001010000101000"; -- -0.12744020482197174
	pesos_i(20143) := b"0000000000000000_0000000000000000_0000011010001010_1010011110101001"; -- 0.02555320626563298
	pesos_i(20144) := b"0000000000000000_0000000000000000_0001110001111000_1101110101011110"; -- 0.11121924928400566
	pesos_i(20145) := b"0000000000000000_0000000000000000_0000000000000011_0100100010101011"; -- 5.010781495157338e-05
	pesos_i(20146) := b"1111111111111111_1111111111111111_1101100110000110_1001010100100001"; -- -0.15029018340559525
	pesos_i(20147) := b"0000000000000000_0000000000000000_0000101011001100_1111100110100101"; -- 0.04219017293924512
	pesos_i(20148) := b"0000000000000000_0000000000000000_0000100111001010_1101001001011100"; -- 0.03825106382100142
	pesos_i(20149) := b"1111111111111111_1111111111111111_1111000110011111_0001100000101011"; -- -0.056166161910290294
	pesos_i(20150) := b"1111111111111111_1111111111111111_1110001110011101_1110001000110010"; -- -0.11087213793912098
	pesos_i(20151) := b"0000000000000000_0000000000000000_0010000100110110_1000101011101001"; -- 0.12973850421769398
	pesos_i(20152) := b"1111111111111111_1111111111111111_1111011110011101_1001110111101110"; -- -0.032751206785952246
	pesos_i(20153) := b"0000000000000000_0000000000000000_0001001010110111_1111000100011000"; -- 0.07311922861925686
	pesos_i(20154) := b"1111111111111111_1111111111111111_1101111100001111_0101100111010110"; -- -0.12867201357366817
	pesos_i(20155) := b"0000000000000000_0000000000000000_0000111010000011_1101000110100100"; -- 0.05669889691235472
	pesos_i(20156) := b"0000000000000000_0000000000000000_0000011011110111_0101111000010000"; -- 0.027212027510968535
	pesos_i(20157) := b"1111111111111111_1111111111111111_1101101011101001_1111110011111010"; -- -0.14486712348400016
	pesos_i(20158) := b"1111111111111111_1111111111111111_1110000101000011_0010100110100111"; -- -0.12006892848494685
	pesos_i(20159) := b"0000000000000000_0000000000000000_0010001110010000_1010011011010110"; -- 0.13892595975464106
	pesos_i(20160) := b"1111111111111111_1111111111111111_1110111000000001_1111100110101011"; -- -0.07028235974007913
	pesos_i(20161) := b"1111111111111111_1111111111111111_1111110101101100_1111100101100111"; -- -0.010055935266107553
	pesos_i(20162) := b"0000000000000000_0000000000000000_0000111111010011_0001010110000001"; -- 0.06181463623773669
	pesos_i(20163) := b"1111111111111111_1111111111111111_1111101011000011_1110000111101001"; -- -0.020448570878991327
	pesos_i(20164) := b"0000000000000000_0000000000000000_0001111100011000_0000101110110101"; -- 0.12146065881457399
	pesos_i(20165) := b"1111111111111111_1111111111111111_1111110100111100_0011111110101001"; -- -0.010799428160781737
	pesos_i(20166) := b"1111111111111111_1111111111111111_1110000011100001_1100010000111011"; -- -0.12155507611574969
	pesos_i(20167) := b"1111111111111111_1111111111111111_1101100011101101_0001011110010010"; -- -0.15263226215754755
	pesos_i(20168) := b"0000000000000000_0000000000000000_0000000000101111_0100101100111100"; -- 0.0007216474305519055
	pesos_i(20169) := b"0000000000000000_0000000000000000_0001101110111101_0111110101000100"; -- 0.10836012748223313
	pesos_i(20170) := b"0000000000000000_0000000000000000_0000001111010011_1001111110111101"; -- 0.014947875549505399
	pesos_i(20171) := b"1111111111111111_1111111111111111_1111010010100010_1010100011100100"; -- -0.04439300942454158
	pesos_i(20172) := b"1111111111111111_1111111111111111_1101110111101101_0100011001111011"; -- -0.1330982160443943
	pesos_i(20173) := b"1111111111111111_1111111111111111_1110100101100100_0111000000100000"; -- -0.08831118786047165
	pesos_i(20174) := b"0000000000000000_0000000000000000_0010010011100110_1001011011010101"; -- 0.1441435116652928
	pesos_i(20175) := b"0000000000000000_0000000000000000_0010000110010110_0000110101111011"; -- 0.13119587190098145
	pesos_i(20176) := b"0000000000000000_0000000000000000_0001000111010110_1011111000111001"; -- 0.06968296901855177
	pesos_i(20177) := b"1111111111111111_1111111111111111_1110100001101101_0111011010010101"; -- -0.09207972396003195
	pesos_i(20178) := b"1111111111111111_1111111111111111_1110001100110010_1110110110110010"; -- -0.11250414291211229
	pesos_i(20179) := b"0000000000000000_0000000000000000_0001000100000010_0010001001100010"; -- 0.06643881706774325
	pesos_i(20180) := b"0000000000000000_0000000000000000_0000101110000111_0110000111000100"; -- 0.04503451371577707
	pesos_i(20181) := b"0000000000000000_0000000000000000_0000111011011101_0101000001111110"; -- 0.058064489983274806
	pesos_i(20182) := b"0000000000000000_0000000000000000_0010011101000100_0111100110101011"; -- 0.15338859974870053
	pesos_i(20183) := b"1111111111111111_1111111111111111_1101111001101001_1001100001011101"; -- -0.13120124562114158
	pesos_i(20184) := b"0000000000000000_0000000000000000_0001010011101011_1100011010011110"; -- 0.08172265382857222
	pesos_i(20185) := b"1111111111111111_1111111111111111_1111110111001101_0001111100100110"; -- -0.008588841662739866
	pesos_i(20186) := b"0000000000000000_0000000000000000_0000111001111011_1111110111111100"; -- 0.05657946969986106
	pesos_i(20187) := b"1111111111111111_1111111111111111_1110010011101111_1000011110010111"; -- -0.10572006764153874
	pesos_i(20188) := b"0000000000000000_0000000000000000_0000000011010000_1101110101000000"; -- 0.0031870155382438315
	pesos_i(20189) := b"1111111111111111_1111111111111111_1111111110100110_0001001100000100"; -- -0.0013721575912229679
	pesos_i(20190) := b"0000000000000000_0000000000000000_0000011110001111_0001000111111010"; -- 0.029526828326519483
	pesos_i(20191) := b"0000000000000000_0000000000000000_0000100011001011_0011000101001100"; -- 0.03435047251873554
	pesos_i(20192) := b"1111111111111111_1111111111111111_1110011000111011_0110001110010010"; -- -0.10065629670282107
	pesos_i(20193) := b"0000000000000000_0000000000000000_0001101110000111_0010010000100100"; -- 0.10753084069869576
	pesos_i(20194) := b"1111111111111111_1111111111111111_1111110110000100_1011011010010011"; -- -0.009693707568525542
	pesos_i(20195) := b"0000000000000000_0000000000000000_0001011001111000_1010111111010000"; -- 0.08777903383117766
	pesos_i(20196) := b"0000000000000000_0000000000000000_0000100111110011_1000101010000000"; -- 0.03887239098444208
	pesos_i(20197) := b"1111111111111111_1111111111111111_1110000111010110_1001110111010111"; -- -0.1178189611947811
	pesos_i(20198) := b"0000000000000000_0000000000000000_0000101000100110_1011111111011000"; -- 0.039653768688917033
	pesos_i(20199) := b"1111111111111111_1111111111111111_1111011100010101_0101110010100100"; -- -0.03483029360319738
	pesos_i(20200) := b"1111111111111111_1111111111111111_1110001111101010_1000111110011000"; -- -0.10970213455709152
	pesos_i(20201) := b"0000000000000000_0000000000000000_0010000100111111_1101110001110111"; -- 0.1298806944248077
	pesos_i(20202) := b"0000000000000000_0000000000000000_0000010010101001_0000110110101011"; -- 0.01820455013375877
	pesos_i(20203) := b"0000000000000000_0000000000000000_0000100100100111_1011010001100101"; -- 0.035762095224211025
	pesos_i(20204) := b"1111111111111111_1111111111111111_1111010101010101_1110001011101100"; -- -0.041658227328158076
	pesos_i(20205) := b"1111111111111111_1111111111111111_1111010010110010_0110001101000111"; -- -0.0441530181548185
	pesos_i(20206) := b"1111111111111111_1111111111111111_1110111111110000_0111010101110101"; -- -0.06273713964238387
	pesos_i(20207) := b"1111111111111111_1111111111111111_1111011001010100_0100101001010101"; -- -0.03777633124543209
	pesos_i(20208) := b"1111111111111111_1111111111111111_1110010111001111_1101111101100001"; -- -0.10229686621493178
	pesos_i(20209) := b"1111111111111111_1111111111111111_1111000011100000_0111100000000000"; -- -0.059074878740023914
	pesos_i(20210) := b"1111111111111111_1111111111111111_1111100010111100_0100110001011001"; -- -0.028376796874736068
	pesos_i(20211) := b"1111111111111111_1111111111111111_1110001011110111_1111101000000001"; -- -0.11340367763645041
	pesos_i(20212) := b"0000000000000000_0000000000000000_0000000001111111_1001111110011101"; -- 0.0019473798826597733
	pesos_i(20213) := b"0000000000000000_0000000000000000_0010010000100101_0101011001010001"; -- 0.1411947201028736
	pesos_i(20214) := b"0000000000000000_0000000000000000_0010001000111010_1101100110010010"; -- 0.13371047794902205
	pesos_i(20215) := b"1111111111111111_1111111111111111_1110100011110001_0011100011101011"; -- -0.09006923927494474
	pesos_i(20216) := b"0000000000000000_0000000000000000_0000101100100111_0011000001010111"; -- 0.0435667239600088
	pesos_i(20217) := b"1111111111111111_1111111111111111_1110000000111111_0000010011101110"; -- -0.12403840236071673
	pesos_i(20218) := b"0000000000000000_0000000000000000_0001010011100101_0001101000011111"; -- 0.0816208195436167
	pesos_i(20219) := b"0000000000000000_0000000000000000_0001111100111110_0011011001110101"; -- 0.12204304077309382
	pesos_i(20220) := b"1111111111111111_1111111111111111_1111110001010101_1101000110101000"; -- -0.014315506466487124
	pesos_i(20221) := b"1111111111111111_1111111111111111_1101011111100111_0100001001010111"; -- -0.15662751557880877
	pesos_i(20222) := b"1111111111111111_1111111111111111_1110001011010101_1101111111011010"; -- -0.11392403542829041
	pesos_i(20223) := b"0000000000000000_0000000000000000_0000101011000111_0001100101011000"; -- 0.04210050953106362
	pesos_i(20224) := b"1111111111111111_1111111111111111_1110101100011011_0111110011011010"; -- -0.08161182092917478
	pesos_i(20225) := b"1111111111111111_1111111111111111_1110110001001010_1101111000101100"; -- -0.07698260704238108
	pesos_i(20226) := b"1111111111111111_1111111111111111_1111100010000001_0000111111001110"; -- -0.029280674269705025
	pesos_i(20227) := b"1111111111111111_1111111111111111_1101101111110111_1010001100100001"; -- -0.14075260589385521
	pesos_i(20228) := b"0000000000000000_0000000000000000_0001100010000110_1010101011100101"; -- 0.09580486387303663
	pesos_i(20229) := b"0000000000000000_0000000000000000_0000100100101001_1111110000000100"; -- 0.03579688161749781
	pesos_i(20230) := b"0000000000000000_0000000000000000_0000101111000001_0111111111101011"; -- 0.045921320801542924
	pesos_i(20231) := b"0000000000000000_0000000000000000_0001010110011001_0111011100010100"; -- 0.08437294237854694
	pesos_i(20232) := b"1111111111111111_1111111111111111_1110011000011101_0000111010001101"; -- -0.10111912775126497
	pesos_i(20233) := b"0000000000000000_0000000000000000_0001001011101011_1110101000011101"; -- 0.07391226970420212
	pesos_i(20234) := b"1111111111111111_1111111111111111_1110101010010011_0101001101110010"; -- -0.08368948430632991
	pesos_i(20235) := b"0000000000000000_0000000000000000_0000101001001110_0100011010111010"; -- 0.04025690124711701
	pesos_i(20236) := b"1111111111111111_1111111111111111_1101101101000000_0111101101011101"; -- -0.14354733456028348
	pesos_i(20237) := b"1111111111111111_1111111111111111_1110001111010101_1011010000111111"; -- -0.11002038448305829
	pesos_i(20238) := b"1111111111111111_1111111111111111_1111001100001010_1011101110011110"; -- -0.050617479199186584
	pesos_i(20239) := b"0000000000000000_0000000000000000_0000100000001010_0001111010110010"; -- 0.0314044173591509
	pesos_i(20240) := b"1111111111111111_1111111111111111_1111000100001011_0111100110001001"; -- -0.058418659181610134
	pesos_i(20241) := b"0000000000000000_0000000000000000_0010000011111011_1001110111111010"; -- 0.1288393722665427
	pesos_i(20242) := b"0000000000000000_0000000000000000_0010001011000010_0100000010100001"; -- 0.1357765572827261
	pesos_i(20243) := b"0000000000000000_0000000000000000_0000000100100000_1110100101110101"; -- 0.004408446413532316
	pesos_i(20244) := b"1111111111111111_1111111111111111_1110101011010111_1111101100101100"; -- -0.08264188927658773
	pesos_i(20245) := b"0000000000000000_0000000000000000_0000000111110100_0101011010011000"; -- 0.0076345559788908645
	pesos_i(20246) := b"0000000000000000_0000000000000000_0001101011010110_0101110000100010"; -- 0.10483337235446334
	pesos_i(20247) := b"0000000000000000_0000000000000000_0010011010010100_1100010111010100"; -- 0.15070759216217824
	pesos_i(20248) := b"0000000000000000_0000000000000000_0010000001100001_0100000110011010"; -- 0.12648401258892777
	pesos_i(20249) := b"0000000000000000_0000000000000000_0001110000001010_0100101110010001"; -- 0.10953209189955407
	pesos_i(20250) := b"1111111111111111_1111111111111111_1101101001100110_1011110011001010"; -- -0.1468698507901532
	pesos_i(20251) := b"1111111111111111_1111111111111111_1110110100101111_0000011011101101"; -- -0.07350117403786519
	pesos_i(20252) := b"0000000000000000_0000000000000000_0001100101110010_0011010111111011"; -- 0.09939896933552489
	pesos_i(20253) := b"1111111111111111_1111111111111111_1110100000101001_1110001111100001"; -- -0.09311080703411563
	pesos_i(20254) := b"0000000000000000_0000000000000000_0001011001100101_0001001011000010"; -- 0.08747975585355112
	pesos_i(20255) := b"1111111111111111_1111111111111111_1110111111100100_0110000101110010"; -- -0.0629214379959892
	pesos_i(20256) := b"1111111111111111_1111111111111111_1101111110000100_1000110010001001"; -- -0.12688371320120548
	pesos_i(20257) := b"1111111111111111_1111111111111111_1111100011100111_1001100111100001"; -- -0.02771604782723275
	pesos_i(20258) := b"1111111111111111_1111111111111111_1101101000010001_0111011110100010"; -- -0.14817096998108126
	pesos_i(20259) := b"1111111111111111_1111111111111111_1110011011101001_0111101101101010"; -- -0.09799984619681071
	pesos_i(20260) := b"0000000000000000_0000000000000000_0000010101111010_1000101011111100"; -- 0.021401106494171453
	pesos_i(20261) := b"1111111111111111_1111111111111111_1110101110001101_0000100010101110"; -- -0.07987924342494863
	pesos_i(20262) := b"0000000000000000_0000000000000000_0001001001110010_0000101011000010"; -- 0.07205264328136679
	pesos_i(20263) := b"0000000000000000_0000000000000000_0000101000011001_1111010100000000"; -- 0.039458572858703286
	pesos_i(20264) := b"1111111111111111_1111111111111111_1111100110001100_0111100001101001"; -- -0.025200342626269457
	pesos_i(20265) := b"1111111111111111_1111111111111111_1110110110010100_0100101110101010"; -- -0.07195593925386104
	pesos_i(20266) := b"0000000000000000_0000000000000000_0001100001111000_0001101110001111"; -- 0.09558269741208308
	pesos_i(20267) := b"0000000000000000_0000000000000000_0000111100001101_0000001010010111"; -- 0.05879226861815848
	pesos_i(20268) := b"0000000000000000_0000000000000000_0001101110110110_1100111100111100"; -- 0.1082582016489192
	pesos_i(20269) := b"1111111111111111_1111111111111111_1110000101001110_0001011000100000"; -- -0.11990224564097945
	pesos_i(20270) := b"1111111111111111_1111111111111111_1110100001100010_1110101000001011"; -- -0.09224068867286407
	pesos_i(20271) := b"0000000000000000_0000000000000000_0000011101000000_1111010000110000"; -- 0.028334867100913062
	pesos_i(20272) := b"0000000000000000_0000000000000000_0001011101001001_1011010101000010"; -- 0.09096844547462943
	pesos_i(20273) := b"0000000000000000_0000000000000000_0000101011111110_0010101010010101"; -- 0.04294077041175182
	pesos_i(20274) := b"1111111111111111_1111111111111111_1111100001100101_0010101111110001"; -- -0.029706243099309488
	pesos_i(20275) := b"1111111111111111_1111111111111111_1111100111110110_0000001110001001"; -- -0.023589877082466914
	pesos_i(20276) := b"1111111111111111_1111111111111111_1111111000011010_0010101001100001"; -- -0.007413245511080772
	pesos_i(20277) := b"0000000000000000_0000000000000000_0000000110101000_0000010000001011"; -- 0.006469967595734354
	pesos_i(20278) := b"0000000000000000_0000000000000000_0010010110110101_0101011000100011"; -- 0.14729822506890852
	pesos_i(20279) := b"1111111111111111_1111111111111111_1110001110111111_1111000001101011"; -- -0.11035249115676375
	pesos_i(20280) := b"0000000000000000_0000000000000000_0001000011000100_0101110011100111"; -- 0.0654962600994216
	pesos_i(20281) := b"1111111111111111_1111111111111111_1110110111101110_0001000101101010"; -- -0.07058612016302622
	pesos_i(20282) := b"1111111111111111_1111111111111111_1111010100001110_0100010001101101"; -- -0.04275104857303798
	pesos_i(20283) := b"1111111111111111_1111111111111111_1110001011110101_1100011110100011"; -- -0.11343719733741914
	pesos_i(20284) := b"0000000000000000_0000000000000000_0000110001000101_0011111011010110"; -- 0.0479316018718186
	pesos_i(20285) := b"0000000000000000_0000000000000000_0000100111011111_0011111001110111"; -- 0.03856268304093804
	pesos_i(20286) := b"1111111111111111_1111111111111111_1111110110101011_1011100000100100"; -- -0.009098521371483754
	pesos_i(20287) := b"1111111111111111_1111111111111111_1110000001101111_0001001111110010"; -- -0.12330508566405912
	pesos_i(20288) := b"1111111111111111_1111111111111111_1110001001010010_0100111110011110"; -- -0.11593153370308958
	pesos_i(20289) := b"1111111111111111_1111111111111111_1111101111100100_1000101011010100"; -- -0.016043971265515378
	pesos_i(20290) := b"0000000000000000_0000000000000000_0001110000110100_0101111111110000"; -- 0.11017417530236782
	pesos_i(20291) := b"1111111111111111_1111111111111111_1111111101101011_0011101100011111"; -- -0.0022700356312331284
	pesos_i(20292) := b"1111111111111111_1111111111111111_1110101100000001_1111111010100101"; -- -0.08200081318464764
	pesos_i(20293) := b"1111111111111111_1111111111111111_1110101111011111_0010110001101100"; -- -0.07862589231617854
	pesos_i(20294) := b"0000000000000000_0000000000000000_0010000111000000_1111101101000000"; -- 0.1318509130954257
	pesos_i(20295) := b"0000000000000000_0000000000000000_0000000010001000_0011000111000000"; -- 0.0020781606175199387
	pesos_i(20296) := b"0000000000000000_0000000000000000_0000011101100001_0111001111101111"; -- 0.028830762677574843
	pesos_i(20297) := b"0000000000000000_0000000000000000_0010001110110011_0100111000010011"; -- 0.13945472694050956
	pesos_i(20298) := b"1111111111111111_1111111111111111_1110110001011000_1111101000001010"; -- -0.07676732299149737
	pesos_i(20299) := b"1111111111111111_1111111111111111_1111100001001001_1001111100010101"; -- -0.03012662641325412
	pesos_i(20300) := b"0000000000000000_0000000000000000_0001111010110010_1100011001010111"; -- 0.11991538642492451
	pesos_i(20301) := b"0000000000000000_0000000000000000_0000010001011011_0011010101110010"; -- 0.017016735425811287
	pesos_i(20302) := b"1111111111111111_1111111111111111_1110010111111100_1011111010101011"; -- -0.10161217044323534
	pesos_i(20303) := b"0000000000000000_0000000000000000_0001001011101111_0110100111001111"; -- 0.07396565729767059
	pesos_i(20304) := b"1111111111111111_1111111111111111_1110110110011110_1001011000000011"; -- -0.07179892002799036
	pesos_i(20305) := b"1111111111111111_1111111111111111_1111101011111100_0000010100101110"; -- -0.01959197634380737
	pesos_i(20306) := b"1111111111111111_1111111111111111_1110011110101001_0110111000110110"; -- -0.09507094548915952
	pesos_i(20307) := b"1111111111111111_1111111111111111_1110011101000011_0110110010101110"; -- -0.0966274333406839
	pesos_i(20308) := b"0000000000000000_0000000000000000_0000000011110101_1101111100101011"; -- 0.0037517051180724955
	pesos_i(20309) := b"1111111111111111_1111111111111111_1110001000000001_1011000100000010"; -- -0.1171616907658463
	pesos_i(20310) := b"0000000000000000_0000000000000000_0010000001011111_0101000100110101"; -- 0.12645442519299127
	pesos_i(20311) := b"1111111111111111_1111111111111111_1110101000000001_1011110110010101"; -- -0.08591094114189803
	pesos_i(20312) := b"0000000000000000_0000000000000000_0001001111010111_0011001000010101"; -- 0.07750237486121142
	pesos_i(20313) := b"0000000000000000_0000000000000000_0001001100101011_0101110010101111"; -- 0.07488040237545734
	pesos_i(20314) := b"0000000000000000_0000000000000000_0001111010101111_1110111101101111"; -- 0.11987205944781346
	pesos_i(20315) := b"1111111111111111_1111111111111111_1111000101010100_0110111001010101"; -- -0.05730543545559714
	pesos_i(20316) := b"0000000000000000_0000000000000000_0000110001001011_1100001001011001"; -- 0.048030993300094034
	pesos_i(20317) := b"1111111111111111_1111111111111111_1110101010000000_0001110011100100"; -- -0.08398265293036178
	pesos_i(20318) := b"0000000000000000_0000000000000000_0001100000100100_1110010101001010"; -- 0.09431298301001269
	pesos_i(20319) := b"0000000000000000_0000000000000000_0000110010111011_1000101101101100"; -- 0.04973670374239343
	pesos_i(20320) := b"1111111111111111_1111111111111111_1101101101101101_0101001111101011"; -- -0.1428630400076909
	pesos_i(20321) := b"1111111111111111_1111111111111111_1111101000000100_1100100000111001"; -- -0.02336453073230121
	pesos_i(20322) := b"1111111111111111_1111111111111111_1111001011000111_0010000101111001"; -- -0.05164900591202729
	pesos_i(20323) := b"0000000000000000_0000000000000000_0001111111011010_0111111100011101"; -- 0.12442774249451174
	pesos_i(20324) := b"0000000000000000_0000000000000000_0000001101110011_0011010000011001"; -- 0.013476616093681658
	pesos_i(20325) := b"0000000000000000_0000000000000000_0001010100011100_0000001110110011"; -- 0.08245871668976013
	pesos_i(20326) := b"0000000000000000_0000000000000000_0000000110101110_0010001100000111"; -- 0.006563367107688978
	pesos_i(20327) := b"1111111111111111_1111111111111111_1110110001101101_1010111000011111"; -- -0.07645141366164417
	pesos_i(20328) := b"1111111111111111_1111111111111111_1110010111001101_0010100011011110"; -- -0.10233826231633772
	pesos_i(20329) := b"1111111111111111_1111111111111111_1101100110010000_0110010111000101"; -- -0.15014041832477362
	pesos_i(20330) := b"1111111111111111_1111111111111111_1110111010101101_1010000001000011"; -- -0.06766317716269353
	pesos_i(20331) := b"1111111111111111_1111111111111111_1101101111101110_1000001011000110"; -- -0.14089186341653165
	pesos_i(20332) := b"1111111111111111_1111111111111111_1111100110011001_1111111001010100"; -- -0.02499399620028827
	pesos_i(20333) := b"1111111111111111_1111111111111111_1111101101111011_1011000011001011"; -- -0.017643881327965787
	pesos_i(20334) := b"1111111111111111_1111111111111111_1110101000101100_0001000110000010"; -- -0.08526506982695951
	pesos_i(20335) := b"0000000000000000_0000000000000000_0000111101001001_0011001110101001"; -- 0.05971072070926271
	pesos_i(20336) := b"1111111111111111_1111111111111111_1110111010110101_1010101011101010"; -- -0.06754047194311275
	pesos_i(20337) := b"0000000000000000_0000000000000000_0010000010101000_0000010010000001"; -- 0.12756374498828923
	pesos_i(20338) := b"1111111111111111_1111111111111111_1110010011000011_0000111000000000"; -- -0.10639870155557977
	pesos_i(20339) := b"0000000000000000_0000000000000000_0010001100101010_1011001000101001"; -- 0.13737023839338816
	pesos_i(20340) := b"1111111111111111_1111111111111111_1111101101111000_0001000011111010"; -- -0.01769918339576111
	pesos_i(20341) := b"0000000000000000_0000000000000000_0000110011000101_0011010011011010"; -- 0.04988413168780921
	pesos_i(20342) := b"1111111111111111_1111111111111111_1110101100010110_0100010010011110"; -- -0.08169146669541077
	pesos_i(20343) := b"0000000000000000_0000000000000000_0010000100010000_1111101000011111"; -- 0.1291652989124422
	pesos_i(20344) := b"0000000000000000_0000000000000000_0000000101100110_1101111011100110"; -- 0.005475932261352494
	pesos_i(20345) := b"0000000000000000_0000000000000000_0000010000110101_1011001110000011"; -- 0.016444415581718982
	pesos_i(20346) := b"0000000000000000_0000000000000000_0010001110100010_1100111000100010"; -- 0.13920296031766402
	pesos_i(20347) := b"1111111111111111_1111111111111111_1111010001001011_0001000100001000"; -- -0.04572957575069213
	pesos_i(20348) := b"1111111111111111_1111111111111111_1111101001001100_1001000000110101"; -- -0.022269236553835593
	pesos_i(20349) := b"0000000000000000_0000000000000000_0010010100111000_0110110111101010"; -- 0.1453922936783422
	pesos_i(20350) := b"1111111111111111_1111111111111111_1111000011111010_0110010000101110"; -- -0.05867933147063881
	pesos_i(20351) := b"1111111111111111_1111111111111111_1111001011111011_0010010101111101"; -- -0.050855309542460814
	pesos_i(20352) := b"0000000000000000_0000000000000000_0001000100010100_0001001110011001"; -- 0.06671259391273322
	pesos_i(20353) := b"0000000000000000_0000000000000000_0000100010001010_0111011011111010"; -- 0.033362804370120375
	pesos_i(20354) := b"1111111111111111_1111111111111111_1101110000111111_1010000100001011"; -- -0.13965409742792656
	pesos_i(20355) := b"0000000000000000_0000000000000000_0001001110110110_1010110100101100"; -- 0.07700617137089441
	pesos_i(20356) := b"1111111111111111_1111111111111111_1101101111000111_1001000111101100"; -- -0.14148605329582395
	pesos_i(20357) := b"0000000000000000_0000000000000000_0001010001110100_0100110011110110"; -- 0.07989960664721195
	pesos_i(20358) := b"1111111111111111_1111111111111111_1110011001010101_1010011000000110"; -- -0.10025560720005533
	pesos_i(20359) := b"0000000000000000_0000000000000000_0010001010000001_1011101101101000"; -- 0.13479205411298012
	pesos_i(20360) := b"0000000000000000_0000000000000000_0001010111000010_0011011110001011"; -- 0.08499476571203976
	pesos_i(20361) := b"0000000000000000_0000000000000000_0001100000010111_0110010011001100"; -- 0.0941069600889547
	pesos_i(20362) := b"0000000000000000_0000000000000000_0010100101101010_1010000010110010"; -- 0.1617832598262784
	pesos_i(20363) := b"0000000000000000_0000000000000000_0000000001011011_1110001111111110"; -- 0.0014021391364374264
	pesos_i(20364) := b"0000000000000000_0000000000000000_0000111001011111_1101001001100010"; -- 0.05614962466147938
	pesos_i(20365) := b"0000000000000000_0000000000000000_0001111011111110_0001011011111100"; -- 0.12106460246222403
	pesos_i(20366) := b"0000000000000000_0000000000000000_0000010110110101_0010010100010110"; -- 0.02229530138198838
	pesos_i(20367) := b"1111111111111111_1111111111111111_1110100001011101_0001001111110101"; -- -0.09232974302128086
	pesos_i(20368) := b"1111111111111111_1111111111111111_1110111110100000_1101111000010111"; -- -0.06395160606062625
	pesos_i(20369) := b"0000000000000000_0000000000000000_0001100010010101_0001110000100100"; -- 0.0960252369985053
	pesos_i(20370) := b"0000000000000000_0000000000000000_0001100100001110_1111110011001010"; -- 0.09788494033711415
	pesos_i(20371) := b"0000000000000000_0000000000000000_0001010000101000_1101100101110010"; -- 0.07874831224710116
	pesos_i(20372) := b"1111111111111111_1111111111111111_1111001110001011_1111110101010001"; -- -0.04864517939395011
	pesos_i(20373) := b"0000000000000000_0000000000000000_0001100111100111_0100111010000101"; -- 0.10118571050107456
	pesos_i(20374) := b"0000000000000000_0000000000000000_0000000010011011_0100001001000010"; -- 0.0023690616141178677
	pesos_i(20375) := b"1111111111111111_1111111111111111_1111010111010000_0100010011101011"; -- -0.03979081406922316
	pesos_i(20376) := b"1111111111111111_1111111111111111_1101111001001101_0111000110101101"; -- -0.1316307975753662
	pesos_i(20377) := b"0000000000000000_0000000000000000_0000101100001010_1000001000010100"; -- 0.04312909118116993
	pesos_i(20378) := b"0000000000000000_0000000000000000_0010010101010101_0100001110000100"; -- 0.1458322713379676
	pesos_i(20379) := b"1111111111111111_1111111111111111_1111011000011000_0010000110101011"; -- -0.038694282254231625
	pesos_i(20380) := b"1111111111111111_1111111111111111_1101111111000110_1101011000110001"; -- -0.12587224292487106
	pesos_i(20381) := b"1111111111111111_1111111111111111_1110000101001101_0110100100110001"; -- -0.11991255329682038
	pesos_i(20382) := b"0000000000000000_0000000000000000_0000101110000011_1001010001010110"; -- 0.04497649281357962
	pesos_i(20383) := b"1111111111111111_1111111111111111_1110001101001011_0011101001100100"; -- -0.11213336036481146
	pesos_i(20384) := b"1111111111111111_1111111111111111_1111100000000101_0001101111110011"; -- -0.03117204010228964
	pesos_i(20385) := b"1111111111111111_1111111111111111_1111111011010010_1101010100011110"; -- -0.004595451537950708
	pesos_i(20386) := b"0000000000000000_0000000000000000_0000010101110100_1100110001010001"; -- 0.021313447737822077
	pesos_i(20387) := b"1111111111111111_1111111111111111_1101011111011001_0101110010100100"; -- -0.1568395710285335
	pesos_i(20388) := b"1111111111111111_1111111111111111_1110011100000010_0111111100000000"; -- -0.09761816271805754
	pesos_i(20389) := b"1111111111111111_1111111111111111_1111011001100111_1100001110111001"; -- -0.0374791787450478
	pesos_i(20390) := b"1111111111111111_1111111111111111_1110000010110011_0010100001010100"; -- -0.12226627307090987
	pesos_i(20391) := b"1111111111111111_1111111111111111_1110000011000010_0110011100001010"; -- -0.12203365326513739
	pesos_i(20392) := b"1111111111111111_1111111111111111_1110010111101011_0011100001000000"; -- -0.10187958186437637
	pesos_i(20393) := b"0000000000000000_0000000000000000_0001110010101110_0111110100011010"; -- 0.11203748591472087
	pesos_i(20394) := b"0000000000000000_0000000000000000_0000000010101111_1101010011001011"; -- 0.002682971581984489
	pesos_i(20395) := b"1111111111111111_1111111111111111_1101111010010001_1101111100011100"; -- -0.13058667719311046
	pesos_i(20396) := b"0000000000000000_0000000000000000_0000101101110111_1101101101011110"; -- 0.04479762110934836
	pesos_i(20397) := b"1111111111111111_1111111111111111_1111101100111110_0100001010010110"; -- -0.018581236262395783
	pesos_i(20398) := b"1111111111111111_1111111111111111_1111100010101001_1110001100111110"; -- -0.02865772006772085
	pesos_i(20399) := b"0000000000000000_0000000000000000_0000010111000000_1101101111110010"; -- 0.022474047316592624
	pesos_i(20400) := b"0000000000000000_0000000000000000_0001100101101001_1010010011001111"; -- 0.09926824617915446
	pesos_i(20401) := b"1111111111111111_1111111111111111_1111010101000111_1011010001000000"; -- -0.041874632211126105
	pesos_i(20402) := b"0000000000000000_0000000000000000_0000010010000110_1101010111001010"; -- 0.017682420442612038
	pesos_i(20403) := b"1111111111111111_1111111111111111_1111100111100101_1101001001101100"; -- -0.02383694523703622
	pesos_i(20404) := b"1111111111111111_1111111111111111_1110110110011110_0100111111111000"; -- -0.07180309488452578
	pesos_i(20405) := b"0000000000000000_0000000000000000_0000101001000111_1001100011011010"; -- 0.04015498469350299
	pesos_i(20406) := b"1111111111111111_1111111111111111_1101111111001001_0010110101001101"; -- -0.12583653319544713
	pesos_i(20407) := b"1111111111111111_1111111111111111_1111101100110010_1011010010110000"; -- -0.018757540842023534
	pesos_i(20408) := b"1111111111111111_1111111111111111_1110100011010110_0110011101010100"; -- -0.0904784602239121
	pesos_i(20409) := b"0000000000000000_0000000000000000_0000110000111011_0100001100100001"; -- 0.04777926975745326
	pesos_i(20410) := b"0000000000000000_0000000000000000_0001001001110111_0011110111101011"; -- 0.07213198651772826
	pesos_i(20411) := b"1111111111111111_1111111111111111_1111110011000001_1000000101101111"; -- -0.012672338878277957
	pesos_i(20412) := b"1111111111111111_1111111111111111_1101101100111010_1111001101000001"; -- -0.14363174113214394
	pesos_i(20413) := b"1111111111111111_1111111111111111_1101100011111100_0111111001001111"; -- -0.152397256491812
	pesos_i(20414) := b"1111111111111111_1111111111111111_1111001100110000_0100111110110000"; -- -0.05004407844441958
	pesos_i(20415) := b"0000000000000000_0000000000000000_0000111000101010_0011100100101010"; -- 0.055331776430968496
	pesos_i(20416) := b"0000000000000000_0000000000000000_0001000001101010_1010010010001011"; -- 0.06412723926890512
	pesos_i(20417) := b"1111111111111111_1111111111111111_1111000000101000_1101010110110101"; -- -0.06187691040363837
	pesos_i(20418) := b"0000000000000000_0000000000000000_0000110101000101_0011011101001001"; -- 0.051837401671854556
	pesos_i(20419) := b"1111111111111111_1111111111111111_1111001001011000_1101100111100001"; -- -0.053331739854486256
	pesos_i(20420) := b"1111111111111111_1111111111111111_1101110010001001_0110001000100010"; -- -0.13852869679128568
	pesos_i(20421) := b"0000000000000000_0000000000000000_0001001100000100_0000001000100010"; -- 0.07427991223015509
	pesos_i(20422) := b"1111111111111111_1111111111111111_1111000010000111_0010010011011100"; -- -0.060437866396264604
	pesos_i(20423) := b"1111111111111111_1111111111111111_1111010001101001_1101110001100110"; -- -0.04525969046393436
	pesos_i(20424) := b"1111111111111111_1111111111111111_1110110000000100_1111100011001110"; -- -0.07804913494693959
	pesos_i(20425) := b"1111111111111111_1111111111111111_1111111001101110_0100010101111001"; -- -0.006129892230854289
	pesos_i(20426) := b"1111111111111111_1111111111111111_1111011110111111_1111010000111000"; -- -0.03222726466549863
	pesos_i(20427) := b"0000000000000000_0000000000000000_0010000110000110_1001001011101111"; -- 0.1309596855472731
	pesos_i(20428) := b"1111111111111111_1111111111111111_1111000100101101_0111011110110110"; -- -0.05789996927928896
	pesos_i(20429) := b"1111111111111111_1111111111111111_1110010110011010_1011111110011011"; -- -0.10310747580091592
	pesos_i(20430) := b"1111111111111111_1111111111111111_1111010010111111_1001000101010100"; -- -0.04395190913719
	pesos_i(20431) := b"0000000000000000_0000000000000000_0001110101111101_0001011110001101"; -- 0.11519000247749557
	pesos_i(20432) := b"1111111111111111_1111111111111111_1111010011001111_0010101011011011"; -- -0.043713876190450356
	pesos_i(20433) := b"0000000000000000_0000000000000000_0001011010111101_0101000110001110"; -- 0.08882627208487813
	pesos_i(20434) := b"0000000000000000_0000000000000000_0001111101000010_0010000110110101"; -- 0.12210283910744077
	pesos_i(20435) := b"0000000000000000_0000000000000000_0001010001000000_0101100001010100"; -- 0.07910682726572905
	pesos_i(20436) := b"0000000000000000_0000000000000000_0001010000110011_0100011110111110"; -- 0.07890747440220876
	pesos_i(20437) := b"1111111111111111_1111111111111111_1101110100111010_1001100110100111"; -- -0.1358245817565094
	pesos_i(20438) := b"0000000000000000_0000000000000000_0001001111000101_0011011110101010"; -- 0.07722804924871467
	pesos_i(20439) := b"1111111111111111_1111111111111111_1101111100011111_0010010111010001"; -- -0.12843097350778201
	pesos_i(20440) := b"1111111111111111_1111111111111111_1110111111001100_0100011011101001"; -- -0.06328923045345913
	pesos_i(20441) := b"1111111111111111_1111111111111111_1110011100001000_0101110101001100"; -- -0.09752861874055829
	pesos_i(20442) := b"0000000000000000_0000000000000000_0000000101000011_1001110100100111"; -- 0.004937955830497676
	pesos_i(20443) := b"1111111111111111_1111111111111111_1110001011110011_1011111100001010"; -- -0.11346822734357803
	pesos_i(20444) := b"1111111111111111_1111111111111111_1111001100111010_1100101011010011"; -- -0.04988415087025359
	pesos_i(20445) := b"1111111111111111_1111111111111111_1110110011110100_1011011111000001"; -- -0.07439090278830965
	pesos_i(20446) := b"0000000000000000_0000000000000000_0001011000111101_1010001001011000"; -- 0.08687796261975458
	pesos_i(20447) := b"1111111111111111_1111111111111111_1110111100110111_1110101101101100"; -- -0.06555298437500931
	pesos_i(20448) := b"0000000000000000_0000000000000000_0000100000110000_0111000011001011"; -- 0.03198914490127707
	pesos_i(20449) := b"1111111111111111_1111111111111111_1110110000101011_0110100100101110"; -- -0.07746260293227379
	pesos_i(20450) := b"1111111111111111_1111111111111111_1101110111101101_0010010100111100"; -- -0.13310019758342076
	pesos_i(20451) := b"0000000000000000_0000000000000000_0001001010001111_1000110100001001"; -- 0.07250291309936324
	pesos_i(20452) := b"1111111111111111_1111111111111111_1110101101111011_0110100111001100"; -- -0.0801481130398459
	pesos_i(20453) := b"0000000000000000_0000000000000000_0001111110101001_0001011100100010"; -- 0.12367386427517175
	pesos_i(20454) := b"1111111111111111_1111111111111111_1111001000100101_1100011101011100"; -- -0.05411104199869368
	pesos_i(20455) := b"0000000000000000_0000000000000000_0000100110000111_1101100010000100"; -- 0.037229091876368615
	pesos_i(20456) := b"1111111111111111_1111111111111111_1110110110101100_0111000111000110"; -- -0.07158745682175212
	pesos_i(20457) := b"0000000000000000_0000000000000000_0010001011010011_0111000101100110"; -- 0.13603886364514733
	pesos_i(20458) := b"1111111111111111_1111111111111111_1101100110011100_1000100001101111"; -- -0.14995524673826297
	pesos_i(20459) := b"0000000000000000_0000000000000000_0000011110111001_0010110111110100"; -- 0.030169365105748504
	pesos_i(20460) := b"1111111111111111_1111111111111111_1110101111101000_1100010000110011"; -- -0.07847951646582368
	pesos_i(20461) := b"0000000000000000_0000000000000000_0001010000001101_1101011001001010"; -- 0.07833613680542817
	pesos_i(20462) := b"0000000000000000_0000000000000000_0000010001001011_1101010010000011"; -- 0.016782075756145026
	pesos_i(20463) := b"0000000000000000_0000000000000000_0001001011010111_0011011110000111"; -- 0.07359644930746276
	pesos_i(20464) := b"0000000000000000_0000000000000000_0001000000001110_1110111011000110"; -- 0.06272785511200323
	pesos_i(20465) := b"0000000000000000_0000000000000000_0000111101010000_0011000110110000"; -- 0.059817414730959126
	pesos_i(20466) := b"0000000000000000_0000000000000000_0001111010000000_1010000001100011"; -- 0.11915018484368758
	pesos_i(20467) := b"0000000000000000_0000000000000000_0001010011111111_1110011101100001"; -- 0.08202978246151928
	pesos_i(20468) := b"0000000000000000_0000000000000000_0001101100001111_0111111000101000"; -- 0.10570515131537174
	pesos_i(20469) := b"0000000000000000_0000000000000000_0001111110000111_1101011100000011"; -- 0.12316650222498667
	pesos_i(20470) := b"1111111111111111_1111111111111111_1111010100001011_1011011111001011"; -- -0.04278994834013898
	pesos_i(20471) := b"0000000000000000_0000000000000000_0001011111110100_0001101001101101"; -- 0.09356846957909705
	pesos_i(20472) := b"1111111111111111_1111111111111111_1111110111010101_0100010100001110"; -- -0.008464511835967204
	pesos_i(20473) := b"0000000000000000_0000000000000000_0001111111100110_1010010010110100"; -- 0.12461308845120134
	pesos_i(20474) := b"0000000000000000_0000000000000000_0000011110110011_0001011110110000"; -- 0.03007648510903135
	pesos_i(20475) := b"0000000000000000_0000000000000000_0010001000011011_1110101000111101"; -- 0.1332384489926526
	pesos_i(20476) := b"0000000000000000_0000000000000000_0001111110101101_0111110110110100"; -- 0.12374101297856115
	pesos_i(20477) := b"1111111111111111_1111111111111111_1111111110001111_1111100001110111"; -- -0.0017094334377258423
	pesos_i(20478) := b"1111111111111111_1111111111111111_1111000101111110_1011101010111100"; -- -0.05666001224965539
	pesos_i(20479) := b"1111111111111111_1111111111111111_1111001111101110_0100110100001000"; -- -0.04714506686633845
	pesos_i(20480) := b"0000000000000000_0000000000000000_0000101000001101_1010000000000110"; -- 0.03927040235318779
	pesos_i(20481) := b"0000000000000000_0000000000000000_0000000111100111_0110111011100010"; -- 0.007437639425348867
	pesos_i(20482) := b"1111111111111111_1111111111111111_1111101100000011_0111000111010000"; -- -0.019478689920582975
	pesos_i(20483) := b"1111111111111111_1111111111111111_1101101101001100_1000000000100111"; -- -0.14336394360261395
	pesos_i(20484) := b"1111111111111111_1111111111111111_1110001000010110_0010110100010110"; -- -0.11684911927494605
	pesos_i(20485) := b"0000000000000000_0000000000000000_0010000101100110_1101000111000010"; -- 0.13047514899392781
	pesos_i(20486) := b"1111111111111111_1111111111111111_1111011111000011_0001110100111001"; -- -0.03217904439800744
	pesos_i(20487) := b"1111111111111111_1111111111111111_1111110000111000_0011111100100011"; -- -0.0147667444981123
	pesos_i(20488) := b"1111111111111111_1111111111111111_1111110011100101_0000111001010111"; -- -0.012129882660769017
	pesos_i(20489) := b"0000000000000000_0000000000000000_0001101010010010_1000110001010110"; -- 0.10379864784534143
	pesos_i(20490) := b"0000000000000000_0000000000000000_0000110010010101_0001100101111010"; -- 0.04915007797698185
	pesos_i(20491) := b"0000000000000000_0000000000000000_0010001000110010_0000110010000010"; -- 0.13357618487725884
	pesos_i(20492) := b"1111111111111111_1111111111111111_1111001101011000_1110101111000011"; -- -0.04942442412591154
	pesos_i(20493) := b"1111111111111111_1111111111111111_1110010010110011_1101111101110110"; -- -0.10663035752644269
	pesos_i(20494) := b"1111111111111111_1111111111111111_1110110011000101_0110101010000111"; -- -0.07511266897148611
	pesos_i(20495) := b"0000000000000000_0000000000000000_0000110001000111_1010010010011001"; -- 0.04796818486397235
	pesos_i(20496) := b"1111111111111111_1111111111111111_1110111101010011_1110001100001010"; -- -0.06512623796509616
	pesos_i(20497) := b"1111111111111111_1111111111111111_1110010010110010_0110100100111100"; -- -0.10665266314711837
	pesos_i(20498) := b"0000000000000000_0000000000000000_0000011010111011_1001000010000100"; -- 0.02629950729350152
	pesos_i(20499) := b"1111111111111111_1111111111111111_1111111101001001_1011101110011111"; -- -0.002781175372252075
	pesos_i(20500) := b"1111111111111111_1111111111111111_1110110011111011_1000000010000100"; -- -0.07428738370354011
	pesos_i(20501) := b"0000000000000000_0000000000000000_0010001011011001_1010001111100111"; -- 0.13613342648268562
	pesos_i(20502) := b"1111111111111111_1111111111111111_1110000110110110_0111101110100100"; -- -0.11830928083614994
	pesos_i(20503) := b"0000000000000000_0000000000000000_0000101010101101_0100010010000010"; -- 0.04170635400128674
	pesos_i(20504) := b"1111111111111111_1111111111111111_1110000111011111_0011010000101011"; -- -0.11768793068481442
	pesos_i(20505) := b"0000000000000000_0000000000000000_0000111100000001_1010011010110100"; -- 0.05861894499422969
	pesos_i(20506) := b"1111111111111111_1111111111111111_1110011111110010_0000001001111111"; -- -0.09396347417480506
	pesos_i(20507) := b"0000000000000000_0000000000000000_0010001010110001_0100011111001101"; -- 0.13551758526064417
	pesos_i(20508) := b"1111111111111111_1111111111111111_1111100111010110_1111110101000101"; -- -0.024063273120406008
	pesos_i(20509) := b"0000000000000000_0000000000000000_0001101000111011_1011001011100011"; -- 0.10247343098044848
	pesos_i(20510) := b"0000000000000000_0000000000000000_0001011100100011_0001110011010010"; -- 0.09037952554014048
	pesos_i(20511) := b"1111111111111111_1111111111111111_1110111101011001_0011010110001111"; -- -0.06504502536089178
	pesos_i(20512) := b"0000000000000000_0000000000000000_0000010010000111_0110011001110111"; -- 0.017691043880713225
	pesos_i(20513) := b"0000000000000000_0000000000000000_0000101011011101_1110111101010100"; -- 0.04244895752345206
	pesos_i(20514) := b"0000000000000000_0000000000000000_0010001000000011_1010010010110001"; -- 0.13286809274204225
	pesos_i(20515) := b"0000000000000000_0000000000000000_0000101010100010_1101101101011110"; -- 0.04154749916831547
	pesos_i(20516) := b"0000000000000000_0000000000000000_0000000110100010_0010001111101001"; -- 0.006380314331231187
	pesos_i(20517) := b"0000000000000000_0000000000000000_0001011011111111_0110100001111000"; -- 0.08983471805773562
	pesos_i(20518) := b"1111111111111111_1111111111111111_1101110011010101_0110111100101000"; -- -0.13736825254466872
	pesos_i(20519) := b"0000000000000000_0000000000000000_0010000101101010_0100100010011011"; -- 0.13052800934913014
	pesos_i(20520) := b"0000000000000000_0000000000000000_0000101100110001_1111111101111011"; -- 0.04373165857498047
	pesos_i(20521) := b"1111111111111111_1111111111111111_1111010001010100_1101101100010010"; -- -0.04558020416008959
	pesos_i(20522) := b"0000000000000000_0000000000000000_0001011010011100_1110000001000010"; -- 0.088331237799689
	pesos_i(20523) := b"0000000000000000_0000000000000000_0001000110110100_0110001101010110"; -- 0.06915875296401697
	pesos_i(20524) := b"1111111111111111_1111111111111111_1110010000110000_1011011000100110"; -- -0.10863172122661913
	pesos_i(20525) := b"1111111111111111_1111111111111111_1110100101001110_0000101010001100"; -- -0.08865293590763448
	pesos_i(20526) := b"0000000000000000_0000000000000000_0001110100111001_0110010011101110"; -- 0.11415701682193265
	pesos_i(20527) := b"1111111111111111_1111111111111111_1110100100110100_0100000110100101"; -- -0.08904638024010231
	pesos_i(20528) := b"1111111111111111_1111111111111111_1110010001011011_0101110100110101"; -- -0.10798089462252948
	pesos_i(20529) := b"1111111111111111_1111111111111111_1111100000110001_0010011010011100"; -- -0.030500018090286914
	pesos_i(20530) := b"0000000000000000_0000000000000000_0001011000011100_1000100001001011"; -- 0.08637286987526467
	pesos_i(20531) := b"0000000000000000_0000000000000000_0010000110101111_0011111100001001"; -- 0.1315802952028338
	pesos_i(20532) := b"0000000000000000_0000000000000000_0000111100011100_1011111010100001"; -- 0.05903235849222639
	pesos_i(20533) := b"0000000000000000_0000000000000000_0010010101010110_0111100111001011"; -- 0.1458507651905957
	pesos_i(20534) := b"0000000000000000_0000000000000000_0001111111000001_1001101100100000"; -- 0.12404794247820065
	pesos_i(20535) := b"1111111111111111_1111111111111111_1111011111001100_0011110010100000"; -- -0.03203984354124678
	pesos_i(20536) := b"1111111111111111_1111111111111111_1110000111011010_0001010100101101"; -- -0.11776607172882783
	pesos_i(20537) := b"0000000000000000_0000000000000000_0000010011010111_0010001111011101"; -- 0.01890777718369341
	pesos_i(20538) := b"0000000000000000_0000000000000000_0000100110010011_0010100001001111"; -- 0.03740169465139078
	pesos_i(20539) := b"1111111111111111_1111111111111111_1111000010101011_0111011101010111"; -- -0.059883633836879474
	pesos_i(20540) := b"0000000000000000_0000000000000000_0000110000011011_1101100101001100"; -- 0.04729993920434233
	pesos_i(20541) := b"0000000000000000_0000000000000000_0000001111101100_0110001011001101"; -- 0.015325713212930319
	pesos_i(20542) := b"0000000000000000_0000000000000000_0001001000111100_1100001101001100"; -- 0.07123966787781327
	pesos_i(20543) := b"1111111111111111_1111111111111111_1101110111101000_0100001110011110"; -- -0.13317468061653692
	pesos_i(20544) := b"1111111111111111_1111111111111111_1110111000001000_0011110011001001"; -- -0.07018680660606302
	pesos_i(20545) := b"0000000000000000_0000000000000000_0001001100100010_0111111011100110"; -- 0.07474511261093252
	pesos_i(20546) := b"0000000000000000_0000000000000000_0001100111110111_1101100101011010"; -- 0.10143812600180453
	pesos_i(20547) := b"1111111111111111_1111111111111111_1111110101101110_0011111110001011"; -- -0.010036495727092172
	pesos_i(20548) := b"0000000000000000_0000000000000000_0000001011011101_1010010100111101"; -- 0.011194541420813772
	pesos_i(20549) := b"1111111111111111_1111111111111111_1110010010110100_0101011101001000"; -- -0.10662321569064415
	pesos_i(20550) := b"0000000000000000_0000000000000000_0001100011110010_1111111100111110"; -- 0.09745784055297817
	pesos_i(20551) := b"1111111111111111_1111111111111111_1111111111111011_1001011011001001"; -- -6.73063631736693e-05
	pesos_i(20552) := b"0000000000000000_0000000000000000_0001011111101111_1101110111011101"; -- 0.09350382457860655
	pesos_i(20553) := b"1111111111111111_1111111111111111_1110001100011010_1110000110101011"; -- -0.1128710705449828
	pesos_i(20554) := b"1111111111111111_1111111111111111_1101110111001110_0110100000001011"; -- -0.13356923792081488
	pesos_i(20555) := b"0000000000000000_0000000000000000_0000101110001100_0010000011100110"; -- 0.04510694137174822
	pesos_i(20556) := b"0000000000000000_0000000000000000_0010001101011111_0000111100111100"; -- 0.1381692430982177
	pesos_i(20557) := b"1111111111111111_1111111111111111_1111100001110010_0101101010101101"; -- -0.02950509333771348
	pesos_i(20558) := b"0000000000000000_0000000000000000_0010000010000111_0001111010100011"; -- 0.12706176267408276
	pesos_i(20559) := b"0000000000000000_0000000000000000_0010010100010100_0101101010001100"; -- 0.14484182284535974
	pesos_i(20560) := b"1111111111111111_1111111111111111_1111001100100110_1110101100101000"; -- -0.05018739949693691
	pesos_i(20561) := b"1111111111111111_1111111111111111_1110000110100011_0000100100001001"; -- -0.11860602895176639
	pesos_i(20562) := b"1111111111111111_1111111111111111_1111001111011100_0111100010001000"; -- -0.04741713217004626
	pesos_i(20563) := b"0000000000000000_0000000000000000_0001000001000000_1100110000101110"; -- 0.06348873253576917
	pesos_i(20564) := b"1111111111111111_1111111111111111_1111101111001111_1100010110111001"; -- -0.01636089545638212
	pesos_i(20565) := b"1111111111111111_1111111111111111_1111011110011000_0111010001110100"; -- -0.03282997287771887
	pesos_i(20566) := b"0000000000000000_0000000000000000_0001010100010001_0100001000100001"; -- 0.08229459093795466
	pesos_i(20567) := b"0000000000000000_0000000000000000_0010000010100110_1011011111000011"; -- 0.12754391208754956
	pesos_i(20568) := b"1111111111111111_1111111111111111_1110010001101100_0110000101001010"; -- -0.10772125201468292
	pesos_i(20569) := b"0000000000000000_0000000000000000_0000111011000010_1101001101111111"; -- 0.05766031114324677
	pesos_i(20570) := b"1111111111111111_1111111111111111_1110001111010100_1101010101100100"; -- -0.11003366764642177
	pesos_i(20571) := b"1111111111111111_1111111111111111_1110010101101100_0000001111010000"; -- -0.10382057350701843
	pesos_i(20572) := b"0000000000000000_0000000000000000_0010001101101000_1001000010000000"; -- 0.13831427692352238
	pesos_i(20573) := b"1111111111111111_1111111111111111_1111010000000011_1011001110111101"; -- -0.04681851043977268
	pesos_i(20574) := b"1111111111111111_1111111111111111_1110100010010000_0000110100111000"; -- -0.09155194657171489
	pesos_i(20575) := b"0000000000000000_0000000000000000_0000011110010000_0111000110100001"; -- 0.02954778840378909
	pesos_i(20576) := b"0000000000000000_0000000000000000_0010000110001001_1100110000011101"; -- 0.1310088700868629
	pesos_i(20577) := b"0000000000000000_0000000000000000_0001101001101000_0100101110101111"; -- 0.10315392507686397
	pesos_i(20578) := b"1111111111111111_1111111111111111_1101111110100011_1000111001110110"; -- -0.12641057595877295
	pesos_i(20579) := b"1111111111111111_1111111111111111_1111010110100011_0000011101110001"; -- -0.040481123814498254
	pesos_i(20580) := b"1111111111111111_1111111111111111_1111000011000111_0101100011101111"; -- -0.059458200214942934
	pesos_i(20581) := b"0000000000000000_0000000000000000_0001100010101001_0011110010110010"; -- 0.09633235299305631
	pesos_i(20582) := b"0000000000000000_0000000000000000_0001101010101000_0101000010000101"; -- 0.10413077586384858
	pesos_i(20583) := b"0000000000000000_0000000000000000_0001011111001101_0000100000000111"; -- 0.0929722802496253
	pesos_i(20584) := b"0000000000000000_0000000000000000_0001001100111111_1001001111010110"; -- 0.07518886533568259
	pesos_i(20585) := b"0000000000000000_0000000000000000_0001100110110010_1111011101110011"; -- 0.10038706346534172
	pesos_i(20586) := b"1111111111111111_1111111111111111_1110101101110000_1000010110010110"; -- -0.08031430333482782
	pesos_i(20587) := b"0000000000000000_0000000000000000_0000011011000110_0001000101100011"; -- 0.026459776663706747
	pesos_i(20588) := b"1111111111111111_1111111111111111_1110100010100110_1010111000110000"; -- -0.09120665861520609
	pesos_i(20589) := b"1111111111111111_1111111111111111_1110101001110110_1101010111010011"; -- -0.08412421798808764
	pesos_i(20590) := b"0000000000000000_0000000000000000_0001110110111010_1000011110001101"; -- 0.11612746414873054
	pesos_i(20591) := b"1111111111111111_1111111111111111_1101100100110011_1011010001101010"; -- -0.15155479828845275
	pesos_i(20592) := b"0000000000000000_0000000000000000_0000010101000001_0000100001110101"; -- 0.02052357548109143
	pesos_i(20593) := b"0000000000000000_0000000000000000_0010100110101011_0010000101000101"; -- 0.1627674860400663
	pesos_i(20594) := b"1111111111111111_1111111111111111_1110011111011010_1010111101000101"; -- -0.09431938717132778
	pesos_i(20595) := b"0000000000000000_0000000000000000_0000110010111000_0011000001100100"; -- 0.049685501398668015
	pesos_i(20596) := b"0000000000000000_0000000000000000_0000001110011011_0111011010111100"; -- 0.01409093938670287
	pesos_i(20597) := b"1111111111111111_1111111111111111_1111110000111000_1000111110001101"; -- -0.01476195150627687
	pesos_i(20598) := b"1111111111111111_1111111111111111_1111111001011000_0011110010001001"; -- -0.006466118272027174
	pesos_i(20599) := b"1111111111111111_1111111111111111_1110101011001110_0011101011011000"; -- -0.08279068220313408
	pesos_i(20600) := b"0000000000000000_0000000000000000_0001010010001100_0100101001011001"; -- 0.08026566192227247
	pesos_i(20601) := b"1111111111111111_1111111111111111_1110100101000001_1010000110111110"; -- -0.08884228808386707
	pesos_i(20602) := b"1111111111111111_1111111111111111_1110110101111100_1100101110010110"; -- -0.07231452554306853
	pesos_i(20603) := b"0000000000000000_0000000000000000_0010000010110101_1110110111010001"; -- 0.1277760158466023
	pesos_i(20604) := b"1111111111111111_1111111111111111_1111010100001011_0110010111011010"; -- -0.04279483250304627
	pesos_i(20605) := b"0000000000000000_0000000000000000_0000100101011100_1101100011000111"; -- 0.036572979449678654
	pesos_i(20606) := b"1111111111111111_1111111111111111_1110101101010010_0000001001100011"; -- -0.08077988714019377
	pesos_i(20607) := b"0000000000000000_0000000000000000_0010000100100001_0001111010001000"; -- 0.1294116097360898
	pesos_i(20608) := b"1111111111111111_1111111111111111_1111100000100010_1000101011110100"; -- -0.03072291901545106
	pesos_i(20609) := b"1111111111111111_1111111111111111_1110001111010110_1001100111011011"; -- -0.11000669855849667
	pesos_i(20610) := b"0000000000000000_0000000000000000_0001011100011111_0101111100010110"; -- 0.09032243995147025
	pesos_i(20611) := b"1111111111111111_1111111111111111_1111001101000000_1001111110001100"; -- -0.04979517786991253
	pesos_i(20612) := b"0000000000000000_0000000000000000_0000001010000011_1010001010111010"; -- 0.009821100619230957
	pesos_i(20613) := b"0000000000000000_0000000000000000_0001011100100110_1101111110001100"; -- 0.09043690841279704
	pesos_i(20614) := b"1111111111111111_1111111111111111_1110000110000010_0110101001010101"; -- -0.11910376965033095
	pesos_i(20615) := b"0000000000000000_0000000000000000_0001011101000111_1111110001011111"; -- 0.09094216641132609
	pesos_i(20616) := b"1111111111111111_1111111111111111_1110101001101100_0000001110111100"; -- -0.08428932826228264
	pesos_i(20617) := b"0000000000000000_0000000000000000_0001000010101000_0110010011011110"; -- 0.06506948867000766
	pesos_i(20618) := b"1111111111111111_1111111111111111_1111001011000101_1100001110100110"; -- -0.05166985693874523
	pesos_i(20619) := b"0000000000000000_0000000000000000_0001011010000000_0100111001100001"; -- 0.08789529673768084
	pesos_i(20620) := b"0000000000000000_0000000000000000_0000011100000100_1001101011100100"; -- 0.02741401745004575
	pesos_i(20621) := b"0000000000000000_0000000000000000_0001011110000000_1110000010001100"; -- 0.09181025902529953
	pesos_i(20622) := b"1111111111111111_1111111111111111_1110111100011110_0000111111000001"; -- -0.06594754728262314
	pesos_i(20623) := b"0000000000000000_0000000000000000_0001000001000001_1010101100011110"; -- 0.0635020206403343
	pesos_i(20624) := b"0000000000000000_0000000000000000_0010011001011111_1001001110110001"; -- 0.14989588816248245
	pesos_i(20625) := b"1111111111111111_1111111111111111_1101110110100000_1000101100101111"; -- -0.1342690478698389
	pesos_i(20626) := b"1111111111111111_1111111111111111_1111000101110111_1111100001000100"; -- -0.05676315624844635
	pesos_i(20627) := b"1111111111111111_1111111111111111_1101101111011110_0011011010000101"; -- -0.1411405491595063
	pesos_i(20628) := b"0000000000000000_0000000000000000_0010010001001110_1011011010110001"; -- 0.14182607482979417
	pesos_i(20629) := b"1111111111111111_1111111111111111_1111000000001100_1110000010100111"; -- -0.06230350415175485
	pesos_i(20630) := b"0000000000000000_0000000000000000_0001100000001101_0111101111101111"; -- 0.09395575136187351
	pesos_i(20631) := b"1111111111111111_1111111111111111_1110100110010110_1110010111010110"; -- -0.08754123227347776
	pesos_i(20632) := b"0000000000000000_0000000000000000_0000000110010011_0011000110011011"; -- 0.006152248735162454
	pesos_i(20633) := b"0000000000000000_0000000000000000_0000011110110110_1010100000110111"; -- 0.030130876088644
	pesos_i(20634) := b"0000000000000000_0000000000000000_0001110001001101_1010111001011110"; -- 0.11056031984806021
	pesos_i(20635) := b"0000000000000000_0000000000000000_0010011100011111_0010100011010111"; -- 0.15281920663372026
	pesos_i(20636) := b"1111111111111111_1111111111111111_1101110101000001_0111001100011001"; -- -0.13572006846963447
	pesos_i(20637) := b"1111111111111111_1111111111111111_1101100111111101_1010111110010001"; -- -0.14847281188085465
	pesos_i(20638) := b"0000000000000000_0000000000000000_0001011011000110_1001000101010010"; -- 0.08896740210584761
	pesos_i(20639) := b"1111111111111111_1111111111111111_1111011110010011_1000111101010010"; -- -0.03290466538273893
	pesos_i(20640) := b"0000000000000000_0000000000000000_0000110011001100_0010101010111100"; -- 0.04999034020822525
	pesos_i(20641) := b"1111111111111111_1111111111111111_1110000101011000_1101011100100011"; -- -0.11973815348618505
	pesos_i(20642) := b"1111111111111111_1111111111111111_1111101101000101_1010010011011110"; -- -0.018468566702479705
	pesos_i(20643) := b"1111111111111111_1111111111111111_1111001100001101_0100110000010001"; -- -0.050578351873371286
	pesos_i(20644) := b"0000000000000000_0000000000000000_0000111010011101_0000011001001100"; -- 0.05708350515687556
	pesos_i(20645) := b"1111111111111111_1111111111111111_1111010001010111_1100111110100100"; -- -0.04553510905329435
	pesos_i(20646) := b"1111111111111111_1111111111111111_1111010111010100_0101011100011110"; -- -0.03972869414391844
	pesos_i(20647) := b"0000000000000000_0000000000000000_0001001110001000_0111011011111110"; -- 0.07630103782766211
	pesos_i(20648) := b"0000000000000000_0000000000000000_0000010110111001_0100011110100000"; -- 0.022358395158332135
	pesos_i(20649) := b"0000000000000000_0000000000000000_0001010111110111_0100011000011110"; -- 0.08580435009972194
	pesos_i(20650) := b"0000000000000000_0000000000000000_0010010011111100_0100100001000111"; -- 0.14447452282650644
	pesos_i(20651) := b"0000000000000000_0000000000000000_0000111000100000_0000111100000000"; -- 0.05517667524415804
	pesos_i(20652) := b"1111111111111111_1111111111111111_1111001001001011_1010000010010001"; -- -0.053533520223102135
	pesos_i(20653) := b"1111111111111111_1111111111111111_1101110110111100_1111100000000001"; -- -0.13383531541384724
	pesos_i(20654) := b"0000000000000000_0000000000000000_0010001101001110_1010110011001110"; -- 0.137919235411846
	pesos_i(20655) := b"1111111111111111_1111111111111111_1111100000100011_0011011001100101"; -- -0.030712700330371708
	pesos_i(20656) := b"0000000000000000_0000000000000000_0001010110011110_0000111001100000"; -- 0.08444299544594788
	pesos_i(20657) := b"1111111111111111_1111111111111111_1110010000110101_1000100111001101"; -- -0.10855807058467382
	pesos_i(20658) := b"0000000000000000_0000000000000000_0001110101000111_0111010010100101"; -- 0.11437157647108526
	pesos_i(20659) := b"1111111111111111_1111111111111111_1101100111111100_1110110101110111"; -- -0.1484843810603167
	pesos_i(20660) := b"1111111111111111_1111111111111111_1111101100100110_1000011001001101"; -- -0.01894341107129789
	pesos_i(20661) := b"0000000000000000_0000000000000000_0000111101011001_1011011101111001"; -- 0.059962718090907766
	pesos_i(20662) := b"0000000000000000_0000000000000000_0001101010100011_1101011001101010"; -- 0.1040624627038186
	pesos_i(20663) := b"1111111111111111_1111111111111111_1110101000001000_1010001000001111"; -- -0.08580577017885037
	pesos_i(20664) := b"1111111111111111_1111111111111111_1110110001100011_1100110101001011"; -- -0.07660214357790987
	pesos_i(20665) := b"1111111111111111_1111111111111111_1110100111101011_0011111111001001"; -- -0.08625413257523672
	pesos_i(20666) := b"1111111111111111_1111111111111111_1111111101010110_0010100101111110"; -- -0.002591521118616715
	pesos_i(20667) := b"0000000000000000_0000000000000000_0001001010001011_0100000000011001"; -- 0.07243729218388477
	pesos_i(20668) := b"0000000000000000_0000000000000000_0001011010110100_1100110010101110"; -- 0.08869628184064217
	pesos_i(20669) := b"1111111111111111_1111111111111111_1111111001010011_1100011100101000"; -- -0.006534149923971356
	pesos_i(20670) := b"1111111111111111_1111111111111111_1110010011000011_0101101011100001"; -- -0.10639411936964975
	pesos_i(20671) := b"0000000000000000_0000000000000000_0010001000010001_0100000100110010"; -- 0.13307578530037825
	pesos_i(20672) := b"1111111111111111_1111111111111111_1111000011000110_1100111110000010"; -- -0.059466391339752046
	pesos_i(20673) := b"1111111111111111_1111111111111111_1111111110010101_1001011011110010"; -- -0.0016236933215907595
	pesos_i(20674) := b"0000000000000000_0000000000000000_0000000010100110_0100111101000000"; -- 0.0025376825688467044
	pesos_i(20675) := b"1111111111111111_1111111111111111_1101110111111000_0000011110010110"; -- -0.1329341182703217
	pesos_i(20676) := b"1111111111111111_1111111111111111_1101110100100011_1000111111111010"; -- -0.1361761106622313
	pesos_i(20677) := b"1111111111111111_1111111111111111_1110110001110101_1010011111001111"; -- -0.07632971946213897
	pesos_i(20678) := b"0000000000000000_0000000000000000_0000100011111010_1111011101000011"; -- 0.035079435172382246
	pesos_i(20679) := b"1111111111111111_1111111111111111_1110000110111101_0100100011110001"; -- -0.11820549133699014
	pesos_i(20680) := b"0000000000000000_0000000000000000_0001101101100000_1011100101011000"; -- 0.10694464110422452
	pesos_i(20681) := b"0000000000000000_0000000000000000_0001011110011111_1111011101110001"; -- 0.09228464607998083
	pesos_i(20682) := b"0000000000000000_0000000000000000_0000100010001100_1100010010000001"; -- 0.033397942949954386
	pesos_i(20683) := b"1111111111111111_1111111111111111_1110001010011010_1000000011001010"; -- -0.11482997003244273
	pesos_i(20684) := b"1111111111111111_1111111111111111_1110000110010010_0000000110000101"; -- -0.11886587632545861
	pesos_i(20685) := b"1111111111111111_1111111111111111_1111101110001101_1011011100011000"; -- -0.017368847455895894
	pesos_i(20686) := b"1111111111111111_1111111111111111_1101111010101101_1000001111010001"; -- -0.13016487261853835
	pesos_i(20687) := b"0000000000000000_0000000000000000_0000000001001110_1001011011100010"; -- 0.0011991789539858731
	pesos_i(20688) := b"1111111111111111_1111111111111111_1110110110110010_1110110011101000"; -- -0.07148856479357558
	pesos_i(20689) := b"0000000000000000_0000000000000000_0001110011100000_0101101011100001"; -- 0.11279838549435384
	pesos_i(20690) := b"1111111111111111_1111111111111111_1111101100011100_0011111001010100"; -- -0.019100288897474667
	pesos_i(20691) := b"0000000000000000_0000000000000000_0001101000101111_1101010111111101"; -- 0.10229241777025824
	pesos_i(20692) := b"0000000000000000_0000000000000000_0000111000010100_1111011110101001"; -- 0.05500743752094615
	pesos_i(20693) := b"1111111111111111_1111111111111111_1110001111101011_1111100101011001"; -- -0.10968057232868057
	pesos_i(20694) := b"1111111111111111_1111111111111111_1101111111100111_1010100101100110"; -- -0.12537137271599963
	pesos_i(20695) := b"1111111111111111_1111111111111111_1101111101111000_0111111000100101"; -- -0.12706767643448236
	pesos_i(20696) := b"1111111111111111_1111111111111111_1110101000111100_1001111111010011"; -- -0.08501244630554071
	pesos_i(20697) := b"0000000000000000_0000000000000000_0000000010100111_1100011000010000"; -- 0.0025600231415561885
	pesos_i(20698) := b"1111111111111111_1111111111111111_1111001011011001_1100110110110101"; -- -0.05136408158594394
	pesos_i(20699) := b"0000000000000000_0000000000000000_0010001110010111_1000110011100101"; -- 0.13903122517330038
	pesos_i(20700) := b"0000000000000000_0000000000000000_0000110011101010_0100001001100010"; -- 0.05044951345103599
	pesos_i(20701) := b"0000000000000000_0000000000000000_0001111001001110_1111011111011111"; -- 0.11839245978374249
	pesos_i(20702) := b"0000000000000000_0000000000000000_0001110101111010_0101011100110101"; -- 0.11514802030495358
	pesos_i(20703) := b"1111111111111111_1111111111111111_1111111011010111_1000100101101000"; -- -0.0045236703899658795
	pesos_i(20704) := b"1111111111111111_1111111111111111_1111011000000011_1101010100010111"; -- -0.03900402245506196
	pesos_i(20705) := b"1111111111111111_1111111111111111_1111000000010011_0111100000110010"; -- -0.062202918835192605
	pesos_i(20706) := b"1111111111111111_1111111111111111_1101110011100100_0101111101101111"; -- -0.13714030782719042
	pesos_i(20707) := b"0000000000000000_0000000000000000_0001000111000000_1100101110000111"; -- 0.06934806870231465
	pesos_i(20708) := b"1111111111111111_1111111111111111_1110110000110010_0010101100111111"; -- -0.07735948276303621
	pesos_i(20709) := b"1111111111111111_1111111111111111_1110111001000111_1011110101101100"; -- -0.06921783555071485
	pesos_i(20710) := b"1111111111111111_1111111111111111_1111011111110111_0101111010010011"; -- -0.031381691949492405
	pesos_i(20711) := b"0000000000000000_0000000000000000_0000100011101100_1011000100010010"; -- 0.03486162848664296
	pesos_i(20712) := b"0000000000000000_0000000000000000_0001010101111011_1011010001010111"; -- 0.0839188301207992
	pesos_i(20713) := b"0000000000000000_0000000000000000_0010010111101010_0111011101101001"; -- 0.1481089240165407
	pesos_i(20714) := b"1111111111111111_1111111111111111_1101111011110011_0110111000100000"; -- -0.12909805032442057
	pesos_i(20715) := b"1111111111111111_1111111111111111_1101110010110010_0111000011001101"; -- -0.13790221206759876
	pesos_i(20716) := b"0000000000000000_0000000000000000_0001000011111010_1100111000100000"; -- 0.06632698326231976
	pesos_i(20717) := b"0000000000000000_0000000000000000_0000001100110001_1000100001010001"; -- 0.012474555762342911
	pesos_i(20718) := b"1111111111111111_1111111111111111_1110111111010111_0010100000111111"; -- -0.06312321155479446
	pesos_i(20719) := b"0000000000000000_0000000000000000_0000110011111111_1100011111000000"; -- 0.050777897275470114
	pesos_i(20720) := b"1111111111111111_1111111111111111_1110110110001101_0011010010100000"; -- -0.07206412405033052
	pesos_i(20721) := b"1111111111111111_1111111111111111_1111101101101101_0110000010001001"; -- -0.017862288151719925
	pesos_i(20722) := b"0000000000000000_0000000000000000_0000011100000100_0011001001111100"; -- 0.027407794334204497
	pesos_i(20723) := b"1111111111111111_1111111111111111_1110100000111110_1111110010000010"; -- -0.09278890434284111
	pesos_i(20724) := b"0000000000000000_0000000000000000_0000011010101100_0010000010110101"; -- 0.026063961203976947
	pesos_i(20725) := b"1111111111111111_1111111111111111_1111011101010010_0011001000111000"; -- -0.033902035987400436
	pesos_i(20726) := b"1111111111111111_1111111111111111_1111111101100111_1101110100100100"; -- -0.0023214136412354983
	pesos_i(20727) := b"1111111111111111_1111111111111111_1111000110001101_0110100111110000"; -- -0.05643594632151642
	pesos_i(20728) := b"0000000000000000_0000000000000000_0000011011000110_1100001101000111"; -- 0.026470379768628767
	pesos_i(20729) := b"0000000000000000_0000000000000000_0010000111111011_1100101100111001"; -- 0.13274831896779737
	pesos_i(20730) := b"1111111111111111_1111111111111111_1110101110011010_1110111110001101"; -- -0.07966711817970519
	pesos_i(20731) := b"0000000000000000_0000000000000000_0001010000000010_1110101001000100"; -- 0.07816948086054025
	pesos_i(20732) := b"1111111111111111_1111111111111111_1111011000110001_1110000000101101"; -- -0.03830145744475438
	pesos_i(20733) := b"0000000000000000_0000000000000000_0000110101001111_0011101000001000"; -- 0.05199015319473696
	pesos_i(20734) := b"0000000000000000_0000000000000000_0000111111011101_1000110000000101"; -- 0.06197428811577075
	pesos_i(20735) := b"1111111111111111_1111111111111111_1111110101001000_1011100011100110"; -- -0.010609096493677177
	pesos_i(20736) := b"1111111111111111_1111111111111111_1101100110110001_0111110111101011"; -- -0.14963543904195778
	pesos_i(20737) := b"1111111111111111_1111111111111111_1111011010010100_1110010100001001"; -- -0.03679054773131286
	pesos_i(20738) := b"0000000000000000_0000000000000000_0010100101100111_1010111001100101"; -- 0.16173829990844535
	pesos_i(20739) := b"0000000000000000_0000000000000000_0000010011001111_1011100101101011"; -- 0.018794621010040383
	pesos_i(20740) := b"0000000000000000_0000000000000000_0001110110101100_1111110111101101"; -- 0.1159208968874347
	pesos_i(20741) := b"1111111111111111_1111111111111111_1111010110010110_1110111011110000"; -- -0.040665689877546145
	pesos_i(20742) := b"0000000000000000_0000000000000000_0010001000100110_1101010000111110"; -- 0.1334049847075401
	pesos_i(20743) := b"1111111111111111_1111111111111111_1111011100011000_1101011001110101"; -- -0.03477725641813904
	pesos_i(20744) := b"1111111111111111_1111111111111111_1110011011000111_1101010001000011"; -- -0.09851334907613166
	pesos_i(20745) := b"1111111111111111_1111111111111111_1110011101001011_1100100101001110"; -- -0.09649984210085216
	pesos_i(20746) := b"0000000000000000_0000000000000000_0000101000010110_0110100011110101"; -- 0.039404449285504545
	pesos_i(20747) := b"0000000000000000_0000000000000000_0001011001010111_0001001101011101"; -- 0.0872661687538373
	pesos_i(20748) := b"0000000000000000_0000000000000000_0000000100100011_0010011011001001"; -- 0.004442619411864625
	pesos_i(20749) := b"1111111111111111_1111111111111111_1110001111011111_0010001001111100"; -- -0.1098764846291033
	pesos_i(20750) := b"1111111111111111_1111111111111111_1101111101100010_0010110100001110"; -- -0.12740820319614093
	pesos_i(20751) := b"0000000000000000_0000000000000000_0000111110010001_1100101101001001"; -- 0.060818391173666345
	pesos_i(20752) := b"0000000000000000_0000000000000000_0001010111101110_1000010110001001"; -- 0.08567080113991402
	pesos_i(20753) := b"0000000000000000_0000000000000000_0000000000000000_1011111000111011"; -- 1.1338710813356809e-05
	pesos_i(20754) := b"0000000000000000_0000000000000000_0001011000111010_1011101110111111"; -- 0.08683370036600432
	pesos_i(20755) := b"1111111111111111_1111111111111111_1111001100011111_1111101101100011"; -- -0.05029324364367314
	pesos_i(20756) := b"1111111111111111_1111111111111111_1110101001101001_0100011010111011"; -- -0.08433111123939502
	pesos_i(20757) := b"1111111111111111_1111111111111111_1110010000011010_1101000001010010"; -- -0.1089658545578218
	pesos_i(20758) := b"0000000000000000_0000000000000000_0000001011100101_1011110000011100"; -- 0.011317974897629868
	pesos_i(20759) := b"0000000000000000_0000000000000000_0000111000010010_1010000100001100"; -- 0.05497175724012746
	pesos_i(20760) := b"1111111111111111_1111111111111111_1101110010110010_1001100000101000"; -- -0.13789986643798874
	pesos_i(20761) := b"1111111111111111_1111111111111111_1111010001110100_1100011010110100"; -- -0.04509313674772553
	pesos_i(20762) := b"0000000000000000_0000000000000000_0001000011100111_1001000001111010"; -- 0.06603339176244467
	pesos_i(20763) := b"0000000000000000_0000000000000000_0010000010000111_1100000111000101"; -- 0.12707148603079427
	pesos_i(20764) := b"0000000000000000_0000000000000000_0010000100001101_0110011111011001"; -- 0.12911080411911155
	pesos_i(20765) := b"1111111111111111_1111111111111111_1111100011110111_1110111100110010"; -- -0.02746682195394535
	pesos_i(20766) := b"1111111111111111_1111111111111111_1111100100001101_0100100010001011"; -- -0.027141061913206383
	pesos_i(20767) := b"1111111111111111_1111111111111111_1111010101100111_1001000101010001"; -- -0.04138843329891923
	pesos_i(20768) := b"1111111111111111_1111111111111111_1110100000011110_1010110011110100"; -- -0.09328192762473204
	pesos_i(20769) := b"0000000000000000_0000000000000000_0001101000110111_1111001111100111"; -- 0.10241627118953636
	pesos_i(20770) := b"1111111111111111_1111111111111111_1110001000100001_1101101011101100"; -- -0.11667091115206743
	pesos_i(20771) := b"1111111111111111_1111111111111111_1110001010101000_0111011010110010"; -- -0.11461694865286252
	pesos_i(20772) := b"1111111111111111_1111111111111111_1111001000010000_0100011110000111"; -- -0.054439096001605194
	pesos_i(20773) := b"0000000000000000_0000000000000000_0000011011000101_1100011110100001"; -- 0.02645538024070614
	pesos_i(20774) := b"1111111111111111_1111111111111111_1111010011111011_1000110111001110"; -- -0.04303659178494617
	pesos_i(20775) := b"1111111111111111_1111111111111111_1110001111010101_1001110001101111"; -- -0.11002180365150038
	pesos_i(20776) := b"1111111111111111_1111111111111111_1111000001010101_1110000110101001"; -- -0.06118955261144646
	pesos_i(20777) := b"0000000000000000_0000000000000000_0010001101111110_0000100011101001"; -- 0.13864188848071904
	pesos_i(20778) := b"1111111111111111_1111111111111111_1111011110111011_0011010111101100"; -- -0.03229964247439529
	pesos_i(20779) := b"1111111111111111_1111111111111111_1111111101100101_0111011011000001"; -- -0.002358034045744157
	pesos_i(20780) := b"1111111111111111_1111111111111111_1110010000011010_0011110101000110"; -- -0.10897461937004087
	pesos_i(20781) := b"0000000000000000_0000000000000000_0001011000101100_0110011111000011"; -- 0.08661507131681995
	pesos_i(20782) := b"1111111111111111_1111111111111111_1111000100100111_1010001100111011"; -- -0.057988927983132106
	pesos_i(20783) := b"1111111111111111_1111111111111111_1110100101000110_0100000000101010"; -- -0.08877181024404096
	pesos_i(20784) := b"1111111111111111_1111111111111111_1110100011111010_1000001001111001"; -- -0.08992752601223838
	pesos_i(20785) := b"0000000000000000_0000000000000000_0000111001011101_1110111011110100"; -- 0.05612080998467361
	pesos_i(20786) := b"0000000000000000_0000000000000000_0001100110000110_1100101100110101"; -- 0.09971303983270033
	pesos_i(20787) := b"0000000000000000_0000000000000000_0001111011110101_0011000100010011"; -- 0.12092882841928122
	pesos_i(20788) := b"0000000000000000_0000000000000000_0000001001001101_0001101101100111"; -- 0.00898906017031454
	pesos_i(20789) := b"1111111111111111_1111111111111111_1110111100110010_1101111000110000"; -- -0.06563006705784354
	pesos_i(20790) := b"1111111111111111_1111111111111111_1111011111000000_1100000011010101"; -- -0.03221506886392299
	pesos_i(20791) := b"1111111111111111_1111111111111111_1110011110001000_1101110001111100"; -- -0.09556791272435945
	pesos_i(20792) := b"0000000000000000_0000000000000000_0001000011100111_1110011001100110"; -- 0.0660385132034502
	pesos_i(20793) := b"1111111111111111_1111111111111111_1101110001001001_0111111100110101"; -- -0.13950352636659125
	pesos_i(20794) := b"1111111111111111_1111111111111111_1111101101101001_0101101000001100"; -- -0.017923709874386292
	pesos_i(20795) := b"0000000000000000_0000000000000000_0001100100011101_1011111111110000"; -- 0.09811019524604815
	pesos_i(20796) := b"1111111111111111_1111111111111111_1111110111010010_1000100101000100"; -- -0.00850622253585329
	pesos_i(20797) := b"0000000000000000_0000000000000000_0000000101100010_1110110111010111"; -- 0.005415787689133011
	pesos_i(20798) := b"0000000000000000_0000000000000000_0000000001100010_1011000101000010"; -- 0.0015059266405669115
	pesos_i(20799) := b"0000000000000000_0000000000000000_0001100111000101_0001000001101100"; -- 0.10066321030645319
	pesos_i(20800) := b"1111111111111111_1111111111111111_1111010100011011_0001100001100110"; -- -0.042555308411308154
	pesos_i(20801) := b"0000000000000000_0000000000000000_0000111101101110_0001011111001110"; -- 0.06027363564821106
	pesos_i(20802) := b"1111111111111111_1111111111111111_1111110001000001_1001001011101110"; -- -0.014624421094532498
	pesos_i(20803) := b"1111111111111111_1111111111111111_1101100000011101_1000001100001000"; -- -0.15579968515479042
	pesos_i(20804) := b"1111111111111111_1111111111111111_1110001100111110_1111011100000001"; -- -0.11232048255734098
	pesos_i(20805) := b"0000000000000000_0000000000000000_0001011110111100_1001010011101011"; -- 0.09272127843580012
	pesos_i(20806) := b"0000000000000000_0000000000000000_0001111100111001_0110101000000100"; -- 0.1219698199897727
	pesos_i(20807) := b"0000000000000000_0000000000000000_0001000010000100_1100010010010110"; -- 0.0645258775957325
	pesos_i(20808) := b"1111111111111111_1111111111111111_1110111011000010_0100100110100001"; -- -0.0673479062558596
	pesos_i(20809) := b"1111111111111111_1111111111111111_1111101110010101_1110000110000100"; -- -0.017244248665269902
	pesos_i(20810) := b"1111111111111111_1111111111111111_1111001011111001_0101001000110000"; -- -0.050883162831564924
	pesos_i(20811) := b"1111111111111111_1111111111111111_1110101000111101_0110000110100011"; -- -0.08500089429387592
	pesos_i(20812) := b"1111111111111111_1111111111111111_1110110011111000_1011101011001001"; -- -0.0743296870270525
	pesos_i(20813) := b"0000000000000000_0000000000000000_0000010001011001_0100011100101100"; -- 0.016987274515629095
	pesos_i(20814) := b"0000000000000000_0000000000000000_0000000010111011_1101001111111100"; -- 0.0028660287801324734
	pesos_i(20815) := b"0000000000000000_0000000000000000_0000101111110101_1000100010101001"; -- 0.046715298795130755
	pesos_i(20816) := b"0000000000000000_0000000000000000_0001011001111000_1111100101110000"; -- 0.08778342228351887
	pesos_i(20817) := b"1111111111111111_1111111111111111_1111001100010001_0100011001010100"; -- -0.05051765871870663
	pesos_i(20818) := b"0000000000000000_0000000000000000_0000101000011010_0101000000010011"; -- 0.039464001277622354
	pesos_i(20819) := b"0000000000000000_0000000000000000_0000110000111100_1101101101100101"; -- 0.04780360423359391
	pesos_i(20820) := b"1111111111111111_1111111111111111_1111101110001110_0011011001111111"; -- -0.01736125383454272
	pesos_i(20821) := b"0000000000000000_0000000000000000_0000010111011110_0100100010101010"; -- 0.022923032216699803
	pesos_i(20822) := b"1111111111111111_1111111111111111_1111000110001001_1100011011110010"; -- -0.05649143784079816
	pesos_i(20823) := b"1111111111111111_1111111111111111_1111101111100110_0111111100010100"; -- -0.01601415397090136
	pesos_i(20824) := b"1111111111111111_1111111111111111_1111110100001011_1011100111011001"; -- -0.011539825847183114
	pesos_i(20825) := b"1111111111111111_1111111111111111_1111111101110000_0001010011001110"; -- -0.002196025680315937
	pesos_i(20826) := b"0000000000000000_0000000000000000_0001011011110110_0010011101100100"; -- 0.08969351004491377
	pesos_i(20827) := b"0000000000000000_0000000000000000_0000111100001000_1011111101010001"; -- 0.058727223689488274
	pesos_i(20828) := b"0000000000000000_0000000000000000_0000001011010000_0001000110100111"; -- 0.010987380292594717
	pesos_i(20829) := b"1111111111111111_1111111111111111_1110101010000000_0011011000101000"; -- -0.08398114704690382
	pesos_i(20830) := b"0000000000000000_0000000000000000_0001010111011000_0010100111010110"; -- 0.08532964194395147
	pesos_i(20831) := b"1111111111111111_1111111111111111_1101101010101011_0001110101010101"; -- -0.1458264986732647
	pesos_i(20832) := b"1111111111111111_1111111111111111_1101101011011001_1000011110110111"; -- -0.1451182535505667
	pesos_i(20833) := b"0000000000000000_0000000000000000_0001011111011111_0101011101000110"; -- 0.09325166180392362
	pesos_i(20834) := b"1111111111111111_1111111111111111_1110010000011110_1001100111001010"; -- -0.10890806978802556
	pesos_i(20835) := b"0000000000000000_0000000000000000_0000111110100100_1011001111010000"; -- 0.06110690902674782
	pesos_i(20836) := b"1111111111111111_1111111111111111_1111010001011000_0101011100011010"; -- -0.0455270349389961
	pesos_i(20837) := b"0000000000000000_0000000000000000_0000101001110010_0001011111001000"; -- 0.04080341942348429
	pesos_i(20838) := b"1111111111111111_1111111111111111_1110000000110010_0111010101101000"; -- -0.12423006265660125
	pesos_i(20839) := b"0000000000000000_0000000000000000_0001100001111100_1001010110011111"; -- 0.09565100801724685
	pesos_i(20840) := b"1111111111111111_1111111111111111_1111111010111001_1111101010111111"; -- -0.0049746784433747976
	pesos_i(20841) := b"0000000000000000_0000000000000000_0010001110010111_1110110100010101"; -- 0.13903695833789462
	pesos_i(20842) := b"1111111111111111_1111111111111111_1101011001000010_1110100000010100"; -- -0.1630415870526903
	pesos_i(20843) := b"1111111111111111_1111111111111111_1110010111101011_0001100000100000"; -- -0.10188149657954487
	pesos_i(20844) := b"0000000000000000_0000000000000000_0000000110101001_0111000000011011"; -- 0.006491667399378754
	pesos_i(20845) := b"0000000000000000_0000000000000000_0001111000100001_0010111011110100"; -- 0.11769383875927596
	pesos_i(20846) := b"1111111111111111_1111111111111111_1101100011011111_0101010011101101"; -- -0.15284222812920933
	pesos_i(20847) := b"1111111111111111_1111111111111111_1111000000000011_1100100110011100"; -- -0.06244220679664795
	pesos_i(20848) := b"0000000000000000_0000000000000000_0010001111011001_0010001111100101"; -- 0.14003204681232811
	pesos_i(20849) := b"0000000000000000_0000000000000000_0001011111100001_1101101111010101"; -- 0.09329008053100428
	pesos_i(20850) := b"1111111111111111_1111111111111111_1110111111110110_1001001110001011"; -- -0.06264379359927323
	pesos_i(20851) := b"0000000000000000_0000000000000000_0010011000100010_0100000111010001"; -- 0.1489602216769371
	pesos_i(20852) := b"0000000000000000_0000000000000000_0001000110011110_1000110010000000"; -- 0.06882551320165016
	pesos_i(20853) := b"0000000000000000_0000000000000000_0001000111001100_0100011101011001"; -- 0.06952329561329078
	pesos_i(20854) := b"1111111111111111_1111111111111111_1101111010011001_0101111011011111"; -- -0.13047225061311882
	pesos_i(20855) := b"0000000000000000_0000000000000000_0000011001010000_0111001111100111"; -- 0.024665111444996633
	pesos_i(20856) := b"0000000000000000_0000000000000000_0000100111100010_1001001001100100"; -- 0.0386134619983154
	pesos_i(20857) := b"0000000000000000_0000000000000000_0000010000111110_0100011001001111"; -- 0.016575235706129003
	pesos_i(20858) := b"0000000000000000_0000000000000000_0010001011010111_0001110011111111"; -- 0.13609486790749165
	pesos_i(20859) := b"1111111111111111_1111111111111111_1110010100001000_1110000110011110"; -- -0.1053332318792613
	pesos_i(20860) := b"1111111111111111_1111111111111111_1111011101101101_1100011100100101"; -- -0.033481172047694845
	pesos_i(20861) := b"1111111111111111_1111111111111111_1101100100011101_1001010000100011"; -- -0.15189241550681662
	pesos_i(20862) := b"1111111111111111_1111111111111111_1111100111001111_1001111111000010"; -- -0.024175658324960127
	pesos_i(20863) := b"0000000000000000_0000000000000000_0000100110000000_1100010001101011"; -- 0.03712108244729809
	pesos_i(20864) := b"0000000000000000_0000000000000000_0000010110110111_1110100000111011"; -- 0.0223374504279803
	pesos_i(20865) := b"1111111111111111_1111111111111111_1101100001100110_0010101000100000"; -- -0.1546910926972398
	pesos_i(20866) := b"0000000000000000_0000000000000000_0001010000100111_1000000011110011"; -- 0.0787277787437301
	pesos_i(20867) := b"0000000000000000_0000000000000000_0000011011101000_0011100011101110"; -- 0.026980932340220965
	pesos_i(20868) := b"0000000000000000_0000000000000000_0001001100011110_1000100001011001"; -- 0.07468464067806753
	pesos_i(20869) := b"1111111111111111_1111111111111111_1110011011110010_0001010101000111"; -- -0.09786860486383375
	pesos_i(20870) := b"1111111111111111_1111111111111111_1111100110111101_1001011011100111"; -- -0.024450844371632967
	pesos_i(20871) := b"0000000000000000_0000000000000000_0000101011101000_0100100111111011"; -- 0.042606948699982515
	pesos_i(20872) := b"0000000000000000_0000000000000000_0001011110011011_0111101101100000"; -- 0.09221621605958275
	pesos_i(20873) := b"0000000000000000_0000000000000000_0001010110100011_1000101111001001"; -- 0.08452676454426836
	pesos_i(20874) := b"1111111111111111_1111111111111111_1110011000111011_1101011010010001"; -- -0.10064944221390054
	pesos_i(20875) := b"0000000000000000_0000000000000000_0001000111111101_0011110000110110"; -- 0.07027031237200003
	pesos_i(20876) := b"1111111111111111_1111111111111111_1111101111110011_1101001101010111"; -- -0.015810767384926594
	pesos_i(20877) := b"1111111111111111_1111111111111111_1111111000011000_1011010011000000"; -- -0.007435515556969109
	pesos_i(20878) := b"1111111111111111_1111111111111111_1101100011110011_0000111111011101"; -- -0.15254116866945236
	pesos_i(20879) := b"0000000000000000_0000000000000000_0000101010100111_1100000110111110"; -- 0.041622265604345766
	pesos_i(20880) := b"1111111111111111_1111111111111111_1111000000100110_0100111000100010"; -- -0.06191550894718964
	pesos_i(20881) := b"1111111111111111_1111111111111111_1111101000110000_1000100101101111"; -- -0.022696886460538714
	pesos_i(20882) := b"0000000000000000_0000000000000000_0000111011011101_0111111001000010"; -- 0.05806721793573474
	pesos_i(20883) := b"0000000000000000_0000000000000000_0001100100010101_1110001000101110"; -- 0.09799016594004971
	pesos_i(20884) := b"0000000000000000_0000000000000000_0001101010001001_1001000000011001"; -- 0.1036615430717251
	pesos_i(20885) := b"1111111111111111_1111111111111111_1110001011010000_0011101000001011"; -- -0.11401021235465512
	pesos_i(20886) := b"0000000000000000_0000000000000000_0001111110010110_0010000001101001"; -- 0.12338450027037658
	pesos_i(20887) := b"0000000000000000_0000000000000000_0001101011011000_0001000100100111"; -- 0.10485942084073852
	pesos_i(20888) := b"1111111111111111_1111111111111111_1110001110000101_0010011110011110"; -- -0.11124946961834159
	pesos_i(20889) := b"0000000000000000_0000000000000000_0001001010000000_1011101011000100"; -- 0.07227675719456306
	pesos_i(20890) := b"1111111111111111_1111111111111111_1111100001111101_1111010100110110"; -- -0.029328035746634614
	pesos_i(20891) := b"0000000000000000_0000000000000000_0010011011000111_0001011111000001"; -- 0.15147541491881625
	pesos_i(20892) := b"0000000000000000_0000000000000000_0010001011111011_1011010110111111"; -- 0.13665328899600046
	pesos_i(20893) := b"1111111111111111_1111111111111111_1110111001111110_0110111011100100"; -- -0.068383282949337
	pesos_i(20894) := b"0000000000000000_0000000000000000_0000001100010011_0110000101111110"; -- 0.012014477965067959
	pesos_i(20895) := b"1111111111111111_1111111111111111_1110100001111011_1110001011000001"; -- -0.09185965330692734
	pesos_i(20896) := b"0000000000000000_0000000000000000_0010001011100111_1010001000010101"; -- 0.13634694107133502
	pesos_i(20897) := b"0000000000000000_0000000000000000_0000001101111010_0110101101100111"; -- 0.013586724031976494
	pesos_i(20898) := b"0000000000000000_0000000000000000_0010001101110101_0110110101100011"; -- 0.13851054828514775
	pesos_i(20899) := b"1111111111111111_1111111111111111_1111110110110000_1001001011110001"; -- -0.009024444670193504
	pesos_i(20900) := b"1111111111111111_1111111111111111_1111101110110100_0001111100011010"; -- -0.016782814203221565
	pesos_i(20901) := b"1111111111111111_1111111111111111_1110110011110101_0011011000110100"; -- -0.07438336595866205
	pesos_i(20902) := b"1111111111111111_1111111111111111_1101100111010101_1110100010100001"; -- -0.1490797620694509
	pesos_i(20903) := b"1111111111111111_1111111111111111_1110111111110000_1111010011010111"; -- -0.06272954709321281
	pesos_i(20904) := b"1111111111111111_1111111111111111_1110101110000011_0111011011101110"; -- -0.08002525980579674
	pesos_i(20905) := b"1111111111111111_1111111111111111_1111011001111010_1001110111101101"; -- -0.03719151465553043
	pesos_i(20906) := b"1111111111111111_1111111111111111_1111000000110101_1110000101110010"; -- -0.06167784652802087
	pesos_i(20907) := b"0000000000000000_0000000000000000_0000010111010111_1001000101011101"; -- 0.02282055398174459
	pesos_i(20908) := b"1111111111111111_1111111111111111_1111111100010101_0111100101100111"; -- -0.0035785791970218226
	pesos_i(20909) := b"1111111111111111_1111111111111111_1111001011001001_0011101101100011"; -- -0.05161694361230158
	pesos_i(20910) := b"1111111111111111_1111111111111111_1101110011010101_0011001001101110"; -- -0.137371872112978
	pesos_i(20911) := b"0000000000000000_0000000000000000_0001110110101010_0011010010111100"; -- 0.11587838736681134
	pesos_i(20912) := b"0000000000000000_0000000000000000_0000111011100010_1011110110101111"; -- 0.05814729237698724
	pesos_i(20913) := b"1111111111111111_1111111111111111_1101111111011100_1001010011000111"; -- -0.12554044861189145
	pesos_i(20914) := b"1111111111111111_1111111111111111_1110001111111100_0110110001010001"; -- -0.10942957902051492
	pesos_i(20915) := b"1111111111111111_1111111111111111_1101101101000011_1100011000101011"; -- -0.143497099368354
	pesos_i(20916) := b"0000000000000000_0000000000000000_0010001100101011_1001000111111000"; -- 0.13738357838488
	pesos_i(20917) := b"1111111111111111_1111111111111111_1101101001100010_0110001110001111"; -- -0.14693620450268424
	pesos_i(20918) := b"0000000000000000_0000000000000000_0001001100000100_1001110111010011"; -- 0.07428919228639533
	pesos_i(20919) := b"0000000000000000_0000000000000000_0000111100010110_0010111001001100"; -- 0.058932202813584356
	pesos_i(20920) := b"0000000000000000_0000000000000000_0001001001100110_1110101011101011"; -- 0.0718828986167003
	pesos_i(20921) := b"0000000000000000_0000000000000000_0000000001010100_0110011111000001"; -- 0.0012879225812266885
	pesos_i(20922) := b"0000000000000000_0000000000000000_0010001010001101_0100001110011100"; -- 0.13496801917019055
	pesos_i(20923) := b"1111111111111111_1111111111111111_1110001111011000_0111101101001111"; -- -0.10997800174650527
	pesos_i(20924) := b"1111111111111111_1111111111111111_1110101011001001_1111011110111100"; -- -0.08285571737437016
	pesos_i(20925) := b"0000000000000000_0000000000000000_0001001011100010_1001100101110010"; -- 0.07377013226896237
	pesos_i(20926) := b"1111111111111111_1111111111111111_1101110001000101_0010010100000101"; -- -0.1395699369208977
	pesos_i(20927) := b"1111111111111111_1111111111111111_1110111101101000_0010010000000100"; -- -0.06481718932318901
	pesos_i(20928) := b"0000000000000000_0000000000000000_0000110010101000_1001011100010111"; -- 0.04944748223239147
	pesos_i(20929) := b"0000000000000000_0000000000000000_0000000010100111_0100000100100100"; -- 0.0025521005148978885
	pesos_i(20930) := b"1111111111111111_1111111111111111_1110111111010011_1101101011110011"; -- -0.06317359512026938
	pesos_i(20931) := b"1111111111111111_1111111111111111_1101110000101001_1000000100000000"; -- -0.13999170066779426
	pesos_i(20932) := b"0000000000000000_0000000000000000_0000010101000111_0101011101000111"; -- 0.020619826199280298
	pesos_i(20933) := b"1111111111111111_1111111111111111_1110100000111001_1100000010010000"; -- -0.0928687714127018
	pesos_i(20934) := b"1111111111111111_1111111111111111_1110011010001000_1010101000100100"; -- -0.09947716351582257
	pesos_i(20935) := b"0000000000000000_0000000000000000_0001000010000011_0101001001100001"; -- 0.06450381159229655
	pesos_i(20936) := b"0000000000000000_0000000000000000_0001110110010001_1111101010111010"; -- 0.1155087188531256
	pesos_i(20937) := b"1111111111111111_1111111111111111_1111010110000100_1000000100011100"; -- -0.04094689431544918
	pesos_i(20938) := b"1111111111111111_1111111111111111_1101011011011100_1001000100110010"; -- -0.1606969121772285
	pesos_i(20939) := b"1111111111111111_1111111111111111_1110100000000110_0010111011011101"; -- -0.09365565392214635
	pesos_i(20940) := b"0000000000000000_0000000000000000_0001110001110100_1111010001001001"; -- 0.11115958005759162
	pesos_i(20941) := b"0000000000000000_0000000000000000_0001101000100010_0001001110100111"; -- 0.1020824702188012
	pesos_i(20942) := b"1111111111111111_1111111111111111_1101101111000101_0111111011100000"; -- -0.14151770623104723
	pesos_i(20943) := b"1111111111111111_1111111111111111_1111000110011111_0111010011110000"; -- -0.05616063256725214
	pesos_i(20944) := b"0000000000000000_0000000000000000_0001001010001000_0010101001000101"; -- 0.07239021487958032
	pesos_i(20945) := b"0000000000000000_0000000000000000_0010001110111011_1101111000101100"; -- 0.13958538597659326
	pesos_i(20946) := b"0000000000000000_0000000000000000_0000001000011111_1100110000111101"; -- 0.008297696120997218
	pesos_i(20947) := b"1111111111111111_1111111111111111_1101110101101000_1011101111100011"; -- -0.13512063702030847
	pesos_i(20948) := b"1111111111111111_1111111111111111_1110101111000011_0010000011101110"; -- -0.0790538233321511
	pesos_i(20949) := b"0000000000000000_0000000000000000_0000001010100100_0011111001001001"; -- 0.010318653924720483
	pesos_i(20950) := b"0000000000000000_0000000000000000_0001010011010000_1011011110011011"; -- 0.08130977186409676
	pesos_i(20951) := b"1111111111111111_1111111111111111_1110100011111001_1010000110011010"; -- -0.08994092936604366
	pesos_i(20952) := b"0000000000000000_0000000000000000_0001111111010010_1110110111101111"; -- 0.12431227758750621
	pesos_i(20953) := b"1111111111111111_1111111111111111_1110011111010010_0111001110011110"; -- -0.0944450130068111
	pesos_i(20954) := b"1111111111111111_1111111111111111_1110110110001101_0011110110001111"; -- -0.0720635915978189
	pesos_i(20955) := b"0000000000000000_0000000000000000_0000000100000010_1111010101100100"; -- 0.003951393932792449
	pesos_i(20956) := b"0000000000000000_0000000000000000_0000001101111011_1110011101011000"; -- 0.013609370328058288
	pesos_i(20957) := b"1111111111111111_1111111111111111_1111110101100010_0011001010111000"; -- -0.010220365485008374
	pesos_i(20958) := b"1111111111111111_1111111111111111_1110110010100111_1011001011110110"; -- -0.07556611525123837
	pesos_i(20959) := b"1111111111111111_1111111111111111_1101110101100010_0101111000111010"; -- -0.13521777230095988
	pesos_i(20960) := b"0000000000000000_0000000000000000_0010000001101001_0110110100000001"; -- 0.12660866992483935
	pesos_i(20961) := b"0000000000000000_0000000000000000_0001100111100101_0111000101011010"; -- 0.10115726886648022
	pesos_i(20962) := b"1111111111111111_1111111111111111_1110000000010111_0011001011010010"; -- -0.12464601863947355
	pesos_i(20963) := b"0000000000000000_0000000000000000_0010000001011000_0001011011010000"; -- 0.12634413305749978
	pesos_i(20964) := b"1111111111111111_1111111111111111_1111000100000000_0010011011111111"; -- -0.058591425768027824
	pesos_i(20965) := b"0000000000000000_0000000000000000_0000001001000101_0111010111110000"; -- 0.008872386043511739
	pesos_i(20966) := b"0000000000000000_0000000000000000_0000111011000111_1100000101111111"; -- 0.057735532304758974
	pesos_i(20967) := b"1111111111111111_1111111111111111_1101111111101010_1100111011010001"; -- -0.12532336607050612
	pesos_i(20968) := b"1111111111111111_1111111111111111_1111010101010000_1101011100010001"; -- -0.04173522793844828
	pesos_i(20969) := b"0000000000000000_0000000000000000_0000000111100001_0101100101100101"; -- 0.00734480591120133
	pesos_i(20970) := b"1111111111111111_1111111111111111_1111110100100011_1110001100000101"; -- -0.011171160972522626
	pesos_i(20971) := b"1111111111111111_1111111111111111_1111100000001110_0110010000000010"; -- -0.031030415940429365
	pesos_i(20972) := b"0000000000000000_0000000000000000_0001100001011000_1111101110100101"; -- 0.09510777258805835
	pesos_i(20973) := b"1111111111111111_1111111111111111_1101101011100110_0101100110101000"; -- -0.14492263469280628
	pesos_i(20974) := b"0000000000000000_0000000000000000_0010000110101110_0000101110110111"; -- 0.13156197748419143
	pesos_i(20975) := b"0000000000000000_0000000000000000_0001111100000111_1100111001100110"; -- 0.12121286374898885
	pesos_i(20976) := b"0000000000000000_0000000000000000_0000101011110010_0001111001101100"; -- 0.0427569402521995
	pesos_i(20977) := b"1111111111111111_1111111111111111_1110001010110111_0110101011101111"; -- -0.11438876792806937
	pesos_i(20978) := b"0000000000000000_0000000000000000_0001111011111010_0010000011101111"; -- 0.1210041603119113
	pesos_i(20979) := b"1111111111111111_1111111111111111_1110011010000010_1101100100110100"; -- -0.09956591109565324
	pesos_i(20980) := b"0000000000000000_0000000000000000_0000000011011110_1111010001011111"; -- 0.0034020167366678603
	pesos_i(20981) := b"0000000000000000_0000000000000000_0000001101000101_0111001011110011"; -- 0.012778458015266444
	pesos_i(20982) := b"0000000000000000_0000000000000000_0001111101111001_0111000110110101"; -- 0.12294684082918657
	pesos_i(20983) := b"1111111111111111_1111111111111111_1111110010110110_1000101010000100"; -- -0.01283964414144575
	pesos_i(20984) := b"0000000000000000_0000000000000000_0001010000001101_1001000000101011"; -- 0.07833195745175361
	pesos_i(20985) := b"0000000000000000_0000000000000000_0001010100000011_1111001000010111"; -- 0.08209145596365111
	pesos_i(20986) := b"0000000000000000_0000000000000000_0001111100100000_1001000010000101"; -- 0.12159064520129012
	pesos_i(20987) := b"1111111111111111_1111111111111111_1110000101100110_0100000100000001"; -- -0.11953347901410043
	pesos_i(20988) := b"0000000000000000_0000000000000000_0001100000111011_1101100011000011"; -- 0.0946631886615166
	pesos_i(20989) := b"1111111111111111_1111111111111111_1101111110001010_0101110000101010"; -- -0.12679504362380267
	pesos_i(20990) := b"1111111111111111_1111111111111111_1111000110011011_1101110111011110"; -- -0.05621541330066724
	pesos_i(20991) := b"1111111111111111_1111111111111111_1101100111010110_1101100100011111"; -- -0.14906542767496098
	pesos_i(20992) := b"1111111111111111_1111111111111111_1110011001110000_0100111100011000"; -- -0.09984880128203791
	pesos_i(20993) := b"1111111111111111_1111111111111111_1111010100000010_1010101010001011"; -- -0.04292806728361824
	pesos_i(20994) := b"1111111111111111_1111111111111111_1110000110111110_1101100100100000"; -- -0.11818163832692045
	pesos_i(20995) := b"0000000000000000_0000000000000000_0001111010100111_0101101100011000"; -- 0.11974114745136857
	pesos_i(20996) := b"1111111111111111_1111111111111111_1110100001011001_1110011110001110"; -- -0.09237816594421237
	pesos_i(20997) := b"1111111111111111_1111111111111111_1110001000111101_1100000011100101"; -- -0.11624521643462513
	pesos_i(20998) := b"1111111111111111_1111111111111111_1101111000111000_0010001000010110"; -- -0.1319559760863157
	pesos_i(20999) := b"1111111111111111_1111111111111111_1101101111100100_0110101111001101"; -- -0.14104582056396525
	pesos_i(21000) := b"1111111111111111_1111111111111111_1110010111010011_1000010110101100"; -- -0.10224117812730926
	pesos_i(21001) := b"0000000000000000_0000000000000000_0000100011101011_1010000001001000"; -- 0.03484536885655913
	pesos_i(21002) := b"1111111111111111_1111111111111111_1110111011011110_1111000011111111"; -- -0.06691068437087827
	pesos_i(21003) := b"1111111111111111_1111111111111111_1101101100101110_0000110000011001"; -- -0.14382862460807821
	pesos_i(21004) := b"1111111111111111_1111111111111111_1111101110111100_0111100001001010"; -- -0.016655427872116244
	pesos_i(21005) := b"0000000000000000_0000000000000000_0000011000111001_1000011000100001"; -- 0.02431524564163161
	pesos_i(21006) := b"0000000000000000_0000000000000000_0000110101010111_0110110100001010"; -- 0.052115263811952875
	pesos_i(21007) := b"0000000000000000_0000000000000000_0000001100001100_1100000000110110"; -- 0.011913312059931921
	pesos_i(21008) := b"0000000000000000_0000000000000000_0001111001000111_0000111011000011"; -- 0.11827175390884968
	pesos_i(21009) := b"1111111111111111_1111111111111111_1110101111000000_0011100101110101"; -- -0.07909813784055478
	pesos_i(21010) := b"1111111111111111_1111111111111111_1111101101101000_1110101111011011"; -- -0.017930277753739038
	pesos_i(21011) := b"1111111111111111_1111111111111111_1111111010001100_1110000110110001"; -- -0.005662817321260817
	pesos_i(21012) := b"1111111111111111_1111111111111111_1110011111111110_1000010001100011"; -- -0.0937726267806666
	pesos_i(21013) := b"1111111111111111_1111111111111111_1111000000101011_1000111101010001"; -- -0.0618353296616725
	pesos_i(21014) := b"1111111111111111_1111111111111111_1111010100110101_0001000101010101"; -- -0.04215900104450372
	pesos_i(21015) := b"0000000000000000_0000000000000000_0000010111000000_0001010001000100"; -- 0.022462145448217157
	pesos_i(21016) := b"0000000000000000_0000000000000000_0001001101100010_1011100001010100"; -- 0.07572509814597893
	pesos_i(21017) := b"1111111111111111_1111111111111111_1110111101011110_0101011111101110"; -- -0.06496668291989086
	pesos_i(21018) := b"1111111111111111_1111111111111111_1110001100101111_0110100100001101"; -- -0.11255782543716887
	pesos_i(21019) := b"1111111111111111_1111111111111111_1111011101100110_0011000011100010"; -- -0.03359693984056157
	pesos_i(21020) := b"1111111111111111_1111111111111111_1110101100110011_0010001001011010"; -- -0.08125100415691894
	pesos_i(21021) := b"0000000000000000_0000000000000000_0001111011010001_1110000100010011"; -- 0.12039000244159763
	pesos_i(21022) := b"1111111111111111_1111111111111111_1101110000010000_1100100111111001"; -- -0.14036882085339838
	pesos_i(21023) := b"1111111111111111_1111111111111111_1101111010110011_0000001000000001"; -- -0.13008105736854333
	pesos_i(21024) := b"1111111111111111_1111111111111111_1110001101001111_1001111100101111"; -- -0.11206631756444055
	pesos_i(21025) := b"1111111111111111_1111111111111111_1111101011011010_1010100100110001"; -- -0.020100999415267776
	pesos_i(21026) := b"1111111111111111_1111111111111111_1110000010001010_0101111011110100"; -- -0.12288862741335228
	pesos_i(21027) := b"0000000000000000_0000000000000000_0000000000001001_0111110000010011"; -- 0.00014472445960028805
	pesos_i(21028) := b"0000000000000000_0000000000000000_0001111001001111_1010001010000100"; -- 0.11840263100322819
	pesos_i(21029) := b"1111111111111111_1111111111111111_1111010100111010_1000000111011100"; -- -0.04207600004699854
	pesos_i(21030) := b"1111111111111111_1111111111111111_1101011000111011_0110110011111101"; -- -0.16315573514169038
	pesos_i(21031) := b"1111111111111111_1111111111111111_1110000101011111_0001011001111111"; -- -0.11964282412784612
	pesos_i(21032) := b"0000000000000000_0000000000000000_0010001101110010_0000110000100100"; -- 0.1384589755639605
	pesos_i(21033) := b"0000000000000000_0000000000000000_0001101110111110_1011100010010000"; -- 0.1083789207141287
	pesos_i(21034) := b"0000000000000000_0000000000000000_0000000001100000_1111100111000010"; -- 0.001479730423821034
	pesos_i(21035) := b"1111111111111111_1111111111111111_1110011011111100_1111000100111010"; -- -0.09770290698603244
	pesos_i(21036) := b"1111111111111111_1111111111111111_1110100111010101_0110111001111000"; -- -0.08658704343421264
	pesos_i(21037) := b"1111111111111111_1111111111111111_1101100111110111_0111111000110001"; -- -0.14856730740308585
	pesos_i(21038) := b"1111111111111111_1111111111111111_1110000111000110_1100101000111011"; -- -0.1180604559942365
	pesos_i(21039) := b"1111111111111111_1111111111111111_1101110010000011_1101001110010000"; -- -0.13861348848871033
	pesos_i(21040) := b"0000000000000000_0000000000000000_0000101000101100_1010000100110100"; -- 0.03974349524537485
	pesos_i(21041) := b"1111111111111111_1111111111111111_1101110011000101_0000010110110110"; -- -0.1376186781259174
	pesos_i(21042) := b"0000000000000000_0000000000000000_0010000000100000_1001001001111010"; -- 0.1254970119058033
	pesos_i(21043) := b"0000000000000000_0000000000000000_0000000101010100_0111110110110111"; -- 0.005195481478000739
	pesos_i(21044) := b"0000000000000000_0000000000000000_0001001110111110_1001100101100000"; -- 0.07712706189283745
	pesos_i(21045) := b"0000000000000000_0000000000000000_0000000101011101_1001110001111011"; -- 0.0053346444434788694
	pesos_i(21046) := b"1111111111111111_1111111111111111_1111011000010001_1100110001101000"; -- -0.038790917037292025
	pesos_i(21047) := b"1111111111111111_1111111111111111_1110101110111101_0011100010011110"; -- -0.07914396415585065
	pesos_i(21048) := b"1111111111111111_1111111111111111_1111010001101010_1011010100100110"; -- -0.045246771077394034
	pesos_i(21049) := b"1111111111111111_1111111111111111_1111100000001110_0011001000011000"; -- -0.031033391204031216
	pesos_i(21050) := b"0000000000000000_0000000000000000_0010010000000011_1000110101011000"; -- 0.1406792012237505
	pesos_i(21051) := b"1111111111111111_1111111111111111_1110001011100101_1110100101000101"; -- -0.11367933344323893
	pesos_i(21052) := b"0000000000000000_0000000000000000_0010001010011100_1000101010011110"; -- 0.13520113338758438
	pesos_i(21053) := b"0000000000000000_0000000000000000_0001001100001110_0110010000000011"; -- 0.07443833409923167
	pesos_i(21054) := b"0000000000000000_0000000000000000_0001110000110010_0000110100011010"; -- 0.11013872041817802
	pesos_i(21055) := b"0000000000000000_0000000000000000_0000111101111111_1111100000110111"; -- 0.06054641095793761
	pesos_i(21056) := b"0000000000000000_0000000000000000_0010001010000110_0110000100011000"; -- 0.1348629649783774
	pesos_i(21057) := b"1111111111111111_1111111111111111_1110110001010110_1110001110000001"; -- -0.07679918382480479
	pesos_i(21058) := b"1111111111111111_1111111111111111_1111110111110101_1110000110100000"; -- -0.00796689829145264
	pesos_i(21059) := b"0000000000000000_0000000000000000_0001101000010100_0110100101000011"; -- 0.10187394988301944
	pesos_i(21060) := b"1111111111111111_1111111111111111_1111111111110111_0011011010011111"; -- -0.0001340734865379573
	pesos_i(21061) := b"1111111111111111_1111111111111111_1111001101001110_1001001110000010"; -- -0.049582272315665255
	pesos_i(21062) := b"0000000000000000_0000000000000000_0000010011001010_0001011011000001"; -- 0.018708631536389218
	pesos_i(21063) := b"0000000000000000_0000000000000000_0000000011110010_1010001010011001"; -- 0.0037023185220783003
	pesos_i(21064) := b"1111111111111111_1111111111111111_1110001011000101_1110010110001110"; -- -0.11416783596761455
	pesos_i(21065) := b"0000000000000000_0000000000000000_0000110111100000_0010111101000000"; -- 0.054202035112448116
	pesos_i(21066) := b"1111111111111111_1111111111111111_1111111000001101_0000001110100101"; -- -0.0076139184706832995
	pesos_i(21067) := b"0000000000000000_0000000000000000_0010011000001100_0011100001011111"; -- 0.14862396545605933
	pesos_i(21068) := b"0000000000000000_0000000000000000_0001001111000111_1000101001000101"; -- 0.07726349047099676
	pesos_i(21069) := b"1111111111111111_1111111111111111_1110001010101110_0110101000010100"; -- -0.11452614799316277
	pesos_i(21070) := b"1111111111111111_1111111111111111_1111100111111010_0101100111110111"; -- -0.023523690361023135
	pesos_i(21071) := b"1111111111111111_1111111111111111_1110001111001011_0100101001100101"; -- -0.11017928153519135
	pesos_i(21072) := b"0000000000000000_0000000000000000_0000100010000000_0100101111001001"; -- 0.03320764217569012
	pesos_i(21073) := b"0000000000000000_0000000000000000_0010000111101100_1101000010000001"; -- 0.1325197519548105
	pesos_i(21074) := b"0000000000000000_0000000000000000_0001000010111001_1000101111011010"; -- 0.06533121179423662
	pesos_i(21075) := b"1111111111111111_1111111111111111_1111010111101100_0101100110010110"; -- -0.039362336101919936
	pesos_i(21076) := b"1111111111111111_1111111111111111_1110001011010100_0111011111010101"; -- -0.11394549409192817
	pesos_i(21077) := b"1111111111111111_1111111111111111_1110011000100100_0111110011011010"; -- -0.10100574194115713
	pesos_i(21078) := b"1111111111111111_1111111111111111_1110001001010000_1111001010001100"; -- -0.11595233988380331
	pesos_i(21079) := b"0000000000000000_0000000000000000_0010000101111100_0100110000100001"; -- 0.13080287747450917
	pesos_i(21080) := b"0000000000000000_0000000000000000_0010000000110001_0111111100101010"; -- 0.12575526019139457
	pesos_i(21081) := b"0000000000000000_0000000000000000_0001100110101010_1001111011101010"; -- 0.10025971611033607
	pesos_i(21082) := b"1111111111111111_1111111111111111_1110001110001010_1001110001010110"; -- -0.11116621884957024
	pesos_i(21083) := b"1111111111111111_1111111111111111_1110111000111100_1001111100110110"; -- -0.06938748288348154
	pesos_i(21084) := b"0000000000000000_0000000000000000_0000110100010101_0101111110001010"; -- 0.051107379246502486
	pesos_i(21085) := b"1111111111111111_1111111111111111_1101110000110101_0100111011101000"; -- -0.13981158108975364
	pesos_i(21086) := b"0000000000000000_0000000000000000_0001010001100011_0000111010111001"; -- 0.07963649762000585
	pesos_i(21087) := b"0000000000000000_0000000000000000_0010001001101111_1111011010010110"; -- 0.13452092321363032
	pesos_i(21088) := b"0000000000000000_0000000000000000_0000001010101000_0100111110101011"; -- 0.010380725138163861
	pesos_i(21089) := b"0000000000000000_0000000000000000_0001001000000111_1100011001010100"; -- 0.07043113276911776
	pesos_i(21090) := b"0000000000000000_0000000000000000_0000011000110010_1011101011101011"; -- 0.02421158071171014
	pesos_i(21091) := b"1111111111111111_1111111111111111_1110000001010111_1111001000000101"; -- -0.12365805993228003
	pesos_i(21092) := b"0000000000000000_0000000000000000_0000011101101010_0101111111011001"; -- 0.02896689463307201
	pesos_i(21093) := b"1111111111111111_1111111111111111_1101100101010100_0111110100100110"; -- -0.15105455230962103
	pesos_i(21094) := b"0000000000000000_0000000000000000_0001011100010100_0110100101001100"; -- 0.0901552020392833
	pesos_i(21095) := b"1111111111111111_1111111111111111_1101110110010100_0100110011000101"; -- -0.13445587341218854
	pesos_i(21096) := b"1111111111111111_1111111111111111_1110100000001101_0101110010110101"; -- -0.09354610996181613
	pesos_i(21097) := b"0000000000000000_0000000000000000_0000010111101110_1111000101011000"; -- 0.023177226916501772
	pesos_i(21098) := b"1111111111111111_1111111111111111_1110111101001001_0011100000101100"; -- -0.06528901023286969
	pesos_i(21099) := b"1111111111111111_1111111111111111_1110110111110101_1110000001000010"; -- -0.07046697987268873
	pesos_i(21100) := b"0000000000000000_0000000000000000_0000011110111010_1011110111100110"; -- 0.030193203637265423
	pesos_i(21101) := b"0000000000000000_0000000000000000_0001010000011011_1101110100000101"; -- 0.07855016104453202
	pesos_i(21102) := b"1111111111111111_1111111111111111_1111010000011100_0001000101010110"; -- -0.04644672064259902
	pesos_i(21103) := b"1111111111111111_1111111111111111_1101110001110011_1010001010100110"; -- -0.13886054470406603
	pesos_i(21104) := b"0000000000000000_0000000000000000_0010001001010011_0101001101000101"; -- 0.13408394267389226
	pesos_i(21105) := b"0000000000000000_0000000000000000_0000000011000101_0010001011100111"; -- 0.003008061894643198
	pesos_i(21106) := b"1111111111111111_1111111111111111_1110100000001111_1011101111101010"; -- -0.09350991763576047
	pesos_i(21107) := b"0000000000000000_0000000000000000_0001110110111111_0100101101010100"; -- 0.11620016859242843
	pesos_i(21108) := b"0000000000000000_0000000000000000_0010000000101011_1111010110110101"; -- 0.12567077320738493
	pesos_i(21109) := b"1111111111111111_1111111111111111_1101001011011000_0001011000110011"; -- -0.17639027840023194
	pesos_i(21110) := b"0000000000000000_0000000000000000_0001010111000010_0111001111100000"; -- 0.0849983617144504
	pesos_i(21111) := b"1111111111111111_1111111111111111_1111001100101011_0111001111110111"; -- -0.05011820996568223
	pesos_i(21112) := b"1111111111111111_1111111111111111_1110101100111011_1010001011010001"; -- -0.08112127674744138
	pesos_i(21113) := b"1111111111111111_1111111111111111_1111101110101101_0010010110111010"; -- -0.016889230761741654
	pesos_i(21114) := b"0000000000000000_0000000000000000_0001111100110000_1101011110001100"; -- 0.12183901957540906
	pesos_i(21115) := b"0000000000000000_0000000000000000_0001010011011001_0101010101101000"; -- 0.08144124773281569
	pesos_i(21116) := b"0000000000000000_0000000000000000_0001100100000101_0000111001101111"; -- 0.09773340436732549
	pesos_i(21117) := b"0000000000000000_0000000000000000_0010001010010110_1100110011011011"; -- 0.13511352880517657
	pesos_i(21118) := b"1111111111111111_1111111111111111_1111111001110000_0001011111011001"; -- -0.006102094128486646
	pesos_i(21119) := b"1111111111111111_1111111111111111_1111011000001001_1001110101101110"; -- -0.0389157872798881
	pesos_i(21120) := b"0000000000000000_0000000000000000_0000110001001100_1000111100010111"; -- 0.04804319690257442
	pesos_i(21121) := b"0000000000000000_0000000000000000_0001011111011110_0111111011001011"; -- 0.09323875863734159
	pesos_i(21122) := b"0000000000000000_0000000000000000_0001100100111010_0110011000111011"; -- 0.09854735316353896
	pesos_i(21123) := b"1111111111111111_1111111111111111_1110011000110000_1000111011101110"; -- -0.10082155892922876
	pesos_i(21124) := b"0000000000000000_0000000000000000_0001000011010011_1100010110000110"; -- 0.06573137791256178
	pesos_i(21125) := b"0000000000000000_0000000000000000_0001010001100000_1000001100000011"; -- 0.07959765277212832
	pesos_i(21126) := b"1111111111111111_1111111111111111_1111001010001000_0011011011100010"; -- -0.05260903349674788
	pesos_i(21127) := b"1111111111111111_1111111111111111_1101111000101111_1111111000111000"; -- -0.1320801841812608
	pesos_i(21128) := b"0000000000000000_0000000000000000_0001111101010101_1110000110111010"; -- 0.12240420133409606
	pesos_i(21129) := b"1111111111111111_1111111111111111_1101100110100010_0100100101110101"; -- -0.14986744786519773
	pesos_i(21130) := b"0000000000000000_0000000000000000_0000001110001111_0101010101000101"; -- 0.013905839225864443
	pesos_i(21131) := b"0000000000000000_0000000000000000_0001101010010010_1011100000110111"; -- 0.10380126323418634
	pesos_i(21132) := b"0000000000000000_0000000000000000_0001101100100111_0000010010000011"; -- 0.10606411167255528
	pesos_i(21133) := b"0000000000000000_0000000000000000_0001100110111111_0101100000000001"; -- 0.10057592405076594
	pesos_i(21134) := b"1111111111111111_1111111111111111_1110111111011101_0011101100110101"; -- -0.06303052851054136
	pesos_i(21135) := b"1111111111111111_1111111111111111_1111010000011111_0101111101001011"; -- -0.04639629755861248
	pesos_i(21136) := b"1111111111111111_1111111111111111_1111101001101100_0111110100101101"; -- -0.02178208962074643
	pesos_i(21137) := b"1111111111111111_1111111111111111_1111111111011000_0110011110010111"; -- -0.0006041770528730213
	pesos_i(21138) := b"0000000000000000_0000000000000000_0010101100000011_1101011011000000"; -- 0.1680273264381317
	pesos_i(21139) := b"0000000000000000_0000000000000000_0000111101010111_1111111000110101"; -- 0.059936416628844476
	pesos_i(21140) := b"1111111111111111_1111111111111111_1110111110111101_1110101001110011"; -- -0.06350836448909372
	pesos_i(21141) := b"1111111111111111_1111111111111111_1111011101100100_0011000100111101"; -- -0.0336274361831719
	pesos_i(21142) := b"1111111111111111_1111111111111111_1111111000001000_1110110110100001"; -- -0.007676265956774306
	pesos_i(21143) := b"0000000000000000_0000000000000000_0001100011001100_0100000001011101"; -- 0.0968666293653174
	pesos_i(21144) := b"1111111111111111_1111111111111111_1101011001010000_0001010011010111"; -- -0.16284055473438339
	pesos_i(21145) := b"0000000000000000_0000000000000000_0001111000100010_1010100000001110"; -- 0.11771631569557299
	pesos_i(21146) := b"1111111111111111_1111111111111111_1101111001100111_1001111101101001"; -- -0.13123134319368704
	pesos_i(21147) := b"0000000000000000_0000000000000000_0010010100111111_1010011000010000"; -- 0.1455024517138838
	pesos_i(21148) := b"0000000000000000_0000000000000000_0000110101001001_1000111110011010"; -- 0.051903700956295484
	pesos_i(21149) := b"1111111111111111_1111111111111111_1110001111001000_0100101010100110"; -- -0.11022504290834895
	pesos_i(21150) := b"1111111111111111_1111111111111111_1111111100011110_0101101110101010"; -- -0.003443022727056566
	pesos_i(21151) := b"0000000000000000_0000000000000000_0001011000100000_0110101000010011"; -- 0.08643210386995832
	pesos_i(21152) := b"1111111111111111_1111111111111111_1111100010110111_1111000010010000"; -- -0.028443302954057014
	pesos_i(21153) := b"0000000000000000_0000000000000000_0000011000010000_0111101100010011"; -- 0.023688976412158114
	pesos_i(21154) := b"1111111111111111_1111111111111111_1110001110001110_1000101010100010"; -- -0.11110623888287918
	pesos_i(21155) := b"0000000000000000_0000000000000000_0001001001000000_0011101100110110"; -- 0.07129259178848342
	pesos_i(21156) := b"1111111111111111_1111111111111111_1101111010000011_0111001110000011"; -- -0.13080671353659892
	pesos_i(21157) := b"0000000000000000_0000000000000000_0000110100011110_1101001111110110"; -- 0.05125164757264627
	pesos_i(21158) := b"0000000000000000_0000000000000000_0001011010011110_1111010111001100"; -- 0.08836303931552357
	pesos_i(21159) := b"1111111111111111_1111111111111111_1110111110010011_1101101110001010"; -- -0.06415012257015652
	pesos_i(21160) := b"0000000000000000_0000000000000000_0010001100111111_1101111010101111"; -- 0.1376933266628019
	pesos_i(21161) := b"1111111111111111_1111111111111111_1111010000010111_1001111111010100"; -- -0.04651452145069371
	pesos_i(21162) := b"0000000000000000_0000000000000000_0001101000000110_0010011111110111"; -- 0.10165643478713643
	pesos_i(21163) := b"0000000000000000_0000000000000000_0001011010101001_0101011110011011"; -- 0.08852145693140964
	pesos_i(21164) := b"0000000000000000_0000000000000000_0000101001001101_0101111010010110"; -- 0.04024306449331184
	pesos_i(21165) := b"1111111111111111_1111111111111111_1110111110011101_0101011111100010"; -- -0.06400538183869729
	pesos_i(21166) := b"1111111111111111_1111111111111111_1101100111011111_1101000111100000"; -- -0.14892853062885317
	pesos_i(21167) := b"1111111111111111_1111111111111111_1111100111111011_1100001010001011"; -- -0.023502198187936557
	pesos_i(21168) := b"1111111111111111_1111111111111111_1111111001000011_1001110101101110"; -- -0.006780777532474871
	pesos_i(21169) := b"1111111111111111_1111111111111111_1101111101100001_1101001010110011"; -- -0.12741358888544072
	pesos_i(21170) := b"1111111111111111_1111111111111111_1101110011010101_1010010100111001"; -- -0.1373650298936707
	pesos_i(21171) := b"0000000000000000_0000000000000000_0001001000000100_1000110110010011"; -- 0.07038197374708094
	pesos_i(21172) := b"0000000000000000_0000000000000000_0001110111110111_1001100011000001"; -- 0.1170592757584426
	pesos_i(21173) := b"1111111111111111_1111111111111111_1110111100110101_1011011110001111"; -- -0.06558659322607235
	pesos_i(21174) := b"0000000000000000_0000000000000000_0000001001111101_0011000000010101"; -- 0.009722714516152375
	pesos_i(21175) := b"1111111111111111_1111111111111111_1101111000000000_1011000100110101"; -- -0.1328019376954165
	pesos_i(21176) := b"0000000000000000_0000000000000000_0001101110110001_0001111101010100"; -- 0.10817142298030506
	pesos_i(21177) := b"0000000000000000_0000000000000000_0001100001110001_0110111000111000"; -- 0.0954808126733747
	pesos_i(21178) := b"1111111111111111_1111111111111111_1110101100111010_1110011100111000"; -- -0.08113245843512167
	pesos_i(21179) := b"0000000000000000_0000000000000000_0001000000100010_1011111001111011"; -- 0.06303015232652948
	pesos_i(21180) := b"1111111111111111_1111111111111111_1111110000000011_0110100011010000"; -- -0.01557297625124552
	pesos_i(21181) := b"0000000000000000_0000000000000000_0001010100111100_0100110011001001"; -- 0.08295135413343863
	pesos_i(21182) := b"1111111111111111_1111111111111111_1110100101110100_0001100011011011"; -- -0.08807224899734475
	pesos_i(21183) := b"1111111111111111_1111111111111111_1110101101000000_0101110110110110"; -- -0.0810491018989731
	pesos_i(21184) := b"0000000000000000_0000000000000000_0001100100010111_0010001011000100"; -- 0.09800927429910057
	pesos_i(21185) := b"1111111111111111_1111111111111111_1110001110111001_1011101011010110"; -- -0.11044723782731403
	pesos_i(21186) := b"0000000000000000_0000000000000000_0010000010000101_0011010110111010"; -- 0.12703262139401097
	pesos_i(21187) := b"1111111111111111_1111111111111111_1101100111111011_0011010010010110"; -- -0.14851065946860795
	pesos_i(21188) := b"1111111111111111_1111111111111111_1111101100010100_0000000010010010"; -- -0.01922604023051007
	pesos_i(21189) := b"0000000000000000_0000000000000000_0000101100100111_1100010000110111"; -- 0.04357553819315985
	pesos_i(21190) := b"1111111111111111_1111111111111111_1110010110000100_0111001110011111"; -- -0.10344769839945678
	pesos_i(21191) := b"1111111111111111_1111111111111111_1111011001100110_0101111000010010"; -- -0.0375004964053933
	pesos_i(21192) := b"0000000000000000_0000000000000000_0000011111100000_0110001010001111"; -- 0.030767593361253887
	pesos_i(21193) := b"0000000000000000_0000000000000000_0010100001101110_0100010000001000"; -- 0.15793252167883745
	pesos_i(21194) := b"1111111111111111_1111111111111111_1111010111100110_0000001000000101"; -- -0.03945910807155653
	pesos_i(21195) := b"1111111111111111_1111111111111111_1111111111010110_0100011010011111"; -- -0.0006366597223186571
	pesos_i(21196) := b"0000000000000000_0000000000000000_0001101111101101_1010001001111011"; -- 0.1090947675159928
	pesos_i(21197) := b"1111111111111111_1111111111111111_1110111100010100_0001001111100000"; -- -0.06609988968992898
	pesos_i(21198) := b"1111111111111111_1111111111111111_1111001001000000_0011101110000110"; -- -0.053707389562820444
	pesos_i(21199) := b"1111111111111111_1111111111111111_1101100011110010_1010000011001011"; -- -0.15254778908808278
	pesos_i(21200) := b"0000000000000000_0000000000000000_0000100100100001_1010111010100101"; -- 0.03567019963553456
	pesos_i(21201) := b"0000000000000000_0000000000000000_0000010101110010_0101100001100110"; -- 0.02127602091678579
	pesos_i(21202) := b"1111111111111111_1111111111111111_1110101110011000_1011011110010101"; -- -0.07970097174864885
	pesos_i(21203) := b"1111111111111111_1111111111111111_1111011110010110_0111010100110001"; -- -0.032860446448659514
	pesos_i(21204) := b"1111111111111111_1111111111111111_1111101000110010_0000010110001010"; -- -0.022674230336580736
	pesos_i(21205) := b"0000000000000000_0000000000000000_0010001101101101_0011110100011111"; -- 0.13838560116269574
	pesos_i(21206) := b"1111111111111111_1111111111111111_1101110111101101_0010110011110010"; -- -0.13309973793210086
	pesos_i(21207) := b"1111111111111111_1111111111111111_1110110101010110_0010101010100010"; -- -0.07290395291163071
	pesos_i(21208) := b"1111111111111111_1111111111111111_1110011000100111_1000111110010101"; -- -0.10095884899841259
	pesos_i(21209) := b"1111111111111111_1111111111111111_1111001011000000_0000010010101000"; -- -0.05175753496557106
	pesos_i(21210) := b"1111111111111111_1111111111111111_1101101100100100_0100111110111011"; -- -0.1439771811957442
	pesos_i(21211) := b"0000000000000000_0000000000000000_0010101010110010_1000011101010111"; -- 0.16678663144130332
	pesos_i(21212) := b"1111111111111111_1111111111111111_1111001100010110_0111101010011000"; -- -0.050438249375509364
	pesos_i(21213) := b"1111111111111111_1111111111111111_1110010000100011_1101010001000101"; -- -0.10882829019443072
	pesos_i(21214) := b"0000000000000000_0000000000000000_0001110001000100_1001000110111010"; -- 0.11042128352692214
	pesos_i(21215) := b"0000000000000000_0000000000000000_0001010001110010_1110111011000100"; -- 0.07987873353941394
	pesos_i(21216) := b"1111111111111111_1111111111111111_1110100111001001_1111110111111010"; -- -0.08676159510314191
	pesos_i(21217) := b"1111111111111111_1111111111111111_1101110001001100_0001100100000000"; -- -0.13946384187057137
	pesos_i(21218) := b"1111111111111111_1111111111111111_1110001010110010_0110110000111010"; -- -0.11446498479381992
	pesos_i(21219) := b"1111111111111111_1111111111111111_1101111001010111_0001000110001101"; -- -0.13148393916103995
	pesos_i(21220) := b"0000000000000000_0000000000000000_0001100111001110_0110000101101000"; -- 0.10080536641748752
	pesos_i(21221) := b"0000000000000000_0000000000000000_0000101110010010_0110110001101010"; -- 0.04520299511669371
	pesos_i(21222) := b"0000000000000000_0000000000000000_0000110000001110_0000010101011111"; -- 0.04708894323030532
	pesos_i(21223) := b"0000000000000000_0000000000000000_0001111011111101_1101010010001001"; -- 0.1210606417225851
	pesos_i(21224) := b"0000000000000000_0000000000000000_0010011000011111_1011000011010100"; -- 0.14892106230302216
	pesos_i(21225) := b"1111111111111111_1111111111111111_1110101001011101_1010100000100111"; -- -0.0845084099780791
	pesos_i(21226) := b"0000000000000000_0000000000000000_0001110110011100_1010011010000010"; -- 0.11567154562117732
	pesos_i(21227) := b"0000000000000000_0000000000000000_0000001000110101_0100111001101100"; -- 0.008625890039521607
	pesos_i(21228) := b"0000000000000000_0000000000000000_0000010110110110_1100001110011101"; -- 0.02232000899453147
	pesos_i(21229) := b"1111111111111111_1111111111111111_1111100101100100_1010011011001110"; -- -0.025807928826703085
	pesos_i(21230) := b"1111111111111111_1111111111111111_1110001100100011_1000111100101001"; -- -0.11273865937840608
	pesos_i(21231) := b"1111111111111111_1111111111111111_1111100010110000_0100110111100101"; -- -0.02855981028818843
	pesos_i(21232) := b"1111111111111111_1111111111111111_1101111011001110_1110010011010000"; -- -0.12965555116185942
	pesos_i(21233) := b"0000000000000000_0000000000000000_0010000101000101_1100000110010101"; -- 0.12997064491528246
	pesos_i(21234) := b"0000000000000000_0000000000000000_0000101011110100_1101010001100001"; -- 0.042798303251745676
	pesos_i(21235) := b"0000000000000000_0000000000000000_0010011110001101_0110110111111010"; -- 0.15450179439405373
	pesos_i(21236) := b"0000000000000000_0000000000000000_0001101011100100_0110000100111010"; -- 0.10504729904323121
	pesos_i(21237) := b"1111111111111111_1111111111111111_1110110110001010_0111101110101111"; -- -0.07210566500489896
	pesos_i(21238) := b"0000000000000000_0000000000000000_0010000000011101_0111010011100011"; -- 0.12544947187474428
	pesos_i(21239) := b"0000000000000000_0000000000000000_0000110101100101_1110010111111011"; -- 0.05233609571157247
	pesos_i(21240) := b"0000000000000000_0000000000000000_0000011100011101_0000010110101100"; -- 0.027786592923092518
	pesos_i(21241) := b"0000000000000000_0000000000000000_0000101100110111_1111010110111101"; -- 0.04382263055785892
	pesos_i(21242) := b"1111111111111111_1111111111111111_1101111000101001_0100001001101100"; -- -0.1321829304880556
	pesos_i(21243) := b"0000000000000000_0000000000000000_0001010010100010_0011011100001011"; -- 0.08060020471342652
	pesos_i(21244) := b"1111111111111111_1111111111111111_1110010010011010_1000101001000010"; -- -0.10701690560729119
	pesos_i(21245) := b"0000000000000000_0000000000000000_0001111000001100_0111100011111111"; -- 0.11737781745394216
	pesos_i(21246) := b"0000000000000000_0000000000000000_0001010111111001_1010000011100000"; -- 0.08584027748569961
	pesos_i(21247) := b"0000000000000000_0000000000000000_0001101101000111_1101100010000111"; -- 0.10656503000067429
	pesos_i(21248) := b"1111111111111111_1111111111111111_1110001011111011_1010101101101000"; -- -0.1133473273707008
	pesos_i(21249) := b"1111111111111111_1111111111111111_1111010001100011_1111110011110100"; -- -0.04534930267736335
	pesos_i(21250) := b"0000000000000000_0000000000000000_0000010111010110_1010001010010110"; -- 0.022806321821210587
	pesos_i(21251) := b"0000000000000000_0000000000000000_0000001000100000_0100000011011000"; -- 0.008304646325943051
	pesos_i(21252) := b"1111111111111111_1111111111111111_1111100111100111_1001110110101011"; -- -0.02380957208800427
	pesos_i(21253) := b"0000000000000000_0000000000000000_0000110000111000_0011010110101001"; -- 0.04773269068777427
	pesos_i(21254) := b"0000000000000000_0000000000000000_0000110001100101_1110101000011010"; -- 0.048430091313514056
	pesos_i(21255) := b"1111111111111111_1111111111111111_1101100011011110_1100111000110111"; -- -0.1528502574692385
	pesos_i(21256) := b"1111111111111111_1111111111111111_1111000010100101_1100110100011001"; -- -0.0599700749917893
	pesos_i(21257) := b"0000000000000000_0000000000000000_0000000110000011_1101000001100001"; -- 0.0059175717264808025
	pesos_i(21258) := b"0000000000000000_0000000000000000_0010001000111100_0000101001000001"; -- 0.13372863841259625
	pesos_i(21259) := b"1111111111111111_1111111111111111_1101110100100000_1111001100100110"; -- -0.13621597598532412
	pesos_i(21260) := b"0000000000000000_0000000000000000_0000101101110100_1001010111101000"; -- 0.044747704682791066
	pesos_i(21261) := b"0000000000000000_0000000000000000_0001110111001110_0001101011110101"; -- 0.11642616725944385
	pesos_i(21262) := b"0000000000000000_0000000000000000_0000011001101011_0111111001001111"; -- 0.025077718949358667
	pesos_i(21263) := b"1111111111111111_1111111111111111_1101101110100000_0111011101110011"; -- -0.14208272398137564
	pesos_i(21264) := b"1111111111111111_1111111111111111_1101101001111100_0100011101011001"; -- -0.14654115757183653
	pesos_i(21265) := b"1111111111111111_1111111111111111_1111010101001011_1101001010000110"; -- -0.04181179258873133
	pesos_i(21266) := b"1111111111111111_1111111111111111_1110100101111101_0101011101000010"; -- -0.08793120040995735
	pesos_i(21267) := b"1111111111111111_1111111111111111_1101101010011110_1111111110000001"; -- -0.14601138201045696
	pesos_i(21268) := b"1111111111111111_1111111111111111_1101101110001010_1000111001101110"; -- -0.14241704767163524
	pesos_i(21269) := b"1111111111111111_1111111111111111_1111111001100011_1000111110101001"; -- -0.006293317048161218
	pesos_i(21270) := b"1111111111111111_1111111111111111_1110100000101010_0111111001110000"; -- -0.09310159468986347
	pesos_i(21271) := b"1111111111111111_1111111111111111_1101110001111111_1010001101111111"; -- -0.13867738870825094
	pesos_i(21272) := b"1111111111111111_1111111111111111_1111001011110011_0001000110111000"; -- -0.05097855811753171
	pesos_i(21273) := b"1111111111111111_1111111111111111_1110110100111000_0101101011000110"; -- -0.07335884738883841
	pesos_i(21274) := b"0000000000000000_0000000000000000_0001010001100110_0010100001110011"; -- 0.07968380754058084
	pesos_i(21275) := b"1111111111111111_1111111111111111_1111011101101011_0110010100011100"; -- -0.033517532891834595
	pesos_i(21276) := b"1111111111111111_1111111111111111_1110111000010010_1000101101011000"; -- -0.07002953621269063
	pesos_i(21277) := b"0000000000000000_0000000000000000_0001100111001110_1101000011111001"; -- 0.10081201637564866
	pesos_i(21278) := b"1111111111111111_1111111111111111_1110010011001001_1110010000101100"; -- -0.10629438326606241
	pesos_i(21279) := b"0000000000000000_0000000000000000_0001010011100001_1101100010110111"; -- 0.08157114482981526
	pesos_i(21280) := b"1111111111111111_1111111111111111_1101110100010000_0100100111101111"; -- -0.13647020267158924
	pesos_i(21281) := b"0000000000000000_0000000000000000_0000110010101110_0011110001010100"; -- 0.04953362519320367
	pesos_i(21282) := b"0000000000000000_0000000000000000_0000101110101010_1011100101101101"; -- 0.04557379649139124
	pesos_i(21283) := b"0000000000000000_0000000000000000_0001101111000110_0100000111011011"; -- 0.10849391563974031
	pesos_i(21284) := b"0000000000000000_0000000000000000_0001000011110000_1111100101111010"; -- 0.06617697930650279
	pesos_i(21285) := b"0000000000000000_0000000000000000_0000101000011110_1000101111100101"; -- 0.03952860210454216
	pesos_i(21286) := b"0000000000000000_0000000000000000_0001100101101001_0011010110100001"; -- 0.09926161949443385
	pesos_i(21287) := b"0000000000000000_0000000000000000_0000100000000011_1101010101110110"; -- 0.03130849974009887
	pesos_i(21288) := b"1111111111111111_1111111111111111_1111000011111001_0010111011101011"; -- -0.058697764917039104
	pesos_i(21289) := b"1111111111111111_1111111111111111_1110000000100001_1110110100011101"; -- -0.12448232692826211
	pesos_i(21290) := b"0000000000000000_0000000000000000_0000011010100110_0100100110101111"; -- 0.025974850883392072
	pesos_i(21291) := b"1111111111111111_1111111111111111_1111111011001100_0011101010101100"; -- -0.004696210016771211
	pesos_i(21292) := b"0000000000000000_0000000000000000_0001001011100011_1111100011010011"; -- 0.07379107629269335
	pesos_i(21293) := b"1111111111111111_1111111111111111_1110110110001011_1110011010001011"; -- -0.07208403689188833
	pesos_i(21294) := b"0000000000000000_0000000000000000_0010000000101011_1101010101111000"; -- 0.12566885155937205
	pesos_i(21295) := b"1111111111111111_1111111111111111_1110111100001111_0000011011001101"; -- -0.06617696279555994
	pesos_i(21296) := b"1111111111111111_1111111111111111_1110000000111000_1110000010100111"; -- -0.124132117566368
	pesos_i(21297) := b"1111111111111111_1111111111111111_1110011011110011_0010101011100100"; -- -0.0978520577495677
	pesos_i(21298) := b"0000000000000000_0000000000000000_0000011111110101_0010100000011100"; -- 0.031084544127222332
	pesos_i(21299) := b"0000000000000000_0000000000000000_0010011001001101_0100110101101010"; -- 0.1496170408802201
	pesos_i(21300) := b"0000000000000000_0000000000000000_0001111011001111_0000000010011011"; -- 0.12034610542158022
	pesos_i(21301) := b"0000000000000000_0000000000000000_0000000001111100_0100000000001000"; -- 0.001895906516118643
	pesos_i(21302) := b"0000000000000000_0000000000000000_0001010011011001_1010101110110101"; -- 0.08144639173329488
	pesos_i(21303) := b"0000000000000000_0000000000000000_0000010001001111_1101001111010001"; -- 0.016843069491413544
	pesos_i(21304) := b"1111111111111111_1111111111111111_1110101100110100_0010101101100111"; -- -0.08123520595073427
	pesos_i(21305) := b"1111111111111111_1111111111111111_1111110010110001_1111000100001100"; -- -0.01290982691008944
	pesos_i(21306) := b"0000000000000000_0000000000000000_0001111101100011_1001010100111010"; -- 0.12261326460188526
	pesos_i(21307) := b"1111111111111111_1111111111111111_1111000101011000_0001110001001101"; -- -0.05724928972149144
	pesos_i(21308) := b"1111111111111111_1111111111111111_1110011101011101_1001100110001101"; -- -0.0962280302794706
	pesos_i(21309) := b"0000000000000000_0000000000000000_0001010010001110_0001011000110001"; -- 0.08029307069625674
	pesos_i(21310) := b"0000000000000000_0000000000000000_0000000011011000_1001110101000110"; -- 0.003305272744496688
	pesos_i(21311) := b"0000000000000000_0000000000000000_0000100101000010_1100101101111010"; -- 0.03617545831735303
	pesos_i(21312) := b"1111111111111111_1111111111111111_1110010000011000_1101000111000010"; -- -0.10899628657808909
	pesos_i(21313) := b"0000000000000000_0000000000000000_0001001010000010_1011000001001101"; -- 0.0723066508110393
	pesos_i(21314) := b"1111111111111111_1111111111111111_1111110100100100_0100111110111011"; -- -0.011164681177545684
	pesos_i(21315) := b"1111111111111111_1111111111111111_1111101101001101_1011011101100100"; -- -0.018345392245248275
	pesos_i(21316) := b"1111111111111111_1111111111111111_1101101100100001_0111110110110011"; -- -0.14402021779389504
	pesos_i(21317) := b"1111111111111111_1111111111111111_1101101000101101_0010001000001011"; -- -0.14774882532646083
	pesos_i(21318) := b"1111111111111111_1111111111111111_1111010011101000_0000001100101010"; -- -0.043334772430237374
	pesos_i(21319) := b"1111111111111111_1111111111111111_1111001111010001_1011110001100010"; -- -0.04758093457879921
	pesos_i(21320) := b"1111111111111111_1111111111111111_1101101010001111_1000110010011001"; -- -0.14624711287007325
	pesos_i(21321) := b"0000000000000000_0000000000000000_0000001101010100_1101011111101100"; -- 0.013013358126614482
	pesos_i(21322) := b"1111111111111111_1111111111111111_1110010100000100_1110001101010010"; -- -0.10539416554643967
	pesos_i(21323) := b"0000000000000000_0000000000000000_0001001100010000_0101000100111011"; -- 0.07446773223859175
	pesos_i(21324) := b"0000000000000000_0000000000000000_0001101110010100_0110010001100111"; -- 0.1077330351186164
	pesos_i(21325) := b"1111111111111111_1111111111111111_1111010000000011_0100011000010001"; -- -0.04682504726177249
	pesos_i(21326) := b"0000000000000000_0000000000000000_0010010101010110_1010100010001110"; -- 0.14585355261601768
	pesos_i(21327) := b"0000000000000000_0000000000000000_0000001110100100_1001011111110101"; -- 0.014230248855578422
	pesos_i(21328) := b"1111111111111111_1111111111111111_1101100101110110_1110111100101100"; -- -0.1505289571334295
	pesos_i(21329) := b"1111111111111111_1111111111111111_1110110110000110_0111011010001100"; -- -0.07216700624972401
	pesos_i(21330) := b"1111111111111111_1111111111111111_1110110111100111_1111110101011110"; -- -0.07067886781400885
	pesos_i(21331) := b"0000000000000000_0000000000000000_0001011010010000_0110110111111001"; -- 0.08814132042905855
	pesos_i(21332) := b"1111111111111111_1111111111111111_1111011111010110_0100011100101001"; -- -0.03188662757237954
	pesos_i(21333) := b"1111111111111111_1111111111111111_1110100010011110_1001100100111111"; -- -0.09132997717158123
	pesos_i(21334) := b"1111111111111111_1111111111111111_1110110111011011_0111110101011001"; -- -0.07086960381570738
	pesos_i(21335) := b"1111111111111111_1111111111111111_1111101010011100_0011001011001000"; -- -0.021054102029295394
	pesos_i(21336) := b"0000000000000000_0000000000000000_0000011001100101_1101000100011001"; -- 0.02499110085740196
	pesos_i(21337) := b"0000000000000000_0000000000000000_0010000110101110_1001000101000111"; -- 0.13156993848636758
	pesos_i(21338) := b"0000000000000000_0000000000000000_0001111100001111_0101101000000010"; -- 0.12132799673965869
	pesos_i(21339) := b"0000000000000000_0000000000000000_0001101111110000_0110011010000000"; -- 0.10913696874361672
	pesos_i(21340) := b"1111111111111111_1111111111111111_1111010010000110_0100011111100000"; -- -0.04482603812649885
	pesos_i(21341) := b"0000000000000000_0000000000000000_0000000011000001_0011010011100101"; -- 0.002948098944962433
	pesos_i(21342) := b"1111111111111111_1111111111111111_1111001110110000_1000111111111101"; -- -0.04808712082625312
	pesos_i(21343) := b"0000000000000000_0000000000000000_0001001000001110_0111001000110100"; -- 0.07053293004217527
	pesos_i(21344) := b"1111111111111111_1111111111111111_1110000001011010_0010100011101011"; -- -0.1236242701606042
	pesos_i(21345) := b"1111111111111111_1111111111111111_1110101111111000_1000011100100110"; -- -0.07823901474223728
	pesos_i(21346) := b"0000000000000000_0000000000000000_0001100110001111_0001011110010110"; -- 0.09983966269694024
	pesos_i(21347) := b"0000000000000000_0000000000000000_0001100111000011_1001110011000000"; -- 0.10064105698137599
	pesos_i(21348) := b"0000000000000000_0000000000000000_0000101101011100_1001100110110110"; -- 0.044381720586107086
	pesos_i(21349) := b"0000000000000000_0000000000000000_0001010110111101_0111001101010010"; -- 0.08492203482643298
	pesos_i(21350) := b"0000000000000000_0000000000000000_0000000011010111_0010101111100000"; -- 0.0032832547251812993
	pesos_i(21351) := b"0000000000000000_0000000000000000_0010001101110001_1110101101000110"; -- 0.13845701663480192
	pesos_i(21352) := b"1111111111111111_1111111111111111_1111110101010001_0111101101010101"; -- -0.010475436924248563
	pesos_i(21353) := b"1111111111111111_1111111111111111_1111101110111001_1100010100100100"; -- -0.01669662341479161
	pesos_i(21354) := b"1111111111111111_1111111111111111_1101110001111101_1001100000010100"; -- -0.13870858670169864
	pesos_i(21355) := b"1111111111111111_1111111111111111_1110010100110100_1001011101101100"; -- -0.1046662675537968
	pesos_i(21356) := b"0000000000000000_0000000000000000_0000011101110101_1100010001111010"; -- 0.02914073915777957
	pesos_i(21357) := b"0000000000000000_0000000000000000_0001010110001100_1111101100011101"; -- 0.0841824480629358
	pesos_i(21358) := b"1111111111111111_1111111111111111_1111000011101110_1011011001100100"; -- -0.05885753684311535
	pesos_i(21359) := b"0000000000000000_0000000000000000_0001110101111011_0110010010101110"; -- 0.11516408211738605
	pesos_i(21360) := b"0000000000000000_0000000000000000_0010001111111000_1111101011000011"; -- 0.1405178763634709
	pesos_i(21361) := b"0000000000000000_0000000000000000_0000100101010011_1110010010011110"; -- 0.03643635615257173
	pesos_i(21362) := b"0000000000000000_0000000000000000_0001010110101011_1110010101010000"; -- 0.08465417091383892
	pesos_i(21363) := b"1111111111111111_1111111111111111_1110110100111111_1100010111000010"; -- -0.07324565891089511
	pesos_i(21364) := b"1111111111111111_1111111111111111_1111110110000011_1100110011101000"; -- -0.009707635244984811
	pesos_i(21365) := b"0000000000000000_0000000000000000_0000000111011101_0100101101100110"; -- 0.007282936471370643
	pesos_i(21366) := b"1111111111111111_1111111111111111_1101101011000100_1101001000001001"; -- -0.14543425837682952
	pesos_i(21367) := b"1111111111111111_1111111111111111_1111110110000110_1110000100111101"; -- -0.00966064699891973
	pesos_i(21368) := b"1111111111111111_1111111111111111_1111001010000001_0110101110010000"; -- -0.05271270488361271
	pesos_i(21369) := b"0000000000000000_0000000000000000_0000100011000110_1101111001110011"; -- 0.034284499238688065
	pesos_i(21370) := b"0000000000000000_0000000000000000_0001100110000110_1011110010110101"; -- 0.09971217554744533
	pesos_i(21371) := b"0000000000000000_0000000000000000_0000101010000111_1101001100100101"; -- 0.041135021815895324
	pesos_i(21372) := b"1111111111111111_1111111111111111_1111111011111000_1100001011011011"; -- -0.004016705920773391
	pesos_i(21373) := b"1111111111111111_1111111111111111_1101101100111101_1011100011011001"; -- -0.14358944598566645
	pesos_i(21374) := b"1111111111111111_1111111111111111_1111111000000001_1100001011110000"; -- -0.007785622071020136
	pesos_i(21375) := b"0000000000000000_0000000000000000_0001011100111100_1000101010111010"; -- 0.09076754611080493
	pesos_i(21376) := b"1111111111111111_1111111111111111_1111101011001010_0101010000110011"; -- -0.020350205870247166
	pesos_i(21377) := b"1111111111111111_1111111111111111_1110110000100000_1101111000100010"; -- -0.07762347860089572
	pesos_i(21378) := b"1111111111111111_1111111111111111_1101011111000100_1111011100110010"; -- -0.15715079344959362
	pesos_i(21379) := b"0000000000000000_0000000000000000_0000010111100101_0100101101101000"; -- 0.023030007226975336
	pesos_i(21380) := b"1111111111111111_1111111111111111_1110101110001010_1111101111101001"; -- -0.07991052198022337
	pesos_i(21381) := b"1111111111111111_1111111111111111_1110001001001010_0111100100111101"; -- -0.11605112315969601
	pesos_i(21382) := b"1111111111111111_1111111111111111_1101101001000001_1000000111001100"; -- -0.14743794230819782
	pesos_i(21383) := b"0000000000000000_0000000000000000_0001110001100010_1011001011000110"; -- 0.11088101709919027
	pesos_i(21384) := b"0000000000000000_0000000000000000_0001001011111000_1010111101000111"; -- 0.07410712704891789
	pesos_i(21385) := b"1111111111111111_1111111111111111_1110011100011011_1010100000000001"; -- -0.09723424878051767
	pesos_i(21386) := b"0000000000000000_0000000000000000_0010001010100101_0100010101101101"; -- 0.13533433827550595
	pesos_i(21387) := b"0000000000000000_0000000000000000_0000011101010111_1011101000110011"; -- 0.02868236288397285
	pesos_i(21388) := b"1111111111111111_1111111111111111_1111011011000000_1011111000101100"; -- -0.03612147732055585
	pesos_i(21389) := b"0000000000000000_0000000000000000_0000000010011001_0111111101111010"; -- 0.00234219283867329
	pesos_i(21390) := b"1111111111111111_1111111111111111_1111010110100110_1100010101001000"; -- -0.04042403210752598
	pesos_i(21391) := b"0000000000000000_0000000000000000_0001110000100111_0011100110110011"; -- 0.1099735319678931
	pesos_i(21392) := b"0000000000000000_0000000000000000_0001010001010000_1001101011111000"; -- 0.07935494005250489
	pesos_i(21393) := b"1111111111111111_1111111111111111_1101111111011100_0100101100001010"; -- -0.12554484372030203
	pesos_i(21394) := b"1111111111111111_1111111111111111_1111110000110011_0001000001101100"; -- -0.014845822889449248
	pesos_i(21395) := b"0000000000000000_0000000000000000_0001111101111001_0011010011100101"; -- 0.12294321620374667
	pesos_i(21396) := b"1111111111111111_1111111111111111_1110001000110010_1101001000100001"; -- -0.11641203592718714
	pesos_i(21397) := b"0000000000000000_0000000000000000_0000001000111100_1011110000111010"; -- 0.008739246555565431
	pesos_i(21398) := b"1111111111111111_1111111111111111_1110010000111001_0010101100101010"; -- -0.10850267633744563
	pesos_i(21399) := b"1111111111111111_1111111111111111_1110000110111000_1001100010001000"; -- -0.11827704129061911
	pesos_i(21400) := b"0000000000000000_0000000000000000_0010101000000111_1011010101011001"; -- 0.16418012076448277
	pesos_i(21401) := b"0000000000000000_0000000000000000_0001000100010111_0110111110010100"; -- 0.0667638528139748
	pesos_i(21402) := b"1111111111111111_1111111111111111_1101101011010111_0001100001011100"; -- -0.14515540838118948
	pesos_i(21403) := b"1111111111111111_1111111111111111_1111100001101111_0011111100001000"; -- -0.02955251752528504
	pesos_i(21404) := b"1111111111111111_1111111111111111_1110110001001110_0101011111101001"; -- -0.07692957456559295
	pesos_i(21405) := b"0000000000000000_0000000000000000_0000100110100011_1101010011101010"; -- 0.037656123275981335
	pesos_i(21406) := b"0000000000000000_0000000000000000_0001110110000111_0011001110101010"; -- 0.11534426600062019
	pesos_i(21407) := b"1111111111111111_1111111111111111_1101111101001011_1100010100111001"; -- -0.12775008547444075
	pesos_i(21408) := b"1111111111111111_1111111111111111_1111010110110010_0111011100001001"; -- -0.04024559046443557
	pesos_i(21409) := b"1111111111111111_1111111111111111_1101111000011100_1001011111111101"; -- -0.13237619460248054
	pesos_i(21410) := b"1111111111111111_1111111111111111_1101100001101001_0010001110011001"; -- -0.1546457053993192
	pesos_i(21411) := b"1111111111111111_1111111111111111_1111010111101011_0111100101011010"; -- -0.03937570145768641
	pesos_i(21412) := b"1111111111111111_1111111111111111_1110000100011101_1110001111100011"; -- -0.12063766198407538
	pesos_i(21413) := b"0000000000000000_0000000000000000_0000101011000010_0100100010011110"; -- 0.04202703333165799
	pesos_i(21414) := b"0000000000000000_0000000000000000_0010011011000110_0110011000101101"; -- 0.15146483029642874
	pesos_i(21415) := b"1111111111111111_1111111111111111_1110011010110010_0111000101001010"; -- -0.09883968298492062
	pesos_i(21416) := b"1111111111111111_1111111111111111_1111001111110001_0011100111111010"; -- -0.04710042612601246
	pesos_i(21417) := b"1111111111111111_1111111111111111_1101101100100111_0110010011101000"; -- -0.14393014269530263
	pesos_i(21418) := b"0000000000000000_0000000000000000_0010000111101010_1100001010000010"; -- 0.13248840020686453
	pesos_i(21419) := b"0000000000000000_0000000000000000_0010101010110001_0010010000111111"; -- 0.1667654660973818
	pesos_i(21420) := b"1111111111111111_1111111111111111_1111110111010011_0011101010101111"; -- -0.008495647700350774
	pesos_i(21421) := b"0000000000000000_0000000000000000_0000000100110101_0011100110000101"; -- 0.004718394139275772
	pesos_i(21422) := b"0000000000000000_0000000000000000_0000000110001000_1111100000100000"; -- 0.005996234774633974
	pesos_i(21423) := b"0000000000000000_0000000000000000_0000100001110000_1001111111000111"; -- 0.032968507954158156
	pesos_i(21424) := b"1111111111111111_1111111111111111_1111011000010010_0010100000011011"; -- -0.038785451414723275
	pesos_i(21425) := b"1111111111111111_1111111111111111_1111010001010101_0101110001011110"; -- -0.04557249746216671
	pesos_i(21426) := b"1111111111111111_1111111111111111_1111011110000100_1101010101000111"; -- -0.0331293774218826
	pesos_i(21427) := b"1111111111111111_1111111111111111_1111001000010010_0110110110010101"; -- -0.05440631028454863
	pesos_i(21428) := b"1111111111111111_1111111111111111_1111000100010011_0011010011100101"; -- -0.058300680208867556
	pesos_i(21429) := b"1111111111111111_1111111111111111_1110101101010000_0101001111110100"; -- -0.08080554290302135
	pesos_i(21430) := b"0000000000000000_0000000000000000_0011001011001011_0111011110101110"; -- 0.1984171675757534
	pesos_i(21431) := b"0000000000000000_0000000000000000_0000011001110011_1001011001010010"; -- 0.02520122049216406
	pesos_i(21432) := b"1111111111111111_1111111111111111_1101111110001111_1011000011001000"; -- -0.12671370614444252
	pesos_i(21433) := b"0000000000000000_0000000000000000_0000000101110010_1001110110010011"; -- 0.005655144159543237
	pesos_i(21434) := b"1111111111111111_1111111111111111_1101111001000111_1010010001101000"; -- -0.1317193265575804
	pesos_i(21435) := b"1111111111111111_1111111111111111_1110101110100101_1010010010011001"; -- -0.07950373910466416
	pesos_i(21436) := b"1111111111111111_1111111111111111_1101101100101000_1101011010101101"; -- -0.14390810271493915
	pesos_i(21437) := b"0000000000000000_0000000000000000_0001111010010100_1100000000010100"; -- 0.11945724944263754
	pesos_i(21438) := b"1111111111111111_1111111111111111_1111010000011011_1101010001100110"; -- -0.04645035286952089
	pesos_i(21439) := b"1111111111111111_1111111111111111_1101100100110011_0111011000011000"; -- -0.1515585127810358
	pesos_i(21440) := b"0000000000000000_0000000000000000_0000110011111111_0001010100000000"; -- 0.05076724287700812
	pesos_i(21441) := b"0000000000000000_0000000000000000_0001011110110011_1010111000100001"; -- 0.09258545206627805
	pesos_i(21442) := b"0000000000000000_0000000000000000_0001001101101001_1111010010100110"; -- 0.07583550495085836
	pesos_i(21443) := b"0000000000000000_0000000000000000_0001101110110010_0000011101001010"; -- 0.10818524881975349
	pesos_i(21444) := b"0000000000000000_0000000000000000_0010010010001101_0101011110011100"; -- 0.14278171128525158
	pesos_i(21445) := b"0000000000000000_0000000000000000_0000110010010010_1100001110101100"; -- 0.049114446094850106
	pesos_i(21446) := b"0000000000000000_0000000000000000_0000010011101100_1111101000000000"; -- 0.01924097526730937
	pesos_i(21447) := b"0000000000000000_0000000000000000_0000010010110101_0110100000010100"; -- 0.018393044456887213
	pesos_i(21448) := b"0000000000000000_0000000000000000_0000101111111001_1011010010010101"; -- 0.04677895201695329
	pesos_i(21449) := b"1111111111111111_1111111111111111_1110110011001101_0000100110010110"; -- -0.0749963769675049
	pesos_i(21450) := b"1111111111111111_1111111111111111_1110010000101111_0110100110111100"; -- -0.10865153467575882
	pesos_i(21451) := b"0000000000000000_0000000000000000_0000011010010001_1010010010110000"; -- 0.025659840502963743
	pesos_i(21452) := b"0000000000000000_0000000000000000_0001100010100001_1101110000001110"; -- 0.0962197812640244
	pesos_i(21453) := b"1111111111111111_1111111111111111_1111110000010010_0101010010101011"; -- -0.015345295145036866
	pesos_i(21454) := b"0000000000000000_0000000000000000_0001101100100100_1111111001001001"; -- 0.10603322296880906
	pesos_i(21455) := b"1111111111111111_1111111111111111_1111011111001101_1001000101110001"; -- -0.03201952918265639
	pesos_i(21456) := b"1111111111111111_1111111111111111_1110111000100001_0101000011101010"; -- -0.0698041371313089
	pesos_i(21457) := b"1111111111111111_1111111111111111_1111001011001111_0011100000101001"; -- -0.051525583319569745
	pesos_i(21458) := b"1111111111111111_1111111111111111_1110110011111011_1010010101111000"; -- -0.07428518116230533
	pesos_i(21459) := b"0000000000000000_0000000000000000_0000101110101001_1111010011001001"; -- 0.045562075611156036
	pesos_i(21460) := b"1111111111111111_1111111111111111_1111001100010100_1011111000010110"; -- -0.05046474427255924
	pesos_i(21461) := b"0000000000000000_0000000000000000_0001000111010000_1101011101111101"; -- 0.06959292222736829
	pesos_i(21462) := b"0000000000000000_0000000000000000_0001111011110110_0101010101110001"; -- 0.1209462548680451
	pesos_i(21463) := b"0000000000000000_0000000000000000_0010000110001110_1101111101000101"; -- 0.1310863058756062
	pesos_i(21464) := b"1111111111111111_1111111111111111_1101100101110011_1011101101110100"; -- -0.1505778161782591
	pesos_i(21465) := b"0000000000000000_0000000000000000_0000000111010101_0110101110100110"; -- 0.007162788382245375
	pesos_i(21466) := b"1111111111111111_1111111111111111_1110111101010100_0001010011010101"; -- -0.06512327004286896
	pesos_i(21467) := b"1111111111111111_1111111111111111_1110001110100000_0100110110101100"; -- -0.11083521403838369
	pesos_i(21468) := b"1111111111111111_1111111111111111_1111101011001000_1001111101000011"; -- -0.02037624946737228
	pesos_i(21469) := b"1111111111111111_1111111111111111_1110000110000001_0001000000111101"; -- -0.11912439841326583
	pesos_i(21470) := b"1111111111111111_1111111111111111_1110011010011001_1100000010111111"; -- -0.09921641677355175
	pesos_i(21471) := b"0000000000000000_0000000000000000_0010000000100111_1100000001110101"; -- 0.1256065641738312
	pesos_i(21472) := b"1111111111111111_1111111111111111_1111100010011111_0010010101110111"; -- -0.028821619498281405
	pesos_i(21473) := b"0000000000000000_0000000000000000_0001011001101011_1000010101001100"; -- 0.08757813547313735
	pesos_i(21474) := b"0000000000000000_0000000000000000_0010001100101111_0101001100101010"; -- 0.1374408700073513
	pesos_i(21475) := b"1111111111111111_1111111111111111_1110111101111101_1011110100000001"; -- -0.06448763584455411
	pesos_i(21476) := b"0000000000000000_0000000000000000_0001011110011110_0110011011010100"; -- 0.09226076768759146
	pesos_i(21477) := b"0000000000000000_0000000000000000_0001111110001000_0011101011111100"; -- 0.1231724611661593
	pesos_i(21478) := b"0000000000000000_0000000000000000_0001111010001000_1010010111110110"; -- 0.11927258728845028
	pesos_i(21479) := b"1111111111111111_1111111111111111_1111001111101010_0110111111011001"; -- -0.04720402681868727
	pesos_i(21480) := b"1111111111111111_1111111111111111_1110011100000000_1101101001000001"; -- -0.09764324110531596
	pesos_i(21481) := b"0000000000000000_0000000000000000_0001010111010010_0010111111110001"; -- 0.0852384532587912
	pesos_i(21482) := b"0000000000000000_0000000000000000_0001000011011110_0110010111100101"; -- 0.06589352454963239
	pesos_i(21483) := b"0000000000000000_0000000000000000_0000011101111101_0110010010011000"; -- 0.029257094431080467
	pesos_i(21484) := b"0000000000000000_0000000000000000_0000000111100101_1100100110000111"; -- 0.007412524549295944
	pesos_i(21485) := b"0000000000000000_0000000000000000_0000010010100110_1111100011111001"; -- 0.018172798973401023
	pesos_i(21486) := b"0000000000000000_0000000000000000_0000110010111110_1011100100011001"; -- 0.04978520255057876
	pesos_i(21487) := b"1111111111111111_1111111111111111_1111100011111011_0110111100101101"; -- -0.027413417333917025
	pesos_i(21488) := b"1111111111111111_1111111111111111_1111000011101001_1010000110110011"; -- -0.05893506416138697
	pesos_i(21489) := b"1111111111111111_1111111111111111_1111000010001101_0000001101101010"; -- -0.060348307359698594
	pesos_i(21490) := b"1111111111111111_1111111111111111_1111010000000001_1101011000111001"; -- -0.04684697255832832
	pesos_i(21491) := b"0000000000000000_0000000000000000_0001010011110111_1100110001010001"; -- 0.08190609909252534
	pesos_i(21492) := b"1111111111111111_1111111111111111_1111111010101100_1100110000001101"; -- -0.005175825903079077
	pesos_i(21493) := b"0000000000000000_0000000000000000_0000101111011110_1001101001110001"; -- 0.04636540668986603
	pesos_i(21494) := b"0000000000000000_0000000000000000_0000011001001010_0101000101000110"; -- 0.024571494773344763
	pesos_i(21495) := b"1111111111111111_1111111111111111_1110101000110100_0100101001011111"; -- -0.0851396099911927
	pesos_i(21496) := b"1111111111111111_1111111111111111_1110001000001110_1100000011010101"; -- -0.11696238326575756
	pesos_i(21497) := b"1111111111111111_1111111111111111_1101111111110101_0111000001110111"; -- -0.12516114324909428
	pesos_i(21498) := b"1111111111111111_1111111111111111_1101011000101011_0110011010001011"; -- -0.16340025991808863
	pesos_i(21499) := b"1111111111111111_1111111111111111_1111000100101011_1011010101111111"; -- -0.05792680415774783
	pesos_i(21500) := b"1111111111111111_1111111111111111_1110010101100011_0001000010000011"; -- -0.10395714573150051
	pesos_i(21501) := b"1111111111111111_1111111111111111_1110101001001000_1111001101011001"; -- -0.08482436253538739
	pesos_i(21502) := b"0000000000000000_0000000000000000_0001111001001000_0000000101101000"; -- 0.1182862166077444
	pesos_i(21503) := b"0000000000000000_0000000000000000_0001011001111110_0100100011001011"; -- 0.0878644461279982
	pesos_i(21504) := b"1111111111111111_1111111111111111_1110110011110010_1100101001001110"; -- -0.07442031479179248
	pesos_i(21505) := b"1111111111111111_1111111111111111_1111101101100000_1101111101101011"; -- -0.01805308956124098
	pesos_i(21506) := b"0000000000000000_0000000000000000_0001110100001000_0101100101111011"; -- 0.11340865379350129
	pesos_i(21507) := b"0000000000000000_0000000000000000_0000101111111110_1001101100110111"; -- 0.04685373402831459
	pesos_i(21508) := b"0000000000000000_0000000000000000_0000100000011000_1111001010111101"; -- 0.03163067936308322
	pesos_i(21509) := b"0000000000000000_0000000000000000_0000100101001011_1010001010101000"; -- 0.0363103541778187
	pesos_i(21510) := b"0000000000000000_0000000000000000_0010010001111101_0110000111010111"; -- 0.1425381804297811
	pesos_i(21511) := b"0000000000000000_0000000000000000_0000100110101000_0001101000010010"; -- 0.037721280435378285
	pesos_i(21512) := b"1111111111111111_1111111111111111_1111011111110100_0100111100010010"; -- -0.031428392599526116
	pesos_i(21513) := b"1111111111111111_1111111111111111_1110011001111011_1001100000001011"; -- -0.09967660656910443
	pesos_i(21514) := b"1111111111111111_1111111111111111_1111110011101010_0111100010000110"; -- -0.012047259611225623
	pesos_i(21515) := b"1111111111111111_1111111111111111_1111010111110010_0110010001100000"; -- -0.03927014023515996
	pesos_i(21516) := b"1111111111111111_1111111111111111_1110001000001100_1000111110011101"; -- -0.11699583452596214
	pesos_i(21517) := b"1111111111111111_1111111111111111_1101100111111010_0101001100010011"; -- -0.14852410102399144
	pesos_i(21518) := b"0000000000000000_0000000000000000_0001011010110101_1011010110010101"; -- 0.08871016404702127
	pesos_i(21519) := b"1111111111111111_1111111111111111_1101101011110011_1011110011000110"; -- -0.144718362420693
	pesos_i(21520) := b"1111111111111111_1111111111111111_1101111100001101_1000011101010011"; -- -0.12869981982315307
	pesos_i(21521) := b"0000000000000000_0000000000000000_0000111110011111_1100000000001101"; -- 0.06103134450971553
	pesos_i(21522) := b"0000000000000000_0000000000000000_0000000001000010_0100100000001001"; -- 0.0010113736177544588
	pesos_i(21523) := b"0000000000000000_0000000000000000_0001000001111110_0011111010111111"; -- 0.06442634726972815
	pesos_i(21524) := b"0000000000000000_0000000000000000_0000110001110000_1101000100110111"; -- 0.04859645455024563
	pesos_i(21525) := b"0000000000000000_0000000000000000_0010010000010001_0010001010100110"; -- 0.1408864646882864
	pesos_i(21526) := b"1111111111111111_1111111111111111_1110100111110110_1011010101101011"; -- -0.08607927442438348
	pesos_i(21527) := b"0000000000000000_0000000000000000_0001110011011010_0101101110001010"; -- 0.11270687221088754
	pesos_i(21528) := b"0000000000000000_0000000000000000_0010101011111111_0100111011110010"; -- 0.16795819682412125
	pesos_i(21529) := b"0000000000000000_0000000000000000_0000110101111000_1011111010100111"; -- 0.05262366849850293
	pesos_i(21530) := b"1111111111111111_1111111111111111_1110111010101111_0001110101100110"; -- -0.06764045954637558
	pesos_i(21531) := b"1111111111111111_1111111111111111_1111010111011011_0001000101001110"; -- -0.03962604376195009
	pesos_i(21532) := b"0000000000000000_0000000000000000_0000010111000001_0001000101111010"; -- 0.022477238081475108
	pesos_i(21533) := b"0000000000000000_0000000000000000_0001111110100111_0110001010110010"; -- 0.12364785036122806
	pesos_i(21534) := b"0000000000000000_0000000000000000_0000001011010111_0010111000111011"; -- 0.01109589509394404
	pesos_i(21535) := b"0000000000000000_0000000000000000_0000111000111110_0100001010001011"; -- 0.05563751110052927
	pesos_i(21536) := b"0000000000000000_0000000000000000_0000101001001100_0101011110101100"; -- 0.040227393701788836
	pesos_i(21537) := b"1111111111111111_1111111111111111_1111101101111100_0011100100111010"; -- -0.017635749212166558
	pesos_i(21538) := b"1111111111111111_1111111111111111_1101101001001010_1010001010100110"; -- -0.14729865490155974
	pesos_i(21539) := b"0000000000000000_0000000000000000_0000011111011101_0000110101011000"; -- 0.03071673773496408
	pesos_i(21540) := b"1111111111111111_1111111111111111_1101111001010001_0111111011011110"; -- -0.13156897612479013
	pesos_i(21541) := b"1111111111111111_1111111111111111_1111011100001111_0101000111101011"; -- -0.03492248556863707
	pesos_i(21542) := b"0000000000000000_0000000000000000_0001111010010100_1111100000000101"; -- 0.11946058388806491
	pesos_i(21543) := b"0000000000000000_0000000000000000_0010000101000111_0101010000100000"; -- 0.12999463836182631
	pesos_i(21544) := b"1111111111111111_1111111111111111_1110110000000010_0111011101011001"; -- -0.07808736876557851
	pesos_i(21545) := b"0000000000000000_0000000000000000_0000011110001101_0111101000000110"; -- 0.029502512526325336
	pesos_i(21546) := b"1111111111111111_1111111111111111_1101111110101111_0000110000001000"; -- -0.12623524475595232
	pesos_i(21547) := b"1111111111111111_1111111111111111_1110101110000000_0010111110000100"; -- -0.080075292732592
	pesos_i(21548) := b"0000000000000000_0000000000000000_0001010010100001_1011110110001101"; -- 0.08059296320043251
	pesos_i(21549) := b"1111111111111111_1111111111111111_1111010011100100_1010001001100010"; -- -0.04338631725367659
	pesos_i(21550) := b"1111111111111111_1111111111111111_1111101101000101_0101110110101001"; -- -0.01847281091021862
	pesos_i(21551) := b"0000000000000000_0000000000000000_0000101100100011_1110011001011000"; -- 0.04351653715065097
	pesos_i(21552) := b"0000000000000000_0000000000000000_0000011001110001_1101001000011001"; -- 0.025174266052955082
	pesos_i(21553) := b"1111111111111111_1111111111111111_1101111000111011_1001010010000011"; -- -0.13190337937576346
	pesos_i(21554) := b"0000000000000000_0000000000000000_0001000111100101_1010100011100001"; -- 0.06991057863888855
	pesos_i(21555) := b"1111111111111111_1111111111111111_1101101101000111_1000011101101101"; -- -0.14343980391790745
	pesos_i(21556) := b"1111111111111111_1111111111111111_1111101001001100_0000101100111111"; -- -0.022277161619298675
	pesos_i(21557) := b"0000000000000000_0000000000000000_0001010101011110_0011000000110100"; -- 0.08346844921531824
	pesos_i(21558) := b"0000000000000000_0000000000000000_0010100110011010_1000010010010000"; -- 0.16251400486054882
	pesos_i(21559) := b"1111111111111111_1111111111111111_1111100001110011_0110001000010001"; -- -0.02948939393713995
	pesos_i(21560) := b"0000000000000000_0000000000000000_0000011001011001_0100110100100101"; -- 0.024800130494871266
	pesos_i(21561) := b"0000000000000000_0000000000000000_0001101101101100_0001101011001001"; -- 0.10711829563145364
	pesos_i(21562) := b"0000000000000000_0000000000000000_0000000001101001_0000101101111000"; -- 0.0016028563356216055
	pesos_i(21563) := b"0000000000000000_0000000000000000_0000110101000010_1011010101100111"; -- 0.05179914250619449
	pesos_i(21564) := b"1111111111111111_1111111111111111_1101100000010000_0101000111101011"; -- -0.15600097675378216
	pesos_i(21565) := b"1111111111111111_1111111111111111_1110101101000001_1000110010100011"; -- -0.08103104609785705
	pesos_i(21566) := b"1111111111111111_1111111111111111_1111010011100101_0001011111110001"; -- -0.043379310171954594
	pesos_i(21567) := b"0000000000000000_0000000000000000_0010011010001000_1100000010001001"; -- 0.15052417122591055
	pesos_i(21568) := b"0000000000000000_0000000000000000_0010010011101100_1101011011110010"; -- 0.14423888592199702
	pesos_i(21569) := b"0000000000000000_0000000000000000_0010001100110000_1010101101000001"; -- 0.13746137931034214
	pesos_i(21570) := b"0000000000000000_0000000000000000_0000110011101110_0001101001111001"; -- 0.05050816965667492
	pesos_i(21571) := b"1111111111111111_1111111111111111_1111111000010101_1010000100011111"; -- -0.0074824617802855126
	pesos_i(21572) := b"1111111111111111_1111111111111111_1101110110010000_0111110000010111"; -- -0.13451408809164306
	pesos_i(21573) := b"1111111111111111_1111111111111111_1101101111000101_1111101000010111"; -- -0.1415103619497865
	pesos_i(21574) := b"0000000000000000_0000000000000000_0010001111101011_1001000001000011"; -- 0.1403131640702978
	pesos_i(21575) := b"1111111111111111_1111111111111111_1111011111111010_1010100001010010"; -- -0.03133152003941489
	pesos_i(21576) := b"0000000000000000_0000000000000000_0000110101101010_0110111100101101"; -- 0.05240530820572224
	pesos_i(21577) := b"1111111111111111_1111111111111111_1111011011100010_1101000000110101"; -- -0.03560160358569585
	pesos_i(21578) := b"0000000000000000_0000000000000000_0001110101000110_0000010100010111"; -- 0.11434966851502418
	pesos_i(21579) := b"0000000000000000_0000000000000000_0000010001001100_1111101000100011"; -- 0.016799577254554703
	pesos_i(21580) := b"1111111111111111_1111111111111111_1101110110001000_0001001000001110"; -- -0.13464247865753667
	pesos_i(21581) := b"0000000000000000_0000000000000000_0010100011100010_1000100110101010"; -- 0.159706691816947
	pesos_i(21582) := b"1111111111111111_1111111111111111_1110100011110011_1000001101100100"; -- -0.09003428271567211
	pesos_i(21583) := b"1111111111111111_1111111111111111_1111011110100100_0100110100110110"; -- -0.0326492063891662
	pesos_i(21584) := b"0000000000000000_0000000000000000_0001100001110001_0100101001110101"; -- 0.09547868117821828
	pesos_i(21585) := b"0000000000000000_0000000000000000_0000100101111011_1001001011000110"; -- 0.03704182938361135
	pesos_i(21586) := b"0000000000000000_0000000000000000_0000111100000001_0011100110110110"; -- 0.05861244857579562
	pesos_i(21587) := b"1111111111111111_1111111111111111_1111110001100010_1100110011001010"; -- -0.014117432372700916
	pesos_i(21588) := b"0000000000000000_0000000000000000_0010001010111111_0000110000000110"; -- 0.13572764525380077
	pesos_i(21589) := b"0000000000000000_0000000000000000_0010001011011101_0110010110011001"; -- 0.1361907480593685
	pesos_i(21590) := b"1111111111111111_1111111111111111_1110011001101111_1000110110100101"; -- -0.09986033179068436
	pesos_i(21591) := b"1111111111111111_1111111111111111_1110100100001100_1001111111111011"; -- -0.08965110892514153
	pesos_i(21592) := b"0000000000000000_0000000000000000_0000001101101111_0001101111001100"; -- 0.01341413235955814
	pesos_i(21593) := b"0000000000000000_0000000000000000_0000011011011100_1111100100100100"; -- 0.026809283644677374
	pesos_i(21594) := b"0000000000000000_0000000000000000_0010000011100101_0011110001111110"; -- 0.1284978682951899
	pesos_i(21595) := b"0000000000000000_0000000000000000_0001110001001110_0110110111011001"; -- 0.11057173292288339
	pesos_i(21596) := b"0000000000000000_0000000000000000_0001110100000110_1011101101010110"; -- 0.11338396877222573
	pesos_i(21597) := b"1111111111111111_1111111111111111_1111010101001010_0110010100001001"; -- -0.04183357751537401
	pesos_i(21598) := b"1111111111111111_1111111111111111_1111011000100000_1100110010001110"; -- -0.03856202636540441
	pesos_i(21599) := b"1111111111111111_1111111111111111_1110000000000000_0000000111100110"; -- -0.12499988694625024
	pesos_i(21600) := b"0000000000000000_0000000000000000_0001110011100111_0111001011101010"; -- 0.11290662970410943
	pesos_i(21601) := b"0000000000000000_0000000000000000_0000001100011101_0011110101011001"; -- 0.012164911468993978
	pesos_i(21602) := b"1111111111111111_1111111111111111_1110001111010100_0110011110110010"; -- -0.11004020601246478
	pesos_i(21603) := b"0000000000000000_0000000000000000_0001000011010100_1101001000010001"; -- 0.0657473841590628
	pesos_i(21604) := b"1111111111111111_1111111111111111_1110111110010110_1101101001000100"; -- -0.06410442203271491
	pesos_i(21605) := b"0000000000000000_0000000000000000_0010001000111011_0011000001101011"; -- 0.13371565444704464
	pesos_i(21606) := b"1111111111111111_1111111111111111_1110110111101000_0011110011001001"; -- -0.07067508774855356
	pesos_i(21607) := b"0000000000000000_0000000000000000_0001010110001100_0111010001000101"; -- 0.08417441061811763
	pesos_i(21608) := b"1111111111111111_1111111111111111_1110111011000001_1010110001111000"; -- -0.06735727388106029
	pesos_i(21609) := b"1111111111111111_1111111111111111_1111110100111000_1110001000110011"; -- -0.01085077537100382
	pesos_i(21610) := b"1111111111111111_1111111111111111_1101111010110010_1001110000100010"; -- -0.13008712929130944
	pesos_i(21611) := b"1111111111111111_1111111111111111_1111101000111110_0001010110110001"; -- -0.022490162275291804
	pesos_i(21612) := b"1111111111111111_1111111111111111_1111010111001101_1000111111011111"; -- -0.03983212296040748
	pesos_i(21613) := b"0000000000000000_0000000000000000_0000011000111000_0110110110100110"; -- 0.024298527669572113
	pesos_i(21614) := b"1111111111111111_1111111111111111_1111101010000100_0110000101101001"; -- -0.021417533691910653
	pesos_i(21615) := b"0000000000000000_0000000000000000_0000000000001101_1010111110111001"; -- 0.00020883817356270713
	pesos_i(21616) := b"0000000000000000_0000000000000000_0001001001110111_1001000100011100"; -- 0.07213694510811221
	pesos_i(21617) := b"1111111111111111_1111111111111111_1110101010100110_0010010010110100"; -- -0.08340235322795529
	pesos_i(21618) := b"1111111111111111_1111111111111111_1110110011101110_0000110001011001"; -- -0.0744926721755381
	pesos_i(21619) := b"1111111111111111_1111111111111111_1111011101010010_1001000100111111"; -- -0.03389637192206162
	pesos_i(21620) := b"1111111111111111_1111111111111111_1110011100011110_1001111011000111"; -- -0.09718902248233136
	pesos_i(21621) := b"1111111111111111_1111111111111111_1111010101100100_1111100011101001"; -- -0.04142803491891796
	pesos_i(21622) := b"1111111111111111_1111111111111111_1111010110000011_1010000010101101"; -- -0.040960271600405655
	pesos_i(21623) := b"1111111111111111_1111111111111111_1110111111101101_0011100011111100"; -- -0.06278652049086085
	pesos_i(21624) := b"1111111111111111_1111111111111111_1110010101111000_1101001010001011"; -- -0.10362514591919446
	pesos_i(21625) := b"0000000000000000_0000000000000000_0000010011010100_1011010111010011"; -- 0.0188707008699528
	pesos_i(21626) := b"1111111111111111_1111111111111111_1111100110011111_1000011110010001"; -- -0.024909522144524656
	pesos_i(21627) := b"1111111111111111_1111111111111111_1110101001010000_0000111100101010"; -- -0.08471589311396487
	pesos_i(21628) := b"1111111111111111_1111111111111111_1110000111001100_0001101000100101"; -- -0.11797939864621733
	pesos_i(21629) := b"1111111111111111_1111111111111111_1111010011010101_0101010000011100"; -- -0.04361986466268573
	pesos_i(21630) := b"1111111111111111_1111111111111111_1101100001101111_0001101000101111"; -- -0.1545547137428278
	pesos_i(21631) := b"0000000000000000_0000000000000000_0001001010111010_1111100101111011"; -- 0.07316550488345819
	pesos_i(21632) := b"1111111111111111_1111111111111111_1111101100100111_1010000000111111"; -- -0.018926605753271524
	pesos_i(21633) := b"0000000000000000_0000000000000000_0010000000011001_1101100111001011"; -- 0.12539445114535575
	pesos_i(21634) := b"0000000000000000_0000000000000000_0000000111000010_0001000001001111"; -- 0.0068674272624475365
	pesos_i(21635) := b"0000000000000000_0000000000000000_0001101111000000_1110100000000111"; -- 0.10841226737882788
	pesos_i(21636) := b"1111111111111111_1111111111111111_1111000110111110_0110101100000011"; -- -0.055688201645756906
	pesos_i(21637) := b"0000000000000000_0000000000000000_0000110011110010_0101000011001110"; -- 0.050572443345876475
	pesos_i(21638) := b"1111111111111111_1111111111111111_1111011000110100_0111111110000111"; -- -0.03826144182575688
	pesos_i(21639) := b"0000000000000000_0000000000000000_0010001111111101_0101011111111010"; -- 0.14058446747939154
	pesos_i(21640) := b"1111111111111111_1111111111111111_1110000011100101_1001111101100111"; -- -0.12149623618087389
	pesos_i(21641) := b"1111111111111111_1111111111111111_1111010010111101_0001001100001001"; -- -0.04398995430724383
	pesos_i(21642) := b"1111111111111111_1111111111111111_1110111111001010_1000001111011100"; -- -0.06331611519180554
	pesos_i(21643) := b"0000000000000000_0000000000000000_0001100001001100_1100110011100101"; -- 0.09492188061763263
	pesos_i(21644) := b"1111111111111111_1111111111111111_1101110001000001_0101001100100110"; -- -0.13962822264583893
	pesos_i(21645) := b"0000000000000000_0000000000000000_0010010010111100_1100011101001011"; -- 0.14350553112453632
	pesos_i(21646) := b"1111111111111111_1111111111111111_1110010000000000_0011010111000001"; -- -0.10937179596653174
	pesos_i(21647) := b"0000000000000000_0000000000000000_0000110001111000_0001001011101010"; -- 0.048707181961700236
	pesos_i(21648) := b"0000000000000000_0000000000000000_0000010011101001_0101101000111011"; -- 0.01918567611401049
	pesos_i(21649) := b"0000000000000000_0000000000000000_0000110001001011_1000100110110100"; -- 0.048027617000378074
	pesos_i(21650) := b"1111111111111111_1111111111111111_1111010111100111_0110101001101010"; -- -0.039437627026523245
	pesos_i(21651) := b"1111111111111111_1111111111111111_1110010100110001_1100101101111001"; -- -0.1047089413901455
	pesos_i(21652) := b"1111111111111111_1111111111111111_1111001101001101_0111110000010010"; -- -0.049598928067659205
	pesos_i(21653) := b"1111111111111111_1111111111111111_1101110110010000_1100010111101110"; -- -0.13450968674625188
	pesos_i(21654) := b"1111111111111111_1111111111111111_1110111111110010_0111000000111111"; -- -0.06270693275107453
	pesos_i(21655) := b"1111111111111111_1111111111111111_1110011000010011_1111010001101101"; -- -0.10125801403078037
	pesos_i(21656) := b"1111111111111111_1111111111111111_1111010001111000_0010010101111100"; -- -0.04504171117999079
	pesos_i(21657) := b"1111111111111111_1111111111111111_1111001111110011_1000011101010111"; -- -0.04706529735130878
	pesos_i(21658) := b"0000000000000000_0000000000000000_0010001011111010_0010001010110111"; -- 0.13662926633352143
	pesos_i(21659) := b"1111111111111111_1111111111111111_1111101101000110_0001111111110010"; -- -0.018461230596927516
	pesos_i(21660) := b"1111111111111111_1111111111111111_1111000100111010_0001101001001011"; -- -0.05770717303580783
	pesos_i(21661) := b"0000000000000000_0000000000000000_0000011100011000_0000110111100001"; -- 0.027710788197199448
	pesos_i(21662) := b"0000000000000000_0000000000000000_0001001010011100_1001010011100000"; -- 0.07270174482560927
	pesos_i(21663) := b"0000000000000000_0000000000000000_0001101100110110_0011110000101100"; -- 0.10629631114614231
	pesos_i(21664) := b"0000000000000000_0000000000000000_0000110100111101_0111000011001100"; -- 0.051718759301345715
	pesos_i(21665) := b"0000000000000000_0000000000000000_0000101000011110_1111101101111101"; -- 0.03953525355332191
	pesos_i(21666) := b"0000000000000000_0000000000000000_0000111010110001_1100010101111011"; -- 0.05740007644024883
	pesos_i(21667) := b"0000000000000000_0000000000000000_0000011111011001_0001101111001110"; -- 0.03065656444424602
	pesos_i(21668) := b"0000000000000000_0000000000000000_0000111000110001_1110010100111010"; -- 0.05544884358699426
	pesos_i(21669) := b"0000000000000000_0000000000000000_0001101100110001_0110000110001101"; -- 0.10622224521855692
	pesos_i(21670) := b"1111111111111111_1111111111111111_1110111101110000_0111010100110110"; -- -0.06469027934792841
	pesos_i(21671) := b"1111111111111111_1111111111111111_1111101100110111_0100110010110011"; -- -0.018687444972779223
	pesos_i(21672) := b"1111111111111111_1111111111111111_1110110111000001_1001001101111000"; -- -0.0712650138648803
	pesos_i(21673) := b"1111111111111111_1111111111111111_1111010010000111_1111100001011111"; -- -0.044800259299560004
	pesos_i(21674) := b"0000000000000000_0000000000000000_0000110001111111_0010111110001000"; -- 0.04881569918997901
	pesos_i(21675) := b"0000000000000000_0000000000000000_0001011101001000_1110111111111010"; -- 0.09095668650557243
	pesos_i(21676) := b"1111111111111111_1111111111111111_1111111010111011_1100010101000010"; -- -0.004947349007081133
	pesos_i(21677) := b"0000000000000000_0000000000000000_0000001001010010_1100010100101011"; -- 0.00907547276894636
	pesos_i(21678) := b"1111111111111111_1111111111111111_1101100100110001_1001100110110100"; -- -0.1515869078068664
	pesos_i(21679) := b"0000000000000000_0000000000000000_0000111011011001_1001110010011000"; -- 0.05800799103408969
	pesos_i(21680) := b"1111111111111111_1111111111111111_1111010001111100_1111110000001100"; -- -0.044967886905913725
	pesos_i(21681) := b"0000000000000000_0000000000000000_0000110110011001_1100110100100011"; -- 0.053128071766963214
	pesos_i(21682) := b"1111111111111111_1111111111111111_1111000000100100_1110110100010001"; -- -0.06193655334304897
	pesos_i(21683) := b"1111111111111111_1111111111111111_1111001110001111_0100110110011001"; -- -0.04859461798001421
	pesos_i(21684) := b"1111111111111111_1111111111111111_1110010111011001_0111101101000010"; -- -0.10215024607637652
	pesos_i(21685) := b"0000000000000000_0000000000000000_0001110110111111_0101000101000010"; -- 0.11620052199642875
	pesos_i(21686) := b"1111111111111111_1111111111111111_1101110010000110_0111111001010110"; -- -0.13857279199494385
	pesos_i(21687) := b"0000000000000000_0000000000000000_0000010100010101_0011110111010100"; -- 0.019855369846569746
	pesos_i(21688) := b"0000000000000000_0000000000000000_0000011011011001_0010101011011110"; -- 0.026751212371588114
	pesos_i(21689) := b"0000000000000000_0000000000000000_0000111100001111_0001010100111011"; -- 0.05882389736859453
	pesos_i(21690) := b"0000000000000000_0000000000000000_0001000101011010_0000001111110010"; -- 0.0677797762037857
	pesos_i(21691) := b"0000000000000000_0000000000000000_0000010011100111_0100011001100111"; -- 0.019153976475491316
	pesos_i(21692) := b"0000000000000000_0000000000000000_0001111111101101_0111101111101100"; -- 0.12471746943315296
	pesos_i(21693) := b"0000000000000000_0000000000000000_0001001001000010_0111001101011100"; -- 0.0713264559970532
	pesos_i(21694) := b"0000000000000000_0000000000000000_0000111011101000_1111000100100111"; -- 0.05824191294518094
	pesos_i(21695) := b"0000000000000000_0000000000000000_0000010100001010_1001001101100000"; -- 0.019692622147271695
	pesos_i(21696) := b"0000000000000000_0000000000000000_0001110010000110_1011101100011001"; -- 0.11143082972832591
	pesos_i(21697) := b"1111111111111111_1111111111111111_1101101110101110_0010011101000111"; -- -0.14187387952116895
	pesos_i(21698) := b"1111111111111111_1111111111111111_1110001101000100_0111100101010100"; -- -0.11223642057432759
	pesos_i(21699) := b"1111111111111111_1111111111111111_1110110111110011_1110000101100101"; -- -0.07049742975476465
	pesos_i(21700) := b"0000000000000000_0000000000000000_0010011001010010_1001111001000011"; -- 0.14969815384040952
	pesos_i(21701) := b"0000000000000000_0000000000000000_0000111101110011_1000110000011110"; -- 0.06035686232488588
	pesos_i(21702) := b"0000000000000000_0000000000000000_0001100000101010_1011100001101101"; -- 0.0944018618261687
	pesos_i(21703) := b"1111111111111111_1111111111111111_1101110110000111_0111010111010111"; -- -0.13465178973128086
	pesos_i(21704) := b"0000000000000000_0000000000000000_0001000101011010_1100011000001110"; -- 0.06779134609163555
	pesos_i(21705) := b"1111111111111111_1111111111111111_1110011111000011_0000101110100111"; -- -0.09468009168109554
	pesos_i(21706) := b"0000000000000000_0000000000000000_0000101101110100_0010011000110001"; -- 0.044741045919230386
	pesos_i(21707) := b"1111111111111111_1111111111111111_1110111110010111_0011000001111000"; -- -0.06409928377476257
	pesos_i(21708) := b"1111111111111111_1111111111111111_1110011110110011_0001111111101010"; -- -0.0949230245191905
	pesos_i(21709) := b"0000000000000000_0000000000000000_0001101110101100_1101010101110001"; -- 0.10810598382027109
	pesos_i(21710) := b"0000000000000000_0000000000000000_0000101111100010_0010100010110001"; -- 0.046419661810654975
	pesos_i(21711) := b"1111111111111111_1111111111111111_1111110001101001_1111111110001110"; -- -0.014007595005214542
	pesos_i(21712) := b"0000000000000000_0000000000000000_0010000011100111_0001110101101000"; -- 0.12852653294934188
	pesos_i(21713) := b"0000000000000000_0000000000000000_0001101010000001_1101101111000001"; -- 0.10354398204636091
	pesos_i(21714) := b"0000000000000000_0000000000000000_0001110001010111_1111101000100100"; -- 0.11071742421532028
	pesos_i(21715) := b"1111111111111111_1111111111111111_1111110101011010_1111110000111110"; -- -0.01033042415566458
	pesos_i(21716) := b"0000000000000000_0000000000000000_0001001010001000_0001101011111000"; -- 0.07238930272626037
	pesos_i(21717) := b"1111111111111111_1111111111111111_1110011101101010_0001001011100110"; -- -0.09603769200279698
	pesos_i(21718) := b"1111111111111111_1111111111111111_1110001001100111_0110001010101101"; -- -0.11560996312122306
	pesos_i(21719) := b"0000000000000000_0000000000000000_0001011010010111_1110101100000100"; -- 0.0882555851781781
	pesos_i(21720) := b"1111111111111111_1111111111111111_1110110100100000_1001110011100101"; -- -0.07372111710227
	pesos_i(21721) := b"0000000000000000_0000000000000000_0001111111110010_1000111010000000"; -- 0.12479487066888853
	pesos_i(21722) := b"1111111111111111_1111111111111111_1110110111101011_0101001101101111"; -- -0.07062796146935799
	pesos_i(21723) := b"1111111111111111_1111111111111111_1110101001111101_1010101100011100"; -- -0.08401995246058162
	pesos_i(21724) := b"0000000000000000_0000000000000000_0000011011111111_1010001101110101"; -- 0.027338234099279147
	pesos_i(21725) := b"0000000000000000_0000000000000000_0010001000010111_1000100001010010"; -- 0.1331715775434484
	pesos_i(21726) := b"1111111111111111_1111111111111111_1110011011100101_1011000101010000"; -- -0.09805766866453526
	pesos_i(21727) := b"0000000000000000_0000000000000000_0001110011101110_1000001100100001"; -- 0.11301440775414957
	pesos_i(21728) := b"1111111111111111_1111111111111111_1111101000101000_0101110110110010"; -- -0.022821563824462845
	pesos_i(21729) := b"1111111111111111_1111111111111111_1111100100100001_1010001000100010"; -- -0.026830545977369908
	pesos_i(21730) := b"0000000000000000_0000000000000000_0001100010111110_0100111001011111"; -- 0.09665384108935235
	pesos_i(21731) := b"1111111111111111_1111111111111111_1101101011100101_1011000000010000"; -- -0.14493274309211251
	pesos_i(21732) := b"1111111111111111_1111111111111111_1110100000001000_1010001011000110"; -- -0.09361822758012349
	pesos_i(21733) := b"0000000000000000_0000000000000000_0000101001010100_0101111111100111"; -- 0.040349954408000405
	pesos_i(21734) := b"1111111111111111_1111111111111111_1111001101111111_0011110100100110"; -- -0.048839739152410674
	pesos_i(21735) := b"1111111111111111_1111111111111111_1111000010010001_1100101000011110"; -- -0.0602754284829568
	pesos_i(21736) := b"0000000000000000_0000000000000000_0000101010001110_1001111111100001"; -- 0.04123877762859204
	pesos_i(21737) := b"0000000000000000_0000000000000000_0001100101001001_1100110010101111"; -- 0.09878234175852395
	pesos_i(21738) := b"1111111111111111_1111111111111111_1101110111010110_0001010011110111"; -- -0.13345211945775434
	pesos_i(21739) := b"1111111111111111_1111111111111111_1110100010000010_1110010000001111"; -- -0.09175276417344269
	pesos_i(21740) := b"1111111111111111_1111111111111111_1110111101011011_1011110100111011"; -- -0.06500642109487731
	pesos_i(21741) := b"1111111111111111_1111111111111111_1110110100101100_0001000011011100"; -- -0.073546358302887
	pesos_i(21742) := b"1111111111111111_1111111111111111_1110100100000001_1011101110111010"; -- -0.08981730180552104
	pesos_i(21743) := b"1111111111111111_1111111111111111_1111001001101011_1111001101000101"; -- -0.05304030962331417
	pesos_i(21744) := b"1111111111111111_1111111111111111_1101110000110110_0011010101100000"; -- -0.1397978440076021
	pesos_i(21745) := b"0000000000000000_0000000000000000_0000000011011001_1101111001010011"; -- 0.003324408800200435
	pesos_i(21746) := b"0000000000000000_0000000000000000_0010010010111101_1101000100001110"; -- 0.1435213718441431
	pesos_i(21747) := b"1111111111111111_1111111111111111_1111110000100100_1101110001111000"; -- -0.015062542659718306
	pesos_i(21748) := b"1111111111111111_1111111111111111_1110011000110010_0101100010011010"; -- -0.10079427954726837
	pesos_i(21749) := b"1111111111111111_1111111111111111_1110100010101101_1100011111011101"; -- -0.09109831659732265
	pesos_i(21750) := b"0000000000000000_0000000000000000_0000001001011111_0100000100110100"; -- 0.009265971473763172
	pesos_i(21751) := b"0000000000000000_0000000000000000_0001101111010010_0101000011010111"; -- 0.1086779140255216
	pesos_i(21752) := b"0000000000000000_0000000000000000_0010000110011101_1011001100111101"; -- 0.13131256323544124
	pesos_i(21753) := b"1111111111111111_1111111111111111_1101110010110111_0101011001100110"; -- -0.13782749180205692
	pesos_i(21754) := b"1111111111111111_1111111111111111_1111001000001000_0110001011111111"; -- -0.05455952900254237
	pesos_i(21755) := b"0000000000000000_0000000000000000_0010010111011001_1100111000000111"; -- 0.14785468733867468
	pesos_i(21756) := b"1111111111111111_1111111111111111_1111001011000000_0100100110100110"; -- -0.05175342271391995
	pesos_i(21757) := b"1111111111111111_1111111111111111_1111111000001110_1111100001101110"; -- -0.007584069462091815
	pesos_i(21758) := b"1111111111111111_1111111111111111_1111010110110110_1111010111001001"; -- -0.040177000461909154
	pesos_i(21759) := b"1111111111111111_1111111111111111_1101111110111010_0101110001110111"; -- -0.12606260381811668
	pesos_i(21760) := b"1111111111111111_1111111111111111_1101101001011001_0110001111110110"; -- -0.14707350954183115
	pesos_i(21761) := b"0000000000000000_0000000000000000_0000101011000101_1001010011100110"; -- 0.04207735646509536
	pesos_i(21762) := b"0000000000000000_0000000000000000_0001111010001101_0100100011011110"; -- 0.1193433324872822
	pesos_i(21763) := b"0000000000000000_0000000000000000_0001000100111100_0000100101101110"; -- 0.06732233928595924
	pesos_i(21764) := b"1111111111111111_1111111111111111_1110000000110111_1111111100001010"; -- -0.12414556507122555
	pesos_i(21765) := b"0000000000000000_0000000000000000_0001101101010000_1101000111101001"; -- 0.10670196470011248
	pesos_i(21766) := b"1111111111111111_1111111111111111_1111010001100101_1111001000100110"; -- -0.04531942919135606
	pesos_i(21767) := b"0000000000000000_0000000000000000_0001000001000111_1011111101010110"; -- 0.06359477852286821
	pesos_i(21768) := b"1111111111111111_1111111111111111_1111000010110000_1000110010011110"; -- -0.05980607162286396
	pesos_i(21769) := b"0000000000000000_0000000000000000_0001101001010010_0110111111000000"; -- 0.10282038150357109
	pesos_i(21770) := b"0000000000000000_0000000000000000_0000101001000011_1110101001111100"; -- 0.040098815341100574
	pesos_i(21771) := b"0000000000000000_0000000000000000_0001010100101001_1101110011010100"; -- 0.08267002281040996
	pesos_i(21772) := b"0000000000000000_0000000000000000_0001101000101001_1101000010100100"; -- 0.10220054624196434
	pesos_i(21773) := b"0000000000000000_0000000000000000_0010011011010011_0100111100000000"; -- 0.1516618132206455
	pesos_i(21774) := b"1111111111111111_1111111111111111_1101111110111111_1111000001010011"; -- -0.12597749696374413
	pesos_i(21775) := b"0000000000000000_0000000000000000_0000000101010100_0100110010010000"; -- 0.005192551872253608
	pesos_i(21776) := b"1111111111111111_1111111111111111_1111001000111001_0000110011101100"; -- -0.05381697890231081
	pesos_i(21777) := b"0000000000000000_0000000000000000_0001100001110100_1100010000010100"; -- 0.09553170661644786
	pesos_i(21778) := b"1111111111111111_1111111111111111_1111110011111100_0001100100011101"; -- -0.011778288271689192
	pesos_i(21779) := b"1111111111111111_1111111111111111_1110101111111100_0110100001001000"; -- -0.07817981961350343
	pesos_i(21780) := b"1111111111111111_1111111111111111_1101011110111011_1100001101011110"; -- -0.15729121166136742
	pesos_i(21781) := b"0000000000000000_0000000000000000_0001001010100100_0111111100111011"; -- 0.07282252489760657
	pesos_i(21782) := b"0000000000000000_0000000000000000_0000010000100110_1111111111101110"; -- 0.016220088656750713
	pesos_i(21783) := b"1111111111111111_1111111111111111_1110010000100010_0000001101110001"; -- -0.10885599595062817
	pesos_i(21784) := b"1111111111111111_1111111111111111_1111111110010101_0000011000111101"; -- -0.001632318602153231
	pesos_i(21785) := b"0000000000000000_0000000000000000_0010011111010000_0101001110010110"; -- 0.15552256028383357
	pesos_i(21786) := b"0000000000000000_0000000000000000_0000101110011000_0010010000110110"; -- 0.04529024427963185
	pesos_i(21787) := b"1111111111111111_1111111111111111_1110001000000001_0101111000011110"; -- -0.11716663141089033
	pesos_i(21788) := b"1111111111111111_1111111111111111_1111011000100100_0101000000111111"; -- -0.03850840065738775
	pesos_i(21789) := b"0000000000000000_0000000000000000_0001010010010100_1101000110011011"; -- 0.08039579429502348
	pesos_i(21790) := b"0000000000000000_0000000000000000_0010000010111011_1001011000111011"; -- 0.12786234809435504
	pesos_i(21791) := b"1111111111111111_1111111111111111_1111100001011111_0110000000100001"; -- -0.029794685379641264
	pesos_i(21792) := b"0000000000000000_0000000000000000_0010001100010010_1110011100010000"; -- 0.13700718070251444
	pesos_i(21793) := b"1111111111111111_1111111111111111_1110010101101010_1000011000111101"; -- -0.10384331703811828
	pesos_i(21794) := b"1111111111111111_1111111111111111_1110111001110111_1100100110001000"; -- -0.06848469189220349
	pesos_i(21795) := b"1111111111111111_1111111111111111_1110101011111100_0110011111000011"; -- -0.08208610047807925
	pesos_i(21796) := b"0000000000000000_0000000000000000_0000100100101100_1001011000110101"; -- 0.03583658985710053
	pesos_i(21797) := b"0000000000000000_0000000000000000_0010010111010011_1010010001100010"; -- 0.14776065248210504
	pesos_i(21798) := b"1111111111111111_1111111111111111_1101100000000001_0011100001110110"; -- -0.15623137583434749
	pesos_i(21799) := b"1111111111111111_1111111111111111_1111111000101000_1001000010011001"; -- -0.007193529782269775
	pesos_i(21800) := b"1111111111111111_1111111111111111_1111011101010110_1011100110100001"; -- -0.0338329299012918
	pesos_i(21801) := b"1111111111111111_1111111111111111_1111011000010000_0000001110111101"; -- -0.03881813657601698
	pesos_i(21802) := b"0000000000000000_0000000000000000_0010100100000101_1001101010110000"; -- 0.16024176395419332
	pesos_i(21803) := b"1111111111111111_1111111111111111_1110011011110110_1110111110011000"; -- -0.09779455692387379
	pesos_i(21804) := b"0000000000000000_0000000000000000_0001000011001000_1111110000111001"; -- 0.06556679145735084
	pesos_i(21805) := b"1111111111111111_1111111111111111_1101010111000001_1011001010001001"; -- -0.16501316208711425
	pesos_i(21806) := b"0000000000000000_0000000000000000_0001010001000111_0100100001111110"; -- 0.07921269493249875
	pesos_i(21807) := b"1111111111111111_1111111111111111_1111100000011010_1001101110111000"; -- -0.030843989873096347
	pesos_i(21808) := b"0000000000000000_0000000000000000_0010011001111001_1010001001001011"; -- 0.1502934869479581
	pesos_i(21809) := b"1111111111111111_1111111111111111_1110100011010111_0100100010011111"; -- -0.09046503184093324
	pesos_i(21810) := b"1111111111111111_1111111111111111_1111000011010101_0101101001100011"; -- -0.05924449039801077
	pesos_i(21811) := b"1111111111111111_1111111111111111_1110011101000101_1101101110010110"; -- -0.09659030530653255
	pesos_i(21812) := b"1111111111111111_1111111111111111_1111011010010011_0111010111011111"; -- -0.036812432350269854
	pesos_i(21813) := b"1111111111111111_1111111111111111_1111000001011110_0000011100011110"; -- -0.06106524969730073
	pesos_i(21814) := b"0000000000000000_0000000000000000_0000101010101100_1111011100001011"; -- 0.04170173668567443
	pesos_i(21815) := b"1111111111111111_1111111111111111_1110100001101111_0001001101111001"; -- -0.09205511366744827
	pesos_i(21816) := b"0000000000000000_0000000000000000_0001011110010110_0110010001000000"; -- 0.09213854369469923
	pesos_i(21817) := b"1111111111111111_1111111111111111_1111100000100100_1010101000010000"; -- -0.030690547122461456
	pesos_i(21818) := b"0000000000000000_0000000000000000_0000111011000011_0010101000100101"; -- 0.0576654758141261
	pesos_i(21819) := b"0000000000000000_0000000000000000_0000101110110000_1000001100011010"; -- 0.045662111054697446
	pesos_i(21820) := b"0000000000000000_0000000000000000_0010100010100101_1110001000010001"; -- 0.15878117486815804
	pesos_i(21821) := b"0000000000000000_0000000000000000_0000100101010011_1101101110110101"; -- 0.03643582498923201
	pesos_i(21822) := b"1111111111111111_1111111111111111_1111101111101010_0010110100010000"; -- -0.015958007362685624
	pesos_i(21823) := b"0000000000000000_0000000000000000_0001110101100011_0000001011101111"; -- 0.1147920449060681
	pesos_i(21824) := b"1111111111111111_1111111111111111_1110001110000100_1010010110010101"; -- -0.11125722030280243
	pesos_i(21825) := b"0000000000000000_0000000000000000_0010001001001110_0001111110011101"; -- 0.1340045697489882
	pesos_i(21826) := b"1111111111111111_1111111111111111_1111010001100011_0111110010111111"; -- -0.04535694434926833
	pesos_i(21827) := b"0000000000000000_0000000000000000_0001000100000111_1010110110111000"; -- 0.06652341603469179
	pesos_i(21828) := b"0000000000000000_0000000000000000_0001000111101111_0011001000110010"; -- 0.0700560924591699
	pesos_i(21829) := b"1111111111111111_1111111111111111_1110110010101111_1011110101100100"; -- -0.07544342342223079
	pesos_i(21830) := b"0000000000000000_0000000000000000_0000110100010010_0101010011100100"; -- 0.05106096817452614
	pesos_i(21831) := b"1111111111111111_1111111111111111_1111111100000011_1000101001011010"; -- -0.0038522271821939927
	pesos_i(21832) := b"1111111111111111_1111111111111111_1110101011000100_1111000110111000"; -- -0.08293236985318984
	pesos_i(21833) := b"0000000000000000_0000000000000000_0010100000011111_1100101111010111"; -- 0.15673517219517108
	pesos_i(21834) := b"1111111111111111_1111111111111111_1110011101010100_1101101010000000"; -- -0.09636148802448877
	pesos_i(21835) := b"1111111111111111_1111111111111111_1111110110001101_1100001010100111"; -- -0.0095556586181217
	pesos_i(21836) := b"0000000000000000_0000000000000000_0010000111000001_1001010100110100"; -- 0.1318600894928474
	pesos_i(21837) := b"0000000000000000_0000000000000000_0010000000011011_1101000100100111"; -- 0.12542445375428105
	pesos_i(21838) := b"0000000000000000_0000000000000000_0010010100111001_1111111110010000"; -- 0.14541623374940915
	pesos_i(21839) := b"0000000000000000_0000000000000000_0000101001000001_1110010101001001"; -- 0.04006798773095087
	pesos_i(21840) := b"0000000000000000_0000000000000000_0010100100111000_0001000011010000"; -- 0.16101174430938123
	pesos_i(21841) := b"0000000000000000_0000000000000000_0000101100111010_0110110000000001"; -- 0.043860197195660776
	pesos_i(21842) := b"0000000000000000_0000000000000000_0000000111100011_1100100010000100"; -- 0.007381946766821455
	pesos_i(21843) := b"1111111111111111_1111111111111111_1111000001000011_0010111000100100"; -- -0.06147491103447409
	pesos_i(21844) := b"0000000000000000_0000000000000000_0000000001001101_0100001000010111"; -- 0.00117886602411113
	pesos_i(21845) := b"0000000000000000_0000000000000000_0000000001100011_1010110001000010"; -- 0.0015208874510146562
	pesos_i(21846) := b"0000000000000000_0000000000000000_0000011111110010_1111111110001010"; -- 0.031051608359081027
	pesos_i(21847) := b"1111111111111111_1111111111111111_1111000111100100_0110000001110110"; -- -0.05510899657777336
	pesos_i(21848) := b"0000000000000000_0000000000000000_0001000011001011_1000001110100110"; -- 0.06560538108864639
	pesos_i(21849) := b"1111111111111111_1111111111111111_1111111000101110_1111100000111000"; -- -0.007095800728689976
	pesos_i(21850) := b"1111111111111111_1111111111111111_1101110111101110_1110101101011011"; -- -0.13307312986782185
	pesos_i(21851) := b"0000000000000000_0000000000000000_0000010100010010_0011111110100010"; -- 0.019809700950266695
	pesos_i(21852) := b"1111111111111111_1111111111111111_1101111111010101_1110100100001111"; -- -0.1256422365821377
	pesos_i(21853) := b"1111111111111111_1111111111111111_1111011010100010_1101100010000000"; -- -0.03657767167040652
	pesos_i(21854) := b"1111111111111111_1111111111111111_1110101001001001_1101010110101001"; -- -0.08481087331749058
	pesos_i(21855) := b"1111111111111111_1111111111111111_1111100001110111_1011111011100011"; -- -0.02942282637517992
	pesos_i(21856) := b"0000000000000000_0000000000000000_0000100001011001_1110101110011001"; -- 0.03262207502465554
	pesos_i(21857) := b"1111111111111111_1111111111111111_1111010000111110_0001000000001110"; -- -0.045927998251501755
	pesos_i(21858) := b"0000000000000000_0000000000000000_0001000000011010_0110101101001101"; -- 0.06290312416352356
	pesos_i(21859) := b"0000000000000000_0000000000000000_0001000001111110_0000010010001101"; -- 0.0644228787832892
	pesos_i(21860) := b"1111111111111111_1111111111111111_1111011011001001_1010100110011000"; -- -0.03598537483100614
	pesos_i(21861) := b"1111111111111111_1111111111111111_1101101010111110_0011100010010000"; -- -0.14553495866940894
	pesos_i(21862) := b"0000000000000000_0000000000000000_0010100010111011_1001010010011000"; -- 0.15911225049488942
	pesos_i(21863) := b"0000000000000000_0000000000000000_0000111001001001_0101010111100111"; -- 0.05580651175503362
	pesos_i(21864) := b"1111111111111111_1111111111111111_1110100100101000_0101001000010110"; -- -0.0892285057851608
	pesos_i(21865) := b"0000000000000000_0000000000000000_0010100000000111_1000101110011010"; -- 0.15636513235512586
	pesos_i(21866) := b"0000000000000000_0000000000000000_0001000001100111_1010000110000011"; -- 0.06408128212094491
	pesos_i(21867) := b"1111111111111111_1111111111111111_1111110011100000_1010001000101101"; -- -0.012197364826696082
	pesos_i(21868) := b"1111111111111111_1111111111111111_1111000010010011_0001000101101011"; -- -0.06025591985042225
	pesos_i(21869) := b"0000000000000000_0000000000000000_0000110100011010_0000111010011000"; -- 0.051178848370325936
	pesos_i(21870) := b"0000000000000000_0000000000000000_0001110000111100_1010001001001111"; -- 0.11030020172650437
	pesos_i(21871) := b"0000000000000000_0000000000000000_0001001100011100_0001101111001010"; -- 0.07464765233459668
	pesos_i(21872) := b"1111111111111111_1111111111111111_1111000011100010_1101111110010011"; -- -0.05903818763522376
	pesos_i(21873) := b"0000000000000000_0000000000000000_0001010011110101_0101001111100100"; -- 0.0818684037003995
	pesos_i(21874) := b"1111111111111111_1111111111111111_1111110001110011_1000101110110010"; -- -0.013861912731440086
	pesos_i(21875) := b"1111111111111111_1111111111111111_1111110100101001_1101000111011100"; -- -0.011080631170533685
	pesos_i(21876) := b"1111111111111111_1111111111111111_1111000111010101_0100010000100101"; -- -0.055339566091648425
	pesos_i(21877) := b"1111111111111111_1111111111111111_1111001110000110_0110111100111001"; -- -0.04872994297586476
	pesos_i(21878) := b"0000000000000000_0000000000000000_0001101110101010_0100000111110111"; -- 0.10806667594342506
	pesos_i(21879) := b"1111111111111111_1111111111111111_1110010010110000_0111000010000111"; -- -0.10668274599737462
	pesos_i(21880) := b"1111111111111111_1111111111111111_1111111101111101_0110000001110001"; -- -0.0019931529277203474
	pesos_i(21881) := b"1111111111111111_1111111111111111_1111011100110011_0000011110100111"; -- -0.03437759562207403
	pesos_i(21882) := b"1111111111111111_1111111111111111_1110011101110001_1011100100010011"; -- -0.09592097550160399
	pesos_i(21883) := b"0000000000000000_0000000000000000_0000001001101101_0001101010000001"; -- 0.009477287674370193
	pesos_i(21884) := b"0000000000000000_0000000000000000_0001000110111001_0001110111111010"; -- 0.06923091276712982
	pesos_i(21885) := b"1111111111111111_1111111111111111_1110101010001011_0111011010110010"; -- -0.08380945346872348
	pesos_i(21886) := b"1111111111111111_1111111111111111_1110010110110011_0000000011011100"; -- -0.10273737553545288
	pesos_i(21887) := b"0000000000000000_0000000000000000_0001110101010101_0111000100110011"; -- 0.11458499417163022
	pesos_i(21888) := b"1111111111111111_1111111111111111_1101110000101010_0111100110110011"; -- -0.139976876964293
	pesos_i(21889) := b"0000000000000000_0000000000000000_0001000010011110_1011110100100001"; -- 0.06492216174550362
	pesos_i(21890) := b"0000000000000000_0000000000000000_0001000101100001_1001100000101101"; -- 0.06789542303569333
	pesos_i(21891) := b"0000000000000000_0000000000000000_0001110111111011_1010111001100001"; -- 0.11712159981107845
	pesos_i(21892) := b"1111111111111111_1111111111111111_1111100000011010_0110100101001100"; -- -0.03084699533752545
	pesos_i(21893) := b"1111111111111111_1111111111111111_1111110000011011_0001100100011011"; -- -0.015211516214346769
	pesos_i(21894) := b"0000000000000000_0000000000000000_0001111010000100_0011011111110101"; -- 0.11920499536135469
	pesos_i(21895) := b"0000000000000000_0000000000000000_0000101110011100_0010001001000011"; -- 0.04535116317696912
	pesos_i(21896) := b"1111111111111111_1111111111111111_1101110000010000_0101010101010011"; -- -0.14037577362144582
	pesos_i(21897) := b"1111111111111111_1111111111111111_1111100001010000_0010001011100011"; -- -0.030027217465260506
	pesos_i(21898) := b"1111111111111111_1111111111111111_1111000010110001_0111101010011010"; -- -0.059791886763220684
	pesos_i(21899) := b"0000000000000000_0000000000000000_0000110011000100_0100000000110011"; -- 0.04986954924250372
	pesos_i(21900) := b"1111111111111111_1111111111111111_1110101110111101_1000100110001000"; -- -0.07913914132248825
	pesos_i(21901) := b"1111111111111111_1111111111111111_1110001011011110_1100101000101000"; -- -0.11378799934108551
	pesos_i(21902) := b"0000000000000000_0000000000000000_0010011000100110_0000011100101111"; -- 0.14901776220885699
	pesos_i(21903) := b"1111111111111111_1111111111111111_1110101010011101_0111101111010111"; -- -0.08353448866133828
	pesos_i(21904) := b"1111111111111111_1111111111111111_1110111101011100_1000001010001101"; -- -0.06499466008551406
	pesos_i(21905) := b"1111111111111111_1111111111111111_1110011001111101_1001110101110011"; -- -0.09964576665763643
	pesos_i(21906) := b"0000000000000000_0000000000000000_0001000110000010_1000110110010011"; -- 0.06839833116149376
	pesos_i(21907) := b"0000000000000000_0000000000000000_0010000100100011_1001100101111101"; -- 0.12944945622021764
	pesos_i(21908) := b"0000000000000000_0000000000000000_0010001101001100_0100010011000100"; -- 0.13788251666300938
	pesos_i(21909) := b"0000000000000000_0000000000000000_0000110100101100_0001111001000111"; -- 0.051454441314546344
	pesos_i(21910) := b"1111111111111111_1111111111111111_1111000001101101_0001001011010010"; -- -0.06083567029956425
	pesos_i(21911) := b"0000000000000000_0000000000000000_0001111111000000_1110100010110110"; -- 0.1240373081656043
	pesos_i(21912) := b"0000000000000000_0000000000000000_0001011100001110_0000000010010100"; -- 0.09005740760345783
	pesos_i(21913) := b"1111111111111111_1111111111111111_1110011010111000_0110111011101110"; -- -0.09874827095834615
	pesos_i(21914) := b"0000000000000000_0000000000000000_0001100111111110_0100110010101011"; -- 0.10153655222700832
	pesos_i(21915) := b"1111111111111111_1111111111111111_1101100110100100_1001001000010110"; -- -0.14983260115638214
	pesos_i(21916) := b"1111111111111111_1111111111111111_1110101010001010_0010111110000000"; -- -0.08382895599563664
	pesos_i(21917) := b"1111111111111111_1111111111111111_1101101011110111_1000111101000010"; -- -0.14466004036947055
	pesos_i(21918) := b"0000000000000000_0000000000000000_0010010001010111_1111001111100011"; -- 0.1419670515128682
	pesos_i(21919) := b"1111111111111111_1111111111111111_1111110110010111_0001101110001010"; -- -0.009413031310904634
	pesos_i(21920) := b"0000000000000000_0000000000000000_0001110010011110_1000100000111000"; -- 0.11179400795028568
	pesos_i(21921) := b"1111111111111111_1111111111111111_1110101110010000_0100100100011110"; -- -0.07982962618876235
	pesos_i(21922) := b"0000000000000000_0000000000000000_0001111100100001_1010101111111000"; -- 0.12160754009484485
	pesos_i(21923) := b"1111111111111111_1111111111111111_1111010101100011_0111111000000000"; -- -0.041450619674360166
	pesos_i(21924) := b"0000000000000000_0000000000000000_0001000111010110_0001010001101110"; -- 0.06967284864233653
	pesos_i(21925) := b"0000000000000000_0000000000000000_0010001011111111_1110101011101011"; -- 0.1367174933797299
	pesos_i(21926) := b"0000000000000000_0000000000000000_0010000010110100_1101110011111110"; -- 0.12775975414732707
	pesos_i(21927) := b"1111111111111111_1111111111111111_1111010000001001_1001110101111100"; -- -0.04672828402697687
	pesos_i(21928) := b"1111111111111111_1111111111111111_1101111110011101_0110101001011010"; -- -0.12650428113456358
	pesos_i(21929) := b"1111111111111111_1111111111111111_1110011110001101_1110101000101000"; -- -0.09549080403075576
	pesos_i(21930) := b"0000000000000000_0000000000000000_0001110001101101_0101001001101001"; -- 0.11104312010343553
	pesos_i(21931) := b"0000000000000000_0000000000000000_0000011101110101_0001101100101000"; -- 0.029130646919286185
	pesos_i(21932) := b"1111111111111111_1111111111111111_1111000000000111_1110111110010011"; -- -0.062378908748632306
	pesos_i(21933) := b"0000000000000000_0000000000000000_0010000111001000_1111010100011010"; -- 0.13197261696233387
	pesos_i(21934) := b"0000000000000000_0000000000000000_0000000100000011_0011100011111011"; -- 0.003955422732750606
	pesos_i(21935) := b"0000000000000000_0000000000000000_0001011100100101_1000110000100011"; -- 0.09041667796101446
	pesos_i(21936) := b"0000000000000000_0000000000000000_0000000011010000_0110010001010000"; -- 0.0031798073201046453
	pesos_i(21937) := b"1111111111111111_1111111111111111_1101110101010101_0111111101101101"; -- -0.1354141578380217
	pesos_i(21938) := b"0000000000000000_0000000000000000_0010010000000001_0000011001110100"; -- 0.1406406433684745
	pesos_i(21939) := b"1111111111111111_1111111111111111_1111000110101100_1111001110111100"; -- -0.05595471060579087
	pesos_i(21940) := b"1111111111111111_1111111111111111_1101011110101111_0010110111110000"; -- -0.15748322372252005
	pesos_i(21941) := b"1111111111111111_1111111111111111_1111101101111000_1110011000010000"; -- -0.017686482459914894
	pesos_i(21942) := b"1111111111111111_1111111111111111_1111101100010011_0101111001100010"; -- -0.019235707419402184
	pesos_i(21943) := b"0000000000000000_0000000000000000_0001101010010010_1000010010100100"; -- 0.10379818912963948
	pesos_i(21944) := b"0000000000000000_0000000000000000_0010010001001111_1101101000111001"; -- 0.1418434513773906
	pesos_i(21945) := b"0000000000000000_0000000000000000_0001101101001000_0111111011111110"; -- 0.10657495205395585
	pesos_i(21946) := b"0000000000000000_0000000000000000_0010000010001101_1011111100010111"; -- 0.12716287916246877
	pesos_i(21947) := b"0000000000000000_0000000000000000_0010000000000010_1001100010000100"; -- 0.12503960827604593
	pesos_i(21948) := b"1111111111111111_1111111111111111_1110001010111010_0001111111110001"; -- -0.11434746146287257
	pesos_i(21949) := b"1111111111111111_1111111111111111_1110110001001011_1000110111111100"; -- -0.07697212788578864
	pesos_i(21950) := b"1111111111111111_1111111111111111_1110000010011001_0000000000010010"; -- -0.12266540118369006
	pesos_i(21951) := b"1111111111111111_1111111111111111_1101100110100101_1100001110110001"; -- -0.14981438563360713
	pesos_i(21952) := b"1111111111111111_1111111111111111_1111011101110010_1110111000011010"; -- -0.033402556024120594
	pesos_i(21953) := b"0000000000000000_0000000000000000_0001000111010101_1110010110010101"; -- 0.06967005631324884
	pesos_i(21954) := b"0000000000000000_0000000000000000_0001110101110001_1000111010000000"; -- 0.11501398689970387
	pesos_i(21955) := b"1111111111111111_1111111111111111_1101101110111011_1101110100110101"; -- -0.14166467147485762
	pesos_i(21956) := b"0000000000000000_0000000000000000_0000000101011011_1111110111110001"; -- 0.00530993585728599
	pesos_i(21957) := b"1111111111111111_1111111111111111_1110111101101100_0010001001011011"; -- -0.06475625293632005
	pesos_i(21958) := b"1111111111111111_1111111111111111_1111101010100110_0100100000110001"; -- -0.020900238131939815
	pesos_i(21959) := b"0000000000000000_0000000000000000_0000100111001010_1011011011000101"; -- 0.03824941924091884
	pesos_i(21960) := b"1111111111111111_1111111111111111_1110111011101000_0011001001001000"; -- -0.06676946385995759
	pesos_i(21961) := b"1111111111111111_1111111111111111_1110000101100110_0010000101001001"; -- -0.11953536961705565
	pesos_i(21962) := b"1111111111111111_1111111111111111_1101111110100111_0110010111001001"; -- -0.12635196533619064
	pesos_i(21963) := b"0000000000000000_0000000000000000_0000010001000010_1110001001101101"; -- 0.016645576173218705
	pesos_i(21964) := b"1111111111111111_1111111111111111_1110010001101010_1110010011101010"; -- -0.10774392392809141
	pesos_i(21965) := b"0000000000000000_0000000000000000_0000100110110110_1111011111001001"; -- 0.03794811874633992
	pesos_i(21966) := b"0000000000000000_0000000000000000_0000010000011011_0011001011100110"; -- 0.016040021185894586
	pesos_i(21967) := b"0000000000000000_0000000000000000_0000001010110011_1100111101110110"; -- 0.010556188765908286
	pesos_i(21968) := b"0000000000000000_0000000000000000_0000110000101010_1011111000010001"; -- 0.04752719787375989
	pesos_i(21969) := b"0000000000000000_0000000000000000_0001001000101000_0100011011110011"; -- 0.07092708053448969
	pesos_i(21970) := b"0000000000000000_0000000000000000_0001001111010111_1010111010000000"; -- 0.07750979071329639
	pesos_i(21971) := b"0000000000000000_0000000000000000_0000110010000110_1110001111001011"; -- 0.04893325524988674
	pesos_i(21972) := b"1111111111111111_1111111111111111_1110000100001100_1101011011001101"; -- -0.12089784138264212
	pesos_i(21973) := b"1111111111111111_1111111111111111_1110001000100001_0101011010111111"; -- -0.11667878941980864
	pesos_i(21974) := b"0000000000000000_0000000000000000_0001001101100011_1111100111000101"; -- 0.07574425754270882
	pesos_i(21975) := b"0000000000000000_0000000000000000_0001100111001001_1001111011000100"; -- 0.10073272982133417
	pesos_i(21976) := b"0000000000000000_0000000000000000_0010000100101011_1010010010101100"; -- 0.12957219318254662
	pesos_i(21977) := b"0000000000000000_0000000000000000_0000110001001101_1011100001000011"; -- 0.04806090950441555
	pesos_i(21978) := b"1111111111111111_1111111111111111_1111001111010100_1011011100001000"; -- -0.04753547732127706
	pesos_i(21979) := b"1111111111111111_1111111111111111_1110111101101010_0011100101010010"; -- -0.06478540173433092
	pesos_i(21980) := b"1111111111111111_1111111111111111_1101101011000001_1111101011100010"; -- -0.14547760001828963
	pesos_i(21981) := b"0000000000000000_0000000000000000_0000011100011111_1010010011010101"; -- 0.027826597116428042
	pesos_i(21982) := b"0000000000000000_0000000000000000_0001010000010100_0110100011111101"; -- 0.07843643351073928
	pesos_i(21983) := b"1111111111111111_1111111111111111_1110000010011100_0111011110000001"; -- -0.12261250594828615
	pesos_i(21984) := b"1111111111111111_1111111111111111_1110011101110111_0010011010101001"; -- -0.09583814976049525
	pesos_i(21985) := b"1111111111111111_1111111111111111_1111001010101010_0111111101011010"; -- -0.05208591515799203
	pesos_i(21986) := b"0000000000000000_0000000000000000_0010010001101101_1110010001110110"; -- 0.14230182533390756
	pesos_i(21987) := b"0000000000000000_0000000000000000_0000111011011111_1010111011000100"; -- 0.05810062676371297
	pesos_i(21988) := b"0000000000000000_0000000000000000_0010000111101110_1100111100010011"; -- 0.1325501844670949
	pesos_i(21989) := b"1111111111111111_1111111111111111_1110000011111101_1010010001010011"; -- -0.12112973177409803
	pesos_i(21990) := b"0000000000000000_0000000000000000_0001010010110110_1100011111110010"; -- 0.08091401733780355
	pesos_i(21991) := b"1111111111111111_1111111111111111_1111001010010011_1110011000000010"; -- -0.05243074837284921
	pesos_i(21992) := b"1111111111111111_1111111111111111_1110010010110011_0011000000000110"; -- -0.10664081444366795
	pesos_i(21993) := b"1111111111111111_1111111111111111_1110110010010101_1011110011001000"; -- -0.07584018811745132
	pesos_i(21994) := b"0000000000000000_0000000000000000_0000000010101011_1110000101000010"; -- 0.002622679388961479
	pesos_i(21995) := b"0000000000000000_0000000000000000_0000000001111110_0100101010001010"; -- 0.001927050313873677
	pesos_i(21996) := b"0000000000000000_0000000000000000_0000101111010101_0111010001101100"; -- 0.046225811318564645
	pesos_i(21997) := b"0000000000000000_0000000000000000_0000100100001100_0101000010010111"; -- 0.03534415896950843
	pesos_i(21998) := b"1111111111111111_1111111111111111_1111100010001001_1111110110011110"; -- -0.02914442918999248
	pesos_i(21999) := b"0000000000000000_0000000000000000_0000001000010000_0001100111001110"; -- 0.008058178727249662
	pesos_i(22000) := b"1111111111111111_1111111111111111_1111101010010010_0111100101110011"; -- -0.021202477801721877
	pesos_i(22001) := b"1111111111111111_1111111111111111_1110001001111001_1111001001010001"; -- -0.11532674340692564
	pesos_i(22002) := b"1111111111111111_1111111111111111_1101111011101101_1001000110010111"; -- -0.12918748911859956
	pesos_i(22003) := b"1111111111111111_1111111111111111_1111010100011111_0101010110110110"; -- -0.0424906188851565
	pesos_i(22004) := b"0000000000000000_0000000000000000_0000101011111100_1001001000001100"; -- 0.04291641985330496
	pesos_i(22005) := b"0000000000000000_0000000000000000_0001111001101000_1011100010101101"; -- 0.11878542160498173
	pesos_i(22006) := b"1111111111111111_1111111111111111_1110101010110101_0010001000101110"; -- -0.08317362192369104
	pesos_i(22007) := b"0000000000000000_0000000000000000_0001011110001100_0111111010100010"; -- 0.09198752826650852
	pesos_i(22008) := b"0000000000000000_0000000000000000_0000010101010111_0010110000000000"; -- 0.020861387175690388
	pesos_i(22009) := b"0000000000000000_0000000000000000_0000001001110011_0001000001011010"; -- 0.009568235326386365
	pesos_i(22010) := b"1111111111111111_1111111111111111_1110110000001000_0011111011001010"; -- -0.07799918709338706
	pesos_i(22011) := b"0000000000000000_0000000000000000_0000110000111000_1011100110110100"; -- 0.04774056096168074
	pesos_i(22012) := b"1111111111111111_1111111111111111_1111011101111000_1001101011010000"; -- -0.033315967717745434
	pesos_i(22013) := b"0000000000000000_0000000000000000_0000100101111000_1110110101001001"; -- 0.03700144791258136
	pesos_i(22014) := b"1111111111111111_1111111111111111_1111111001011111_0110111000110100"; -- -0.006356346483663541
	pesos_i(22015) := b"0000000000000000_0000000000000000_0000001100011111_0001011101010010"; -- 0.012193162566283895
	pesos_i(22016) := b"1111111111111111_1111111111111111_1101100111101101_0110100011011000"; -- -0.1487211677602698
	pesos_i(22017) := b"1111111111111111_1111111111111111_1110100000000101_1001000100001101"; -- -0.09366506028133889
	pesos_i(22018) := b"1111111111111111_1111111111111111_1111010100101110_1010100011100100"; -- -0.04225677909369994
	pesos_i(22019) := b"0000000000000000_0000000000000000_0001100100100110_1110100011111110"; -- 0.09824997133868518
	pesos_i(22020) := b"0000000000000000_0000000000000000_0001001011010100_0110110011010000"; -- 0.07355384907779036
	pesos_i(22021) := b"1111111111111111_1111111111111111_1110110000000100_1101101011011000"; -- -0.07805092063280848
	pesos_i(22022) := b"1111111111111111_1111111111111111_1110110010010010_0110101110100110"; -- -0.07589080055541074
	pesos_i(22023) := b"0000000000000000_0000000000000000_0000111110111101_1010011010100100"; -- 0.06148759362712025
	pesos_i(22024) := b"1111111111111111_1111111111111111_1110101100011011_1101010001111111"; -- -0.08160659693539295
	pesos_i(22025) := b"1111111111111111_1111111111111111_1110100100010011_1111011111101000"; -- -0.08953905674217373
	pesos_i(22026) := b"1111111111111111_1111111111111111_1101101101110101_1110101101111111"; -- -0.14273193512946905
	pesos_i(22027) := b"0000000000000000_0000000000000000_0000011000100011_1010001011010011"; -- 0.023981262790684046
	pesos_i(22028) := b"1111111111111111_1111111111111111_1111010011000110_1001011101100000"; -- -0.04384473722020271
	pesos_i(22029) := b"1111111111111111_1111111111111111_1111000110000100_0111001011110110"; -- -0.05657273753599659
	pesos_i(22030) := b"0000000000000000_0000000000000000_0010000111100000_0111001011010111"; -- 0.13233106363570554
	pesos_i(22031) := b"1111111111111111_1111111111111111_1101101110000000_1001110000111001"; -- -0.1425688134918223
	pesos_i(22032) := b"0000000000000000_0000000000000000_0010010001101010_1111111010110101"; -- 0.14225761338163367
	pesos_i(22033) := b"1111111111111111_1111111111111111_1111100010101001_1000110000101100"; -- -0.028662909719558455
	pesos_i(22034) := b"0000000000000000_0000000000000000_0001001011000010_0011010101101011"; -- 0.07327588894847878
	pesos_i(22035) := b"1111111111111111_1111111111111111_1111000110111011_0010111000000111"; -- -0.055737612885623275
	pesos_i(22036) := b"0000000000000000_0000000000000000_0001111010101010_0000100011101010"; -- 0.11978202544217433
	pesos_i(22037) := b"0000000000000000_0000000000000000_0000010010101101_0100001000111110"; -- 0.01826871892161355
	pesos_i(22038) := b"1111111111111111_1111111111111111_1110110111100100_0001100010011000"; -- -0.07073828030552308
	pesos_i(22039) := b"1111111111111111_1111111111111111_1111011100000111_0010111111110011"; -- -0.035046580381367085
	pesos_i(22040) := b"0000000000000000_0000000000000000_0000011010000011_0011111101101101"; -- 0.025440181923551807
	pesos_i(22041) := b"1111111111111111_1111111111111111_1110001000100111_1100000100001101"; -- -0.1165809005984851
	pesos_i(22042) := b"1111111111111111_1111111111111111_1111110100000001_1010010010111011"; -- -0.011693672542421499
	pesos_i(22043) := b"0000000000000000_0000000000000000_0010001111001110_0011010001101001"; -- 0.139865184452041
	pesos_i(22044) := b"0000000000000000_0000000000000000_0000101011000001_0100100011010000"; -- 0.04201178614058001
	pesos_i(22045) := b"0000000000000000_0000000000000000_0001100100101000_0111111100101101"; -- 0.0982741817331439
	pesos_i(22046) := b"0000000000000000_0000000000000000_0001010101100001_0010000011100011"; -- 0.0835133127969955
	pesos_i(22047) := b"1111111111111111_1111111111111111_1101101100010010_0011100111011111"; -- -0.14425314251022858
	pesos_i(22048) := b"0000000000000000_0000000000000000_0000000000000010_1010000100001110"; -- 4.0117139772645554e-05
	pesos_i(22049) := b"1111111111111111_1111111111111111_1111101000000010_0010100100110000"; -- -0.023404527528326655
	pesos_i(22050) := b"0000000000000000_0000000000000000_0001111111011101_0100010100011001"; -- 0.12447006095546653
	pesos_i(22051) := b"0000000000000000_0000000000000000_0010011000001110_0111111110111100"; -- 0.14865873653019018
	pesos_i(22052) := b"1111111111111111_1111111111111111_1110100110110001_1010100000100011"; -- -0.08713292252603784
	pesos_i(22053) := b"0000000000000000_0000000000000000_0001110100100010_1001111110101001"; -- 0.11380956533346266
	pesos_i(22054) := b"0000000000000000_0000000000000000_0010010010101000_1101101011010110"; -- 0.14320152024134025
	pesos_i(22055) := b"0000000000000000_0000000000000000_0001000100111001_1100001110110101"; -- 0.06728766596484384
	pesos_i(22056) := b"0000000000000000_0000000000000000_0001010000110001_1110010001010011"; -- 0.07888628989372932
	pesos_i(22057) := b"0000000000000000_0000000000000000_0000111010001011_0001111010111000"; -- 0.056810302653856636
	pesos_i(22058) := b"0000000000000000_0000000000000000_0000111001111100_0011000100011001"; -- 0.056582516178923174
	pesos_i(22059) := b"1111111111111111_1111111111111111_1101010001001101_1111011000100100"; -- -0.17068540204644894
	pesos_i(22060) := b"1111111111111111_1111111111111111_1110011001000011_1110101111100110"; -- -0.10052610043133983
	pesos_i(22061) := b"1111111111111111_1111111111111111_1111100001000001_1100001000001000"; -- -0.03024661349429297
	pesos_i(22062) := b"1111111111111111_1111111111111111_1111000101010111_1000010100111001"; -- -0.05725829463965864
	pesos_i(22063) := b"0000000000000000_0000000000000000_0001100011010011_1001101101010011"; -- 0.09697886248230604
	pesos_i(22064) := b"1111111111111111_1111111111111111_1110000100100100_1001110110110111"; -- -0.12053503308038899
	pesos_i(22065) := b"1111111111111111_1111111111111111_1111011111100100_0010101011000000"; -- -0.0316746978933844
	pesos_i(22066) := b"0000000000000000_0000000000000000_0010000001010111_0000100001000000"; -- 0.12632800631369992
	pesos_i(22067) := b"1111111111111111_1111111111111111_1110001001001100_0000110011011000"; -- -0.11602706638177014
	pesos_i(22068) := b"0000000000000000_0000000000000000_0000101111110000_0100101010111111"; -- 0.04663531451986197
	pesos_i(22069) := b"1111111111111111_1111111111111111_1110010110000010_0101000110010110"; -- -0.10348024451853961
	pesos_i(22070) := b"0000000000000000_0000000000000000_0000100010111101_1100110100010100"; -- 0.034146134739502454
	pesos_i(22071) := b"1111111111111111_1111111111111111_1111110001010000_0101001101001010"; -- -0.014399332379109332
	pesos_i(22072) := b"1111111111111111_1111111111111111_1110110001000101_1100110100111001"; -- -0.07705991122138268
	pesos_i(22073) := b"1111111111111111_1111111111111111_1111111001111010_1111101011011010"; -- -0.005935975777858227
	pesos_i(22074) := b"1111111111111111_1111111111111111_1111011100100001_1111001011000110"; -- -0.03463823942909005
	pesos_i(22075) := b"0000000000000000_0000000000000000_0000101111100010_1100110111101110"; -- 0.04642951071077958
	pesos_i(22076) := b"0000000000000000_0000000000000000_0000010001101111_0110101010101110"; -- 0.017325084278637992
	pesos_i(22077) := b"1111111111111111_1111111111111111_1110101100110001_1100010001101110"; -- -0.08127186126594015
	pesos_i(22078) := b"0000000000000000_0000000000000000_0001001111101101_0100010101011110"; -- 0.07783921761035986
	pesos_i(22079) := b"1111111111111111_1111111111111111_1101111101001100_1110101100010101"; -- -0.12773257001049254
	pesos_i(22080) := b"1111111111111111_1111111111111111_1111011001011000_0101001110011010"; -- -0.037714743507356416
	pesos_i(22081) := b"0000000000000000_0000000000000000_0000100110000001_0101011111000001"; -- 0.03712986436267613
	pesos_i(22082) := b"0000000000000000_0000000000000000_0010100001110000_0101110010100111"; -- 0.15796450691221164
	pesos_i(22083) := b"0000000000000000_0000000000000000_0000110011001111_1001000000000110"; -- 0.050042153847857075
	pesos_i(22084) := b"0000000000000000_0000000000000000_0000001011111111_1110110100101100"; -- 0.011717627749654227
	pesos_i(22085) := b"1111111111111111_1111111111111111_1111111100010110_1000100101001011"; -- -0.0035623733206413396
	pesos_i(22086) := b"1111111111111111_1111111111111111_1101100101101100_1010001101000110"; -- -0.150686068879409
	pesos_i(22087) := b"0000000000000000_0000000000000000_0001001010001111_0011010111011100"; -- 0.07249771700102609
	pesos_i(22088) := b"1111111111111111_1111111111111111_1111010100101001_1110011011111110"; -- -0.04232937148757986
	pesos_i(22089) := b"1111111111111111_1111111111111111_1111010000000100_0110110111000010"; -- -0.04680742276131972
	pesos_i(22090) := b"1111111111111111_1111111111111111_1101100110111110_1110111011001101"; -- -0.14943034635980137
	pesos_i(22091) := b"0000000000000000_0000000000000000_0000101110111010_0010001101100100"; -- 0.04580899412527746
	pesos_i(22092) := b"1111111111111111_1111111111111111_1101110100000110_1100011010010100"; -- -0.13661536119303058
	pesos_i(22093) := b"1111111111111111_1111111111111111_1110111001100111_1011100110010111"; -- -0.06872978277631428
	pesos_i(22094) := b"1111111111111111_1111111111111111_1110101100010011_0111101001010110"; -- -0.08173404121933613
	pesos_i(22095) := b"0000000000000000_0000000000000000_0000100100100010_1001001000011110"; -- 0.035683758104325544
	pesos_i(22096) := b"0000000000000000_0000000000000000_0000110101010001_1011100010110011"; -- 0.052028220868423555
	pesos_i(22097) := b"0000000000000000_0000000000000000_0001111110011001_1011001010100011"; -- 0.1234389924136013
	pesos_i(22098) := b"0000000000000000_0000000000000000_0000111010100111_0010100110011111"; -- 0.057238198531883104
	pesos_i(22099) := b"1111111111111111_1111111111111111_1110001011100000_1110011010101001"; -- -0.11375578286461706
	pesos_i(22100) := b"0000000000000000_0000000000000000_0000011000011001_1110101100000011"; -- 0.023832977563718317
	pesos_i(22101) := b"0000000000000000_0000000000000000_0001100010100111_0001011110011000"; -- 0.09629962412293908
	pesos_i(22102) := b"0000000000000000_0000000000000000_0010000110011101_1010010011010101"; -- 0.13131170452420468
	pesos_i(22103) := b"1111111111111111_1111111111111111_1111001011000010_1011011110101001"; -- -0.05171634795032322
	pesos_i(22104) := b"1111111111111111_1111111111111111_1111000111111000_0011010010000011"; -- -0.05480644037106182
	pesos_i(22105) := b"0000000000000000_0000000000000000_0010010000110101_0010100011100111"; -- 0.14143615372866042
	pesos_i(22106) := b"0000000000000000_0000000000000000_0000000000011111_0011001001010011"; -- 0.0004760220707037877
	pesos_i(22107) := b"1111111111111111_1111111111111111_1111001111111110_1000001101001001"; -- -0.04689769236868458
	pesos_i(22108) := b"1111111111111111_1111111111111111_1101100111101111_0110011101001111"; -- -0.14869074165128568
	pesos_i(22109) := b"0000000000000000_0000000000000000_0000010110110110_1100111000000010"; -- 0.022320628737862787
	pesos_i(22110) := b"1111111111111111_1111111111111111_1111000011101100_0100111010000001"; -- -0.05889424649286574
	pesos_i(22111) := b"1111111111111111_1111111111111111_1101100001010110_0010000100110001"; -- -0.15493576577285229
	pesos_i(22112) := b"0000000000000000_0000000000000000_0010110101001011_0111100101111101"; -- 0.17693290034651826
	pesos_i(22113) := b"1111111111111111_1111111111111111_1111110111000010_0100000110001110"; -- -0.00875463756642253
	pesos_i(22114) := b"1111111111111111_1111111111111111_1111001011001111_0010010110110001"; -- -0.05152668408148201
	pesos_i(22115) := b"1111111111111111_1111111111111111_1110100100000111_0110010001101110"; -- -0.08973095249066872
	pesos_i(22116) := b"0000000000000000_0000000000000000_0000011100101001_1100011011001011"; -- 0.027981209289773473
	pesos_i(22117) := b"0000000000000000_0000000000000000_0001101101010001_0000011101000011"; -- 0.1067051447930453
	pesos_i(22118) := b"1111111111111111_1111111111111111_1111001101001001_1100010101111011"; -- -0.04965558754700887
	pesos_i(22119) := b"1111111111111111_1111111111111111_1110010101000000_1111010110001100"; -- -0.10447755186717238
	pesos_i(22120) := b"1111111111111111_1111111111111111_1101101100010101_1000001001100110"; -- -0.14420304298789433
	pesos_i(22121) := b"1111111111111111_1111111111111111_1110011101001011_0011110101100010"; -- -0.0965081820776826
	pesos_i(22122) := b"0000000000000000_0000000000000000_0000111101111101_0110110101000011"; -- 0.060507611101316486
	pesos_i(22123) := b"1111111111111111_1111111111111111_1111101000000001_1000010000100111"; -- -0.023414364285118693
	pesos_i(22124) := b"1111111111111111_1111111111111111_1111010111001100_0001100011010000"; -- -0.03985447800836147
	pesos_i(22125) := b"1111111111111111_1111111111111111_1111110010001001_1000111011001011"; -- -0.01352603484987912
	pesos_i(22126) := b"1111111111111111_1111111111111111_1111010111100011_1000101111100001"; -- -0.039496667421271364
	pesos_i(22127) := b"1111111111111111_1111111111111111_1111110111101100_0111101010011001"; -- -0.00811036828423803
	pesos_i(22128) := b"0000000000000000_0000000000000000_0001110101110001_1101100000010010"; -- 0.11501837192172316
	pesos_i(22129) := b"1111111111111111_1111111111111111_1110111110011110_1001011000101001"; -- -0.0639864109977593
	pesos_i(22130) := b"0000000000000000_0000000000000000_0000001010011100_1111011010110001"; -- 0.01020757507001309
	pesos_i(22131) := b"0000000000000000_0000000000000000_0010100010000010_1100001110101010"; -- 0.15824530498419404
	pesos_i(22132) := b"0000000000000000_0000000000000000_0010010100100110_1000101111110111"; -- 0.14511942657417473
	pesos_i(22133) := b"1111111111111111_1111111111111111_1110100101010110_1110011001111001"; -- -0.08851775683248257
	pesos_i(22134) := b"1111111111111111_1111111111111111_1110010010111100_1111101111101001"; -- -0.10649133265113772
	pesos_i(22135) := b"0000000000000000_0000000000000000_0001101011001010_1000111011101010"; -- 0.10465329371786186
	pesos_i(22136) := b"0000000000000000_0000000000000000_0000100001111010_1001101111001010"; -- 0.03312085793499062
	pesos_i(22137) := b"0000000000000000_0000000000000000_0000010010010111_0110111001000110"; -- 0.017935649967483147
	pesos_i(22138) := b"1111111111111111_1111111111111111_1111100001000111_0111000011100011"; -- -0.030159897333516872
	pesos_i(22139) := b"1111111111111111_1111111111111111_1111111110011101_1101101110001110"; -- -0.0014975337212506388
	pesos_i(22140) := b"1111111111111111_1111111111111111_1110001111011000_1010010110000010"; -- -0.10997548646101869
	pesos_i(22141) := b"0000000000000000_0000000000000000_0001111000100001_1000010010010010"; -- 0.11769894182349899
	pesos_i(22142) := b"0000000000000000_0000000000000000_0000001111110111_0000111111101110"; -- 0.015488620378049335
	pesos_i(22143) := b"1111111111111111_1111111111111111_1110010100011000_0100110110001010"; -- -0.1050979172781853
	pesos_i(22144) := b"0000000000000000_0000000000000000_0010110111000000_0101110111000110"; -- 0.17871652676401528
	pesos_i(22145) := b"1111111111111111_1111111111111111_1110100101111111_0110100110001011"; -- -0.08789959296739625
	pesos_i(22146) := b"0000000000000000_0000000000000000_0000101000000111_1101011001011111"; -- 0.03918208892217879
	pesos_i(22147) := b"0000000000000000_0000000000000000_0000001111010101_0111101100001111"; -- 0.014976207002546212
	pesos_i(22148) := b"0000000000000000_0000000000000000_0000011001100001_0000110011011010"; -- 0.0249183686468496
	pesos_i(22149) := b"1111111111111111_1111111111111111_1111011001000000_0010000110101011"; -- -0.03808393082185672
	pesos_i(22150) := b"0000000000000000_0000000000000000_0000010100011000_1100001000010000"; -- 0.01990902804354883
	pesos_i(22151) := b"1111111111111111_1111111111111111_1110100100100110_0000101010110011"; -- -0.08926327840174933
	pesos_i(22152) := b"1111111111111111_1111111111111111_1110010010100001_1011111101000010"; -- -0.10690693502664231
	pesos_i(22153) := b"0000000000000000_0000000000000000_0010010100100101_1111010111010000"; -- 0.1451104766647983
	pesos_i(22154) := b"0000000000000000_0000000000000000_0000101110111001_1100110010111100"; -- 0.04580382900262199
	pesos_i(22155) := b"1111111111111111_1111111111111111_1110000110000101_0110111001001000"; -- -0.11905775766935899
	pesos_i(22156) := b"0000000000000000_0000000000000000_0010001010010010_0000000001100011"; -- 0.13504030626869928
	pesos_i(22157) := b"0000000000000000_0000000000000000_0001001111011111_0100110100011001"; -- 0.0776260553794455
	pesos_i(22158) := b"1111111111111111_1111111111111111_1111010110100101_1110010000110101"; -- -0.0404374476154846
	pesos_i(22159) := b"0000000000000000_0000000000000000_0000101111101010_1000000111010100"; -- 0.04654704500273624
	pesos_i(22160) := b"0000000000000000_0000000000000000_0010011101010001_0011010001111111"; -- 0.15358284085777554
	pesos_i(22161) := b"1111111111111111_1111111111111111_1110101110010111_1100110100110000"; -- -0.07971494272993887
	pesos_i(22162) := b"0000000000000000_0000000000000000_0010001110111010_0100010111111100"; -- 0.13956105605966124
	pesos_i(22163) := b"1111111111111111_1111111111111111_1111111110011011_0110001111110110"; -- -0.001535179641110973
	pesos_i(22164) := b"0000000000000000_0000000000000000_0001111111100101_0011111110000110"; -- 0.12459179904230218
	pesos_i(22165) := b"1111111111111111_1111111111111111_1110100110101110_1100000110001111"; -- -0.08717718371218137
	pesos_i(22166) := b"0000000000000000_0000000000000000_0001000010010000_1101000011111111"; -- 0.06470972282376837
	pesos_i(22167) := b"0000000000000000_0000000000000000_0000100011101000_1011100111001110"; -- 0.03480111386091292
	pesos_i(22168) := b"0000000000000000_0000000000000000_0000100110011111_0100101111101000"; -- 0.03758692188996496
	pesos_i(22169) := b"1111111111111111_1111111111111111_1110001111100000_1010000010100000"; -- -0.10985370720650607
	pesos_i(22170) := b"1111111111111111_1111111111111111_1111011010111111_1111001010000000"; -- -0.03613361712680126
	pesos_i(22171) := b"0000000000000000_0000000000000000_0001000100110100_0001001110101101"; -- 0.06720087988523725
	pesos_i(22172) := b"1111111111111111_1111111111111111_1110000001001110_1100010001100101"; -- -0.12379810850610212
	pesos_i(22173) := b"1111111111111111_1111111111111111_1110110101010101_0000101101001101"; -- -0.07292107940649033
	pesos_i(22174) := b"0000000000000000_0000000000000000_0001001001110101_0001100110101001"; -- 0.0720993077832711
	pesos_i(22175) := b"0000000000000000_0000000000000000_0010011110011010_0011000111101100"; -- 0.15469657908951073
	pesos_i(22176) := b"0000000000000000_0000000000000000_0001110101000000_1000101010010110"; -- 0.11426607282906853
	pesos_i(22177) := b"0000000000000000_0000000000000000_0000111000011100_0001011101000110"; -- 0.05511613327472913
	pesos_i(22178) := b"0000000000000000_0000000000000000_0000100111100000_0110010010100010"; -- 0.03858021696671522
	pesos_i(22179) := b"0000000000000000_0000000000000000_0000110110111110_1100011101010101"; -- 0.053692300956616215
	pesos_i(22180) := b"0000000000000000_0000000000000000_0001110010000010_0101100010001011"; -- 0.1113639202255445
	pesos_i(22181) := b"0000000000000000_0000000000000000_0001001011100110_0000101001010011"; -- 0.07382263687020035
	pesos_i(22182) := b"0000000000000000_0000000000000000_0001100001101001_0111110100110111"; -- 0.09535963619636866
	pesos_i(22183) := b"1111111111111111_1111111111111111_1110100110011101_0101010010111111"; -- -0.08744306893266814
	pesos_i(22184) := b"0000000000000000_0000000000000000_0000010010100010_0101111001101011"; -- 0.018102551483154185
	pesos_i(22185) := b"0000000000000000_0000000000000000_0000011010011010_1011110000001110"; -- 0.02579856252831718
	pesos_i(22186) := b"0000000000000000_0000000000000000_0010100000101101_1111010000001100"; -- 0.1569511918302469
	pesos_i(22187) := b"1111111111111111_1111111111111111_1101110010000111_0011011111111010"; -- -0.13856172712686074
	pesos_i(22188) := b"1111111111111111_1111111111111111_1101110110100000_0010111111010111"; -- -0.13427449218861737
	pesos_i(22189) := b"1111111111111111_1111111111111111_1111011000000111_1100001100011100"; -- -0.0389440591602034
	pesos_i(22190) := b"0000000000000000_0000000000000000_0010000000101110_1101111110000000"; -- 0.12571522591830647
	pesos_i(22191) := b"1111111111111111_1111111111111111_1111101110001001_1010011010110000"; -- -0.01743086054835244
	pesos_i(22192) := b"1111111111111111_1111111111111111_1110010111001111_0011010110110100"; -- -0.1023069797100983
	pesos_i(22193) := b"1111111111111111_1111111111111111_1111111000000101_0011010101100001"; -- -0.007733024311239685
	pesos_i(22194) := b"0000000000000000_0000000000000000_0001010011010001_0000100101101000"; -- 0.08131464759588389
	pesos_i(22195) := b"1111111111111111_1111111111111111_1111000110110000_0111111111101100"; -- -0.055900578349392986
	pesos_i(22196) := b"1111111111111111_1111111111111111_1111001011101001_1100110100111001"; -- -0.051119969959234846
	pesos_i(22197) := b"1111111111111111_1111111111111111_1110001001010101_0111000011010001"; -- -0.11588377864116707
	pesos_i(22198) := b"1111111111111111_1111111111111111_1111000111111011_0001001111110011"; -- -0.054762604812894265
	pesos_i(22199) := b"0000000000000000_0000000000000000_0010011001001010_1001101010010000"; -- 0.1495758630919854
	pesos_i(22200) := b"0000000000000000_0000000000000000_0000101110000011_0110111101100001"; -- 0.04497429012631632
	pesos_i(22201) := b"0000000000000000_0000000000000000_0010000011100100_0000111111011001"; -- 0.12847994850072866
	pesos_i(22202) := b"1111111111111111_1111111111111111_1111010111110111_1101011111101110"; -- -0.03918695863682113
	pesos_i(22203) := b"0000000000000000_0000000000000000_0001101110010000_1100110001001001"; -- 0.10767819191159676
	pesos_i(22204) := b"1111111111111111_1111111111111111_1110110101101101_1000111000101000"; -- -0.0725470689255927
	pesos_i(22205) := b"0000000000000000_0000000000000000_0000011010111001_1101001011111010"; -- 0.02627295115592113
	pesos_i(22206) := b"1111111111111111_1111111111111111_1110011001000001_1001001111001001"; -- -0.10056186996212597
	pesos_i(22207) := b"1111111111111111_1111111111111111_1110111011100010_1000011010011101"; -- -0.06685599005103848
	pesos_i(22208) := b"1111111111111111_1111111111111111_1111001010100010_0001111000000101"; -- -0.05221378680924414
	pesos_i(22209) := b"0000000000000000_0000000000000000_0001100010000001_1010110000010011"; -- 0.09572864026758221
	pesos_i(22210) := b"0000000000000000_0000000000000000_0000111011010001_0101000011100010"; -- 0.057881407859949593
	pesos_i(22211) := b"0000000000000000_0000000000000000_0001011100010110_1110001011001111"; -- 0.09019296218486945
	pesos_i(22212) := b"1111111111111111_1111111111111111_1110111101110010_1001010111111001"; -- -0.06465780909415633
	pesos_i(22213) := b"1111111111111111_1111111111111111_1111100001111111_1111100110011111"; -- -0.029297255262751655
	pesos_i(22214) := b"0000000000000000_0000000000000000_0001011100100001_0100111100001011"; -- 0.0903520013092428
	pesos_i(22215) := b"1111111111111111_1111111111111111_1110001110010001_1010010111011100"; -- -0.11105883958274859
	pesos_i(22216) := b"0000000000000000_0000000000000000_0001011110011000_0011001101110010"; -- 0.09216615239752529
	pesos_i(22217) := b"0000000000000000_0000000000000000_0000101000100111_0001011010110010"; -- 0.03965894547860638
	pesos_i(22218) := b"0000000000000000_0000000000000000_0000000101011100_1111010011011011"; -- 0.005324653189223884
	pesos_i(22219) := b"1111111111111111_1111111111111111_1110100111001010_1101011001000011"; -- -0.08674870370821457
	pesos_i(22220) := b"0000000000000000_0000000000000000_0010000111011100_1111100001101011"; -- 0.13227799043476018
	pesos_i(22221) := b"1111111111111111_1111111111111111_1111011101101100_1111101100010011"; -- -0.033493335578616286
	pesos_i(22222) := b"0000000000000000_0000000000000000_0001000000000001_1101001100111100"; -- 0.06252784944560756
	pesos_i(22223) := b"0000000000000000_0000000000000000_0000011010000100_1100001101110110"; -- 0.025463310618456247
	pesos_i(22224) := b"1111111111111111_1111111111111111_1111001100100011_0010101100111001"; -- -0.05024461603582343
	pesos_i(22225) := b"1111111111111111_1111111111111111_1111101010001010_0001111101110101"; -- -0.021329912197148495
	pesos_i(22226) := b"1111111111111111_1111111111111111_1110110010111001_1000010011010110"; -- -0.07529420649287724
	pesos_i(22227) := b"0000000000000000_0000000000000000_0000110010111110_1010010101001110"; -- 0.049784022860898045
	pesos_i(22228) := b"1111111111111111_1111111111111111_1111000111001111_0000110101100000"; -- -0.055434383375108406
	pesos_i(22229) := b"0000000000000000_0000000000000000_0001100111111101_1110100110010111"; -- 0.10153064675933926
	pesos_i(22230) := b"0000000000000000_0000000000000000_0000000001010110_1100001110110001"; -- 0.001323920014037698
	pesos_i(22231) := b"0000000000000000_0000000000000000_0001000101001010_0010000101100110"; -- 0.06753739111392251
	pesos_i(22232) := b"0000000000000000_0000000000000000_0001100111001000_1001101110010011"; -- 0.10071728085189492
	pesos_i(22233) := b"1111111111111111_1111111111111111_1110000101101011_1101110011101010"; -- -0.11944789211407278
	pesos_i(22234) := b"0000000000000000_0000000000000000_0001001111100000_1011000011001001"; -- 0.07764725599202742
	pesos_i(22235) := b"1111111111111111_1111111111111111_1101100101000011_1110010101010000"; -- -0.15130774315288043
	pesos_i(22236) := b"1111111111111111_1111111111111111_1111110001000000_0100111000000001"; -- -0.014643788017040364
	pesos_i(22237) := b"1111111111111111_1111111111111111_1111010100100011_1011110000111001"; -- -0.042423473413313255
	pesos_i(22238) := b"1111111111111111_1111111111111111_1110111100001001_1001010101010001"; -- -0.06626002103091837
	pesos_i(22239) := b"1111111111111111_1111111111111111_1101111011010011_0110101001101011"; -- -0.12958655254059853
	pesos_i(22240) := b"1111111111111111_1111111111111111_1111011010101100_1110101101111111"; -- -0.036423951557339886
	pesos_i(22241) := b"0000000000000000_0000000000000000_0000111110010111_0000001101000000"; -- 0.060898020958233795
	pesos_i(22242) := b"1111111111111111_1111111111111111_1101100100010111_1010101101000111"; -- -0.1519825890050207
	pesos_i(22243) := b"0000000000000000_0000000000000000_0010010100101010_0101001001011101"; -- 0.14517702833381038
	pesos_i(22244) := b"0000000000000000_0000000000000000_0010000001110000_0111011000010010"; -- 0.12671602198176213
	pesos_i(22245) := b"0000000000000000_0000000000000000_0000011110101101_1001001011001111"; -- 0.0299922709259031
	pesos_i(22246) := b"0000000000000000_0000000000000000_0001010101100000_0111001101010110"; -- 0.08350296824574709
	pesos_i(22247) := b"0000000000000000_0000000000000000_0000100000011001_1100001111100001"; -- 0.03164314505862867
	pesos_i(22248) := b"1111111111111111_1111111111111111_1101101000000101_1010110011110111"; -- -0.1483508964839867
	pesos_i(22249) := b"1111111111111111_1111111111111111_1101110011001000_0110110001110110"; -- -0.1375667774153755
	pesos_i(22250) := b"1111111111111111_1111111111111111_1110101110010101_1111010010000000"; -- -0.07974311713866185
	pesos_i(22251) := b"1111111111111111_1111111111111111_1110101101011111_0001010100011001"; -- -0.08058040755131843
	pesos_i(22252) := b"1111111111111111_1111111111111111_1110000000001100_0000000110101001"; -- -0.12481679564709927
	pesos_i(22253) := b"1111111111111111_1111111111111111_1101111001111101_0011110010101001"; -- -0.13090153579286992
	pesos_i(22254) := b"1111111111111111_1111111111111111_1110110101011000_1111011111000110"; -- -0.07286120801795559
	pesos_i(22255) := b"0000000000000000_0000000000000000_0000111000110011_0001001100110010"; -- 0.05546684231352545
	pesos_i(22256) := b"1111111111111111_1111111111111111_1101100000001001_0101010110100000"; -- -0.15610756715925547
	pesos_i(22257) := b"0000000000000000_0000000000000000_0000011010001010_0001101011000110"; -- 0.025544808785134078
	pesos_i(22258) := b"1111111111111111_1111111111111111_1111110101111100_1100101101001000"; -- -0.009814543685475725
	pesos_i(22259) := b"0000000000000000_0000000000000000_0001010100001011_1101100011011111"; -- 0.08221202321286283
	pesos_i(22260) := b"0000000000000000_0000000000000000_0000110001011100_1001000100111011"; -- 0.04828746499457817
	pesos_i(22261) := b"1111111111111111_1111111111111111_1101101101100011_1001000010111000"; -- -0.14301200389837512
	pesos_i(22262) := b"0000000000000000_0000000000000000_0000001000111101_0111010101001111"; -- 0.008750278238184177
	pesos_i(22263) := b"1111111111111111_1111111111111111_1111010001010111_0011010110111010"; -- -0.04554428293526601
	pesos_i(22264) := b"1111111111111111_1111111111111111_1110100001100110_0110010101000110"; -- -0.09218756725831227
	pesos_i(22265) := b"0000000000000000_0000000000000000_0001010101000111_1110011111001110"; -- 0.08312844065039168
	pesos_i(22266) := b"0000000000000000_0000000000000000_0001111111101011_0011001011011110"; -- 0.12468259737334453
	pesos_i(22267) := b"1111111111111111_1111111111111111_1101101001011110_1011011011000001"; -- -0.1469922807794992
	pesos_i(22268) := b"0000000000000000_0000000000000000_0000010010100110_0101101011101010"; -- 0.018163377810018033
	pesos_i(22269) := b"1111111111111111_1111111111111111_1111111111111110_0111111100010010"; -- -2.2943705888817373e-05
	pesos_i(22270) := b"1111111111111111_1111111111111111_1110111111001011_0000111001000010"; -- -0.0633078659659055
	pesos_i(22271) := b"0000000000000000_0000000000000000_0010000001001001_0101001000110010"; -- 0.12611879085924377
	pesos_i(22272) := b"1111111111111111_1111111111111111_1110101111110100_1110011000010110"; -- -0.07829439125898105
	pesos_i(22273) := b"1111111111111111_1111111111111111_1110001011010111_1111111010110101"; -- -0.11389167868839656
	pesos_i(22274) := b"0000000000000000_0000000000000000_0000100011111110_0101110010100011"; -- 0.03513125410529125
	pesos_i(22275) := b"0000000000000000_0000000000000000_0000100010101011_1000000011011010"; -- 0.03386693297057371
	pesos_i(22276) := b"1111111111111111_1111111111111111_1110110100101000_0110101001001000"; -- -0.07360206350247978
	pesos_i(22277) := b"1111111111111111_1111111111111111_1110011110111101_0011010010001011"; -- -0.09476920699324852
	pesos_i(22278) := b"1111111111111111_1111111111111111_1111110010001010_0110100000100111"; -- -0.013513079070203736
	pesos_i(22279) := b"0000000000000000_0000000000000000_0010011001110101_1011001010001110"; -- 0.15023342104610418
	pesos_i(22280) := b"0000000000000000_0000000000000000_0010000001010001_0100011000000000"; -- 0.12624013427575267
	pesos_i(22281) := b"1111111111111111_1111111111111111_1111011110001000_1100110100011110"; -- -0.033068828675027084
	pesos_i(22282) := b"1111111111111111_1111111111111111_1111100101000111_0100111110110111"; -- -0.026255624713907577
	pesos_i(22283) := b"0000000000000000_0000000000000000_0001000110000111_1111001011010010"; -- 0.0684806598106366
	pesos_i(22284) := b"1111111111111111_1111111111111111_1111001011100111_0100001011100111"; -- -0.051158731975929156
	pesos_i(22285) := b"1111111111111111_1111111111111111_1110011111000100_0111001010011011"; -- -0.09465869621349195
	pesos_i(22286) := b"1111111111111111_1111111111111111_1110101010000010_0011110111000011"; -- -0.0839501760699698
	pesos_i(22287) := b"0000000000000000_0000000000000000_0001110010001011_1011110111111000"; -- 0.11150729479342415
	pesos_i(22288) := b"0000000000000000_0000000000000000_0001011101111000_0101011111111111"; -- 0.09168004966898656
	pesos_i(22289) := b"0000000000000000_0000000000000000_0001110100010000_0000100100111010"; -- 0.11352594059993579
	pesos_i(22290) := b"1111111111111111_1111111111111111_1110100101100011_1110100110000010"; -- -0.08831921178972404
	pesos_i(22291) := b"0000000000000000_0000000000000000_0001101001100101_0011000010101011"; -- 0.10310653850746335
	pesos_i(22292) := b"1111111111111111_1111111111111111_1110111010011010_1001000011010001"; -- -0.06795401473231474
	pesos_i(22293) := b"1111111111111111_1111111111111111_1111011000110100_0010101001010101"; -- -0.03826651970908483
	pesos_i(22294) := b"0000000000000000_0000000000000000_0001110110101011_0011000010001000"; -- 0.11589339552913822
	pesos_i(22295) := b"0000000000000000_0000000000000000_0010011010111001_0101100001000101"; -- 0.1512656372535312
	pesos_i(22296) := b"0000000000000000_0000000000000000_0000100010101101_0111011000111101"; -- 0.033896818082890925
	pesos_i(22297) := b"1111111111111111_1111111111111111_1111011010000000_1111110101101011"; -- -0.03709427000673204
	pesos_i(22298) := b"1111111111111111_1111111111111111_1110100100001101_0111001101101001"; -- -0.08963850681852578
	pesos_i(22299) := b"1111111111111111_1111111111111111_1110111010110101_0000110000001011"; -- -0.06754994136497477
	pesos_i(22300) := b"1111111111111111_1111111111111111_1111010110110111_1101100001101011"; -- -0.04016349216883281
	pesos_i(22301) := b"1111111111111111_1111111111111111_1110001011111010_0000010010111001"; -- -0.113372521290958
	pesos_i(22302) := b"1111111111111111_1111111111111111_1111111010110111_1000111110001110"; -- -0.005011584968939478
	pesos_i(22303) := b"0000000000000000_0000000000000000_0000001101011111_0010000101110111"; -- 0.013170329530838505
	pesos_i(22304) := b"0000000000000000_0000000000000000_0001001010110000_0000000110001011"; -- 0.07299813885823493
	pesos_i(22305) := b"1111111111111111_1111111111111111_1111111000000011_1111110111100000"; -- -0.007751591583201279
	pesos_i(22306) := b"0000000000000000_0000000000000000_0001111100010110_1100101101001100"; -- 0.12144156091362786
	pesos_i(22307) := b"1111111111111111_1111111111111111_1110100010010111_1001001001010111"; -- -0.09143720030611299
	pesos_i(22308) := b"1111111111111111_1111111111111111_1111010001011110_0100000101111110"; -- -0.04543677025842304
	pesos_i(22309) := b"0000000000000000_0000000000000000_0001100101101100_0011000010001111"; -- 0.09930709361074935
	pesos_i(22310) := b"0000000000000000_0000000000000000_0000000000011011_0111111011100111"; -- 0.0004195511875850971
	pesos_i(22311) := b"0000000000000000_0000000000000000_0010101110100110_0110001001100110"; -- 0.17050757389242951
	pesos_i(22312) := b"0000000000000000_0000000000000000_0000001011110010_1101110101011000"; -- 0.011518320049502569
	pesos_i(22313) := b"1111111111111111_1111111111111111_1101011000001000_0001100110100000"; -- -0.16393890241360543
	pesos_i(22314) := b"0000000000000000_0000000000000000_0010001010011010_0010001010000111"; -- 0.1351644115681166
	pesos_i(22315) := b"1111111111111111_1111111111111111_1110010001100101_0000001100011000"; -- -0.1078336779345433
	pesos_i(22316) := b"1111111111111111_1111111111111111_1111101001001000_1010000101110101"; -- -0.022329243656276764
	pesos_i(22317) := b"0000000000000000_0000000000000000_0010100000010000_1110110011001011"; -- 0.15650825455254067
	pesos_i(22318) := b"0000000000000000_0000000000000000_0010010001111110_0010111011010111"; -- 0.14255039924847204
	pesos_i(22319) := b"0000000000000000_0000000000000000_0001111000100110_1010000111010011"; -- 0.11777697937250754
	pesos_i(22320) := b"1111111111111111_1111111111111111_1111000110000011_1000100011000000"; -- -0.05658669761766016
	pesos_i(22321) := b"0000000000000000_0000000000000000_0000101001111100_0101010110010011"; -- 0.040959690380996554
	pesos_i(22322) := b"0000000000000000_0000000000000000_0000000001011110_1000000000011000"; -- 0.0014419611932585067
	pesos_i(22323) := b"0000000000000000_0000000000000000_0010010110110000_1010011010110010"; -- 0.14722673270881262
	pesos_i(22324) := b"0000000000000000_0000000000000000_0000010110100001_1000000011010100"; -- 0.02199559383909578
	pesos_i(22325) := b"1111111111111111_1111111111111111_1101010101000010_1011011000001111"; -- -0.16695081846374563
	pesos_i(22326) := b"0000000000000000_0000000000000000_0001001110000100_0100001100111010"; -- 0.07623691725212482
	pesos_i(22327) := b"0000000000000000_0000000000000000_0001001000001011_0101111000101101"; -- 0.07048595996985167
	pesos_i(22328) := b"1111111111111111_1111111111111111_1101101110111110_0000111101011101"; -- -0.14163116445642787
	pesos_i(22329) := b"1111111111111111_1111111111111111_1110111010010111_0011011101010111"; -- -0.06800512433577892
	pesos_i(22330) := b"1111111111111111_1111111111111111_1111001011111011_1000010100000000"; -- -0.050849616586118224
	pesos_i(22331) := b"1111111111111111_1111111111111111_1110011111111000_0111000011001100"; -- -0.09386534712023369
	pesos_i(22332) := b"0000000000000000_0000000000000000_0000001101011100_1000110101110111"; -- 0.013130990449712566
	pesos_i(22333) := b"0000000000000000_0000000000000000_0001110000011111_0001100010000111"; -- 0.10984948451926456
	pesos_i(22334) := b"1111111111111111_1111111111111111_1110011110010000_0101010000011101"; -- -0.09545397089773718
	pesos_i(22335) := b"0000000000000000_0000000000000000_0001101010010000_1011101000011101"; -- 0.1037708587328731
	pesos_i(22336) := b"1111111111111111_1111111111111111_1110100011010111_1001011100110010"; -- -0.09046034833858278
	pesos_i(22337) := b"0000000000000000_0000000000000000_0000011010110101_0001100000111100"; -- 0.026200785279714582
	pesos_i(22338) := b"1111111111111111_1111111111111111_1111000011011000_1010010100101001"; -- -0.05919425724437063
	pesos_i(22339) := b"1111111111111111_1111111111111111_1110110111101001_0100101011010011"; -- -0.07065899234312967
	pesos_i(22340) := b"0000000000000000_0000000000000000_0000101111101111_1110110110100101"; -- 0.04662976536575273
	pesos_i(22341) := b"1111111111111111_1111111111111111_1110001110100011_0101110111101011"; -- -0.11078846944042324
	pesos_i(22342) := b"1111111111111111_1111111111111111_1110101110110110_0110000101011100"; -- -0.0792483473745738
	pesos_i(22343) := b"1111111111111111_1111111111111111_1110011000010101_0010100011011000"; -- -0.10123963104603455
	pesos_i(22344) := b"1111111111111111_1111111111111111_1110110001010110_0010101000011001"; -- -0.07681023482628434
	pesos_i(22345) := b"1111111111111111_1111111111111111_1110101110000010_1011001010011100"; -- -0.08003696142311842
	pesos_i(22346) := b"1111111111111111_1111111111111111_1110110001111000_0100011001100101"; -- -0.07628974938643511
	pesos_i(22347) := b"1111111111111111_1111111111111111_1111011101001110_0100000011100100"; -- -0.03396219678452086
	pesos_i(22348) := b"1111111111111111_1111111111111111_1111101000101010_1110111111111111"; -- -0.022782326043899435
	pesos_i(22349) := b"1111111111111111_1111111111111111_1110011011000001_0000100011001000"; -- -0.09861703021816531
	pesos_i(22350) := b"1111111111111111_1111111111111111_1110110011110111_0010101110101001"; -- -0.07435347675948552
	pesos_i(22351) := b"1111111111111111_1111111111111111_1101111111001010_0011100111011110"; -- -0.1258205253663484
	pesos_i(22352) := b"0000000000000000_0000000000000000_0010001011000111_0000111100110010"; -- 0.1358499048016572
	pesos_i(22353) := b"0000000000000000_0000000000000000_0000001011110000_0110100110111010"; -- 0.011480911066433465
	pesos_i(22354) := b"1111111111111111_1111111111111111_1111111001011100_1011000110111001"; -- -0.006398098253506908
	pesos_i(22355) := b"0000000000000000_0000000000000000_0001101001110001_1100110010001001"; -- 0.10329893429463491
	pesos_i(22356) := b"0000000000000000_0000000000000000_0010001011110110_0111011001100010"; -- 0.13657321817184145
	pesos_i(22357) := b"0000000000000000_0000000000000000_0001010001000110_1001110111010000"; -- 0.07920252167440472
	pesos_i(22358) := b"1111111111111111_1111111111111111_1110010001011010_1011100111110111"; -- -0.10799062463931779
	pesos_i(22359) := b"1111111111111111_1111111111111111_1110101110100100_1001001011100011"; -- -0.07952005338304322
	pesos_i(22360) := b"1111111111111111_1111111111111111_1101011111100100_0101101011110010"; -- -0.15667182530462218
	pesos_i(22361) := b"1111111111111111_1111111111111111_1110000011101101_1111011101101101"; -- -0.12136891920985518
	pesos_i(22362) := b"0000000000000000_0000000000000000_0010001101100000_1000000101110101"; -- 0.13819130993681725
	pesos_i(22363) := b"1111111111111111_1111111111111111_1101101001101001_0010011101101111"; -- -0.14683297678957366
	pesos_i(22364) := b"0000000000000000_0000000000000000_0000010011100010_1111100000111110"; -- 0.019088282676865805
	pesos_i(22365) := b"0000000000000000_0000000000000000_0001111011101100_1000101010100111"; -- 0.12079683843960044
	pesos_i(22366) := b"1111111111111111_1111111111111111_1111100001100010_0110101111011110"; -- -0.029748209312430277
	pesos_i(22367) := b"0000000000000000_0000000000000000_0000101101101111_0000001110110110"; -- 0.0446626967550289
	pesos_i(22368) := b"1111111111111111_1111111111111111_1111001110101110_0001100110111101"; -- -0.048124686597341676
	pesos_i(22369) := b"1111111111111111_1111111111111111_1110000110011111_0101011111110100"; -- -0.11866236002200116
	pesos_i(22370) := b"0000000000000000_0000000000000000_0010000101100111_0000100010010001"; -- 0.1304784157573999
	pesos_i(22371) := b"0000000000000000_0000000000000000_0000001110101100_0011101101010001"; -- 0.014346797310906392
	pesos_i(22372) := b"0000000000000000_0000000000000000_0000011100000011_0110010110111000"; -- 0.027395589228246194
	pesos_i(22373) := b"0000000000000000_0000000000000000_0001101101000100_1111000000010111"; -- 0.10652065808321066
	pesos_i(22374) := b"1111111111111111_1111111111111111_1110111111000011_0100010010111111"; -- -0.06342668852649806
	pesos_i(22375) := b"1111111111111111_1111111111111111_1111111001000011_1000111100001110"; -- -0.006781634442752037
	pesos_i(22376) := b"1111111111111111_1111111111111111_1110000001110011_1101111100011011"; -- -0.12323194102697102
	pesos_i(22377) := b"1111111111111111_1111111111111111_1111110101011011_1001001011101111"; -- -0.010321442318768427
	pesos_i(22378) := b"0000000000000000_0000000000000000_0000110010000111_1100110010110111"; -- 0.048947138515869675
	pesos_i(22379) := b"0000000000000000_0000000000000000_0010001101001001_0111011010000101"; -- 0.13783970597106723
	pesos_i(22380) := b"1111111111111111_1111111111111111_1111100001011101_0110111001110111"; -- -0.02982434846277192
	pesos_i(22381) := b"0000000000000000_0000000000000000_0010001000110111_1010000100010101"; -- 0.13366133460864163
	pesos_i(22382) := b"0000000000000000_0000000000000000_0000101001010011_0111000101100001"; -- 0.04033573734770022
	pesos_i(22383) := b"0000000000000000_0000000000000000_0010100100100110_0100011011011111"; -- 0.16074030816020413
	pesos_i(22384) := b"1111111111111111_1111111111111111_1111000011100000_1111010111001000"; -- -0.05906738151132354
	pesos_i(22385) := b"1111111111111111_1111111111111111_1111000000101010_0011101100111010"; -- -0.061855600567555416
	pesos_i(22386) := b"1111111111111111_1111111111111111_1111010100010011_0011000001100101"; -- -0.04267594844620824
	pesos_i(22387) := b"1111111111111111_1111111111111111_1110000001000101_1110110110100000"; -- -0.1239329799952499
	pesos_i(22388) := b"1111111111111111_1111111111111111_1110100011100010_0100010000000111"; -- -0.09029745890057679
	pesos_i(22389) := b"1111111111111111_1111111111111111_1101001111110111_0111111011010100"; -- -0.17200476960796673
	pesos_i(22390) := b"0000000000000000_0000000000000000_0000110110001010_1100101111101010"; -- 0.05289911713404514
	pesos_i(22391) := b"1111111111111111_1111111111111111_1111111100011000_1011110001110111"; -- -0.0035288055823386073
	pesos_i(22392) := b"1111111111111111_1111111111111111_1111001000110100_0010001000100000"; -- -0.05389200904594596
	pesos_i(22393) := b"0000000000000000_0000000000000000_0001010000111000_0110100111110011"; -- 0.07898580725897046
	pesos_i(22394) := b"0000000000000000_0000000000000000_0001001111100111_0111011111001110"; -- 0.07775067114951621
	pesos_i(22395) := b"1111111111111111_1111111111111111_1101011011100111_0100110000101011"; -- -0.160533179849051
	pesos_i(22396) := b"0000000000000000_0000000000000000_0001111101010100_1011011011100010"; -- 0.12238638892174941
	pesos_i(22397) := b"0000000000000000_0000000000000000_0001001110011001_1000101100110000"; -- 0.07656164090913486
	pesos_i(22398) := b"0000000000000000_0000000000000000_0010001000110101_0010111001110010"; -- 0.1336239842889376
	pesos_i(22399) := b"1111111111111111_1111111111111111_1101010110011111_0000111011001011"; -- -0.16554172091302075
	pesos_i(22400) := b"0000000000000000_0000000000000000_0010000001111010_0101111001110101"; -- 0.12686720227429038
	pesos_i(22401) := b"0000000000000000_0000000000000000_0010000101101111_0111111100000010"; -- 0.13060754589177656
	pesos_i(22402) := b"1111111111111111_1111111111111111_1101011101011010_1001010101001001"; -- -0.158774060945074
	pesos_i(22403) := b"1111111111111111_1111111111111111_1111110100000011_1000011011001001"; -- -0.011664939715546321
	pesos_i(22404) := b"1111111111111111_1111111111111111_1110100000001100_1010011101101110"; -- -0.09355691486249598
	pesos_i(22405) := b"1111111111111111_1111111111111111_1111111001110001_0010001101010000"; -- -0.006086152155575914
	pesos_i(22406) := b"0000000000000000_0000000000000000_0010010000010101_1111111001100011"; -- 0.14096059714683531
	pesos_i(22407) := b"1111111111111111_1111111111111111_1101100001111000_1110100001100010"; -- -0.15440509417983753
	pesos_i(22408) := b"1111111111111111_1111111111111111_1110001110110000_0001010001001010"; -- -0.1105944937449444
	pesos_i(22409) := b"1111111111111111_1111111111111111_1111011111000000_0101100111111000"; -- -0.03222119991777576
	pesos_i(22410) := b"0000000000000000_0000000000000000_0000010111010111_0000101011010111"; -- 0.022812535675459333
	pesos_i(22411) := b"1111111111111111_1111111111111111_1111111010001100_0010110101011000"; -- -0.005673566924926398
	pesos_i(22412) := b"0000000000000000_0000000000000000_0010001111111010_0100100000101001"; -- 0.14053774832269048
	pesos_i(22413) := b"0000000000000000_0000000000000000_0001110111001000_1000001000101010"; -- 0.11634076621711803
	pesos_i(22414) := b"0000000000000000_0000000000000000_0000100111000100_1000100111010110"; -- 0.03815518824270893
	pesos_i(22415) := b"1111111111111111_1111111111111111_1110111111010101_1100111111100010"; -- -0.06314373712015059
	pesos_i(22416) := b"1111111111111111_1111111111111111_1110001000001010_1010000100011111"; -- -0.1170253084616985
	pesos_i(22417) := b"0000000000000000_0000000000000000_0001011011001111_0111110000000100"; -- 0.08910346112896206
	pesos_i(22418) := b"0000000000000000_0000000000000000_0000000110111011_0100011000001110"; -- 0.006763819025691733
	pesos_i(22419) := b"0000000000000000_0000000000000000_0000010000100101_1100010011101011"; -- 0.01620131244543318
	pesos_i(22420) := b"1111111111111111_1111111111111111_1111110101000111_0100110010011101"; -- -0.010630809426252472
	pesos_i(22421) := b"1111111111111111_1111111111111111_1111101001110000_0100010111001111"; -- -0.021724354776959817
	pesos_i(22422) := b"0000000000000000_0000000000000000_0000011001111111_0011101011111011"; -- 0.025378881681272426
	pesos_i(22423) := b"1111111111111111_1111111111111111_1111101000010101_1010100010110001"; -- -0.023107010747055363
	pesos_i(22424) := b"1111111111111111_1111111111111111_1111111111101101_1100111101110101"; -- -0.0002775516133071991
	pesos_i(22425) := b"1111111111111111_1111111111111111_1101100001110001_1100111111100110"; -- -0.1545133650677907
	pesos_i(22426) := b"1111111111111111_1111111111111111_1110111011011101_1010110111010000"; -- -0.0669299475986137
	pesos_i(22427) := b"0000000000000000_0000000000000000_0001011100101100_0111111100010101"; -- 0.0905227114116867
	pesos_i(22428) := b"0000000000000000_0000000000000000_0001101001011000_0111011101010111"; -- 0.10291238653269827
	pesos_i(22429) := b"1111111111111111_1111111111111111_1111000110110010_0110000101010001"; -- -0.05587188510642121
	pesos_i(22430) := b"1111111111111111_1111111111111111_1101111101100010_0100100011110100"; -- -0.12740654033528642
	pesos_i(22431) := b"1111111111111111_1111111111111111_1110011010111000_0111001001100011"; -- -0.0987480647875187
	pesos_i(22432) := b"0000000000000000_0000000000000000_0000101000101001_0101000111010101"; -- 0.03969298799361419
	pesos_i(22433) := b"0000000000000000_0000000000000000_0000010010100100_0101100111010001"; -- 0.018132794885956594
	pesos_i(22434) := b"0000000000000000_0000000000000000_0001100000100101_0100001111000101"; -- 0.09431861467391064
	pesos_i(22435) := b"0000000000000000_0000000000000000_0001000110111110_1111010101100110"; -- 0.06932004680846636
	pesos_i(22436) := b"1111111111111111_1111111111111111_1110011000000101_1011101001110111"; -- -0.10147509194068673
	pesos_i(22437) := b"0000000000000000_0000000000000000_0000001101011111_1110010000001101"; -- 0.013181927928802814
	pesos_i(22438) := b"0000000000000000_0000000000000000_0000100000011110_0001111111001110"; -- 0.03170965945959514
	pesos_i(22439) := b"1111111111111111_1111111111111111_1111111110101001_1000100011110011"; -- -0.0013193517594583025
	pesos_i(22440) := b"1111111111111111_1111111111111111_1111110000100101_0000011001010100"; -- -0.01506004754461394
	pesos_i(22441) := b"1111111111111111_1111111111111111_1101101111010000_1110101100110000"; -- -0.14134340351537986
	pesos_i(22442) := b"1111111111111111_1111111111111111_1111001001111011_0011010110100100"; -- -0.052807471818935525
	pesos_i(22443) := b"0000000000000000_0000000000000000_0010000111100101_0011101001001011"; -- 0.13240398711925583
	pesos_i(22444) := b"1111111111111111_1111111111111111_1111000000011101_0010000000111110"; -- -0.06205557325758182
	pesos_i(22445) := b"1111111111111111_1111111111111111_1110011000100111_1010100100011101"; -- -0.10095732738530627
	pesos_i(22446) := b"1111111111111111_1111111111111111_1110010011001111_0111111100111111"; -- -0.10620884631612888
	pesos_i(22447) := b"0000000000000000_0000000000000000_0001101101101001_1101010101100011"; -- 0.10708364178781245
	pesos_i(22448) := b"0000000000000000_0000000000000000_0001110101001101_0110101010010000"; -- 0.11446252844882869
	pesos_i(22449) := b"0000000000000000_0000000000000000_0000101001000001_0111001011111010"; -- 0.04006117444105752
	pesos_i(22450) := b"0000000000000000_0000000000000000_0000000100001000_1011111000101010"; -- 0.004039655071519179
	pesos_i(22451) := b"1111111111111111_1111111111111111_1111101111000010_1011100101110000"; -- -0.01655999190889951
	pesos_i(22452) := b"0000000000000000_0000000000000000_0010011101000001_0100001001001111"; -- 0.15333952348599703
	pesos_i(22453) := b"1111111111111111_1111111111111111_1110011101011100_1111111110000111"; -- -0.09623721075486188
	pesos_i(22454) := b"1111111111111111_1111111111111111_1110000101010001_0000101010100000"; -- -0.11985715476824964
	pesos_i(22455) := b"0000000000000000_0000000000000000_0001100010011111_0111101111001111"; -- 0.09618352707974438
	pesos_i(22456) := b"0000000000000000_0000000000000000_0000101111000001_0101111100000110"; -- 0.04591936003334796
	pesos_i(22457) := b"0000000000000000_0000000000000000_0000011100000100_0110000100111011"; -- 0.027410580536857198
	pesos_i(22458) := b"1111111111111111_1111111111111111_1111001010111000_1101010101110001"; -- -0.051867160603564305
	pesos_i(22459) := b"0000000000000000_0000000000000000_0001101101000000_1111010000111110"; -- 0.10645987036555225
	pesos_i(22460) := b"0000000000000000_0000000000000000_0010000001111111_1100010001000011"; -- 0.12694956439438285
	pesos_i(22461) := b"1111111111111111_1111111111111111_1111000000010010_0001001000011011"; -- -0.06222426268946392
	pesos_i(22462) := b"1111111111111111_1111111111111111_1111100000111110_1010100100111101"; -- -0.030293867611066297
	pesos_i(22463) := b"0000000000000000_0000000000000000_0000100000100101_1111011100011010"; -- 0.031829303492158297
	pesos_i(22464) := b"0000000000000000_0000000000000000_0000000101001100_1100010010101010"; -- 0.005077639947397377
	pesos_i(22465) := b"0000000000000000_0000000000000000_0010000110001011_0011100001000111"; -- 0.13103057608395421
	pesos_i(22466) := b"1111111111111111_1111111111111111_1111011001101100_1001011010011000"; -- -0.03740557475746056
	pesos_i(22467) := b"1111111111111111_1111111111111111_1110101101110100_1101001100011100"; -- -0.08024864738616604
	pesos_i(22468) := b"0000000000000000_0000000000000000_0000110101010110_1101111000111001"; -- 0.05210675129597627
	pesos_i(22469) := b"0000000000000000_0000000000000000_0000000110100100_0001000011011000"; -- 0.00640969528837689
	pesos_i(22470) := b"0000000000000000_0000000000000000_0001110010110011_0100010011110110"; -- 0.11211043367117969
	pesos_i(22471) := b"0000000000000000_0000000000000000_0000101101110010_1001010000001100"; -- 0.04471707623904956
	pesos_i(22472) := b"1111111111111111_1111111111111111_1111011010000100_0111001000100000"; -- -0.03704153753236203
	pesos_i(22473) := b"0000000000000000_0000000000000000_0001001010111010_0111001101110000"; -- 0.07315751544228413
	pesos_i(22474) := b"0000000000000000_0000000000000000_0010000100100111_1001001110001111"; -- 0.12951013795680044
	pesos_i(22475) := b"1111111111111111_1111111111111111_1110100111101101_0111101111110101"; -- -0.0862200284737198
	pesos_i(22476) := b"0000000000000000_0000000000000000_0010001010110111_0111010001101110"; -- 0.13561179824833833
	pesos_i(22477) := b"0000000000000000_0000000000000000_0000010111010000_1101011101110001"; -- 0.022717919528983676
	pesos_i(22478) := b"1111111111111111_1111111111111111_1110110000000001_0100101011000001"; -- -0.07810528545062619
	pesos_i(22479) := b"1111111111111111_1111111111111111_1111000101110000_1011110000000010"; -- -0.056873559588508586
	pesos_i(22480) := b"0000000000000000_0000000000000000_0010101001111101_1000101110000000"; -- 0.16597816353983544
	pesos_i(22481) := b"1111111111111111_1111111111111111_1111101001101001_0110100010001010"; -- -0.02182909613161674
	pesos_i(22482) := b"0000000000000000_0000000000000000_0001010001110001_0010110001000010"; -- 0.07985188102479707
	pesos_i(22483) := b"1111111111111111_1111111111111111_1111001000010111_0100111011100001"; -- -0.05433184622257621
	pesos_i(22484) := b"1111111111111111_1111111111111111_1110100101101100_1110000111011110"; -- -0.0881823380229071
	pesos_i(22485) := b"0000000000000000_0000000000000000_0001010011110111_0001001101010110"; -- 0.08189507352278567
	pesos_i(22486) := b"0000000000000000_0000000000000000_0000011010100010_0110101010111010"; -- 0.025915785127584173
	pesos_i(22487) := b"1111111111111111_1111111111111111_1111010110011010_0101000000010011"; -- -0.040614123696024726
	pesos_i(22488) := b"1111111111111111_1111111111111111_1111011011100111_1011110110001001"; -- -0.03552642246753161
	pesos_i(22489) := b"1111111111111111_1111111111111111_1110110110011100_1011110101011101"; -- -0.07182709187473209
	pesos_i(22490) := b"1111111111111111_1111111111111111_1101111010110011_0001001010010110"; -- -0.13008006891478507
	pesos_i(22491) := b"0000000000000000_0000000000000000_0000101100100011_1101000000100001"; -- 0.04351521304066346
	pesos_i(22492) := b"1111111111111111_1111111111111111_1110101011110011_0011001110101111"; -- -0.08222653358014388
	pesos_i(22493) := b"0000000000000000_0000000000000000_0001111011001010_0001100000000011"; -- 0.12027120649149545
	pesos_i(22494) := b"1111111111111111_1111111111111111_1110100001011010_1001010011101001"; -- -0.09236783335807015
	pesos_i(22495) := b"0000000000000000_0000000000000000_0001010101110110_0011010010100110"; -- 0.08383492526034048
	pesos_i(22496) := b"0000000000000000_0000000000000000_0000010100001110_1110000011100110"; -- 0.0197582779599872
	pesos_i(22497) := b"1111111111111111_1111111111111111_1110010110011110_0111101011011101"; -- -0.10305053813287429
	pesos_i(22498) := b"1111111111111111_1111111111111111_1110011000000010_0010000100000111"; -- -0.1015300138250597
	pesos_i(22499) := b"1111111111111111_1111111111111111_1110111011100001_0010001010011010"; -- -0.06687721000222567
	pesos_i(22500) := b"0000000000000000_0000000000000000_0010001110011101_0000011111000101"; -- 0.13911484292227194
	pesos_i(22501) := b"1111111111111111_1111111111111111_1111001011010110_1001000110001101"; -- -0.05141344374105169
	pesos_i(22502) := b"0000000000000000_0000000000000000_0000000001001101_1101110101111101"; -- 0.0011881284002985492
	pesos_i(22503) := b"0000000000000000_0000000000000000_0001000001001100_1011101001100100"; -- 0.0636707776179959
	pesos_i(22504) := b"1111111111111111_1111111111111111_1101111011011110_0000100101000111"; -- -0.12942449595221747
	pesos_i(22505) := b"0000000000000000_0000000000000000_0001000000111110_0011101101000111"; -- 0.0634495780397852
	pesos_i(22506) := b"0000000000000000_0000000000000000_0010001010011110_1101000101110101"; -- 0.13523587330773829
	pesos_i(22507) := b"1111111111111111_1111111111111111_1111011010000001_0011101001110010"; -- -0.037090632605014245
	pesos_i(22508) := b"1111111111111111_1111111111111111_1110100001010010_0000111000011110"; -- -0.09249793783293905
	pesos_i(22509) := b"1111111111111111_1111111111111111_1110101001101010_1110011011111111"; -- -0.0843062999491694
	pesos_i(22510) := b"1111111111111111_1111111111111111_1111001001101110_0100110111000110"; -- -0.053004397596218056
	pesos_i(22511) := b"1111111111111111_1111111111111111_1101011001111001_0100111100010010"; -- -0.1622114736642157
	pesos_i(22512) := b"0000000000000000_0000000000000000_0001000010001001_0000110110000011"; -- 0.0645912594137134
	pesos_i(22513) := b"0000000000000000_0000000000000000_0001110100110111_1110000111100101"; -- 0.11413394769930091
	pesos_i(22514) := b"0000000000000000_0000000000000000_0001000001101000_0101111001101000"; -- 0.06409254100483104
	pesos_i(22515) := b"1111111111111111_1111111111111111_1110010101000010_1000111001010011"; -- -0.10445318680636612
	pesos_i(22516) := b"0000000000000000_0000000000000000_0001000001111001_1100100010111000"; -- 0.06435827720139631
	pesos_i(22517) := b"1111111111111111_1111111111111111_1111111001000011_1111110111011110"; -- -0.006775029426845187
	pesos_i(22518) := b"0000000000000000_0000000000000000_0001000101111010_1011101010010100"; -- 0.06827894329480697
	pesos_i(22519) := b"1111111111111111_1111111111111111_1110110111010000_1001010110010111"; -- -0.0710360056965741
	pesos_i(22520) := b"1111111111111111_1111111111111111_1110100110001001_0001100001110100"; -- -0.0877518384941867
	pesos_i(22521) := b"0000000000000000_0000000000000000_0000011000010010_1101000110001111"; -- 0.023724648894015123
	pesos_i(22522) := b"1111111111111111_1111111111111111_1111101001010000_1011001111111011"; -- -0.022206069161620788
	pesos_i(22523) := b"1111111111111111_1111111111111111_1111000110011000_0001011110001011"; -- -0.05627301068880973
	pesos_i(22524) := b"1111111111111111_1111111111111111_1110001110010000_0010011001111101"; -- -0.11108169031432619
	pesos_i(22525) := b"1111111111111111_1111111111111111_1110101010011010_1110000011110000"; -- -0.08357423912510073
	pesos_i(22526) := b"0000000000000000_0000000000000000_0010001100001000_1101100000011000"; -- 0.13685370041262188
	pesos_i(22527) := b"1111111111111111_1111111111111111_1111011000111100_0111011111101111"; -- -0.03813982415765174
	pesos_i(22528) := b"0000000000000000_0000000000000000_0001111101100100_0001000001000000"; -- 0.12262059749568366
	pesos_i(22529) := b"0000000000000000_0000000000000000_0000011010000111_0001111011010100"; -- 0.025499274046770777
	pesos_i(22530) := b"0000000000000000_0000000000000000_0001110111101101_0100100110000010"; -- 0.11690196449994678
	pesos_i(22531) := b"1111111111111111_1111111111111111_1111100000000101_0101101001101111"; -- -0.031168315844007064
	pesos_i(22532) := b"1111111111111111_1111111111111111_1110010111000111_0011100111111001"; -- -0.10242879564210196
	pesos_i(22533) := b"1111111111111111_1111111111111111_1110101001010001_1111100000010000"; -- -0.08468675235904548
	pesos_i(22534) := b"1111111111111111_1111111111111111_1110000000000010_1010100110100110"; -- -0.12495937064568967
	pesos_i(22535) := b"1111111111111111_1111111111111111_1110111100010110_1000010000100010"; -- -0.06606268083854304
	pesos_i(22536) := b"0000000000000000_0000000000000000_0010001010000011_1110000100111111"; -- 0.13482482706812185
	pesos_i(22537) := b"0000000000000000_0000000000000000_0001111001011001_1101000011011111"; -- 0.11855798194900635
	pesos_i(22538) := b"1111111111111111_1111111111111111_1110111000010101_1001101011111010"; -- -0.06998282808881835
	pesos_i(22539) := b"0000000000000000_0000000000000000_0000000101111001_0000011010111001"; -- 0.005752964250996089
	pesos_i(22540) := b"1111111111111111_1111111111111111_1111110001101100_1111010011011101"; -- -0.01396245580941462
	pesos_i(22541) := b"1111111111111111_1111111111111111_1110100111100100_0001101011100001"; -- -0.08636314393754856
	pesos_i(22542) := b"1111111111111111_1111111111111111_1111001111111110_0010100101011010"; -- -0.0469030528919858
	pesos_i(22543) := b"0000000000000000_0000000000000000_0000111110000100_1001010101011101"; -- 0.060616812841097954
	pesos_i(22544) := b"1111111111111111_1111111111111111_1110011000001101_0011111001011000"; -- -0.10136041975298404
	pesos_i(22545) := b"1111111111111111_1111111111111111_1110101001001000_0011101010100000"; -- -0.08483537289068811
	pesos_i(22546) := b"0000000000000000_0000000000000000_0010101001011011_1000000010000101"; -- 0.1654587101703559
	pesos_i(22547) := b"0000000000000000_0000000000000000_0010001110100111_1010110000001110"; -- 0.13927722312678004
	pesos_i(22548) := b"1111111111111111_1111111111111111_1111100111010111_0011000000010011"; -- -0.02406024480663104
	pesos_i(22549) := b"1111111111111111_1111111111111111_1110000010101110_0100101000101101"; -- -0.12234054942640624
	pesos_i(22550) := b"1111111111111111_1111111111111111_1110111000010110_1111011111010111"; -- -0.06996203419073159
	pesos_i(22551) := b"1111111111111111_1111111111111111_1111010101010101_1101100110000010"; -- -0.04165878844233067
	pesos_i(22552) := b"1111111111111111_1111111111111111_1111010101101000_1001001111110100"; -- -0.041373017199472076
	pesos_i(22553) := b"0000000000000000_0000000000000000_0001001100000001_1111101100010101"; -- 0.07424897443436769
	pesos_i(22554) := b"1111111111111111_1111111111111111_1110111001001111_0000001101101110"; -- -0.06910685121654393
	pesos_i(22555) := b"0000000000000000_0000000000000000_0001111101001000_0100001100111000"; -- 0.12219638927528936
	pesos_i(22556) := b"1111111111111111_1111111111111111_1111000011100011_0101110000111001"; -- -0.05903075796195987
	pesos_i(22557) := b"0000000000000000_0000000000000000_0001000011010110_0001011100010111"; -- 0.06576675705551473
	pesos_i(22558) := b"0000000000000000_0000000000000000_0000101011101110_1101110011101101"; -- 0.04270725994369202
	pesos_i(22559) := b"1111111111111111_1111111111111111_1111110011111011_0011111110010101"; -- -0.011791254207715348
	pesos_i(22560) := b"0000000000000000_0000000000000000_0010010000101100_0010000011011111"; -- 0.14129834602116706
	pesos_i(22561) := b"0000000000000000_0000000000000000_0000111001000011_1011001111011100"; -- 0.055720559307383066
	pesos_i(22562) := b"0000000000000000_0000000000000000_0000000011000110_0111001100010011"; -- 0.003028099195215666
	pesos_i(22563) := b"0000000000000000_0000000000000000_0010010000100110_0110000010100010"; -- 0.14121059384085025
	pesos_i(22564) := b"1111111111111111_1111111111111111_1111000000100010_0010001101011101"; -- -0.0619790934094532
	pesos_i(22565) := b"1111111111111111_1111111111111111_1111111101010001_0110100010000111"; -- -0.0026640577179403505
	pesos_i(22566) := b"1111111111111111_1111111111111111_1110110001101001_0011111111110011"; -- -0.07651901536462126
	pesos_i(22567) := b"0000000000000000_0000000000000000_0001011010011101_0100001000010011"; -- 0.0883370681993864
	pesos_i(22568) := b"1111111111111111_1111111111111111_1111100110001011_1111000011010101"; -- -0.025208423584556394
	pesos_i(22569) := b"0000000000000000_0000000000000000_0000011000010001_0001111001111001"; -- 0.02369871566317935
	pesos_i(22570) := b"1111111111111111_1111111111111111_1110110011010001_0011010011110100"; -- -0.07493275691958018
	pesos_i(22571) := b"0000000000000000_0000000000000000_0001110010111000_1011010000110010"; -- 0.11219335772827738
	pesos_i(22572) := b"1111111111111111_1111111111111111_1110001001101010_1001110100001000"; -- -0.11556070861042224
	pesos_i(22573) := b"1111111111111111_1111111111111111_1110000011110001_1000101100010111"; -- -0.12131434146270666
	pesos_i(22574) := b"1111111111111111_1111111111111111_1110100010000001_0100000110011110"; -- -0.09177770515507115
	pesos_i(22575) := b"1111111111111111_1111111111111111_1110100000101101_0010000110001001"; -- -0.09306135561068242
	pesos_i(22576) := b"0000000000000000_0000000000000000_0000001001111001_1001111001110001"; -- 0.009668257399139596
	pesos_i(22577) := b"0000000000000000_0000000000000000_0010000111101101_0001001100100111"; -- 0.13252372462846349
	pesos_i(22578) := b"0000000000000000_0000000000000000_0000110110000100_1100101011111101"; -- 0.05280750930466853
	pesos_i(22579) := b"1111111111111111_1111111111111111_1110100011111100_0011001111111110"; -- -0.08990168623786099
	pesos_i(22580) := b"1111111111111111_1111111111111111_1111011100100111_0110011101011111"; -- -0.03455499580497551
	pesos_i(22581) := b"1111111111111111_1111111111111111_1111011110111010_0100010100100100"; -- -0.03231399417373415
	pesos_i(22582) := b"1111111111111111_1111111111111111_1111111000010000_1100010001101000"; -- -0.007556652719859574
	pesos_i(22583) := b"0000000000000000_0000000000000000_0001001100100010_1100000001011111"; -- 0.07474901500723646
	pesos_i(22584) := b"0000000000000000_0000000000000000_0000011000010000_1110110110111001"; -- 0.023695810012249845
	pesos_i(22585) := b"0000000000000000_0000000000000000_0001010101101011_0011011100010000"; -- 0.08366722235912326
	pesos_i(22586) := b"1111111111111111_1111111111111111_1110110011101011_0100000101010110"; -- -0.0745352903086884
	pesos_i(22587) := b"0000000000000000_0000000000000000_0010000010101001_1010111110000100"; -- 0.1275891970006071
	pesos_i(22588) := b"0000000000000000_0000000000000000_0001001101000101_0011011110000011"; -- 0.07527491514397618
	pesos_i(22589) := b"1111111111111111_1111111111111111_1111110010101010_1110011100010110"; -- -0.0130172319952021
	pesos_i(22590) := b"0000000000000000_0000000000000000_0000010001011110_1010101011100110"; -- 0.01706951253772098
	pesos_i(22591) := b"1111111111111111_1111111111111111_1101111111011010_0110011000101101"; -- -0.12557374377828634
	pesos_i(22592) := b"1111111111111111_1111111111111111_1110010010101101_0111001111000000"; -- -0.10672833014241735
	pesos_i(22593) := b"1111111111111111_1111111111111111_1101111001110010_0110011010010111"; -- -0.13106688322255938
	pesos_i(22594) := b"1111111111111111_1111111111111111_1111101110100000_0001111000110000"; -- -0.017088044348393918
	pesos_i(22595) := b"1111111111111111_1111111111111111_1101111110010010_0111001100000100"; -- -0.1266716114396015
	pesos_i(22596) := b"0000000000000000_0000000000000000_0000001111000000_0111011000000011"; -- 0.01465547158780449
	pesos_i(22597) := b"0000000000000000_0000000000000000_0010001111101100_1010110011110111"; -- 0.14033013383028037
	pesos_i(22598) := b"1111111111111111_1111111111111111_1101111001101100_0010101000100100"; -- -0.13116203906058194
	pesos_i(22599) := b"1111111111111111_1111111111111111_1111110010111110_1110000001101100"; -- -0.01271245343625808
	pesos_i(22600) := b"0000000000000000_0000000000000000_0010000101011000_0111000000001100"; -- 0.13025570202852815
	pesos_i(22601) := b"1111111111111111_1111111111111111_1111001000111010_1000110000000100"; -- -0.05379414458153266
	pesos_i(22602) := b"0000000000000000_0000000000000000_0001000101010001_0110011001001101"; -- 0.0676483096025219
	pesos_i(22603) := b"1111111111111111_1111111111111111_1110010100101101_0100001100100111"; -- -0.10477810179249368
	pesos_i(22604) := b"1111111111111111_1111111111111111_1110110010000110_0111010101000011"; -- -0.07607333283716314
	pesos_i(22605) := b"0000000000000000_0000000000000000_0010100000100001_0100000100101010"; -- 0.15675742407795834
	pesos_i(22606) := b"1111111111111111_1111111111111111_1101110110000101_1100010001101000"; -- -0.1346776243174185
	pesos_i(22607) := b"0000000000000000_0000000000000000_0001110010110000_0101011101001011"; -- 0.11206574997026432
	pesos_i(22608) := b"0000000000000000_0000000000000000_0001011011110001_1110011011101100"; -- 0.08962863224580674
	pesos_i(22609) := b"1111111111111111_1111111111111111_1111110010110011_0000101000001010"; -- -0.012893078295432297
	pesos_i(22610) := b"1111111111111111_1111111111111111_1110000000000100_1101010001011011"; -- -0.12492630744469028
	pesos_i(22611) := b"1111111111111111_1111111111111111_1111101110011011_0010111001011011"; -- -0.01716337477054144
	pesos_i(22612) := b"1111111111111111_1111111111111111_1110101111111100_1101100001000011"; -- -0.0781731449471583
	pesos_i(22613) := b"1111111111111111_1111111111111111_1111110110101101_1110010111010110"; -- -0.009065280296661227
	pesos_i(22614) := b"0000000000000000_0000000000000000_0010011000100101_1001101101110010"; -- 0.14901134039160793
	pesos_i(22615) := b"0000000000000000_0000000000000000_0010010000000111_1110001010000010"; -- 0.14074531235402157
	pesos_i(22616) := b"0000000000000000_0000000000000000_0000111000001010_0001100011010000"; -- 0.05484156680752012
	pesos_i(22617) := b"1111111111111111_1111111111111111_1110011111011111_0001110101101111"; -- -0.09425178564798184
	pesos_i(22618) := b"1111111111111111_1111111111111111_1111111001001110_1001001000011010"; -- -0.006613606096631202
	pesos_i(22619) := b"0000000000000000_0000000000000000_0010000000001001_0010001101000011"; -- 0.12513943077753986
	pesos_i(22620) := b"1111111111111111_1111111111111111_1110110011010001_0110010101000100"; -- -0.07492987723011624
	pesos_i(22621) := b"1111111111111111_1111111111111111_1111111001111111_1101101000101010"; -- -0.005861630131299761
	pesos_i(22622) := b"1111111111111111_1111111111111111_1110010010100001_1101011000011011"; -- -0.1069055732876622
	pesos_i(22623) := b"1111111111111111_1111111111111111_1111110100100000_1100111011100011"; -- -0.011218137383030947
	pesos_i(22624) := b"0000000000000000_0000000000000000_0000000001000101_1101100000111110"; -- 0.0010657454377852905
	pesos_i(22625) := b"1111111111111111_1111111111111111_1111111100101000_1101110111000001"; -- -0.0032826808225427024
	pesos_i(22626) := b"0000000000000000_0000000000000000_0000000110011010_1100100011101000"; -- 0.006268078554501042
	pesos_i(22627) := b"0000000000000000_0000000000000000_0010010111011111_0100001010111110"; -- 0.1479379380856238
	pesos_i(22628) := b"1111111111111111_1111111111111111_1110001011111101_1000100100000111"; -- -0.1133188590120027
	pesos_i(22629) := b"1111111111111111_1111111111111111_1110010101101011_0001001101011101"; -- -0.10383490534674292
	pesos_i(22630) := b"1111111111111111_1111111111111111_1110000101010110_1110111000110111"; -- -0.11976729552380692
	pesos_i(22631) := b"1111111111111111_1111111111111111_1111101111100010_0001101101101110"; -- -0.016081128672766853
	pesos_i(22632) := b"1111111111111111_1111111111111111_1110111111110101_0001101101011011"; -- -0.06266621608076238
	pesos_i(22633) := b"0000000000000000_0000000000000000_0010000110000000_0101001101010100"; -- 0.1308643418576672
	pesos_i(22634) := b"1111111111111111_1111111111111111_1110001010101000_1110100101101101"; -- -0.11461011023384102
	pesos_i(22635) := b"1111111111111111_1111111111111111_1101100011000101_0100100110110100"; -- -0.1532396255893782
	pesos_i(22636) := b"0000000000000000_0000000000000000_0001011010110010_0100001101000001"; -- 0.08865757302102813
	pesos_i(22637) := b"0000000000000000_0000000000000000_0000111011001110_1101011010111011"; -- 0.057843609496199516
	pesos_i(22638) := b"1111111111111111_1111111111111111_1110001001000010_0000001011111001"; -- -0.11618024279662785
	pesos_i(22639) := b"0000000000000000_0000000000000000_0001100111010000_0010111111110000"; -- 0.10083293534960536
	pesos_i(22640) := b"1111111111111111_1111111111111111_1110111011101000_0010010011111110"; -- -0.06677025598208057
	pesos_i(22641) := b"1111111111111111_1111111111111111_1111010100101110_0111100001101000"; -- -0.04225966881575879
	pesos_i(22642) := b"0000000000000000_0000000000000000_0000010111110111_0000110101001111"; -- 0.023300964082890636
	pesos_i(22643) := b"0000000000000000_0000000000000000_0000101110110001_0111010101010011"; -- 0.04567654862769573
	pesos_i(22644) := b"1111111111111111_1111111111111111_1111000001100011_0011010001011110"; -- -0.06098625858856166
	pesos_i(22645) := b"0000000000000000_0000000000000000_0001000100101100_1011001001010000"; -- 0.06708826497081334
	pesos_i(22646) := b"1111111111111111_1111111111111111_1110011001100001_0001001111001001"; -- -0.10008121809689717
	pesos_i(22647) := b"0000000000000000_0000000000000000_0000101100010001_1110111001011011"; -- 0.043242356510423484
	pesos_i(22648) := b"1111111111111111_1111111111111111_1101101001010100_1001101101000011"; -- -0.14714650746454455
	pesos_i(22649) := b"1111111111111111_1111111111111111_1101110101100011_0101001101100100"; -- -0.13520315935118052
	pesos_i(22650) := b"0000000000000000_0000000000000000_0000011001001110_0101100111111010"; -- 0.02463304846381933
	pesos_i(22651) := b"1111111111111111_1111111111111111_1110001000111000_1100100011000100"; -- -0.1163210411780299
	pesos_i(22652) := b"0000000000000000_0000000000000000_0000110111111100_0100010011000110"; -- 0.054630564159103605
	pesos_i(22653) := b"0000000000000000_0000000000000000_0010010101010110_0001101100001111"; -- 0.1458451187523098
	pesos_i(22654) := b"0000000000000000_0000000000000000_0001101010101000_1000100100111001"; -- 0.10413415556704105
	pesos_i(22655) := b"0000000000000000_0000000000000000_0001010000111001_1100100111000001"; -- 0.07900677642654803
	pesos_i(22656) := b"1111111111111111_1111111111111111_1110101110100011_0010011110110110"; -- -0.07954170031992577
	pesos_i(22657) := b"1111111111111111_1111111111111111_1111111100111110_1000001010001010"; -- -0.002952424233491056
	pesos_i(22658) := b"1111111111111111_1111111111111111_1111101001001100_1100110000100101"; -- -0.022265664095421966
	pesos_i(22659) := b"1111111111111111_1111111111111111_1101111001111010_1001111100111001"; -- -0.13094143724217325
	pesos_i(22660) := b"0000000000000000_0000000000000000_0001011101001001_1001001011110011"; -- 0.09096640047882955
	pesos_i(22661) := b"0000000000000000_0000000000000000_0001110010000000_0101010110011110"; -- 0.11133322806871018
	pesos_i(22662) := b"0000000000000000_0000000000000000_0010000101010100_0101100100100000"; -- 0.13019330047650857
	pesos_i(22663) := b"0000000000000000_0000000000000000_0000011000011101_0100011111100010"; -- 0.02388428950043754
	pesos_i(22664) := b"1111111111111111_1111111111111111_1111011110001000_0101111010100010"; -- -0.03307541412451247
	pesos_i(22665) := b"0000000000000000_0000000000000000_0010000000101110_0001101010100100"; -- 0.12570349210561665
	pesos_i(22666) := b"1111111111111111_1111111111111111_1111000101000010_0011001011100000"; -- -0.05758363752797553
	pesos_i(22667) := b"1111111111111111_1111111111111111_1110110111010100_0010011101111010"; -- -0.07098153375287287
	pesos_i(22668) := b"1111111111111111_1111111111111111_1111000001111100_1001100000010010"; -- -0.0605988460364946
	pesos_i(22669) := b"0000000000000000_0000000000000000_0000000111010010_1111010111000111"; -- 0.007125245129587455
	pesos_i(22670) := b"1111111111111111_1111111111111111_1111000111011011_1110100010000100"; -- -0.05523821625909124
	pesos_i(22671) := b"1111111111111111_1111111111111111_1111000000001100_1100011111001000"; -- -0.06230498663390219
	pesos_i(22672) := b"1111111111111111_1111111111111111_1111000101010010_0101011010100100"; -- -0.05733736513277515
	pesos_i(22673) := b"0000000000000000_0000000000000000_0010010110000011_1001111111011000"; -- 0.14653967890410585
	pesos_i(22674) := b"1111111111111111_1111111111111111_1110011110011100_1100011000101000"; -- -0.09526406787362682
	pesos_i(22675) := b"0000000000000000_0000000000000000_0001011111000110_1101100100001111"; -- 0.09287792790982502
	pesos_i(22676) := b"1111111111111111_1111111111111111_1110011000011100_0011000011101000"; -- -0.10113233879951887
	pesos_i(22677) := b"1111111111111111_1111111111111111_1110100000100001_1000000001011011"; -- -0.09323880941232493
	pesos_i(22678) := b"0000000000000000_0000000000000000_0001011111111110_0001110010001110"; -- 0.09372118448008994
	pesos_i(22679) := b"0000000000000000_0000000000000000_0000000110000001_1111011110100011"; -- 0.005889394070296154
	pesos_i(22680) := b"1111111111111111_1111111111111111_1111110101000011_0011111010010100"; -- -0.01069268110238679
	pesos_i(22681) := b"0000000000000000_0000000000000000_0010010000001100_0011001001101101"; -- 0.1408111111863405
	pesos_i(22682) := b"1111111111111111_1111111111111111_1111010100110011_1110001010100111"; -- -0.042177042226978226
	pesos_i(22683) := b"0000000000000000_0000000000000000_0001000101011001_1010100101010100"; -- 0.0677743748783063
	pesos_i(22684) := b"0000000000000000_0000000000000000_0010000000010110_1010011001010101"; -- 0.12534560754221685
	pesos_i(22685) := b"1111111111111111_1111111111111111_1110110010011001_1110000010001010"; -- -0.07577702166643711
	pesos_i(22686) := b"0000000000000000_0000000000000000_0010000000001110_1000110100010100"; -- 0.1252220319030741
	pesos_i(22687) := b"0000000000000000_0000000000000000_0001111111100111_1111111111000111"; -- 0.12463377584232621
	pesos_i(22688) := b"0000000000000000_0000000000000000_0000111111111001_1000011101010101"; -- 0.0624012550012945
	pesos_i(22689) := b"1111111111111111_1111111111111111_1110011010000010_1001011001101111"; -- -0.09956989080145855
	pesos_i(22690) := b"0000000000000000_0000000000000000_0010001111101011_0001111001111010"; -- 0.14030638201470594
	pesos_i(22691) := b"1111111111111111_1111111111111111_1111110100111001_1100001101110101"; -- -0.010837348962423603
	pesos_i(22692) := b"1111111111111111_1111111111111111_1101111011100011_0111000110000001"; -- -0.1293419895793731
	pesos_i(22693) := b"1111111111111111_1111111111111111_1111001011110101_1001100110000000"; -- -0.05093994741423366
	pesos_i(22694) := b"0000000000000000_0000000000000000_0010000000010111_0000100101011111"; -- 0.12535151072684755
	pesos_i(22695) := b"1111111111111111_1111111111111111_1110011110101011_0110010011010111"; -- -0.09504098647957876
	pesos_i(22696) := b"1111111111111111_1111111111111111_1110110010000110_0111000011110001"; -- -0.07607359040095293
	pesos_i(22697) := b"1111111111111111_1111111111111111_1110011001101101_1110001000011101"; -- -0.09988581464841104
	pesos_i(22698) := b"0000000000000000_0000000000000000_0010001011000100_1101111000000000"; -- 0.13581645479088275
	pesos_i(22699) := b"1111111111111111_1111111111111111_1110010101101110_1101010001110111"; -- -0.1037776193116822
	pesos_i(22700) := b"0000000000000000_0000000000000000_0000010111011111_1001100011111101"; -- 0.022943078882862615
	pesos_i(22701) := b"1111111111111111_1111111111111111_1111011001010000_1001000001001100"; -- -0.037833196076086664
	pesos_i(22702) := b"1111111111111111_1111111111111111_1111010000101111_1010101101100001"; -- -0.04614762185376346
	pesos_i(22703) := b"1111111111111111_1111111111111111_1101101010100001_0001101010110111"; -- -0.14597924268922513
	pesos_i(22704) := b"0000000000000000_0000000000000000_0000000001011100_0100000110111001"; -- 0.0014077259829325033
	pesos_i(22705) := b"0000000000000000_0000000000000000_0000011110110001_0101101110000111"; -- 0.030050011031774435
	pesos_i(22706) := b"1111111111111111_1111111111111111_1111111100001001_1011000110100100"; -- -0.0037583327894350174
	pesos_i(22707) := b"1111111111111111_1111111111111111_1110110110110100_0111000010101111"; -- -0.07146545143663263
	pesos_i(22708) := b"1111111111111111_1111111111111111_1111000011110010_0011110010010111"; -- -0.05880376152211324
	pesos_i(22709) := b"0000000000000000_0000000000000000_0001011111010111_0010100111100011"; -- 0.09312688629581829
	pesos_i(22710) := b"1111111111111111_1111111111111111_1101110100010111_1100111111110001"; -- -0.136355403640334
	pesos_i(22711) := b"0000000000000000_0000000000000000_0000011001010101_1110101100111100"; -- 0.024748518047543792
	pesos_i(22712) := b"1111111111111111_1111111111111111_1110000100100100_1111000001101001"; -- -0.12053010407563838
	pesos_i(22713) := b"1111111111111111_1111111111111111_1111001010110000_0111101100011110"; -- -0.05199461481419511
	pesos_i(22714) := b"1111111111111111_1111111111111111_1110100001111101_0010000010110000"; -- -0.09184070300026824
	pesos_i(22715) := b"1111111111111111_1111111111111111_1101100001111110_0001000011111011"; -- -0.15432638049542496
	pesos_i(22716) := b"0000000000000000_0000000000000000_0010001101001111_0011001001101001"; -- 0.13792719898531308
	pesos_i(22717) := b"0000000000000000_0000000000000000_0000111001110110_1011011100001011"; -- 0.05649894739849403
	pesos_i(22718) := b"1111111111111111_1111111111111111_1110101100010110_0100110100100010"; -- -0.08169095908466749
	pesos_i(22719) := b"0000000000000000_0000000000000000_0000010001111100_0011110001100000"; -- 0.017520688469069113
	pesos_i(22720) := b"1111111111111111_1111111111111111_1110110011101010_1110111011101001"; -- -0.07454020325882943
	pesos_i(22721) := b"0000000000000000_0000000000000000_0000100111001001_0110010000010110"; -- 0.03822923229222261
	pesos_i(22722) := b"1111111111111111_1111111111111111_1111111100010001_0001111110010110"; -- -0.0036449680149748614
	pesos_i(22723) := b"0000000000000000_0000000000000000_0000101011111111_1000100111010101"; -- 0.04296170665966744
	pesos_i(22724) := b"1111111111111111_1111111111111111_1110101100010111_1100000000001011"; -- -0.08166885114071425
	pesos_i(22725) := b"1111111111111111_1111111111111111_1111100111111100_0110100100101011"; -- -0.023492266742681206
	pesos_i(22726) := b"0000000000000000_0000000000000000_0001000010101010_1101010011100111"; -- 0.06510668412062505
	pesos_i(22727) := b"1111111111111111_1111111111111111_1101110000110110_1010100011110101"; -- -0.13979095469245206
	pesos_i(22728) := b"0000000000000000_0000000000000000_0001100101111110_1000111010101101"; -- 0.09958736146889904
	pesos_i(22729) := b"1111111111111111_1111111111111111_1111011000110001_1101110100001011"; -- -0.03830164409176721
	pesos_i(22730) := b"0000000000000000_0000000000000000_0001111011101010_0110011000101110"; -- 0.12076414711180371
	pesos_i(22731) := b"1111111111111111_1111111111111111_1111000001110000_1001001000001010"; -- -0.0607823110482828
	pesos_i(22732) := b"1111111111111111_1111111111111111_1110110111110100_1011100011010010"; -- -0.07048458932254874
	pesos_i(22733) := b"0000000000000000_0000000000000000_0001000101101100_0000110111011100"; -- 0.0680550253144164
	pesos_i(22734) := b"0000000000000000_0000000000000000_0001100011101100_1101101010001011"; -- 0.0973641003415986
	pesos_i(22735) := b"0000000000000000_0000000000000000_0001111111011100_1000101011110001"; -- 0.12445896509244707
	pesos_i(22736) := b"1111111111111111_1111111111111111_1111111011100010_0001110110111100"; -- -0.004362241444899277
	pesos_i(22737) := b"0000000000000000_0000000000000000_0000110010111110_1111110111001100"; -- 0.049789297466257446
	pesos_i(22738) := b"0000000000000000_0000000000000000_0010001001101110_1111010110011100"; -- 0.13450560615917506
	pesos_i(22739) := b"1111111111111111_1111111111111111_1101100010100001_1011101101011100"; -- -0.1537821675079068
	pesos_i(22740) := b"1111111111111111_1111111111111111_1110101011111001_1101100100001000"; -- -0.08212512547657702
	pesos_i(22741) := b"1111111111111111_1111111111111111_1111001011111000_0101011101010010"; -- -0.05089811552618863
	pesos_i(22742) := b"1111111111111111_1111111111111111_1111010011001000_0011000101110011"; -- -0.04382029468105803
	pesos_i(22743) := b"1111111111111111_1111111111111111_1110111110101010_0011010101110100"; -- -0.0638090697413403
	pesos_i(22744) := b"0000000000000000_0000000000000000_0000011110110101_1110101011000000"; -- 0.030119583048201365
	pesos_i(22745) := b"0000000000000000_0000000000000000_0000010000101011_1001001001101100"; -- 0.016289855315838327
	pesos_i(22746) := b"0000000000000000_0000000000000000_0000100111001000_1101010110101011"; -- 0.038220743521963925
	pesos_i(22747) := b"0000000000000000_0000000000000000_0001010101010001_0111011101011001"; -- 0.08327432553251882
	pesos_i(22748) := b"1111111111111111_1111111111111111_1110111111111010_1001110101001101"; -- -0.06258217678613366
	pesos_i(22749) := b"0000000000000000_0000000000000000_0001000101000101_0001100101001001"; -- 0.06746061354272233
	pesos_i(22750) := b"1111111111111111_1111111111111111_1111001110011101_1101010110111010"; -- -0.04837288100394317
	pesos_i(22751) := b"0000000000000000_0000000000000000_0001100010011110_1010101010000110"; -- 0.09617105271913345
	pesos_i(22752) := b"1111111111111111_1111111111111111_1110110010000011_0001111000011110"; -- -0.07612430355615321
	pesos_i(22753) := b"1111111111111111_1111111111111111_1111111111000010_1010010111000010"; -- -0.0009361649697357831
	pesos_i(22754) := b"1111111111111111_1111111111111111_1110111111000111_0010001100011110"; -- -0.06336765779474052
	pesos_i(22755) := b"0000000000000000_0000000000000000_0001000111111101_1111111110000101"; -- 0.07028195378584731
	pesos_i(22756) := b"0000000000000000_0000000000000000_0000011010111001_1101010011100001"; -- 0.026273064478095357
	pesos_i(22757) := b"0000000000000000_0000000000000000_0010000101000111_1100001111100010"; -- 0.13000129959809228
	pesos_i(22758) := b"1111111111111111_1111111111111111_1101100110001010_1000100110000000"; -- -0.15022984152854685
	pesos_i(22759) := b"0000000000000000_0000000000000000_0001010101100000_0001010100101100"; -- 0.08349735562249555
	pesos_i(22760) := b"0000000000000000_0000000000000000_0000000110001111_1100011100001010"; -- 0.006100120445523521
	pesos_i(22761) := b"1111111111111111_1111111111111111_1111011011001000_0100110000000001"; -- -0.03600621196312074
	pesos_i(22762) := b"0000000000000000_0000000000000000_0000000101011001_0000000000010111"; -- 0.0052642876386587165
	pesos_i(22763) := b"0000000000000000_0000000000000000_0010001010100000_1111100110001110"; -- 0.1352687807977895
	pesos_i(22764) := b"0000000000000000_0000000000000000_0001100000100111_1101001011100010"; -- 0.09435766239133024
	pesos_i(22765) := b"0000000000000000_0000000000000000_0001010000111010_1110010011001110"; -- 0.07902364767402455
	pesos_i(22766) := b"0000000000000000_0000000000000000_0010011011011100_0110010100011101"; -- 0.1518004604064383
	pesos_i(22767) := b"0000000000000000_0000000000000000_0000010100100011_1010111000010010"; -- 0.02007568301531623
	pesos_i(22768) := b"1111111111111111_1111111111111111_1111100111110000_1010101111111011"; -- -0.023671389843714415
	pesos_i(22769) := b"0000000000000000_0000000000000000_0000001001100101_1001001001111001"; -- 0.009362368167002208
	pesos_i(22770) := b"0000000000000000_0000000000000000_0000011101011110_0111001000101000"; -- 0.028784880299072706
	pesos_i(22771) := b"0000000000000000_0000000000000000_0001101101000110_0001001000101111"; -- 0.10653794901934936
	pesos_i(22772) := b"0000000000000000_0000000000000000_0000100010001000_1100110101001110"; -- 0.033337432358660705
	pesos_i(22773) := b"0000000000000000_0000000000000000_0001000010100010_1000111111110111"; -- 0.0649805047151984
	pesos_i(22774) := b"1111111111111111_1111111111111111_1101110110001011_0111110001011011"; -- -0.13459036615041042
	pesos_i(22775) := b"1111111111111111_1111111111111111_1110110001001001_0100011110010111"; -- -0.0770068413895777
	pesos_i(22776) := b"0000000000000000_0000000000000000_0010000000111111_0101000110110011"; -- 0.12596617342515234
	pesos_i(22777) := b"1111111111111111_1111111111111111_1110010100000001_1101010110110110"; -- -0.10544075303703898
	pesos_i(22778) := b"1111111111111111_1111111111111111_1111110011001011_1111110010010000"; -- -0.012512411885229967
	pesos_i(22779) := b"0000000000000000_0000000000000000_0001000011100010_1110010011001110"; -- 0.06596212423974002
	pesos_i(22780) := b"0000000000000000_0000000000000000_0001001101111001_0110110110000101"; -- 0.07607159133825876
	pesos_i(22781) := b"1111111111111111_1111111111111111_1111001001100001_0001000001000010"; -- -0.05320642850520364
	pesos_i(22782) := b"1111111111111111_1111111111111111_1111000110110101_0001100100000011"; -- -0.05583041827932752
	pesos_i(22783) := b"0000000000000000_0000000000000000_0001101110111000_0110111111011000"; -- 0.10828303368383534
	pesos_i(22784) := b"1111111111111111_1111111111111111_1111100110010011_1111000010000110"; -- -0.025086371742035957
	pesos_i(22785) := b"0000000000000000_0000000000000000_0001111111001011_0011010010010100"; -- 0.1241944179946324
	pesos_i(22786) := b"0000000000000000_0000000000000000_0001101111100111_0111111011100000"; -- 0.10900109269751937
	pesos_i(22787) := b"0000000000000000_0000000000000000_0001110011011000_1100101011010001"; -- 0.11268298734952903
	pesos_i(22788) := b"0000000000000000_0000000000000000_0001101001010010_0101000111101010"; -- 0.10281860324945141
	pesos_i(22789) := b"1111111111111111_1111111111111111_1111111011011011_0000000001110011"; -- -0.0044707984950058035
	pesos_i(22790) := b"0000000000000000_0000000000000000_0000110101001000_1000110111001111"; -- 0.051888335267483314
	pesos_i(22791) := b"0000000000000000_0000000000000000_0001101001000100_0111100011001001"; -- 0.10260729694992439
	pesos_i(22792) := b"1111111111111111_1111111111111111_1111111010110010_0010110000100011"; -- -0.005093804820434346
	pesos_i(22793) := b"1111111111111111_1111111111111111_1110110011000111_1000110100011010"; -- -0.0750800906302105
	pesos_i(22794) := b"0000000000000000_0000000000000000_0010000001011000_0010001111010110"; -- 0.12634490933180503
	pesos_i(22795) := b"0000000000000000_0000000000000000_0000000001101110_0001110010011110"; -- 0.0016801725669544033
	pesos_i(22796) := b"0000000000000000_0000000000000000_0001000011011011_0100000101000001"; -- 0.06584556432880732
	pesos_i(22797) := b"1111111111111111_1111111111111111_1101111000110001_1101011111011101"; -- -0.13205195296735256
	pesos_i(22798) := b"0000000000000000_0000000000000000_0001001110111000_1011000110111001"; -- 0.07703696037390768
	pesos_i(22799) := b"0000000000000000_0000000000000000_0010010111010010_0111001010001111"; -- 0.14774242403361826
	pesos_i(22800) := b"0000000000000000_0000000000000000_0001101100001111_1011001100000110"; -- 0.10570830237754236
	pesos_i(22801) := b"0000000000000000_0000000000000000_0000110011100100_1110101001001101"; -- 0.05036796926183473
	pesos_i(22802) := b"0000000000000000_0000000000000000_0001110101111111_0000000101000100"; -- 0.11521919175433715
	pesos_i(22803) := b"0000000000000000_0000000000000000_0010010101010001_1110100001000100"; -- 0.14578105612119688
	pesos_i(22804) := b"1111111111111111_1111111111111111_1110011100111110_0101110010010001"; -- -0.09670468768253856
	pesos_i(22805) := b"1111111111111111_1111111111111111_1111111110100100_1001111000000111"; -- -0.001394389447895729
	pesos_i(22806) := b"1111111111111111_1111111111111111_1110100000111111_0000110100101111"; -- -0.09278791055628563
	pesos_i(22807) := b"1111111111111111_1111111111111111_1101101100011000_0101110101111000"; -- -0.14415946781774316
	pesos_i(22808) := b"0000000000000000_0000000000000000_0001000010100100_0100110011100000"; -- 0.0650070234935006
	pesos_i(22809) := b"1111111111111111_1111111111111111_1111011001100000_0100110101111000"; -- -0.03759303871225876
	pesos_i(22810) := b"1111111111111111_1111111111111111_1110000011011101_1001010101110111"; -- -0.12161889874098948
	pesos_i(22811) := b"1111111111111111_1111111111111111_1111110001001101_1000011000100110"; -- -0.014442077323887517
	pesos_i(22812) := b"0000000000000000_0000000000000000_0001100000001000_1000010101010110"; -- 0.09388001779383678
	pesos_i(22813) := b"0000000000000000_0000000000000000_0010001011101001_1000011011111100"; -- 0.13637584348854578
	pesos_i(22814) := b"0000000000000000_0000000000000000_0001100110101011_0100100111101101"; -- 0.10026990933729003
	pesos_i(22815) := b"1111111111111111_1111111111111111_1110100101000100_1010101100011100"; -- -0.08879595332034693
	pesos_i(22816) := b"0000000000000000_0000000000000000_0000100000101001_1111110100111010"; -- 0.031890703817461195
	pesos_i(22817) := b"1111111111111111_1111111111111111_1110101110101101_1011101010010011"; -- -0.07938035887972245
	pesos_i(22818) := b"0000000000000000_0000000000000000_0000111100010110_1101000101101011"; -- 0.05894192574612446
	pesos_i(22819) := b"1111111111111111_1111111111111111_1110011001110011_1010011110010100"; -- -0.09979775091582456
	pesos_i(22820) := b"1111111111111111_1111111111111111_1111010000010101_1101000101100011"; -- -0.046542084972900404
	pesos_i(22821) := b"1111111111111111_1111111111111111_1110100000010110_1111011011111010"; -- -0.0933995856359983
	pesos_i(22822) := b"0000000000000000_0000000000000000_0010010000000101_1100100011101100"; -- 0.14071326975998227
	pesos_i(22823) := b"1111111111111111_1111111111111111_1111101100111111_0100010010101010"; -- -0.018565853642771437
	pesos_i(22824) := b"0000000000000000_0000000000000000_0000100100111100_0100110100110100"; -- 0.036076378903927765
	pesos_i(22825) := b"1111111111111111_1111111111111111_1110001101101011_0001011101001111"; -- -0.11164717029364261
	pesos_i(22826) := b"0000000000000000_0000000000000000_0001101011101001_0101000110010110"; -- 0.10512266077113959
	pesos_i(22827) := b"0000000000000000_0000000000000000_0001011000110011_0000000111011101"; -- 0.0867158093950268
	pesos_i(22828) := b"1111111111111111_1111111111111111_1110000101101000_1010001110011111"; -- -0.11949708342179785
	pesos_i(22829) := b"1111111111111111_1111111111111111_1111000011011110_0111110011011011"; -- -0.059105106962648604
	pesos_i(22830) := b"0000000000000000_0000000000000000_0000111001100000_0010100011001011"; -- 0.0561547751212679
	pesos_i(22831) := b"1111111111111111_1111111111111111_1111110011010001_1010110101001110"; -- -0.012425583388550737
	pesos_i(22832) := b"1111111111111111_1111111111111111_1110011101100001_1101110101010011"; -- -0.09616295556442164
	pesos_i(22833) := b"0000000000000000_0000000000000000_0001100101101111_0100100101001000"; -- 0.09935434350501134
	pesos_i(22834) := b"1111111111111111_1111111111111111_1110101101110110_1011010111100101"; -- -0.08021987109963886
	pesos_i(22835) := b"0000000000000000_0000000000000000_0010010101101010_0111110111110101"; -- 0.14615618926745771
	pesos_i(22836) := b"0000000000000000_0000000000000000_0001101001000001_1101111111011101"; -- 0.10256766451741908
	pesos_i(22837) := b"1111111111111111_1111111111111111_1110100000100010_1110010000101011"; -- -0.09321760139460769
	pesos_i(22838) := b"1111111111111111_1111111111111111_1110011010111011_1000001001001101"; -- -0.09870133990120052
	pesos_i(22839) := b"1111111111111111_1111111111111111_1110001010011100_0010010110111100"; -- -0.114804879687381
	pesos_i(22840) := b"0000000000000000_0000000000000000_0001100000100010_0001100110001011"; -- 0.09427032140801421
	pesos_i(22841) := b"1111111111111111_1111111111111111_1111111000110111_1010001010111001"; -- -0.006963567624316379
	pesos_i(22842) := b"1111111111111111_1111111111111111_1111100100100110_0100110111110010"; -- -0.026759270053659787
	pesos_i(22843) := b"0000000000000000_0000000000000000_0001110001101001_0100101100111011"; -- 0.11098165695782322
	pesos_i(22844) := b"1111111111111111_1111111111111111_1111011110011011_1000011000110101"; -- -0.032783138222753756
	pesos_i(22845) := b"0000000000000000_0000000000000000_0001110000011000_0111110101101010"; -- 0.10974868608328389
	pesos_i(22846) := b"1111111111111111_1111111111111111_1101110010001100_1000111000101111"; -- -0.1384802946904398
	pesos_i(22847) := b"1111111111111111_1111111111111111_1101110101100011_1001101010101111"; -- -0.13519890994270484
	pesos_i(22848) := b"0000000000000000_0000000000000000_0000011010101111_1101010011000011"; -- 0.026120469625910327
	pesos_i(22849) := b"1111111111111111_1111111111111111_1110111111100110_0011100001001011"; -- -0.06289337312797073
	pesos_i(22850) := b"1111111111111111_1111111111111111_1110111111001100_1010101110100011"; -- -0.06328322663471801
	pesos_i(22851) := b"0000000000000000_0000000000000000_0000011000000010_0111011101101010"; -- 0.02347513516696062
	pesos_i(22852) := b"1111111111111111_1111111111111111_1101011101100111_0001011101111101"; -- -0.15858319462323894
	pesos_i(22853) := b"1111111111111111_1111111111111111_1111010100000110_1110001100010001"; -- -0.042863663077392034
	pesos_i(22854) := b"1111111111111111_1111111111111111_1111011110110011_1111111110101101"; -- -0.03240968739033253
	pesos_i(22855) := b"0000000000000000_0000000000000000_0010001111010111_1101100010101010"; -- 0.14001230372260806
	pesos_i(22856) := b"1111111111111111_1111111111111111_1110011110011111_1010010101101101"; -- -0.0952202424260722
	pesos_i(22857) := b"1111111111111111_1111111111111111_1101101111111100_0000001011101011"; -- -0.14068586113421602
	pesos_i(22858) := b"0000000000000000_0000000000000000_0001101000100100_0110010101010010"; -- 0.10211785561771289
	pesos_i(22859) := b"1111111111111111_1111111111111111_1111000111101010_1011111100100001"; -- -0.05501180117762656
	pesos_i(22860) := b"1111111111111111_1111111111111111_1101011010100101_1110111001010110"; -- -0.16153059396386005
	pesos_i(22861) := b"1111111111111111_1111111111111111_1111001000100101_0101110001010001"; -- -0.05411742237826535
	pesos_i(22862) := b"0000000000000000_0000000000000000_0001110111100100_1010010010010110"; -- 0.1167700640264197
	pesos_i(22863) := b"0000000000000000_0000000000000000_0001100111000100_1011100101011001"; -- 0.1006580202547244
	pesos_i(22864) := b"0000000000000000_0000000000000000_0001111001101011_1110001010010110"; -- 0.1188336959153688
	pesos_i(22865) := b"1111111111111111_1111111111111111_1101110100001011_1010110001111011"; -- -0.13654062272908063
	pesos_i(22866) := b"1111111111111111_1111111111111111_1111011101101001_1110101111111111"; -- -0.033540010756485744
	pesos_i(22867) := b"0000000000000000_0000000000000000_0001010101010001_1011110100001101"; -- 0.08327848012747609
	pesos_i(22868) := b"0000000000000000_0000000000000000_0010000101010000_0001000001001111"; -- 0.13012792518049174
	pesos_i(22869) := b"0000000000000000_0000000000000000_0001111001111101_1110010000110000"; -- 0.11910844974319529
	pesos_i(22870) := b"0000000000000000_0000000000000000_0001011010111111_0000010101111000"; -- 0.08885225468665447
	pesos_i(22871) := b"0000000000000000_0000000000000000_0010011110000010_0111101100010010"; -- 0.15433472819231325
	pesos_i(22872) := b"0000000000000000_0000000000000000_0000111100110110_1110010101010111"; -- 0.05943139425859082
	pesos_i(22873) := b"0000000000000000_0000000000000000_0010000011011000_0100001110101001"; -- 0.12829993140417953
	pesos_i(22874) := b"1111111111111111_1111111111111111_1110011001111000_1101000001111000"; -- -0.09971901963732947
	pesos_i(22875) := b"1111111111111111_1111111111111111_1101011010101110_1110110111010011"; -- -0.16139329518739434
	pesos_i(22876) := b"1111111111111111_1111111111111111_1111110011110000_0011100110101101"; -- -0.011959452786661492
	pesos_i(22877) := b"1111111111111111_1111111111111111_1111101000100001_0010101100101111"; -- -0.022931385967004576
	pesos_i(22878) := b"1111111111111111_1111111111111111_1111000111111101_1110010110101010"; -- -0.05471958727847048
	pesos_i(22879) := b"1111111111111111_1111111111111111_1111101000010011_0001000111010101"; -- -0.023146520251677127
	pesos_i(22880) := b"0000000000000000_0000000000000000_0000101111001011_0100101010111001"; -- 0.04607073807607377
	pesos_i(22881) := b"1111111111111111_1111111111111111_1111111011000110_1101101000101110"; -- -0.004778255332226534
	pesos_i(22882) := b"1111111111111111_1111111111111111_1110100111000111_1001000100101101"; -- -0.08679859773835637
	pesos_i(22883) := b"1111111111111111_1111111111111111_1110011110101111_0110011110100010"; -- -0.09497978480447043
	pesos_i(22884) := b"0000000000000000_0000000000000000_0010000100101101_1101010001000111"; -- 0.1296055481539418
	pesos_i(22885) := b"1111111111111111_1111111111111111_1110100100010111_0001001000000100"; -- -0.08949172400906243
	pesos_i(22886) := b"1111111111111111_1111111111111111_1101100111101000_1011000011010100"; -- -0.14879317108621293
	pesos_i(22887) := b"1111111111111111_1111111111111111_1101001001010110_0001111100111011"; -- -0.17837338259403376
	pesos_i(22888) := b"1111111111111111_1111111111111111_1110101001000110_1000001010101000"; -- -0.08486159697731309
	pesos_i(22889) := b"1111111111111111_1111111111111111_1101101110000000_0100101110100010"; -- -0.14257361683116884
	pesos_i(22890) := b"0000000000000000_0000000000000000_0000011001111100_1101001010101001"; -- 0.025342146116428696
	pesos_i(22891) := b"1111111111111111_1111111111111111_1101110100101001_0101000011011111"; -- -0.1360883194298387
	pesos_i(22892) := b"0000000000000000_0000000000000000_0010010010000011_0011001011001010"; -- 0.14262692857607184
	pesos_i(22893) := b"0000000000000000_0000000000000000_0000000000010101_0110001001111110"; -- 0.0003263050470227506
	pesos_i(22894) := b"1111111111111111_1111111111111111_1111100010111110_1001001000001101"; -- -0.02834212481604894
	pesos_i(22895) := b"1111111111111111_1111111111111111_1111000000101011_1000111110111010"; -- -0.06183530530002617
	pesos_i(22896) := b"1111111111111111_1111111111111111_1111000111001011_1110101011110011"; -- -0.055482211662814404
	pesos_i(22897) := b"0000000000000000_0000000000000000_0000000000110101_0100101111111000"; -- 0.0008132438820923624
	pesos_i(22898) := b"0000000000000000_0000000000000000_0001010001100010_1000011011111100"; -- 0.07962840697651863
	pesos_i(22899) := b"0000000000000000_0000000000000000_0001111010100100_0111001110111001"; -- 0.11969683909676906
	pesos_i(22900) := b"1111111111111111_1111111111111111_1110011110111011_1100110001010101"; -- -0.09479067723947768
	pesos_i(22901) := b"0000000000000000_0000000000000000_0000101000100010_0010010111001010"; -- 0.03958355129135116
	pesos_i(22902) := b"0000000000000000_0000000000000000_0001100001000000_0000010010110001"; -- 0.09472684201709572
	pesos_i(22903) := b"0000000000000000_0000000000000000_0000010010110011_1110001110001111"; -- 0.018369886727787582
	pesos_i(22904) := b"1111111111111111_1111111111111111_1111101111011000_0001101101010101"; -- -0.01623372240236676
	pesos_i(22905) := b"1111111111111111_1111111111111111_1110110001100011_0001001101010100"; -- -0.076613227898928
	pesos_i(22906) := b"1111111111111111_1111111111111111_1110100101000011_0110001111100100"; -- -0.08881545710249145
	pesos_i(22907) := b"0000000000000000_0000000000000000_0000111101001010_0111110110100100"; -- 0.05973038908774094
	pesos_i(22908) := b"1111111111111111_1111111111111111_1110100000111001_1101110101111001"; -- -0.09286704827158088
	pesos_i(22909) := b"0000000000000000_0000000000000000_0000111010111100_1011111100100001"; -- 0.057567544476300796
	pesos_i(22910) := b"0000000000000000_0000000000000000_0001001111010010_0011111100111100"; -- 0.07742686473765224
	pesos_i(22911) := b"0000000000000000_0000000000000000_0001111101111101_1111010111000010"; -- 0.12301574696869473
	pesos_i(22912) := b"1111111111111111_1111111111111111_1111000010110011_0010000001101001"; -- -0.0597667450710206
	pesos_i(22913) := b"0000000000000000_0000000000000000_0001111100011001_0101010111010010"; -- 0.12148033503070613
	pesos_i(22914) := b"0000000000000000_0000000000000000_0000001011011000_0110001111111111"; -- 0.011114358750770098
	pesos_i(22915) := b"0000000000000000_0000000000000000_0000100010110011_1100111001001110"; -- 0.033993620074919885
	pesos_i(22916) := b"1111111111111111_1111111111111111_1110000100001110_0101001000000100"; -- -0.12087523834400338
	pesos_i(22917) := b"1111111111111111_1111111111111111_1111001110111011_1001100000110011"; -- -0.04791878477251434
	pesos_i(22918) := b"1111111111111111_1111111111111111_1111001110011111_1100011000000111"; -- -0.04834329924749348
	pesos_i(22919) := b"1111111111111111_1111111111111111_1111111111111110_1001010100001100"; -- -2.1633729057367128e-05
	pesos_i(22920) := b"0000000000000000_0000000000000000_0000011100101100_1000111110101011"; -- 0.028023700087031186
	pesos_i(22921) := b"0000000000000000_0000000000000000_0001001111010110_1001010111111101"; -- 0.07749307085196602
	pesos_i(22922) := b"0000000000000000_0000000000000000_0000010100110011_0111110100111001"; -- 0.02031691216281396
	pesos_i(22923) := b"1111111111111111_1111111111111111_1101111100110010_1110100100101011"; -- -0.1281294127370517
	pesos_i(22924) := b"0000000000000000_0000000000000000_0001000000001011_0011110101011111"; -- 0.06267150476481047
	pesos_i(22925) := b"0000000000000000_0000000000000000_0000100011111101_0011100000010111"; -- 0.03511381688387341
	pesos_i(22926) := b"0000000000000000_0000000000000000_0001010011100000_1000110000110111"; -- 0.08155132619103625
	pesos_i(22927) := b"1111111111111111_1111111111111111_1101101001101100_1110110111010000"; -- -0.14677537604483412
	pesos_i(22928) := b"1111111111111111_1111111111111111_1111101101000011_0000100110110001"; -- -0.01850833347835042
	pesos_i(22929) := b"1111111111111111_1111111111111111_1110110111011011_0000111011011011"; -- -0.07087618973778516
	pesos_i(22930) := b"1111111111111111_1111111111111111_1101110011101110_0000111011110011"; -- -0.13699251715264682
	pesos_i(22931) := b"1111111111111111_1111111111111111_1110000010000001_1111011101000100"; -- -0.12301687811728028
	pesos_i(22932) := b"1111111111111111_1111111111111111_1110010011000010_1001011001100011"; -- -0.10640583126134585
	pesos_i(22933) := b"0000000000000000_0000000000000000_0001011011100000_0001100000000101"; -- 0.08935690046666192
	pesos_i(22934) := b"1111111111111111_1111111111111111_1110010100111111_1010111101100110"; -- -0.10449699165387809
	pesos_i(22935) := b"0000000000000000_0000000000000000_0000110011111011_0010100111101001"; -- 0.05070745418138752
	pesos_i(22936) := b"1111111111111111_1111111111111111_1110000101000100_0110010110111101"; -- -0.12005008832599028
	pesos_i(22937) := b"0000000000000000_0000000000000000_0001001010111100_1110111011001111"; -- 0.07319538636956407
	pesos_i(22938) := b"0000000000000000_0000000000000000_0001100000101010_0001100111011000"; -- 0.0943924096159038
	pesos_i(22939) := b"0000000000000000_0000000000000000_0010000101100110_0001100101101000"; -- 0.13046416081409223
	pesos_i(22940) := b"0000000000000000_0000000000000000_0000010100011011_0011000110101111"; -- 0.019946198633938067
	pesos_i(22941) := b"1111111111111111_1111111111111111_1110001011110001_0100010000000000"; -- -0.11350607861573787
	pesos_i(22942) := b"0000000000000000_0000000000000000_0010001110010001_0101111101011111"; -- 0.13893695905370163
	pesos_i(22943) := b"0000000000000000_0000000000000000_0001010100010110_0000010010100110"; -- 0.08236722042298977
	pesos_i(22944) := b"1111111111111111_1111111111111111_1101100000100011_1110110010111010"; -- -0.15570183243236743
	pesos_i(22945) := b"1111111111111111_1111111111111111_1111011111101001_0100111001100001"; -- -0.031596280500849505
	pesos_i(22946) := b"1111111111111111_1111111111111111_1111110100111000_0111100111111110"; -- -0.010856986488614712
	pesos_i(22947) := b"0000000000000000_0000000000000000_0001101111101011_1011101110001001"; -- 0.10906574339723811
	pesos_i(22948) := b"1111111111111111_1111111111111111_1110000111101011_1001101101110110"; -- -0.1174986683168772
	pesos_i(22949) := b"1111111111111111_1111111111111111_1110010010110110_0100001011110001"; -- -0.10659391037030025
	pesos_i(22950) := b"0000000000000000_0000000000000000_0000110010110111_1001011011111100"; -- 0.049676357685912324
	pesos_i(22951) := b"1111111111111111_1111111111111111_1110111010001100_0011111100101000"; -- -0.06817250506120114
	pesos_i(22952) := b"0000000000000000_0000000000000000_0000010110110010_1010100011111011"; -- 0.022257386390926656
	pesos_i(22953) := b"0000000000000000_0000000000000000_0010100011010111_0111000101000110"; -- 0.15953739118448454
	pesos_i(22954) := b"0000000000000000_0000000000000000_0001011101011000_1111000101100101"; -- 0.09120091178075648
	pesos_i(22955) := b"1111111111111111_1111111111111111_1110011001101111_1111100111011110"; -- -0.09985388126292416
	pesos_i(22956) := b"0000000000000000_0000000000000000_0001001111111010_1100010111111100"; -- 0.07804524796134284
	pesos_i(22957) := b"1111111111111111_1111111111111111_1111010001010011_1110110011010111"; -- -0.04559440365989561
	pesos_i(22958) := b"1111111111111111_1111111111111111_1111100010110111_0111100010001111"; -- -0.028450455759062694
	pesos_i(22959) := b"1111111111111111_1111111111111111_1111100000010101_0100100001001110"; -- -0.030925255846113085
	pesos_i(22960) := b"0000000000000000_0000000000000000_0000011110001001_0100111010111001"; -- 0.02943889640560161
	pesos_i(22961) := b"1111111111111111_1111111111111111_1110010111001101_0100101110000001"; -- -0.10233619794332341
	pesos_i(22962) := b"1111111111111111_1111111111111111_1111010000010100_1011001110100010"; -- -0.046559117314813644
	pesos_i(22963) := b"1111111111111111_1111111111111111_1101101010111001_0000111000101111"; -- -0.14561377856187152
	pesos_i(22964) := b"0000000000000000_0000000000000000_0010000100110111_0010000001001111"; -- 0.12974740918375638
	pesos_i(22965) := b"0000000000000000_0000000000000000_0001011010010110_1011000111011100"; -- 0.08823691949035592
	pesos_i(22966) := b"1111111111111111_1111111111111111_1110010101100001_0010010110100110"; -- -0.10398640344915702
	pesos_i(22967) := b"0000000000000000_0000000000000000_0001101001001100_1000011100000111"; -- 0.10273021615297963
	pesos_i(22968) := b"0000000000000000_0000000000000000_0001011001001101_0101100110001000"; -- 0.08711776332771887
	pesos_i(22969) := b"1111111111111111_1111111111111111_1110001011011110_0110011100100110"; -- -0.11379390076581182
	pesos_i(22970) := b"1111111111111111_1111111111111111_1110111110000011_0000100010111001"; -- -0.06440682882886926
	pesos_i(22971) := b"1111111111111111_1111111111111111_1111110100001101_0100000010001101"; -- -0.011516538161599909
	pesos_i(22972) := b"1111111111111111_1111111111111111_1101110010110100_1111010010101110"; -- -0.13786383399492486
	pesos_i(22973) := b"1111111111111111_1111111111111111_1111010101010001_1000001111000110"; -- -0.04172493389270977
	pesos_i(22974) := b"0000000000000000_0000000000000000_0010001110010011_0001000000001000"; -- 0.1389627475981306
	pesos_i(22975) := b"1111111111111111_1111111111111111_1101101101100100_0110011100111111"; -- -0.142999217051775
	pesos_i(22976) := b"0000000000000000_0000000000000000_0000011010101101_1100110011101100"; -- 0.026089484906066402
	pesos_i(22977) := b"0000000000000000_0000000000000000_0010000010000000_1000111100111010"; -- 0.12696166192203065
	pesos_i(22978) := b"1111111111111111_1111111111111111_1111000110001111_0011110011110101"; -- -0.056408109892214134
	pesos_i(22979) := b"0000000000000000_0000000000000000_0000100110111111_0110011010000010"; -- 0.0380767887472941
	pesos_i(22980) := b"0000000000000000_0000000000000000_0001010011000100_1011101111101111"; -- 0.0811269243264436
	pesos_i(22981) := b"0000000000000000_0000000000000000_0000001100101001_0110011000101010"; -- 0.012350449699513813
	pesos_i(22982) := b"0000000000000000_0000000000000000_0001111101001100_1101001011000110"; -- 0.12226598093891428
	pesos_i(22983) := b"1111111111111111_1111111111111111_1110100000110111_0111010100101000"; -- -0.09290378355956364
	pesos_i(22984) := b"1111111111111111_1111111111111111_1111110010001011_0000111100010011"; -- -0.013503129760050515
	pesos_i(22985) := b"1111111111111111_1111111111111111_1110100101100111_0011011111000110"; -- -0.08826877045609378
	pesos_i(22986) := b"1111111111111111_1111111111111111_1110001110000100_1101000010011011"; -- -0.11125465595161757
	pesos_i(22987) := b"1111111111111111_1111111111111111_1111110011101010_1111111001010111"; -- -0.012039283433653201
	pesos_i(22988) := b"0000000000000000_0000000000000000_0010011100000111_0110100001010001"; -- 0.1524567791614096
	pesos_i(22989) := b"1111111111111111_1111111111111111_1110101011110111_0101000000100111"; -- -0.08216380155448674
	pesos_i(22990) := b"0000000000000000_0000000000000000_0000010101110111_0100110011001110"; -- 0.021351623873997944
	pesos_i(22991) := b"0000000000000000_0000000000000000_0000100011011011_1101111001110111"; -- 0.03460493476458007
	pesos_i(22992) := b"0000000000000000_0000000000000000_0000000001101101_1011111001000010"; -- 0.0016745482950924198
	pesos_i(22993) := b"0000000000000000_0000000000000000_0000100010011101_0010111010110001"; -- 0.033648412801585675
	pesos_i(22994) := b"0000000000000000_0000000000000000_0001010100000010_0100111111010111"; -- 0.08206652644063457
	pesos_i(22995) := b"1111111111111111_1111111111111111_1101110011100001_1010001111001001"; -- -0.1371820100292238
	pesos_i(22996) := b"0000000000000000_0000000000000000_0001010111001110_1101001000100110"; -- 0.08518708646510664
	pesos_i(22997) := b"0000000000000000_0000000000000000_0000101001001101_0110100010011111"; -- 0.040243662659329264
	pesos_i(22998) := b"0000000000000000_0000000000000000_0010010101101100_0000001010100100"; -- 0.14617935667259876
	pesos_i(22999) := b"0000000000000000_0000000000000000_0010001101110010_1010110010111011"; -- 0.13846854747906867
	pesos_i(23000) := b"0000000000000000_0000000000000000_0000010101100110_0000100101100111"; -- 0.021088206870115766
	pesos_i(23001) := b"1111111111111111_1111111111111111_1111001010101010_1011001101001011"; -- -0.05208281905975934
	pesos_i(23002) := b"0000000000000000_0000000000000000_0001001111111001_0001100001001110"; -- 0.07801963722214153
	pesos_i(23003) := b"0000000000000000_0000000000000000_0000100110001011_0111010011111100"; -- 0.03728419455529404
	pesos_i(23004) := b"0000000000000000_0000000000000000_0001100000101101_0101000000000101"; -- 0.09444141497313534
	pesos_i(23005) := b"0000000000000000_0000000000000000_0010011000110010_0101011110110010"; -- 0.1492056664574801
	pesos_i(23006) := b"1111111111111111_1111111111111111_1110000101110001_0110011111011001"; -- -0.1193633169345589
	pesos_i(23007) := b"0000000000000000_0000000000000000_0010000101011000_0011000011101011"; -- 0.1302519392343493
	pesos_i(23008) := b"1111111111111111_1111111111111111_1110110100001101_0101011011110010"; -- -0.07401520341277992
	pesos_i(23009) := b"1111111111111111_1111111111111111_1111001111001011_0011001010010110"; -- -0.047680700547123034
	pesos_i(23010) := b"1111111111111111_1111111111111111_1111011011010000_1000011100110110"; -- -0.035880612598363316
	pesos_i(23011) := b"1111111111111111_1111111111111111_1111000100000000_1110000111010101"; -- -0.05858028938555389
	pesos_i(23012) := b"1111111111111111_1111111111111111_1110101110100011_0001111110010100"; -- -0.07954218527289902
	pesos_i(23013) := b"1111111111111111_1111111111111111_1110110111100000_1011010101010001"; -- -0.07078997397749107
	pesos_i(23014) := b"0000000000000000_0000000000000000_0001110111010111_0011110000011001"; -- 0.11656547165014547
	pesos_i(23015) := b"1111111111111111_1111111111111111_1110100011011001_1101011111001010"; -- -0.09042598067477248
	pesos_i(23016) := b"0000000000000000_0000000000000000_0001101001101001_0111010000110100"; -- 0.10317159905009367
	pesos_i(23017) := b"1111111111111111_1111111111111111_1110101000100010_1111001001001010"; -- -0.08540425956810888
	pesos_i(23018) := b"1111111111111111_1111111111111111_1110100110110010_1111010111110010"; -- -0.08711302595290639
	pesos_i(23019) := b"0000000000000000_0000000000000000_0000010110000010_0111000011000000"; -- 0.021521612978205807
	pesos_i(23020) := b"0000000000000000_0000000000000000_0000010000010100_0100011010101001"; -- 0.015934387393469474
	pesos_i(23021) := b"0000000000000000_0000000000000000_0001010110011101_1000010100011101"; -- 0.0844348141467625
	pesos_i(23022) := b"1111111111111111_1111111111111111_1110000111111101_1001101010101000"; -- -0.11722405816023145
	pesos_i(23023) := b"1111111111111111_1111111111111111_1101100101001000_0110011011111110"; -- -0.15123897832827587
	pesos_i(23024) := b"1111111111111111_1111111111111111_1110011101100110_1111010011011111"; -- -0.09608525802426937
	pesos_i(23025) := b"1111111111111111_1111111111111111_1111100110111100_0101010010000011"; -- -0.024470060477530614
	pesos_i(23026) := b"0000000000000000_0000000000000000_0001101010110110_1000010101101110"; -- 0.10434755269321816
	pesos_i(23027) := b"1111111111111111_1111111111111111_1110010101101011_1101110100011011"; -- -0.1038228806342263
	pesos_i(23028) := b"0000000000000000_0000000000000000_0001110101110001_1110001010010000"; -- 0.11501899742182164
	pesos_i(23029) := b"0000000000000000_0000000000000000_0000110011101011_0111100001101100"; -- 0.05046799324667968
	pesos_i(23030) := b"0000000000000000_0000000000000000_0001100100111010_1000111110000010"; -- 0.09854981344565557
	pesos_i(23031) := b"1111111111111111_1111111111111111_1111001111000001_1101000111001010"; -- -0.04782379935231312
	pesos_i(23032) := b"0000000000000000_0000000000000000_0000110011100111_0101100111100001"; -- 0.05040513757034397
	pesos_i(23033) := b"0000000000000000_0000000000000000_0000110001111010_0010011110101011"; -- 0.048738936570242836
	pesos_i(23034) := b"0000000000000000_0000000000000000_0001010100000010_0010101001110110"; -- 0.08206429845119902
	pesos_i(23035) := b"0000000000000000_0000000000000000_0001100110001111_1101111110100001"; -- 0.09985158606044811
	pesos_i(23036) := b"0000000000000000_0000000000000000_0001010110101011_0011001110010000"; -- 0.08464357635450967
	pesos_i(23037) := b"0000000000000000_0000000000000000_0010011100010001_1101011001001000"; -- 0.15261592168583818
	pesos_i(23038) := b"1111111111111111_1111111111111111_1110110111010101_0111011001101110"; -- -0.07096156885430548
	pesos_i(23039) := b"1111111111111111_1111111111111111_1111000001011001_0101011000110010"; -- -0.06113683009952133
	pesos_i(23040) := b"0000000000000000_0000000000000000_0001011110001011_1111011001111010"; -- 0.09197941276136769
	pesos_i(23041) := b"1111111111111111_1111111111111111_1111110100011101_1000110111111011"; -- -0.011267782468023051
	pesos_i(23042) := b"0000000000000000_0000000000000000_0001111100001001_0101001110011110"; -- 0.12123606302961877
	pesos_i(23043) := b"1111111111111111_1111111111111111_1111111101011100_1100110111100011"; -- -0.0024901696166619463
	pesos_i(23044) := b"1111111111111111_1111111111111111_1110000000000011_1110110001110110"; -- -0.1249401294565452
	pesos_i(23045) := b"1111111111111111_1111111111111111_1101100101011000_0011100011111101"; -- -0.15099757986101756
	pesos_i(23046) := b"0000000000000000_0000000000000000_0000011101100010_0111110000101111"; -- 0.028846513285415005
	pesos_i(23047) := b"0000000000000000_0000000000000000_0001000011100110_1011010110100110"; -- 0.06602034859220397
	pesos_i(23048) := b"1111111111111111_1111111111111111_1111110100101111_1100100101101001"; -- -0.010989581940934466
	pesos_i(23049) := b"1111111111111111_1111111111111111_1110010111001011_0100011111011100"; -- -0.10236693264880553
	pesos_i(23050) := b"1111111111111111_1111111111111111_1110000010111010_0011101100001100"; -- -0.1221583457070105
	pesos_i(23051) := b"0000000000000000_0000000000000000_0000011000011011_1101111001011001"; -- 0.023862740349501633
	pesos_i(23052) := b"1111111111111111_1111111111111111_1111101011111010_0011111111001011"; -- -0.01961900034289873
	pesos_i(23053) := b"1111111111111111_1111111111111111_1110000111111100_1101101001011000"; -- -0.11723552085789457
	pesos_i(23054) := b"0000000000000000_0000000000000000_0010010101110001_0111110110001000"; -- 0.14626297546871528
	pesos_i(23055) := b"1111111111111111_1111111111111111_1111011111110001_1000011011001001"; -- -0.03147084807873992
	pesos_i(23056) := b"0000000000000000_0000000000000000_0010001000001111_1011111010100100"; -- 0.13305274489753108
	pesos_i(23057) := b"1111111111111111_1111111111111111_1111011100111011_0010001011000010"; -- -0.03425390968871611
	pesos_i(23058) := b"1111111111111111_1111111111111111_1111000000100101_0011010101101110"; -- -0.061932240036178796
	pesos_i(23059) := b"1111111111111111_1111111111111111_1111010000101000_0011110010101101"; -- -0.04626103188826374
	pesos_i(23060) := b"1111111111111111_1111111111111111_1111011110011101_1111010000011001"; -- -0.032746070797837624
	pesos_i(23061) := b"0000000000000000_0000000000000000_0000111111110101_1000010001000101"; -- 0.06234003711114569
	pesos_i(23062) := b"0000000000000000_0000000000000000_0000110110010010_0110111110110001"; -- 0.05301569061591085
	pesos_i(23063) := b"1111111111111111_1111111111111111_1110110001100000_1000110100101010"; -- -0.07665174213887173
	pesos_i(23064) := b"0000000000000000_0000000000000000_0001010010101010_0101000101011011"; -- 0.08072384320165592
	pesos_i(23065) := b"1111111111111111_1111111111111111_1111011001000001_1101010001111011"; -- -0.038058013822656354
	pesos_i(23066) := b"0000000000000000_0000000000000000_0010001101100111_0011111010111100"; -- 0.13829414446647237
	pesos_i(23067) := b"0000000000000000_0000000000000000_0000111011001101_1000110101100000"; -- 0.05782397839720845
	pesos_i(23068) := b"1111111111111111_1111111111111111_1111111001110000_0100000001011000"; -- -0.00609968051457462
	pesos_i(23069) := b"0000000000000000_0000000000000000_0000100111000100_0110010000001100"; -- 0.03815293583007566
	pesos_i(23070) := b"1111111111111111_1111111111111111_1111001001000101_1000110000111100"; -- -0.05362628487352535
	pesos_i(23071) := b"1111111111111111_1111111111111111_1101100000110010_1010010111101010"; -- -0.15547717141299755
	pesos_i(23072) := b"0000000000000000_0000000000000000_0010010001110100_0010100101100110"; -- 0.1423974871712225
	pesos_i(23073) := b"0000000000000000_0000000000000000_0000010101101011_1111010000100110"; -- 0.021178492727466077
	pesos_i(23074) := b"1111111111111111_1111111111111111_1111101000000100_1101001110000100"; -- -0.023363857478033098
	pesos_i(23075) := b"0000000000000000_0000000000000000_0001001100111101_0111010010001101"; -- 0.07515648317408198
	pesos_i(23076) := b"1111111111111111_1111111111111111_1111110001000010_1011110011101101"; -- -0.014606659061444855
	pesos_i(23077) := b"0000000000000000_0000000000000000_0000001011111111_1110101100000110"; -- 0.011717499665669496
	pesos_i(23078) := b"0000000000000000_0000000000000000_0001101100101100_1110001110001100"; -- 0.10615369957890411
	pesos_i(23079) := b"1111111111111111_1111111111111111_1111111100000000_1111100111010100"; -- -0.003891359064528078
	pesos_i(23080) := b"1111111111111111_1111111111111111_1110101110111000_1000111010010010"; -- -0.07921513501773339
	pesos_i(23081) := b"1111111111111111_1111111111111111_1110110001000101_1010110110110101"; -- -0.07706178989182914
	pesos_i(23082) := b"0000000000000000_0000000000000000_0000011101011010_1111000111101100"; -- 0.02873146078898159
	pesos_i(23083) := b"0000000000000000_0000000000000000_0001101110111101_0101001101000000"; -- 0.10835762316352585
	pesos_i(23084) := b"1111111111111111_1111111111111111_1110010101110010_1110100001110000"; -- -0.10371539361792745
	pesos_i(23085) := b"1111111111111111_1111111111111111_1110111110111000_0111110101000101"; -- -0.06359116617024894
	pesos_i(23086) := b"0000000000000000_0000000000000000_0001001001110011_1101101010011011"; -- 0.07208029055670666
	pesos_i(23087) := b"1111111111111111_1111111111111111_1111001101011001_1111010000001111"; -- -0.04940867081088602
	pesos_i(23088) := b"0000000000000000_0000000000000000_0000001011101111_1101011111100001"; -- 0.011472217963874475
	pesos_i(23089) := b"1111111111111111_1111111111111111_1111000100111001_0110101001001000"; -- -0.05771766418511462
	pesos_i(23090) := b"0000000000000000_0000000000000000_0001110110101000_0100111010101000"; -- 0.11584941495478547
	pesos_i(23091) := b"0000000000000000_0000000000000000_0001111010101001_1110010101101010"; -- 0.11977990938214451
	pesos_i(23092) := b"1111111111111111_1111111111111111_1111001000100010_1001111110101011"; -- -0.05415918422087543
	pesos_i(23093) := b"1111111111111111_1111111111111111_1111001100011010_0110000111001010"; -- -0.05037869291506069
	pesos_i(23094) := b"0000000000000000_0000000000000000_0010110000100111_1111111100001100"; -- 0.1724852948501863
	pesos_i(23095) := b"1111111111111111_1111111111111111_1110101110001100_1011100100011001"; -- -0.07988398694338443
	pesos_i(23096) := b"1111111111111111_1111111111111111_1101110011101011_0110001101110110"; -- -0.13703325633148838
	pesos_i(23097) := b"0000000000000000_0000000000000000_0001010011110101_0010110000100100"; -- 0.08186603436137113
	pesos_i(23098) := b"0000000000000000_0000000000000000_0000111100011110_0000011011111111"; -- 0.05905193056618766
	pesos_i(23099) := b"0000000000000000_0000000000000000_0010001000001101_0110001100011001"; -- 0.13301677091158967
	pesos_i(23100) := b"1111111111111111_1111111111111111_1111000001101111_1101101110001101"; -- -0.06079318812747312
	pesos_i(23101) := b"0000000000000000_0000000000000000_0000000110000111_1011111011100011"; -- 0.005977564371364925
	pesos_i(23102) := b"0000000000000000_0000000000000000_0001000010111111_0111100101111100"; -- 0.0654216697443518
	pesos_i(23103) := b"0000000000000000_0000000000000000_0010001110000000_0110101110111101"; -- 0.13867829663748424
	pesos_i(23104) := b"1111111111111111_1111111111111111_1101100010101001_0100010110001000"; -- -0.15366712027422774
	pesos_i(23105) := b"1111111111111111_1111111111111111_1111100011100101_1110100100011101"; -- -0.02774184277759429
	pesos_i(23106) := b"1111111111111111_1111111111111111_1110001100011011_1001010100011000"; -- -0.11286037593223411
	pesos_i(23107) := b"0000000000000000_0000000000000000_0000000110100101_1000110111101101"; -- 0.0064324096349759755
	pesos_i(23108) := b"1111111111111111_1111111111111111_1101111000101001_1011101100111111"; -- -0.1321757288592264
	pesos_i(23109) := b"1111111111111111_1111111111111111_1110100010010100_1010001111011110"; -- -0.09148193194097383
	pesos_i(23110) := b"1111111111111111_1111111111111111_1110011111000011_1010001100011101"; -- -0.094671063765558
	pesos_i(23111) := b"1111111111111111_1111111111111111_1111001110010110_0111000110011001"; -- -0.0484856607822447
	pesos_i(23112) := b"0000000000000000_0000000000000000_0010101111001100_1001000100010001"; -- 0.17109018966068518
	pesos_i(23113) := b"1111111111111111_1111111111111111_1110111001100010_0001000001100111"; -- -0.06881616110691963
	pesos_i(23114) := b"0000000000000000_0000000000000000_0001100000111110_1110010100110110"; -- 0.09470970687949028
	pesos_i(23115) := b"1111111111111111_1111111111111111_1110110101101101_1000011101010100"; -- -0.07254747581807937
	pesos_i(23116) := b"1111111111111111_1111111111111111_1101111111000111_1001010110100010"; -- -0.1258608322602171
	pesos_i(23117) := b"0000000000000000_0000000000000000_0001101111110101_1111010111110100"; -- 0.10922181331923574
	pesos_i(23118) := b"0000000000000000_0000000000000000_0000011100100100_0101011000010111"; -- 0.02789819779340987
	pesos_i(23119) := b"1111111111111111_1111111111111111_1110001010100100_1010011010000110"; -- -0.11467513299916433
	pesos_i(23120) := b"1111111111111111_1111111111111111_1101111110110111_0100011000001101"; -- -0.12610971614512448
	pesos_i(23121) := b"0000000000000000_0000000000000000_0001111101110001_1000110001110100"; -- 0.12282636489947502
	pesos_i(23122) := b"0000000000000000_0000000000000000_0000100111000000_1001101001010110"; -- 0.03809513661157508
	pesos_i(23123) := b"1111111111111111_1111111111111111_1110010101101011_1000011111101100"; -- -0.10382795791858328
	pesos_i(23124) := b"0000000000000000_0000000000000000_0000000111010100_1111111010100011"; -- 0.007156290716827945
	pesos_i(23125) := b"1111111111111111_1111111111111111_1111111110000101_0001000011111010"; -- -0.001875819176188453
	pesos_i(23126) := b"1111111111111111_1111111111111111_1110111001100011_0101100101110101"; -- -0.06879654783470365
	pesos_i(23127) := b"1111111111111111_1111111111111111_1111011011111101_1001001111001101"; -- -0.03519321679432283
	pesos_i(23128) := b"0000000000000000_0000000000000000_0001010111101011_0010110000100011"; -- 0.08561969618151004
	pesos_i(23129) := b"1111111111111111_1111111111111111_1101111010100111_0010011111111111"; -- -0.1302618982322647
	pesos_i(23130) := b"0000000000000000_0000000000000000_0010011010111110_0011101100101111"; -- 0.15134019747533248
	pesos_i(23131) := b"1111111111111111_1111111111111111_1110101001111100_1100000100000100"; -- -0.08403390561208604
	pesos_i(23132) := b"1111111111111111_1111111111111111_1111110000001010_1011111001111100"; -- -0.015461058288213357
	pesos_i(23133) := b"1111111111111111_1111111111111111_1111011010001110_1011000010001101"; -- -0.03688522880941704
	pesos_i(23134) := b"1111111111111111_1111111111111111_1101111000110010_1100111100011101"; -- -0.13203721559144338
	pesos_i(23135) := b"0000000000000000_0000000000000000_0000000000011100_1101100100010100"; -- 0.00044018493547123616
	pesos_i(23136) := b"1111111111111111_1111111111111111_1110010011101010_1101001111110100"; -- -0.1057918098906596
	pesos_i(23137) := b"1111111111111111_1111111111111111_1110111111011001_1100111100011111"; -- -0.06308274729232821
	pesos_i(23138) := b"1111111111111111_1111111111111111_1110101000110000_0000000100001110"; -- -0.08520501536193192
	pesos_i(23139) := b"1111111111111111_1111111111111111_1110000101100111_1001100110001100"; -- -0.11951294254474053
	pesos_i(23140) := b"1111111111111111_1111111111111111_1110010010100101_0011101100011010"; -- -0.10685377718742624
	pesos_i(23141) := b"0000000000000000_0000000000000000_0001010110100011_1101100111011111"; -- 0.08453141870622348
	pesos_i(23142) := b"0000000000000000_0000000000000000_0010001111011011_1010001100110101"; -- 0.14007015267668918
	pesos_i(23143) := b"0000000000000000_0000000000000000_0001011000111110_0001110111000110"; -- 0.086885319590034
	pesos_i(23144) := b"1111111111111111_1111111111111111_1110101100001001_1010110011100011"; -- -0.08188361599303111
	pesos_i(23145) := b"1111111111111111_1111111111111111_1111111111111001_0001001111101101"; -- -0.00010562392110533288
	pesos_i(23146) := b"1111111111111111_1111111111111111_1110001111101010_1010000100011001"; -- -0.10970109111606917
	pesos_i(23147) := b"1111111111111111_1111111111111111_1101011010100110_0010001100001111"; -- -0.1615274513851822
	pesos_i(23148) := b"0000000000000000_0000000000000000_0001001110010110_0100000111011111"; -- 0.07651149450077067
	pesos_i(23149) := b"1111111111111111_1111111111111111_1110001011100111_1001001101101111"; -- -0.11365393209531909
	pesos_i(23150) := b"1111111111111111_1111111111111111_1101110101011101_1110001110101110"; -- -0.1352861118306708
	pesos_i(23151) := b"1111111111111111_1111111111111111_1110110111010100_1001001001110001"; -- -0.07097515803032806
	pesos_i(23152) := b"0000000000000000_0000000000000000_0000000010000111_0010000100010001"; -- 0.0020619073239623114
	pesos_i(23153) := b"0000000000000000_0000000000000000_0000000011010110_1010110011011100"; -- 0.0032756841518501376
	pesos_i(23154) := b"1111111111111111_1111111111111111_1110111101000001_0010101100100110"; -- -0.0654118568783095
	pesos_i(23155) := b"1111111111111111_1111111111111111_1111001001010001_0110111100010010"; -- -0.053444917700728456
	pesos_i(23156) := b"1111111111111111_1111111111111111_1101100010000000_0000101000101000"; -- -0.15429626970771057
	pesos_i(23157) := b"1111111111111111_1111111111111111_1111010001011111_0011110010111100"; -- -0.04542179490248269
	pesos_i(23158) := b"0000000000000000_0000000000000000_0000011100011011_1000111010101000"; -- 0.02776424023255646
	pesos_i(23159) := b"1111111111111111_1111111111111111_1110111010001000_1011110110000000"; -- -0.068226009705504
	pesos_i(23160) := b"1111111111111111_1111111111111111_1111000000001000_1111000111110010"; -- -0.06236350850758825
	pesos_i(23161) := b"1111111111111111_1111111111111111_1110100011011100_0111101001011001"; -- -0.0903857740017258
	pesos_i(23162) := b"0000000000000000_0000000000000000_0000101000101110_0010111101000001"; -- 0.03976722082630057
	pesos_i(23163) := b"0000000000000000_0000000000000000_0001111010010011_1111101000111010"; -- 0.11944545661916363
	pesos_i(23164) := b"0000000000000000_0000000000000000_0001101001100101_1011011000110010"; -- 0.10311449730980969
	pesos_i(23165) := b"0000000000000000_0000000000000000_0000010011110010_1001001110101101"; -- 0.019326429207312583
	pesos_i(23166) := b"0000000000000000_0000000000000000_0000001001100001_0000101101001100"; -- 0.009293275777920539
	pesos_i(23167) := b"0000000000000000_0000000000000000_0010010001101100_0000001000110101"; -- 0.14227308069269082
	pesos_i(23168) := b"0000000000000000_0000000000000000_0001001000001010_0110110111010001"; -- 0.07047163345242478
	pesos_i(23169) := b"0000000000000000_0000000000000000_0000110111000111_1100111011101001"; -- 0.05383008174788241
	pesos_i(23170) := b"1111111111111111_1111111111111111_1110100101001101_1001001000000110"; -- -0.08866011953747084
	pesos_i(23171) := b"1111111111111111_1111111111111111_1110100001001010_0000110111111100"; -- -0.09262001612370883
	pesos_i(23172) := b"0000000000000000_0000000000000000_0000000100110001_0000000101110110"; -- 0.004654017824080486
	pesos_i(23173) := b"0000000000000000_0000000000000000_0001101111000010_1000000111101000"; -- 0.10843669812573965
	pesos_i(23174) := b"1111111111111111_1111111111111111_1111000000001010_1001110011111000"; -- -0.062338056069773384
	pesos_i(23175) := b"0000000000000000_0000000000000000_0000111011100000_1011111101110111"; -- 0.05811688096970584
	pesos_i(23176) := b"1111111111111111_1111111111111111_1110110111001101_0101110001010111"; -- -0.07108519437078234
	pesos_i(23177) := b"0000000000000000_0000000000000000_0000111001010101_0010111101111010"; -- 0.055987326839443644
	pesos_i(23178) := b"1111111111111111_1111111111111111_1110111101110000_1111100011011010"; -- -0.06468243301271812
	pesos_i(23179) := b"1111111111111111_1111111111111111_1101110110000100_1001010100000110"; -- -0.13469570745796913
	pesos_i(23180) := b"1111111111111111_1111111111111111_1101110110000001_1110101011100111"; -- -0.13473636502801808
	pesos_i(23181) := b"0000000000000000_0000000000000000_0001111111010010_1101011100111111"; -- 0.12431092542155203
	pesos_i(23182) := b"1111111111111111_1111111111111111_1110110000011000_0101000010011100"; -- -0.07775398425830798
	pesos_i(23183) := b"0000000000000000_0000000000000000_0010001010000011_0100010100001010"; -- 0.13481551645272088
	pesos_i(23184) := b"0000000000000000_0000000000000000_0000111011010000_1110001100010001"; -- 0.05787486225125841
	pesos_i(23185) := b"1111111111111111_1111111111111111_1101111110101011_1011000111000100"; -- -0.12628640145173867
	pesos_i(23186) := b"0000000000000000_0000000000000000_0010010101110100_0011100000100000"; -- 0.14630461491505262
	pesos_i(23187) := b"0000000000000000_0000000000000000_0001010011001010_1111101001111001"; -- 0.08122220467628839
	pesos_i(23188) := b"1111111111111111_1111111111111111_1111011011111111_1010111101001010"; -- -0.03516106070807678
	pesos_i(23189) := b"0000000000000000_0000000000000000_0001010100101010_0111011100110110"; -- 0.08267922476252788
	pesos_i(23190) := b"0000000000000000_0000000000000000_0000101110110110_1011100111001100"; -- 0.04575692407251771
	pesos_i(23191) := b"1111111111111111_1111111111111111_1111101011100111_0001011100000001"; -- -0.01991134857117704
	pesos_i(23192) := b"1111111111111111_1111111111111111_1111101100000010_0010011001011100"; -- -0.019498445983626204
	pesos_i(23193) := b"0000000000000000_0000000000000000_0001001001010010_0011010010010011"; -- 0.0715668544349686
	pesos_i(23194) := b"1111111111111111_1111111111111111_1111111000101110_1000110110110110"; -- -0.0071021491078394105
	pesos_i(23195) := b"1111111111111111_1111111111111111_1110000111001100_1011110111011010"; -- -0.11796964104122207
	pesos_i(23196) := b"1111111111111111_1111111111111111_1111111111100111_1001000101001000"; -- -0.00037281029784546195
	pesos_i(23197) := b"0000000000000000_0000000000000000_0001010110101101_0000010111011001"; -- 0.0846713689454345
	pesos_i(23198) := b"0000000000000000_0000000000000000_0000000000001010_0011010101110011"; -- 0.00015577376786270468
	pesos_i(23199) := b"0000000000000000_0000000000000000_0000111110000001_0110110011000101"; -- 0.06056861698492497
	pesos_i(23200) := b"1111111111111111_1111111111111111_1110101110101011_1011100111100011"; -- -0.07941091746940254
	pesos_i(23201) := b"1111111111111111_1111111111111111_1110110010101111_1100110001000001"; -- -0.07544253742016631
	pesos_i(23202) := b"0000000000000000_0000000000000000_0000110000000010_1000110110010000"; -- 0.04691395525041724
	pesos_i(23203) := b"1111111111111111_1111111111111111_1111100111010110_0101001100000000"; -- -0.024073421931280096
	pesos_i(23204) := b"0000000000000000_0000000000000000_0000110100100110_0100101101001011"; -- 0.05136557173685328
	pesos_i(23205) := b"0000000000000000_0000000000000000_0001100111111010_0111011001011110"; -- 0.10147800241975946
	pesos_i(23206) := b"1111111111111111_1111111111111111_1110011011100010_0011110001100000"; -- -0.09811041503715236
	pesos_i(23207) := b"1111111111111111_1111111111111111_1111010001111001_0000001001110111"; -- -0.04502853965551955
	pesos_i(23208) := b"1111111111111111_1111111111111111_1110110000011110_0110000001011110"; -- -0.07766149247355629
	pesos_i(23209) := b"0000000000000000_0000000000000000_0001111100001011_0000101010001101"; -- 0.12126222556777712
	pesos_i(23210) := b"0000000000000000_0000000000000000_0000110101101110_1101100001010001"; -- 0.052472610164172935
	pesos_i(23211) := b"0000000000000000_0000000000000000_0000100000100100_0101100111100000"; -- 0.03180467345612907
	pesos_i(23212) := b"0000000000000000_0000000000000000_0001011000010010_1100100101010100"; -- 0.08622415835833845
	pesos_i(23213) := b"0000000000000000_0000000000000000_0010000101100100_0101111011110100"; -- 0.13043778865928032
	pesos_i(23214) := b"0000000000000000_0000000000000000_0000101111011010_0111110011010110"; -- 0.04630260684211433
	pesos_i(23215) := b"0000000000000000_0000000000000000_0000100100001010_0100101001010110"; -- 0.035313268763592365
	pesos_i(23216) := b"0000000000000000_0000000000000000_0001101101111010_0010111001111011"; -- 0.107333092752073
	pesos_i(23217) := b"1111111111111111_1111111111111111_1111011010101010_1010001111110100"; -- -0.0364587334291388
	pesos_i(23218) := b"1111111111111111_1111111111111111_1110011000001100_0000100011111010"; -- -0.10137885944969002
	pesos_i(23219) := b"0000000000000000_0000000000000000_0010010000110010_1011111000011010"; -- 0.14139927045361644
	pesos_i(23220) := b"1111111111111111_1111111111111111_1111100110110010_0100001011100100"; -- -0.024623698450609986
	pesos_i(23221) := b"0000000000000000_0000000000000000_0001100011110010_0111100000010110"; -- 0.0974497846081843
	pesos_i(23222) := b"1111111111111111_1111111111111111_1101011000101001_0111000001011011"; -- -0.16343019276568863
	pesos_i(23223) := b"0000000000000000_0000000000000000_0001011110110000_0011110001010100"; -- 0.09253289267012497
	pesos_i(23224) := b"0000000000000000_0000000000000000_0001001101001011_0011010111000110"; -- 0.07536636433573426
	pesos_i(23225) := b"1111111111111111_1111111111111111_1111000011101100_1101111001111100"; -- -0.05888566472453368
	pesos_i(23226) := b"1111111111111111_1111111111111111_1110100001001111_0000001111100111"; -- -0.09254432299734554
	pesos_i(23227) := b"1111111111111111_1111111111111111_1110101010110010_0011001101000100"; -- -0.08321837986199412
	pesos_i(23228) := b"1111111111111111_1111111111111111_1110001000001010_1010011000001100"; -- -0.11702501484507057
	pesos_i(23229) := b"1111111111111111_1111111111111111_1111111001110011_1101101100101011"; -- -0.0060446757197053945
	pesos_i(23230) := b"1111111111111111_1111111111111111_1110100110000101_0001011010110010"; -- -0.08781297827813342
	pesos_i(23231) := b"1111111111111111_1111111111111111_1101100110000100_1010010001000000"; -- -0.1503197997322454
	pesos_i(23232) := b"0000000000000000_0000000000000000_0001001010100000_0100101110101100"; -- 0.072758416749949
	pesos_i(23233) := b"1111111111111111_1111111111111111_1111110001011110_1110110011101111"; -- -0.01417655158588811
	pesos_i(23234) := b"1111111111111111_1111111111111111_1111001111001001_1001010110110000"; -- -0.047705311371341284
	pesos_i(23235) := b"0000000000000000_0000000000000000_0000100011100000_1010000000101010"; -- 0.03467751529647212
	pesos_i(23236) := b"1111111111111111_1111111111111111_1111100100101100_1110001110101011"; -- -0.02665879329382994
	pesos_i(23237) := b"1111111111111111_1111111111111111_1111001100101101_0001100101000011"; -- -0.05009309867411795
	pesos_i(23238) := b"0000000000000000_0000000000000000_0001101010011100_0110111010101011"; -- 0.10394946733109492
	pesos_i(23239) := b"1111111111111111_1111111111111111_1111010111110111_1110000000010110"; -- -0.039186472616095154
	pesos_i(23240) := b"0000000000000000_0000000000000000_0000000001011111_0000101000001000"; -- 0.0014501827981140913
	pesos_i(23241) := b"0000000000000000_0000000000000000_0001111110010100_0001100111000001"; -- 0.12335358583432811
	pesos_i(23242) := b"0000000000000000_0000000000000000_0000000011100111_1011111010010111"; -- 0.003536140315987712
	pesos_i(23243) := b"1111111111111111_1111111111111111_1110100101001111_0000111100110111"; -- -0.08863739871201386
	pesos_i(23244) := b"0000000000000000_0000000000000000_0010001110000100_0110001110011100"; -- 0.13873884741137216
	pesos_i(23245) := b"0000000000000000_0000000000000000_0001100010111110_1110001011000100"; -- 0.09666268620505766
	pesos_i(23246) := b"1111111111111111_1111111111111111_1111100001011101_1111101000000111"; -- -0.029816029710803858
	pesos_i(23247) := b"0000000000000000_0000000000000000_0001111111111101_1111101010001001"; -- 0.12496915660119906
	pesos_i(23248) := b"1111111111111111_1111111111111111_1101011111101100_0100000001101011"; -- -0.15655133628318532
	pesos_i(23249) := b"0000000000000000_0000000000000000_0010000110010011_0001101010001010"; -- 0.1311508739070879
	pesos_i(23250) := b"0000000000000000_0000000000000000_0001111110000001_1111100100011001"; -- 0.12307698117342271
	pesos_i(23251) := b"0000000000000000_0000000000000000_0000010010011111_0100101010010010"; -- 0.018055592204951027
	pesos_i(23252) := b"0000000000000000_0000000000000000_0000001001110100_1111001110100011"; -- 0.009597041378127502
	pesos_i(23253) := b"0000000000000000_0000000000000000_0001000001101001_1110000001010000"; -- 0.0641155429797033
	pesos_i(23254) := b"0000000000000000_0000000000000000_0000000101100001_0110101001101100"; -- 0.0053926956867600346
	pesos_i(23255) := b"1111111111111111_1111111111111111_1111001111010011_0001101000101101"; -- -0.04756008533932557
	pesos_i(23256) := b"1111111111111111_1111111111111111_1110011101111001_1001110110100101"; -- -0.0958005400991739
	pesos_i(23257) := b"1111111111111111_1111111111111111_1110001010001010_1001001101011110"; -- -0.11507300344261838
	pesos_i(23258) := b"1111111111111111_1111111111111111_1110010001101101_0100001101100101"; -- -0.10770777498592943
	pesos_i(23259) := b"0000000000000000_0000000000000000_0010001001000101_1110011101010100"; -- 0.13387914476814908
	pesos_i(23260) := b"0000000000000000_0000000000000000_0001000000001000_0000001000001010"; -- 0.06262219178700344
	pesos_i(23261) := b"1111111111111111_1111111111111111_1111111111101000_1010010110011010"; -- -0.0003563403353521978
	pesos_i(23262) := b"1111111111111111_1111111111111111_1110011111100100_1110011010101100"; -- -0.09416349693711258
	pesos_i(23263) := b"1111111111111111_1111111111111111_1111001010010111_1100011111010101"; -- -0.05237151202802911
	pesos_i(23264) := b"1111111111111111_1111111111111111_1111100111101110_1101011011001111"; -- -0.023699354687650418
	pesos_i(23265) := b"1111111111111111_1111111111111111_1110001110011000_0000011110010111"; -- -0.11096146173265982
	pesos_i(23266) := b"0000000000000000_0000000000000000_0001100110010110_1101001011100010"; -- 0.09995763787690234
	pesos_i(23267) := b"0000000000000000_0000000000000000_0001001011101110_1000011100100101"; -- 0.07395214708721605
	pesos_i(23268) := b"0000000000000000_0000000000000000_0001111011101000_0011100100101111"; -- 0.12073094755872733
	pesos_i(23269) := b"1111111111111111_1111111111111111_1111001111010100_0010100001011100"; -- -0.0475439810445257
	pesos_i(23270) := b"1111111111111111_1111111111111111_1111001111000011_1011001010000110"; -- -0.047795145342947716
	pesos_i(23271) := b"0000000000000000_0000000000000000_0000101001111001_0010011111100101"; -- 0.04091119126642011
	pesos_i(23272) := b"0000000000000000_0000000000000000_0000000001111010_1111101011101100"; -- 0.0018765283826467948
	pesos_i(23273) := b"0000000000000000_0000000000000000_0000110111110001_0110001100101110"; -- 0.054464529653634394
	pesos_i(23274) := b"1111111111111111_1111111111111111_1111001001001001_1111111111100111"; -- -0.053558355331928355
	pesos_i(23275) := b"1111111111111111_1111111111111111_1101111011001110_1001100110101101"; -- -0.12966002965222406
	pesos_i(23276) := b"1111111111111111_1111111111111111_1111100000100010_0010010010011100"; -- -0.030729019125499784
	pesos_i(23277) := b"0000000000000000_0000000000000000_0000100111001101_1100001111100101"; -- 0.03829597806510846
	pesos_i(23278) := b"0000000000000000_0000000000000000_0001111001011101_0100000101011100"; -- 0.11861046308689523
	pesos_i(23279) := b"1111111111111111_1111111111111111_1111011001000011_1101000101111110"; -- -0.03802767448588645
	pesos_i(23280) := b"1111111111111111_1111111111111111_1111101110100000_1010100010110011"; -- -0.01707978855690375
	pesos_i(23281) := b"1111111111111111_1111111111111111_1110111111101000_1000110110011110"; -- -0.06285776998755536
	pesos_i(23282) := b"1111111111111111_1111111111111111_1111111111110010_1100101101100101"; -- -0.00020149976368233173
	pesos_i(23283) := b"1111111111111111_1111111111111111_1110111011100100_1111101001100100"; -- -0.06681857159746936
	pesos_i(23284) := b"1111111111111111_1111111111111111_1111110011011010_1100111000001000"; -- -0.012286303676287143
	pesos_i(23285) := b"0000000000000000_0000000000000000_0000001101100000_1011010001011001"; -- 0.013194343244430076
	pesos_i(23286) := b"1111111111111111_1111111111111111_1111111001001111_1110001111110011"; -- -0.006593468878005826
	pesos_i(23287) := b"1111111111111111_1111111111111111_1111001011101001_1111110100010011"; -- -0.05111711768706024
	pesos_i(23288) := b"1111111111111111_1111111111111111_1111000011110111_1010010100111010"; -- -0.05872123084923256
	pesos_i(23289) := b"1111111111111111_1111111111111111_1111000111000001_1011101011110001"; -- -0.05563766114478736
	pesos_i(23290) := b"1111111111111111_1111111111111111_1111101010111011_1110010010011110"; -- -0.020570479890213593
	pesos_i(23291) := b"1111111111111111_1111111111111111_1110010110100001_1110010100001001"; -- -0.10299843343723629
	pesos_i(23292) := b"0000000000000000_0000000000000000_0000101000101000_0000011000100101"; -- 0.03967321773112451
	pesos_i(23293) := b"1111111111111111_1111111111111111_1111100001100111_1001001110000100"; -- -0.029669552038148247
	pesos_i(23294) := b"0000000000000000_0000000000000000_0000100010000101_0100011111011001"; -- 0.03328370150351559
	pesos_i(23295) := b"0000000000000000_0000000000000000_0000110110100011_1010000101010001"; -- 0.05327804782665286
	pesos_i(23296) := b"0000000000000000_0000000000000000_0001010101010001_0110011111011101"; -- 0.08327340275179985
	pesos_i(23297) := b"1111111111111111_1111111111111111_1111101110000110_1101100110111001"; -- -0.017473594923874017
	pesos_i(23298) := b"0000000000000000_0000000000000000_0001111000000001_1011000110000000"; -- 0.11721333867365341
	pesos_i(23299) := b"1111111111111111_1111111111111111_1111010100100111_0000000001101001"; -- -0.04237363281044543
	pesos_i(23300) := b"1111111111111111_1111111111111111_1101111111100101_1010110010101000"; -- -0.12540169611708155
	pesos_i(23301) := b"0000000000000000_0000000000000000_0000001001100001_0101011101111001"; -- 0.00929781621305369
	pesos_i(23302) := b"0000000000000000_0000000000000000_0001000111010100_0010101110110010"; -- 0.06964371780577486
	pesos_i(23303) := b"0000000000000000_0000000000000000_0000110001111011_0110110011101110"; -- 0.048758323687777834
	pesos_i(23304) := b"1111111111111111_1111111111111111_1110101110010011_1001001110010110"; -- -0.0797794112810216
	pesos_i(23305) := b"0000000000000000_0000000000000000_0001101000000101_1010111101000011"; -- 0.1016492403460206
	pesos_i(23306) := b"0000000000000000_0000000000000000_0001101110101011_1101010100010111"; -- 0.10809070398478919
	pesos_i(23307) := b"1111111111111111_1111111111111111_1111111111011011_1000110001101001"; -- -0.0005562060981422229
	pesos_i(23308) := b"0000000000000000_0000000000000000_0001001101101111_1110011001111010"; -- 0.07592621311583507
	pesos_i(23309) := b"0000000000000000_0000000000000000_0001101111110001_1100000100110111"; -- 0.10915763469537576
	pesos_i(23310) := b"0000000000000000_0000000000000000_0000010011111000_0111000010111010"; -- 0.01941589872506283
	pesos_i(23311) := b"0000000000000000_0000000000000000_0010010001000100_1101011000111101"; -- 0.14167536715202925
	pesos_i(23312) := b"0000000000000000_0000000000000000_0001100111101010_1000011001111100"; -- 0.10123482261910234
	pesos_i(23313) := b"1111111111111111_1111111111111111_1111111100011110_0010011001010011"; -- -0.0034462020919224837
	pesos_i(23314) := b"1111111111111111_1111111111111111_1110111000101010_0101100010111100"; -- -0.06966634191945362
	pesos_i(23315) := b"1111111111111111_1111111111111111_1111101111111100_1100000010000100"; -- -0.015674560272586204
	pesos_i(23316) := b"0000000000000000_0000000000000000_0000111110011110_1101000001111100"; -- 0.06101706541354123
	pesos_i(23317) := b"0000000000000000_0000000000000000_0001000111111011_1111000000011110"; -- 0.07025051826462224
	pesos_i(23318) := b"0000000000000000_0000000000000000_0010100001111100_0010100011100101"; -- 0.15814452744495505
	pesos_i(23319) := b"1111111111111111_1111111111111111_1110111011011111_0000100100000000"; -- -0.06690925363326526
	pesos_i(23320) := b"0000000000000000_0000000000000000_0000011100110000_0110100101101111"; -- 0.028082456102841265
	pesos_i(23321) := b"0000000000000000_0000000000000000_0000111001110110_1101110010111000"; -- 0.05650119291644873
	pesos_i(23322) := b"0000000000000000_0000000000000000_0000110000011101_0011001011110100"; -- 0.04732054197744953
	pesos_i(23323) := b"0000000000000000_0000000000000000_0001001001110010_1010001001101101"; -- 0.07206168327292052
	pesos_i(23324) := b"1111111111111111_1111111111111111_1110111100111100_0011111100001011"; -- -0.06548696497000984
	pesos_i(23325) := b"0000000000000000_0000000000000000_0010001001100000_0110100010011111"; -- 0.13428357974067362
	pesos_i(23326) := b"0000000000000000_0000000000000000_0001100110110100_1111100100001101"; -- 0.10041767662706819
	pesos_i(23327) := b"1111111111111111_1111111111111111_1101110011011000_0011001101111101"; -- -0.13732603253276815
	pesos_i(23328) := b"0000000000000000_0000000000000000_0001100000111111_0000100101011001"; -- 0.09471186098147312
	pesos_i(23329) := b"0000000000000000_0000000000000000_0010001011010001_1101000000100110"; -- 0.13601399349165322
	pesos_i(23330) := b"0000000000000000_0000000000000000_0010010111010000_1101110010001110"; -- 0.14771822420357072
	pesos_i(23331) := b"1111111111111111_1111111111111111_1110010111010100_1111100110010101"; -- -0.10221901056270845
	pesos_i(23332) := b"1111111111111111_1111111111111111_1110000001111000_0110100010000111"; -- -0.12316271490757412
	pesos_i(23333) := b"0000000000000000_0000000000000000_0000010110101110_1010011000110111"; -- 0.02219618639330338
	pesos_i(23334) := b"0000000000000000_0000000000000000_0001010110111000_0011110010010111"; -- 0.08484247853878504
	pesos_i(23335) := b"0000000000000000_0000000000000000_0001000000110101_0001000100101000"; -- 0.06330973847301692
	pesos_i(23336) := b"1111111111111111_1111111111111111_1111000011110110_1101000001100011"; -- -0.058733917087231115
	pesos_i(23337) := b"0000000000000000_0000000000000000_0000011001001110_0111100011110100"; -- 0.024634894883794823
	pesos_i(23338) := b"1111111111111111_1111111111111111_1110000110100110_0011011011100110"; -- -0.11855751877077274
	pesos_i(23339) := b"0000000000000000_0000000000000000_0000111010010010_0000011100111110"; -- 0.05691571480077494
	pesos_i(23340) := b"1111111111111111_1111111111111111_1111010010010110_1001110000001010"; -- -0.0445768811023347
	pesos_i(23341) := b"1111111111111111_1111111111111111_1110010010010010_0101001110010000"; -- -0.10714223608576955
	pesos_i(23342) := b"1111111111111111_1111111111111111_1110111110000010_1001000010100110"; -- -0.06441398572577711
	pesos_i(23343) := b"1111111111111111_1111111111111111_1110101011111110_1011110111011010"; -- -0.08205045159939793
	pesos_i(23344) := b"0000000000000000_0000000000000000_0000111010110010_1001111000001101"; -- 0.057412985039643365
	pesos_i(23345) := b"0000000000000000_0000000000000000_0000011010111011_0001101001101001"; -- 0.026292467646259796
	pesos_i(23346) := b"0000000000000000_0000000000000000_0001011011101101_0111010110011001"; -- 0.08956084239704108
	pesos_i(23347) := b"1111111111111111_1111111111111111_1101111000100111_0110011000000000"; -- -0.13221132760168883
	pesos_i(23348) := b"1111111111111111_1111111111111111_1111010011110000_0101000001111111"; -- -0.043208092703775056
	pesos_i(23349) := b"1111111111111111_1111111111111111_1101110101111101_1010001100110000"; -- -0.13480167463273343
	pesos_i(23350) := b"1111111111111111_1111111111111111_1111100111110001_0001100000101000"; -- -0.023664942061338227
	pesos_i(23351) := b"0000000000000000_0000000000000000_0010001011100011_0000100010110010"; -- 0.13627676341793082
	pesos_i(23352) := b"0000000000000000_0000000000000000_0001100110011111_0100000001010010"; -- 0.10008623113967334
	pesos_i(23353) := b"0000000000000000_0000000000000000_0001011100010100_1101011100110001"; -- 0.09016175221991982
	pesos_i(23354) := b"1111111111111111_1111111111111111_1111110010110011_1101100011011000"; -- -0.012880751941437858
	pesos_i(23355) := b"1111111111111111_1111111111111111_1110100101111000_1100100011001101"; -- -0.08800072670907193
	pesos_i(23356) := b"0000000000000000_0000000000000000_0000000111010101_0000010100010110"; -- 0.007156675147496643
	pesos_i(23357) := b"1111111111111111_1111111111111111_1110100101110101_1110001011000100"; -- -0.0880449553350687
	pesos_i(23358) := b"0000000000000000_0000000000000000_0000011110001001_1010001100001010"; -- 0.029443921952141915
	pesos_i(23359) := b"1111111111111111_1111111111111111_1111101011011010_0110001101101011"; -- -0.020105158102668698
	pesos_i(23360) := b"1111111111111111_1111111111111111_1110010000001111_0100000011010010"; -- -0.10914225454256489
	pesos_i(23361) := b"0000000000000000_0000000000000000_0000111100010010_0100111101101011"; -- 0.05887314193733895
	pesos_i(23362) := b"0000000000000000_0000000000000000_0001110000011001_0101000001010100"; -- 0.10976125759242923
	pesos_i(23363) := b"1111111111111111_1111111111111111_1110011101101110_0110111000110010"; -- -0.09597121506584891
	pesos_i(23364) := b"0000000000000000_0000000000000000_0001011010000000_0110010100010100"; -- 0.0878966498229862
	pesos_i(23365) := b"1111111111111111_1111111111111111_1101100011111100_1101111001100011"; -- -0.15239152986674415
	pesos_i(23366) := b"1111111111111111_1111111111111111_1101011111010011_0000011100110011"; -- -0.15693621632870158
	pesos_i(23367) := b"1111111111111111_1111111111111111_1111010100000110_1100011011110101"; -- -0.04286533842410592
	pesos_i(23368) := b"0000000000000000_0000000000000000_0000111011011011_1000010010001101"; -- 0.058037075553196045
	pesos_i(23369) := b"0000000000000000_0000000000000000_0000111101000111_1101110101011001"; -- 0.05969031740577544
	pesos_i(23370) := b"1111111111111111_1111111111111111_1111111011011111_1000111001101010"; -- -0.004401301541126705
	pesos_i(23371) := b"1111111111111111_1111111111111111_1111011101010011_1010110110001001"; -- -0.0338794271001432
	pesos_i(23372) := b"0000000000000000_0000000000000000_0010001110111001_1011111001111110"; -- 0.13955298030178265
	pesos_i(23373) := b"0000000000000000_0000000000000000_0010011100010110_0111010111111001"; -- 0.1526864751407347
	pesos_i(23374) := b"1111111111111111_1111111111111111_1111001111111110_1110100001110101"; -- -0.04689166202714406
	pesos_i(23375) := b"0000000000000000_0000000000000000_0000010011010011_1001001110010000"; -- 0.01885339993018244
	pesos_i(23376) := b"1111111111111111_1111111111111111_1110100000110010_1111101011010110"; -- -0.09297210957112183
	pesos_i(23377) := b"0000000000000000_0000000000000000_0001111000011011_0111011101110100"; -- 0.11760660737689438
	pesos_i(23378) := b"0000000000000000_0000000000000000_0000001000101001_0100100000001000"; -- 0.008442403841963621
	pesos_i(23379) := b"0000000000000000_0000000000000000_0000011101011100_0101101111010111"; -- 0.028753032719690742
	pesos_i(23380) := b"0000000000000000_0000000000000000_0000111100101010_0010011110110011"; -- 0.059236985467492745
	pesos_i(23381) := b"1111111111111111_1111111111111111_1101110011100110_1001101001010000"; -- -0.1371062808459911
	pesos_i(23382) := b"0000000000000000_0000000000000000_0000111001000000_0101011110000100"; -- 0.05566927886222277
	pesos_i(23383) := b"0000000000000000_0000000000000000_0010001100001110_0001011111010100"; -- 0.136933793347581
	pesos_i(23384) := b"0000000000000000_0000000000000000_0001101101000100_0100100001111011"; -- 0.1065106678706881
	pesos_i(23385) := b"1111111111111111_1111111111111111_1111010101110101_0101110000100101"; -- -0.04117797946460472
	pesos_i(23386) := b"0000000000000000_0000000000000000_0000111100000110_1111001010001110"; -- 0.05869976002022581
	pesos_i(23387) := b"0000000000000000_0000000000000000_0000100000011000_0000011000011000"; -- 0.03161657415469651
	pesos_i(23388) := b"0000000000000000_0000000000000000_0001001111111010_1111100110111000"; -- 0.07804833176355429
	pesos_i(23389) := b"0000000000000000_0000000000000000_0010000101011100_0111000011101011"; -- 0.13031678894520576
	pesos_i(23390) := b"1111111111111111_1111111111111111_1101100111000000_1010000000000101"; -- -0.14940452455038672
	pesos_i(23391) := b"1111111111111111_1111111111111111_1110111010011001_1110110111010100"; -- -0.06796372954067276
	pesos_i(23392) := b"0000000000000000_0000000000000000_0010001010111001_0110011110101101"; -- 0.13564155548726015
	pesos_i(23393) := b"1111111111111111_1111111111111111_1110011000010110_1110001001011011"; -- -0.10121331474205114
	pesos_i(23394) := b"1111111111111111_1111111111111111_1110010101010110_0000000001000110"; -- -0.10415647783526037
	pesos_i(23395) := b"0000000000000000_0000000000000000_0000011010010111_1100100001000100"; -- 0.025753513845958666
	pesos_i(23396) := b"1111111111111111_1111111111111111_1111101100011111_1010001001010011"; -- -0.01904855223079512
	pesos_i(23397) := b"1111111111111111_1111111111111111_1101100110100100_0010011010011010"; -- -0.14983900783033957
	pesos_i(23398) := b"1111111111111111_1111111111111111_1111111010001010_0000111101100010"; -- -0.005705870126532847
	pesos_i(23399) := b"0000000000000000_0000000000000000_0001010110000011_1101101101110110"; -- 0.08404323215775668
	pesos_i(23400) := b"0000000000000000_0000000000000000_0000110001011000_1011100011010000"; -- 0.04822878920903927
	pesos_i(23401) := b"0000000000000000_0000000000000000_0000010011101100_0100110001111000"; -- 0.019230632110157103
	pesos_i(23402) := b"0000000000000000_0000000000000000_0001100000110101_1111011101010010"; -- 0.094573457188844
	pesos_i(23403) := b"1111111111111111_1111111111111111_1111110111000111_0001010100100100"; -- -0.008680990905772162
	pesos_i(23404) := b"0000000000000000_0000000000000000_0010001110001001_1110101101100011"; -- 0.1388232343538829
	pesos_i(23405) := b"1111111111111111_1111111111111111_1110000011111100_0110010100101111"; -- -0.12114875403865909
	pesos_i(23406) := b"0000000000000000_0000000000000000_0000010100001000_0010001000110000"; -- 0.019655358051799274
	pesos_i(23407) := b"0000000000000000_0000000000000000_0000010010110110_0011100111010000"; -- 0.018405545423575774
	pesos_i(23408) := b"1111111111111111_1111111111111111_1110111110011101_1011111001010000"; -- -0.06399927664614163
	pesos_i(23409) := b"1111111111111111_1111111111111111_1110110110101011_1011101100100100"; -- -0.07159834252654686
	pesos_i(23410) := b"1111111111111111_1111111111111111_1101100101011001_0010111010011000"; -- -0.15098294064868584
	pesos_i(23411) := b"0000000000000000_0000000000000000_0010000101011111_0100011011010111"; -- 0.13036005731359523
	pesos_i(23412) := b"0000000000000000_0000000000000000_0000100101110000_0001101000101111"; -- 0.03686679507603123
	pesos_i(23413) := b"0000000000000000_0000000000000000_0001100011110010_1011011001111110"; -- 0.09745350439317486
	pesos_i(23414) := b"0000000000000000_0000000000000000_0010011101011001_0000101110000101"; -- 0.15370246890772082
	pesos_i(23415) := b"0000000000000000_0000000000000000_0000000011000010_1000111000011011"; -- 0.002968675191263246
	pesos_i(23416) := b"0000000000000000_0000000000000000_0001011110000000_0010011100000101"; -- 0.09179920063013979
	pesos_i(23417) := b"1111111111111111_1111111111111111_1111000011101111_1101111100011000"; -- -0.058839852072830635
	pesos_i(23418) := b"0000000000000000_0000000000000000_0000100101011000_0101111010101000"; -- 0.03650466527465978
	pesos_i(23419) := b"0000000000000000_0000000000000000_0000110100010000_1110110010110111"; -- 0.0510394998144094
	pesos_i(23420) := b"1111111111111111_1111111111111111_1101110001001011_1100001010111110"; -- -0.13946898322090295
	pesos_i(23421) := b"1111111111111111_1111111111111111_1111100111110010_0111110100101000"; -- -0.02364366323763315
	pesos_i(23422) := b"0000000000000000_0000000000000000_0001110000111001_0000101000100110"; -- 0.11024535586124444
	pesos_i(23423) := b"0000000000000000_0000000000000000_0000000111111001_1110011110010100"; -- 0.007719491582882763
	pesos_i(23424) := b"1111111111111111_1111111111111111_1111111000001010_0101011001010000"; -- -0.007654767484071038
	pesos_i(23425) := b"1111111111111111_1111111111111111_1110101001010100_1111010010011001"; -- -0.08464118261323483
	pesos_i(23426) := b"0000000000000000_0000000000000000_0000111000001101_0101100000011010"; -- 0.05489111562737005
	pesos_i(23427) := b"0000000000000000_0000000000000000_0000101101001111_1100001110001111"; -- 0.044185850570506086
	pesos_i(23428) := b"0000000000000000_0000000000000000_0001110001111100_0010100001110101"; -- 0.11126950133625454
	pesos_i(23429) := b"1111111111111111_1111111111111111_1111011000111011_1110111010110101"; -- -0.03814800336790947
	pesos_i(23430) := b"1111111111111111_1111111111111111_1101110110110000_1011011010110010"; -- -0.13402231352934102
	pesos_i(23431) := b"0000000000000000_0000000000000000_0000000101001000_1110001110110001"; -- 0.00501845428802954
	pesos_i(23432) := b"0000000000000000_0000000000000000_0000111001010100_1101110110111100"; -- 0.05598245479587095
	pesos_i(23433) := b"1111111111111111_1111111111111111_1101101101100110_1010001101100110"; -- -0.14296511425734176
	pesos_i(23434) := b"1111111111111111_1111111111111111_1111010110011110_1101101001000110"; -- -0.040544851224245476
	pesos_i(23435) := b"1111111111111111_1111111111111111_1111011100011010_0000001011001101"; -- -0.03475935460518269
	pesos_i(23436) := b"0000000000000000_0000000000000000_0010001110110011_1010111100010010"; -- 0.13946050822757158
	pesos_i(23437) := b"0000000000000000_0000000000000000_0001000111001010_0101101010000010"; -- 0.06949391999480453
	pesos_i(23438) := b"1111111111111111_1111111111111111_1111110010010001_0100011110100100"; -- -0.013408205558976146
	pesos_i(23439) := b"0000000000000000_0000000000000000_0000100000000010_1010000000100000"; -- 0.0312900617294395
	pesos_i(23440) := b"0000000000000000_0000000000000000_0001010100011100_1110111000111010"; -- 0.082472695612023
	pesos_i(23441) := b"1111111111111111_1111111111111111_1111111110001111_1101010111001000"; -- -0.0017115007982824316
	pesos_i(23442) := b"1111111111111111_1111111111111111_1111110100011001_0101000101100001"; -- -0.0113324296138332
	pesos_i(23443) := b"0000000000000000_0000000000000000_0000010000010011_1111100101100101"; -- 0.01592978211415506
	pesos_i(23444) := b"1111111111111111_1111111111111111_1110010010101100_0110011101011100"; -- -0.10674432754569771
	pesos_i(23445) := b"1111111111111111_1111111111111111_1101111001001001_1000100000011011"; -- -0.1316904959007737
	pesos_i(23446) := b"0000000000000000_0000000000000000_0010011111011101_1011000010001010"; -- 0.15572646485283956
	pesos_i(23447) := b"0000000000000000_0000000000000000_0010011010001001_0101100110100000"; -- 0.15053329619641428
	pesos_i(23448) := b"0000000000000000_0000000000000000_0001000100110000_1010111110011010"; -- 0.0671491386247617
	pesos_i(23449) := b"0000000000000000_0000000000000000_0000100101010000_1110010010101011"; -- 0.03639058287618384
	pesos_i(23450) := b"1111111111111111_1111111111111111_1110110101100101_0100010010100100"; -- -0.07267352090897947
	pesos_i(23451) := b"0000000000000000_0000000000000000_0001011100100101_0110000000001001"; -- 0.09041404935535893
	pesos_i(23452) := b"0000000000000000_0000000000000000_0000000010011011_0001010011011100"; -- 0.0023663556255292505
	pesos_i(23453) := b"0000000000000000_0000000000000000_0000100100001111_0000010111000011"; -- 0.035385475213979584
	pesos_i(23454) := b"0000000000000000_0000000000000000_0001010011100111_0011000101110000"; -- 0.08165272700974813
	pesos_i(23455) := b"1111111111111111_1111111111111111_1110000010101000_0010010101011000"; -- -0.12243429746819652
	pesos_i(23456) := b"1111111111111111_1111111111111111_1110000100111111_1001010111100011"; -- -0.12012351223114193
	pesos_i(23457) := b"1111111111111111_1111111111111111_1111111000000001_1000001010100110"; -- -0.007789454043971994
	pesos_i(23458) := b"1111111111111111_1111111111111111_1110111111001101_1001100010100111"; -- -0.0632690995392911
	pesos_i(23459) := b"0000000000000000_0000000000000000_0001101011000111_0111111111101001"; -- 0.10460662301886994
	pesos_i(23460) := b"0000000000000000_0000000000000000_0000101000001000_1111111100001000"; -- 0.039199771296724674
	pesos_i(23461) := b"0000000000000000_0000000000000000_0001101110011111_1001001010111101"; -- 0.10790364383080447
	pesos_i(23462) := b"1111111111111111_1111111111111111_1110101100000000_1011001010000110"; -- -0.08202060923091783
	pesos_i(23463) := b"1111111111111111_1111111111111111_1110000110000100_1000101101111101"; -- -0.11907127566058699
	pesos_i(23464) := b"0000000000000000_0000000000000000_0000000110110100_0100110100001010"; -- 0.006657424033455629
	pesos_i(23465) := b"0000000000000000_0000000000000000_0000010001011001_0000100110001111"; -- 0.016983601863334072
	pesos_i(23466) := b"0000000000000000_0000000000000000_0000011001001100_0100100111111101"; -- 0.024601578076278132
	pesos_i(23467) := b"1111111111111111_1111111111111111_1111101111111011_1101001100111110"; -- -0.01568870304374956
	pesos_i(23468) := b"0000000000000000_0000000000000000_0010001111111100_0000010101011110"; -- 0.14056428473611873
	pesos_i(23469) := b"1111111111111111_1111111111111111_1110000101011010_1100110110011110"; -- -0.11970820316017117
	pesos_i(23470) := b"1111111111111111_1111111111111111_1111000000010101_1100011111111000"; -- -0.06216764640059615
	pesos_i(23471) := b"1111111111111111_1111111111111111_1111010010011000_0110101000101100"; -- -0.04454933569525278
	pesos_i(23472) := b"1111111111111111_1111111111111111_1111001011010101_1101100001111101"; -- -0.05142447413995268
	pesos_i(23473) := b"0000000000000000_0000000000000000_0000101011110100_0000000000011010"; -- 0.042785650470475986
	pesos_i(23474) := b"1111111111111111_1111111111111111_1101110011000001_0011010011001100"; -- -0.13767690671778668
	pesos_i(23475) := b"0000000000000000_0000000000000000_0010000001001001_1101100110010100"; -- 0.12612686026201897
	pesos_i(23476) := b"1111111111111111_1111111111111111_1111110000000100_1110110101101101"; -- -0.015549813256525172
	pesos_i(23477) := b"1111111111111111_1111111111111111_1110100101000101_0110101110100010"; -- -0.08878447819128114
	pesos_i(23478) := b"1111111111111111_1111111111111111_1111010111110111_0110001001111011"; -- -0.03919395918726114
	pesos_i(23479) := b"1111111111111111_1111111111111111_1110110000011101_0000110110110100"; -- -0.0776816782694524
	pesos_i(23480) := b"1111111111111111_1111111111111111_1110111101111010_0000011001010001"; -- -0.06454430119718702
	pesos_i(23481) := b"1111111111111111_1111111111111111_1110001111100000_0000100101110011"; -- -0.10986271799117055
	pesos_i(23482) := b"1111111111111111_1111111111111111_1110110000110011_0000010111010100"; -- -0.07734645433062512
	pesos_i(23483) := b"1111111111111111_1111111111111111_1110000001111001_0111011101100011"; -- -0.12314657054665708
	pesos_i(23484) := b"0000000000000000_0000000000000000_0000110001110111_1011001011100110"; -- 0.04870145903326964
	pesos_i(23485) := b"1111111111111111_1111111111111111_1111101111100000_0111100001010110"; -- -0.016106108652191614
	pesos_i(23486) := b"0000000000000000_0000000000000000_0000000011000011_0100001111110101"; -- 0.0029795143154505515
	pesos_i(23487) := b"1111111111111111_1111111111111111_1101110001110000_0001000000001111"; -- -0.13891505840929919
	pesos_i(23488) := b"0000000000000000_0000000000000000_0000011000010010_1101011010010000"; -- 0.023724947155762798
	pesos_i(23489) := b"0000000000000000_0000000000000000_0001111100110100_1000011000001100"; -- 0.12189519678111739
	pesos_i(23490) := b"0000000000000000_0000000000000000_0001101011000110_0110001100100101"; -- 0.10458964975844513
	pesos_i(23491) := b"0000000000000000_0000000000000000_0000110110000001_0001000111011111"; -- 0.05275069907922092
	pesos_i(23492) := b"0000000000000000_0000000000000000_0010000111100100_0001101001001010"; -- 0.13238682096805157
	pesos_i(23493) := b"1111111111111111_1111111111111111_1111001001001110_0011110010101100"; -- -0.053493698065359904
	pesos_i(23494) := b"1111111111111111_1111111111111111_1111011111000011_1001110010110111"; -- -0.03217144521121107
	pesos_i(23495) := b"1111111111111111_1111111111111111_1110001110010010_1101001101100010"; -- -0.1110408673319683
	pesos_i(23496) := b"0000000000000000_0000000000000000_0001001010010111_1100100101101100"; -- 0.07262858281215209
	pesos_i(23497) := b"1111111111111111_1111111111111111_1111001101001000_0101010111110111"; -- -0.04967749339462174
	pesos_i(23498) := b"1111111111111111_1111111111111111_1110011001000101_1110101000001111"; -- -0.10049569252277357
	pesos_i(23499) := b"0000000000000000_0000000000000000_0001110001000001_0110110001111001"; -- 0.11037328679350555
	pesos_i(23500) := b"1111111111111111_1111111111111111_1111000001010110_1111101101001111"; -- -0.06117276499274146
	pesos_i(23501) := b"1111111111111111_1111111111111111_1111110101000111_0001110101000101"; -- -0.010633631283499981
	pesos_i(23502) := b"0000000000000000_0000000000000000_0010001001111100_0111010100001000"; -- 0.1347115653488273
	pesos_i(23503) := b"0000000000000000_0000000000000000_0000101100100111_0011100100010100"; -- 0.04356724493876907
	pesos_i(23504) := b"0000000000000000_0000000000000000_0010001101001011_0111011001100101"; -- 0.13787021600144655
	pesos_i(23505) := b"1111111111111111_1111111111111111_1111100110101010_1001010101100110"; -- -0.024740851070625985
	pesos_i(23506) := b"0000000000000000_0000000000000000_0001000110110100_1110010100011011"; -- 0.06916648776009127
	pesos_i(23507) := b"1111111111111111_1111111111111111_1111101110010001_0110000010011110"; -- -0.017312966826782846
	pesos_i(23508) := b"0000000000000000_0000000000000000_0010001001011111_0101100110011000"; -- 0.13426742522920898
	pesos_i(23509) := b"0000000000000000_0000000000000000_0001011001011001_0001001010100110"; -- 0.0872966438712565
	pesos_i(23510) := b"1111111111111111_1111111111111111_1111101110010110_0001010101111111"; -- -0.017241150458941847
	pesos_i(23511) := b"0000000000000000_0000000000000000_0000001110011100_1101001111001110"; -- 0.014111745676419757
	pesos_i(23512) := b"1111111111111111_1111111111111111_1110001100001000_1010000100110110"; -- -0.11314957086691188
	pesos_i(23513) := b"1111111111111111_1111111111111111_1111011110101011_1101100010101010"; -- -0.032534082928946724
	pesos_i(23514) := b"0000000000000000_0000000000000000_0010010110001010_0100100100001111"; -- 0.14664131758794738
	pesos_i(23515) := b"1111111111111111_1111111111111111_1110000010001101_0011110011010101"; -- -0.1228448849621829
	pesos_i(23516) := b"1111111111111111_1111111111111111_1110101010000101_0000000010100100"; -- -0.08390804276491422
	pesos_i(23517) := b"0000000000000000_0000000000000000_0010000100110101_0101101000111110"; -- 0.12972034478841724
	pesos_i(23518) := b"0000000000000000_0000000000000000_0001100111000111_1101101011111100"; -- 0.10070580142350087
	pesos_i(23519) := b"0000000000000000_0000000000000000_0001101010100010_1001111111100010"; -- 0.10404395348511783
	pesos_i(23520) := b"0000000000000000_0000000000000000_0000000101010011_0000100000010100"; -- 0.00517321103223216
	pesos_i(23521) := b"0000000000000000_0000000000000000_0010000011010011_0000101111111010"; -- 0.1282203184495351
	pesos_i(23522) := b"0000000000000000_0000000000000000_0001101101100101_1001010100110100"; -- 0.10701878094061358
	pesos_i(23523) := b"0000000000000000_0000000000000000_0000000101101001_0100110001010000"; -- 0.005512971396492333
	pesos_i(23524) := b"1111111111111111_1111111111111111_1110010011110011_1010011011011111"; -- -0.1056571679443872
	pesos_i(23525) := b"1111111111111111_1111111111111111_1110010101001010_1110100011010011"; -- -0.10432572215447072
	pesos_i(23526) := b"0000000000000000_0000000000000000_0000000110100011_0100111010000001"; -- 0.0063981117116416845
	pesos_i(23527) := b"1111111111111111_1111111111111111_1111011100011111_0000101010001000"; -- -0.03468259980985779
	pesos_i(23528) := b"1111111111111111_1111111111111111_1111101011010101_0001101011010000"; -- -0.020185779728404733
	pesos_i(23529) := b"1111111111111111_1111111111111111_1101111010000111_0100110000110001"; -- -0.13074802204977853
	pesos_i(23530) := b"1111111111111111_1111111111111111_1110110100100000_1100010001011110"; -- -0.07371876439350843
	pesos_i(23531) := b"0000000000000000_0000000000000000_0000100001011011_0101010010001010"; -- 0.03264358877288669
	pesos_i(23532) := b"0000000000000000_0000000000000000_0001000110111011_0111100001011101"; -- 0.06926681786701075
	pesos_i(23533) := b"1111111111111111_1111111111111111_1110110000001011_1111110001111111"; -- -0.0779421034844774
	pesos_i(23534) := b"0000000000000000_0000000000000000_0000101100110010_0000010000101110"; -- 0.04373193854502856
	pesos_i(23535) := b"1111111111111111_1111111111111111_1110101101101001_0010111101000011"; -- -0.08042626005391264
	pesos_i(23536) := b"0000000000000000_0000000000000000_0001010100010000_0000010000100110"; -- 0.08227563787210883
	pesos_i(23537) := b"0000000000000000_0000000000000000_0001001010000111_0110101011100001"; -- 0.07237880695690666
	pesos_i(23538) := b"1111111111111111_1111111111111111_1101101110010011_0001100000111010"; -- -0.14228676392522666
	pesos_i(23539) := b"0000000000000000_0000000000000000_0001111000111101_1001011000110111"; -- 0.11812723963233175
	pesos_i(23540) := b"0000000000000000_0000000000000000_0000000001001011_1100000000011111"; -- 0.0011558604534558875
	pesos_i(23541) := b"0000000000000000_0000000000000000_0001101010111000_0001101000001011"; -- 0.10437166958483714
	pesos_i(23542) := b"0000000000000000_0000000000000000_0001111011100110_0111101000001010"; -- 0.12070429548530456
	pesos_i(23543) := b"1111111111111111_1111111111111111_1110011110101010_0000110011110010"; -- -0.09506148436577588
	pesos_i(23544) := b"1111111111111111_1111111111111111_1111111101000111_0001010111011001"; -- -0.002821573802031371
	pesos_i(23545) := b"0000000000000000_0000000000000000_0000100000111100_0111000010100111"; -- 0.03217224194322577
	pesos_i(23546) := b"0000000000000000_0000000000000000_0001011010111010_1101100100011101"; -- 0.0887885757291699
	pesos_i(23547) := b"1111111111111111_1111111111111111_1110100011011011_0110000110111001"; -- -0.09040250040648816
	pesos_i(23548) := b"0000000000000000_0000000000000000_0001011001000101_0000100101000011"; -- 0.0869909085782606
	pesos_i(23549) := b"0000000000000000_0000000000000000_0001010011100011_0000110110010101"; -- 0.081589554668249
	pesos_i(23550) := b"0000000000000000_0000000000000000_0001010001100110_1010111011001010"; -- 0.07969181469278508
	pesos_i(23551) := b"0000000000000000_0000000000000000_0000001010111110_1000101000010111"; -- 0.010719900654216989
	pesos_i(23552) := b"1111111111111111_1111111111111111_1110100101010001_1011010110001111"; -- -0.08859696645188089
	pesos_i(23553) := b"0000000000000000_0000000000000000_0000111110111100_0011100110100111"; -- 0.06146583873788399
	pesos_i(23554) := b"0000000000000000_0000000000000000_0000110011001110_1011000011101000"; -- 0.05002885492502971
	pesos_i(23555) := b"1111111111111111_1111111111111111_1111001011101010_0010001011011101"; -- -0.051114865310669624
	pesos_i(23556) := b"1111111111111111_1111111111111111_1111100100101111_0001101000110010"; -- -0.02662502547930448
	pesos_i(23557) := b"1111111111111111_1111111111111111_1110101101001111_1100011000111001"; -- -0.08081399057338613
	pesos_i(23558) := b"1111111111111111_1111111111111111_1101110001100100_1001100011110111"; -- -0.13909000371029834
	pesos_i(23559) := b"0000000000000000_0000000000000000_0001010010010111_0100111010111110"; -- 0.08043377048692414
	pesos_i(23560) := b"1111111111111111_1111111111111111_1101111001001010_0010110100010000"; -- -0.13168066364019174
	pesos_i(23561) := b"0000000000000000_0000000000000000_0000110111111110_1111000011111110"; -- 0.054671346786560424
	pesos_i(23562) := b"0000000000000000_0000000000000000_0000110011101100_1101000011001010"; -- 0.050488518906331055
	pesos_i(23563) := b"0000000000000000_0000000000000000_0001011110000111_0001001111100011"; -- 0.09190487182144672
	pesos_i(23564) := b"0000000000000000_0000000000000000_0001111101010001_0000110100001000"; -- 0.12233048860813031
	pesos_i(23565) := b"0000000000000000_0000000000000000_0000010110101000_1010000000011010"; -- 0.02210426935367974
	pesos_i(23566) := b"0000000000000000_0000000000000000_0000000110101001_1000110010101000"; -- 0.006493369087896843
	pesos_i(23567) := b"1111111111111111_1111111111111111_1101111000111101_1001110000111000"; -- -0.1318724024495459
	pesos_i(23568) := b"0000000000000000_0000000000000000_0010001101011111_1001011101011111"; -- 0.13817735740567605
	pesos_i(23569) := b"0000000000000000_0000000000000000_0000111101111100_0011000100000110"; -- 0.060488761842864454
	pesos_i(23570) := b"1111111111111111_1111111111111111_1111001010100000_0111100100011100"; -- -0.05223887512922637
	pesos_i(23571) := b"0000000000000000_0000000000000000_0010010001001011_1110111000000100"; -- 0.14178359608201452
	pesos_i(23572) := b"0000000000000000_0000000000000000_0001001001101111_1001010001011110"; -- 0.07201506896483173
	pesos_i(23573) := b"1111111111111111_1111111111111111_1111100111011110_0101001011110100"; -- -0.023951354420679593
	pesos_i(23574) := b"1111111111111111_1111111111111111_1111000110100101_1001010011101110"; -- -0.05606717285146758
	pesos_i(23575) := b"0000000000000000_0000000000000000_0000100010011000_0011100110011110"; -- 0.03357277027903588
	pesos_i(23576) := b"0000000000000000_0000000000000000_0001111000011111_1010100001011101"; -- 0.11767055761254995
	pesos_i(23577) := b"0000000000000000_0000000000000000_0001001010100101_0011010001111100"; -- 0.07283332841831129
	pesos_i(23578) := b"0000000000000000_0000000000000000_0001111101011000_0011110000001001"; -- 0.12244010179534416
	pesos_i(23579) := b"0000000000000000_0000000000000000_0001101011110001_1010100110101100"; -- 0.1052499813686198
	pesos_i(23580) := b"1111111111111111_1111111111111111_1111000111111110_1011101010001111"; -- -0.05470689780988864
	pesos_i(23581) := b"1111111111111111_1111111111111111_1111001011000010_0110101010001101"; -- -0.05172094389980209
	pesos_i(23582) := b"0000000000000000_0000000000000000_0000000010011011_0101001111001000"; -- 0.0023701061238222587
	pesos_i(23583) := b"1111111111111111_1111111111111111_1101101010110010_1101000100010110"; -- -0.14570897316668738
	pesos_i(23584) := b"1111111111111111_1111111111111111_1111001011101100_1001101001101110"; -- -0.051077221062547674
	pesos_i(23585) := b"1111111111111111_1111111111111111_1111110000101111_1101111111010111"; -- -0.014894494915985422
	pesos_i(23586) := b"1111111111111111_1111111111111111_1111110000111101_1000000001100101"; -- -0.014686560921984242
	pesos_i(23587) := b"1111111111111111_1111111111111111_1111100100001111_1010111000100001"; -- -0.02710448927514332
	pesos_i(23588) := b"0000000000000000_0000000000000000_0000101101001011_0110111101000110"; -- 0.044119791616766935
	pesos_i(23589) := b"0000000000000000_0000000000000000_0000110011011001_0011101110010101"; -- 0.050189708482898526
	pesos_i(23590) := b"1111111111111111_1111111111111111_1111110010110111_1010011010101000"; -- -0.012822708043183462
	pesos_i(23591) := b"1111111111111111_1111111111111111_1111011001111001_0111010011010011"; -- -0.037209223339636235
	pesos_i(23592) := b"0000000000000000_0000000000000000_0010000111000111_0100011111011100"; -- 0.13194703218948925
	pesos_i(23593) := b"1111111111111111_1111111111111111_1110001111000010_0010001111100010"; -- -0.11031890618425996
	pesos_i(23594) := b"1111111111111111_1111111111111111_1110110100011001_1010001111101100"; -- -0.07382750983966725
	pesos_i(23595) := b"0000000000000000_0000000000000000_0000010100010000_0100110111110010"; -- 0.019780036521762776
	pesos_i(23596) := b"1111111111111111_1111111111111111_1101110000011001_0101000000010110"; -- -0.1402387567575032
	pesos_i(23597) := b"0000000000000000_0000000000000000_0001100000001011_1100001100110001"; -- 0.0939294809173666
	pesos_i(23598) := b"1111111111111111_1111111111111111_1111000010100000_0010001101110011"; -- -0.060056480739077024
	pesos_i(23599) := b"1111111111111111_1111111111111111_1111101010111111_0010111100111000"; -- -0.02052025682290391
	pesos_i(23600) := b"0000000000000000_0000000000000000_0000011001010011_0100001000000100"; -- 0.02470791434989174
	pesos_i(23601) := b"1111111111111111_1111111111111111_1111000000010101_1010111111000011"; -- -0.06216908926232138
	pesos_i(23602) := b"0000000000000000_0000000000000000_0000101110001001_0000001111011111"; -- 0.04505943474612232
	pesos_i(23603) := b"1111111111111111_1111111111111111_1101111110100100_1011111100010101"; -- -0.12639241912438065
	pesos_i(23604) := b"0000000000000000_0000000000000000_0010000010010011_1011001001111101"; -- 0.1272536806734302
	pesos_i(23605) := b"1111111111111111_1111111111111111_1110010011101111_0110000111110000"; -- -0.10572231180555554
	pesos_i(23606) := b"1111111111111111_1111111111111111_1101111100000110_0011001001001101"; -- -0.12881169914563967
	pesos_i(23607) := b"1111111111111111_1111111111111111_1111000000011110_0101001101110110"; -- -0.062037261769804765
	pesos_i(23608) := b"0000000000000000_0000000000000000_0001010000011101_1000001100100010"; -- 0.07857532107672188
	pesos_i(23609) := b"0000000000000000_0000000000000000_0001010111000111_1100111011001111"; -- 0.08508007566475967
	pesos_i(23610) := b"0000000000000000_0000000000000000_0000010001001101_0100000001110001"; -- 0.016803767665229317
	pesos_i(23611) := b"0000000000000000_0000000000000000_0010000111001111_0001110101000100"; -- 0.1320665636924862
	pesos_i(23612) := b"1111111111111111_1111111111111111_1110110011011101_0010110111111101"; -- -0.0747500665345985
	pesos_i(23613) := b"1111111111111111_1111111111111111_1110001100010000_0111011000111001"; -- -0.11303006274311457
	pesos_i(23614) := b"1111111111111111_1111111111111111_1110101001100100_0010010100101001"; -- -0.08440940629144666
	pesos_i(23615) := b"0000000000000000_0000000000000000_0001110010010100_0001111000100010"; -- 0.11163509680809243
	pesos_i(23616) := b"1111111111111111_1111111111111111_1111011101110010_0011101000110100"; -- -0.033413278984053475
	pesos_i(23617) := b"0000000000000000_0000000000000000_0010010001010100_0101101100010011"; -- 0.14191216678256313
	pesos_i(23618) := b"0000000000000000_0000000000000000_0001001111001000_1000011011111111"; -- 0.07727855418269455
	pesos_i(23619) := b"0000000000000000_0000000000000000_0001111100110010_1100011011111110"; -- 0.12186855026878556
	pesos_i(23620) := b"1111111111111111_1111111111111111_1111100111101000_0001001100010101"; -- -0.023802573604895547
	pesos_i(23621) := b"0000000000000000_0000000000000000_0000110000000000_0101101111101011"; -- 0.046880478828647716
	pesos_i(23622) := b"0000000000000000_0000000000000000_0001110110010110_0011010011100101"; -- 0.11557322119033801
	pesos_i(23623) := b"1111111111111111_1111111111111111_1101100001001101_0010011001001010"; -- -0.15507279109101224
	pesos_i(23624) := b"0000000000000000_0000000000000000_0000101100001110_1001010101101101"; -- 0.04319127959979424
	pesos_i(23625) := b"1111111111111111_1111111111111111_1111001111001110_1100101100101100"; -- -0.047625829389232384
	pesos_i(23626) := b"0000000000000000_0000000000000000_0000010010100011_0100100110111011"; -- 0.018116577218753024
	pesos_i(23627) := b"1111111111111111_1111111111111111_1110110010101111_1001010001111100"; -- -0.07544586148382651
	pesos_i(23628) := b"1111111111111111_1111111111111111_1110101111100111_1111001101011001"; -- -0.07849196498095212
	pesos_i(23629) := b"0000000000000000_0000000000000000_0001010101010100_1101011001000110"; -- 0.0833257599073371
	pesos_i(23630) := b"1111111111111111_1111111111111111_1110011001010101_0000001100101010"; -- -0.10026531424342762
	pesos_i(23631) := b"1111111111111111_1111111111111111_1101111011010010_1111000000111101"; -- -0.12959383490473422
	pesos_i(23632) := b"0000000000000000_0000000000000000_0001011011011000_1110001001111011"; -- 0.08924689766601748
	pesos_i(23633) := b"0000000000000000_0000000000000000_0001111111010010_1001101101101000"; -- 0.1243073585801256
	pesos_i(23634) := b"1111111111111111_1111111111111111_1111000100011011_0001000011000111"; -- -0.05818076272710996
	pesos_i(23635) := b"0000000000000000_0000000000000000_0010010110101100_1000111101011101"; -- 0.1471643067912539
	pesos_i(23636) := b"0000000000000000_0000000000000000_0000000110111100_1110111110010110"; -- 0.006789182679351583
	pesos_i(23637) := b"0000000000000000_0000000000000000_0001011011111111_1101010011110001"; -- 0.08984118339772197
	pesos_i(23638) := b"0000000000000000_0000000000000000_0000111010010000_0100001111100101"; -- 0.05688881243232422
	pesos_i(23639) := b"0000000000000000_0000000000000000_0000101111101000_0000101000111000"; -- 0.04650939811935403
	pesos_i(23640) := b"1111111111111111_1111111111111111_1110011010000001_0011110011011100"; -- -0.09959048880046453
	pesos_i(23641) := b"1111111111111111_1111111111111111_1101011001000001_0110110000111010"; -- -0.16306422780389587
	pesos_i(23642) := b"0000000000000000_0000000000000000_0010101000110001_1111101001001101"; -- 0.1648250997891423
	pesos_i(23643) := b"0000000000000000_0000000000000000_0000010010111010_0010100011011001"; -- 0.018465569448861144
	pesos_i(23644) := b"0000000000000000_0000000000000000_0001101011100011_1011110001101001"; -- 0.10503747524677269
	pesos_i(23645) := b"0000000000000000_0000000000000000_0001110101011000_1011000110101010"; -- 0.11463461314498101
	pesos_i(23646) := b"1111111111111111_1111111111111111_1101101000100001_1001101011111011"; -- -0.1479247223452714
	pesos_i(23647) := b"0000000000000000_0000000000000000_0000101111101010_0111011011011101"; -- 0.04654639142121076
	pesos_i(23648) := b"0000000000000000_0000000000000000_0001101001001000_1101110010001111"; -- 0.10267427924347475
	pesos_i(23649) := b"1111111111111111_1111111111111111_1110010001011101_1011001101101101"; -- -0.10794523810850802
	pesos_i(23650) := b"1111111111111111_1111111111111111_1101111000001011_0110101010011110"; -- -0.1326382983865043
	pesos_i(23651) := b"1111111111111111_1111111111111111_1101111000001000_1100001000101000"; -- -0.1326788571717789
	pesos_i(23652) := b"1111111111111111_1111111111111111_1111101001100001_0100000101001100"; -- -0.021953505372050965
	pesos_i(23653) := b"0000000000000000_0000000000000000_0001110001000011_1000010101100001"; -- 0.11040528882450132
	pesos_i(23654) := b"0000000000000000_0000000000000000_0001010111000000_1110110010101011"; -- 0.0849750441197296
	pesos_i(23655) := b"0000000000000000_0000000000000000_0000001011011111_1011011110010000"; -- 0.011226151135216147
	pesos_i(23656) := b"1111111111111111_1111111111111111_1111001101010001_1110101111100111"; -- -0.04953122717793971
	pesos_i(23657) := b"0000000000000000_0000000000000000_0000011011010001_0000010101101110"; -- 0.026626910509865036
	pesos_i(23658) := b"0000000000000000_0000000000000000_0010000001000010_0101011110000111"; -- 0.1260122971926337
	pesos_i(23659) := b"0000000000000000_0000000000000000_0000011111011011_0001111111010001"; -- 0.030687321247353717
	pesos_i(23660) := b"0000000000000000_0000000000000000_0000000101010111_1001100000001001"; -- 0.005242826542322012
	pesos_i(23661) := b"0000000000000000_0000000000000000_0000010010110000_0000000111101011"; -- 0.01831066124685429
	pesos_i(23662) := b"0000000000000000_0000000000000000_0001111001001001_0001000101101100"; -- 0.11830243011743433
	pesos_i(23663) := b"1111111111111111_1111111111111111_1101100110001100_0100011001010110"; -- -0.15020332718622403
	pesos_i(23664) := b"1111111111111111_1111111111111111_1110110101001110_1001000110010000"; -- -0.0730198881838807
	pesos_i(23665) := b"1111111111111111_1111111111111111_1110100100111111_0001111010110111"; -- -0.08888061562274642
	pesos_i(23666) := b"0000000000000000_0000000000000000_0000001111011110_1101100101001000"; -- 0.01511915218101483
	pesos_i(23667) := b"1111111111111111_1111111111111111_1111101100100101_1011010101110000"; -- -0.018955860176006475
	pesos_i(23668) := b"0000000000000000_0000000000000000_0000101000010101_1001111011111001"; -- 0.039392410043998155
	pesos_i(23669) := b"1111111111111111_1111111111111111_1110100011010100_0100100000100100"; -- -0.09051083687977117
	pesos_i(23670) := b"1111111111111111_1111111111111111_1101110001011110_0101101010010001"; -- -0.13918527575930545
	pesos_i(23671) := b"1111111111111111_1111111111111111_1110101001001000_0010101000010000"; -- -0.08483636000510399
	pesos_i(23672) := b"1111111111111111_1111111111111111_1110110111101001_0001011110110100"; -- -0.07066203926908733
	pesos_i(23673) := b"0000000000000000_0000000000000000_0001000110011100_1000110110100001"; -- 0.06879506291315057
	pesos_i(23674) := b"0000000000000000_0000000000000000_0000011000100101_1010111101111011"; -- 0.024012534745725615
	pesos_i(23675) := b"0000000000000000_0000000000000000_0001010000001010_0110001000101010"; -- 0.07828343900518829
	pesos_i(23676) := b"0000000000000000_0000000000000000_0001110101000001_1100110111111100"; -- 0.11428534892243213
	pesos_i(23677) := b"1111111111111111_1111111111111111_1110010001011000_1001110001000010"; -- -0.10802291280428515
	pesos_i(23678) := b"1111111111111111_1111111111111111_1110100111000110_0111101010101100"; -- -0.08681519802667337
	pesos_i(23679) := b"0000000000000000_0000000000000000_0001100000011111_0110100010000110"; -- 0.0942292524602415
	pesos_i(23680) := b"1111111111111111_1111111111111111_1111001110011111_0111110101011100"; -- -0.04834763046727301
	pesos_i(23681) := b"0000000000000000_0000000000000000_0000111111111110_1011010100100010"; -- 0.062480278807616814
	pesos_i(23682) := b"1111111111111111_1111111111111111_1110111110001110_1010110011000000"; -- -0.06422920520132279
	pesos_i(23683) := b"1111111111111111_1111111111111111_1111010111111101_0101111110101111"; -- -0.03910257321872832
	pesos_i(23684) := b"0000000000000000_0000000000000000_0000111110101001_1000010010001010"; -- 0.0611803853782646
	pesos_i(23685) := b"1111111111111111_1111111111111111_1111111111101011_0100110100000111"; -- -0.0003158434735462282
	pesos_i(23686) := b"1111111111111111_1111111111111111_1110001100100010_1110111011100000"; -- -0.11274821307272027
	pesos_i(23687) := b"0000000000000000_0000000000000000_0001100011100111_0000110000000011"; -- 0.09727549629977195
	pesos_i(23688) := b"0000000000000000_0000000000000000_0000011010010110_0010101111010111"; -- 0.025728931366218438
	pesos_i(23689) := b"1111111111111111_1111111111111111_1110100000001001_1011011111001111"; -- -0.09360171511137924
	pesos_i(23690) := b"1111111111111111_1111111111111111_1110000010000001_1000010101010111"; -- -0.12302366845596953
	pesos_i(23691) := b"1111111111111111_1111111111111111_1110110011110011_1110011100100101"; -- -0.07440333694816019
	pesos_i(23692) := b"1111111111111111_1111111111111111_1101111100111000_1000001000100011"; -- -0.1280440011252551
	pesos_i(23693) := b"0000000000000000_0000000000000000_0001011111110110_1000111110001111"; -- 0.09360596892633545
	pesos_i(23694) := b"0000000000000000_0000000000000000_0001001101000010_1111101000110111"; -- 0.07524074398568312
	pesos_i(23695) := b"1111111111111111_1111111111111111_1101100101010000_1100000010101010"; -- -0.1511115633021389
	pesos_i(23696) := b"0000000000000000_0000000000000000_0001001111000100_1111010111100101"; -- 0.07722412904437803
	pesos_i(23697) := b"0000000000000000_0000000000000000_0010000100100101_1010000010001010"; -- 0.1294803940180453
	pesos_i(23698) := b"1111111111111111_1111111111111111_1110001000010101_0000000011111100"; -- -0.11686700664025218
	pesos_i(23699) := b"1111111111111111_1111111111111111_1110001111100000_1111000101111100"; -- -0.10984888757852648
	pesos_i(23700) := b"0000000000000000_0000000000000000_0010000010010010_1011011110010110"; -- 0.12723872588179008
	pesos_i(23701) := b"0000000000000000_0000000000000000_0001010010011100_1001011001011000"; -- 0.08051433227071696
	pesos_i(23702) := b"1111111111111111_1111111111111111_1110100000100111_0011101011100101"; -- -0.09315139686924939
	pesos_i(23703) := b"1111111111111111_1111111111111111_1111101010111010_0110111000011111"; -- -0.02059280145196225
	pesos_i(23704) := b"0000000000000000_0000000000000000_0001101100100011_1100100111101110"; -- 0.10601484367900575
	pesos_i(23705) := b"0000000000000000_0000000000000000_0001010100000011_0110010101100011"; -- 0.08208306953797169
	pesos_i(23706) := b"0000000000000000_0000000000000000_0000001101011110_1101000011011100"; -- 0.013165525045510518
	pesos_i(23707) := b"0000000000000000_0000000000000000_0000100011001011_0100000100000000"; -- 0.03435140837109066
	pesos_i(23708) := b"1111111111111111_1111111111111111_1101100110000101_0111111011010001"; -- -0.1503067721834212
	pesos_i(23709) := b"0000000000000000_0000000000000000_0001101101000101_1100110000110100"; -- 0.10653377785211998
	pesos_i(23710) := b"0000000000000000_0000000000000000_0001010000000100_1001111101100000"; -- 0.07819553467971956
	pesos_i(23711) := b"0000000000000000_0000000000000000_0000001100100110_0100110111110011"; -- 0.012303230036097058
	pesos_i(23712) := b"1111111111111111_1111111111111111_1110100110000101_0000110010011000"; -- -0.08781358034796978
	pesos_i(23713) := b"0000000000000000_0000000000000000_0001101100100100_0001100000001110"; -- 0.10601950017526178
	pesos_i(23714) := b"0000000000000000_0000000000000000_0000101000100010_1000101101100110"; -- 0.039589607725089314
	pesos_i(23715) := b"0000000000000000_0000000000000000_0000011011101101_1011010101100001"; -- 0.027064644092253
	pesos_i(23716) := b"0000000000000000_0000000000000000_0001100001001001_1011011000100100"; -- 0.09487474801221603
	pesos_i(23717) := b"1111111111111111_1111111111111111_1101110001101110_0011000110011000"; -- -0.13894357715514066
	pesos_i(23718) := b"1111111111111111_1111111111111111_1111010111101100_1100101101110000"; -- -0.03935555007688869
	pesos_i(23719) := b"0000000000000000_0000000000000000_0001000100000000_0011000100111010"; -- 0.06640918410752927
	pesos_i(23720) := b"1111111111111111_1111111111111111_1110110100100111_1001001000011011"; -- -0.07361494859586228
	pesos_i(23721) := b"1111111111111111_1111111111111111_1110010011000011_1010000101101011"; -- -0.10638991481989894
	pesos_i(23722) := b"0000000000000000_0000000000000000_0001100100001100_1000101001001101"; -- 0.09784759889942092
	pesos_i(23723) := b"0000000000000000_0000000000000000_0010100010111101_1110111011011100"; -- 0.1591481482721637
	pesos_i(23724) := b"0000000000000000_0000000000000000_0000000000011010_1010000110100101"; -- 0.00040636322227093964
	pesos_i(23725) := b"0000000000000000_0000000000000000_0001010000100100_0010101101000011"; -- 0.07867689508916864
	pesos_i(23726) := b"0000000000000000_0000000000000000_0001111110110001_1011011010101010"; -- 0.12380544325686177
	pesos_i(23727) := b"1111111111111111_1111111111111111_1110101100001111_1001011110000100"; -- -0.08179333722920852
	pesos_i(23728) := b"0000000000000000_0000000000000000_0000011100111000_1010111101111110"; -- 0.02820870229135158
	pesos_i(23729) := b"0000000000000000_0000000000000000_0001111100111111_1101001000101000"; -- 0.12206757989179173
	pesos_i(23730) := b"0000000000000000_0000000000000000_0000100011010011_0110001010111100"; -- 0.0344754894947637
	pesos_i(23731) := b"1111111111111111_1111111111111111_1110000101010100_1100100001010001"; -- -0.11980007202615134
	pesos_i(23732) := b"1111111111111111_1111111111111111_1110000010010100_0000010011000000"; -- -0.12274141620797693
	pesos_i(23733) := b"0000000000000000_0000000000000000_0001000011100011_1110001011001001"; -- 0.06597726250326054
	pesos_i(23734) := b"1111111111111111_1111111111111111_1101011011000011_0010010101110011"; -- -0.16108480397452446
	pesos_i(23735) := b"0000000000000000_0000000000000000_0000011011110111_1001010100101111"; -- 0.027215312989234054
	pesos_i(23736) := b"1111111111111111_1111111111111111_1101101000110010_0010110101100101"; -- -0.14767185486383838
	pesos_i(23737) := b"1111111111111111_1111111111111111_1110000010010001_1100110001010001"; -- -0.12277529730990058
	pesos_i(23738) := b"0000000000000000_0000000000000000_0000111110111010_0100011101101010"; -- 0.06143614130175869
	pesos_i(23739) := b"0000000000000000_0000000000000000_0000100010111100_1100000111000000"; -- 0.034130200701799104
	pesos_i(23740) := b"0000000000000000_0000000000000000_0001001000110001_0111000010011111"; -- 0.07106689331437811
	pesos_i(23741) := b"1111111111111111_1111111111111111_1101100000101011_0011100101010111"; -- -0.15559045440870958
	pesos_i(23742) := b"1111111111111111_1111111111111111_1110010011011010_0111111100101110"; -- -0.10604100360064649
	pesos_i(23743) := b"0000000000000000_0000000000000000_0000100101100011_0101010110110010"; -- 0.036671978049649424
	pesos_i(23744) := b"0000000000000000_0000000000000000_0000100100101110_1111100100011011"; -- 0.035873002024960625
	pesos_i(23745) := b"1111111111111111_1111111111111111_1111100011100100_1100111111111110"; -- -0.027758598840975892
	pesos_i(23746) := b"0000000000000000_0000000000000000_0001010101010100_1000100100010110"; -- 0.08332115918206354
	pesos_i(23747) := b"0000000000000000_0000000000000000_0001001000100110_1000100101100101"; -- 0.07090052323318755
	pesos_i(23748) := b"0000000000000000_0000000000000000_0000110111001100_0100011101000011"; -- 0.05389829043812423
	pesos_i(23749) := b"0000000000000000_0000000000000000_0000010111101000_0001011001100011"; -- 0.023072623397676677
	pesos_i(23750) := b"0000000000000000_0000000000000000_0010011100011011_1111111011100100"; -- 0.15277092994636132
	pesos_i(23751) := b"1111111111111111_1111111111111111_1111001100110110_1010001100100011"; -- -0.0499475516071778
	pesos_i(23752) := b"1111111111111111_1111111111111111_1111000011101101_0011111011110100"; -- -0.05887991472502485
	pesos_i(23753) := b"1111111111111111_1111111111111111_1101110111110000_1110001111110111"; -- -0.1330430528910418
	pesos_i(23754) := b"1111111111111111_1111111111111111_1101111011100100_1001110101001000"; -- -0.1293241213712178
	pesos_i(23755) := b"1111111111111111_1111111111111111_1111001100011111_0110101001100010"; -- -0.050301886696734036
	pesos_i(23756) := b"1111111111111111_1111111111111111_1101111111100011_0010100011100110"; -- -0.12544006707682398
	pesos_i(23757) := b"1111111111111111_1111111111111111_1110101100111100_1100001100001011"; -- -0.08110409708179023
	pesos_i(23758) := b"0000000000000000_0000000000000000_0001101110100101_1010111001001000"; -- 0.1079968382015815
	pesos_i(23759) := b"0000000000000000_0000000000000000_0000010010010100_1111100100000110"; -- 0.017898143747142402
	pesos_i(23760) := b"1111111111111111_1111111111111111_1111001001000101_1001110111010010"; -- -0.053625236709440194
	pesos_i(23761) := b"1111111111111111_1111111111111111_1110010011110011_1001101001101010"; -- -0.10565791055286536
	pesos_i(23762) := b"1111111111111111_1111111111111111_1110111000000100_0000000011011001"; -- -0.0702514143145822
	pesos_i(23763) := b"1111111111111111_1111111111111111_1111000000111011_1000111110000010"; -- -0.0615911777930469
	pesos_i(23764) := b"1111111111111111_1111111111111111_1110010110010101_0101110011110101"; -- -0.10318964982780013
	pesos_i(23765) := b"1111111111111111_1111111111111111_1111001011100011_0010100010100111"; -- -0.0512213317343095
	pesos_i(23766) := b"1111111111111111_1111111111111111_1111101110101100_0111010010001110"; -- -0.016899791001829333
	pesos_i(23767) := b"1111111111111111_1111111111111111_1101100101000011_1100100011100011"; -- -0.15130943733902819
	pesos_i(23768) := b"0000000000000000_0000000000000000_0010100001000000_0101101100001110"; -- 0.15723198984765702
	pesos_i(23769) := b"1111111111111111_1111111111111111_1110001001001001_0110110101100111"; -- -0.11606708740495615
	pesos_i(23770) := b"0000000000000000_0000000000000000_0001101000100001_1001011000001100"; -- 0.10207498351679674
	pesos_i(23771) := b"1111111111111111_1111111111111111_1110100101010111_1101010101010110"; -- -0.08850351950711312
	pesos_i(23772) := b"1111111111111111_1111111111111111_1110001001111111_0011011011000000"; -- -0.11524637033629312
	pesos_i(23773) := b"0000000000000000_0000000000000000_0000111111111000_1010101010000001"; -- 0.062388092559781456
	pesos_i(23774) := b"0000000000000000_0000000000000000_0000001011110100_1000110011010000"; -- 0.011544037598714238
	pesos_i(23775) := b"1111111111111111_1111111111111111_1111000011100111_1110000100000010"; -- -0.05896180833192114
	pesos_i(23776) := b"1111111111111111_1111111111111111_1101100111001001_1011000101101010"; -- -0.1492661586994467
	pesos_i(23777) := b"1111111111111111_1111111111111111_1111110001101110_1000011101001101"; -- -0.013938468650333184
	pesos_i(23778) := b"0000000000000000_0000000000000000_0001010100111110_1100111101000111"; -- 0.08298964960977961
	pesos_i(23779) := b"1111111111111111_1111111111111111_1110001101110110_0111001010100000"; -- -0.11147388081876747
	pesos_i(23780) := b"1111111111111111_1111111111111111_1101100001110011_0110011000001110"; -- -0.15448915625193863
	pesos_i(23781) := b"0000000000000000_0000000000000000_0001100001000111_0011101111111011"; -- 0.09483694913416436
	pesos_i(23782) := b"0000000000000000_0000000000000000_0001111110110100_0111110010001100"; -- 0.12384775561320142
	pesos_i(23783) := b"1111111111111111_1111111111111111_1101110000101110_1000010010000001"; -- -0.1399151978401697
	pesos_i(23784) := b"1111111111111111_1111111111111111_1111011001100000_0100001101011110"; -- -0.037593640813331594
	pesos_i(23785) := b"0000000000000000_0000000000000000_0000110000000001_0011011001011100"; -- 0.04689349874958969
	pesos_i(23786) := b"0000000000000000_0000000000000000_0010000011111101_0101101001011000"; -- 0.12886585847865253
	pesos_i(23787) := b"1111111111111111_1111111111111111_1111100000111101_1101000101000111"; -- -0.03030673985260541
	pesos_i(23788) := b"0000000000000000_0000000000000000_0010011000010111_0010001101101100"; -- 0.14879056351035497
	pesos_i(23789) := b"0000000000000000_0000000000000000_0000001001011001_0000110010001110"; -- 0.00917128055813034
	pesos_i(23790) := b"1111111111111111_1111111111111111_1110100100000101_0111110100111100"; -- -0.08975999146107083
	pesos_i(23791) := b"1111111111111111_1111111111111111_1111111110011010_0011110000000011"; -- -0.0015528194057261612
	pesos_i(23792) := b"1111111111111111_1111111111111111_1110111000110110_1000101100110100"; -- -0.06948022818306022
	pesos_i(23793) := b"1111111111111111_1111111111111111_1110101111101101_1110000001011000"; -- -0.07840154496296985
	pesos_i(23794) := b"0000000000000000_0000000000000000_0001100000000110_0101100011100111"; -- 0.09384685179052955
	pesos_i(23795) := b"1111111111111111_1111111111111111_1111101010111000_0000011011011010"; -- -0.020629474452198034
	pesos_i(23796) := b"0000000000000000_0000000000000000_0001100100100111_0101001111010010"; -- 0.09825633882411251
	pesos_i(23797) := b"0000000000000000_0000000000000000_0010010001111111_1000000001111101"; -- 0.1425705247155313
	pesos_i(23798) := b"1111111111111111_1111111111111111_1110001001100110_0010101011101000"; -- -0.1156285462074738
	pesos_i(23799) := b"1111111111111111_1111111111111111_1111000010010011_0011110100011000"; -- -0.060253316541250955
	pesos_i(23800) := b"0000000000000000_0000000000000000_0010001011110000_1100000010001101"; -- 0.1364860864020904
	pesos_i(23801) := b"1111111111111111_1111111111111111_1111110100101100_1000001011001001"; -- -0.011039567913207905
	pesos_i(23802) := b"0000000000000000_0000000000000000_0000011001011011_0010110001100111"; -- 0.02482869633511111
	pesos_i(23803) := b"1111111111111111_1111111111111111_1110011101011011_0000111111011101"; -- -0.09626675463473923
	pesos_i(23804) := b"1111111111111111_1111111111111111_1110010101101000_0000111010000010"; -- -0.10388097125532772
	pesos_i(23805) := b"0000000000000000_0000000000000000_0001110011001101_1000010010010010"; -- 0.11251095346374876
	pesos_i(23806) := b"1111111111111111_1111111111111111_1110001001001111_0110101011011100"; -- -0.11597568638003108
	pesos_i(23807) := b"1111111111111111_1111111111111111_1110001111001101_0101000000000000"; -- -0.11014842984505263
	pesos_i(23808) := b"1111111111111111_1111111111111111_1111011111010111_0110000010010101"; -- -0.031869853597718885
	pesos_i(23809) := b"1111111111111111_1111111111111111_1101110111111111_0010110101000101"; -- -0.1328250604796158
	pesos_i(23810) := b"1111111111111111_1111111111111111_1101010001010100_0110010010000011"; -- -0.17058727086609426
	pesos_i(23811) := b"0000000000000000_0000000000000000_0010000001010111_1010001001011010"; -- 0.12633719157669626
	pesos_i(23812) := b"1111111111111111_1111111111111111_1110010001110000_1000110001010110"; -- -0.1076576509088141
	pesos_i(23813) := b"1111111111111111_1111111111111111_1111001010110101_1101101010111101"; -- -0.0519126212646413
	pesos_i(23814) := b"0000000000000000_0000000000000000_0000000100010110_1110111110110110"; -- 0.004256231228603707
	pesos_i(23815) := b"0000000000000000_0000000000000000_0000111111001011_0101011000111010"; -- 0.061696423658172815
	pesos_i(23816) := b"1111111111111111_1111111111111111_1111001110111110_1100101010101001"; -- -0.04787000062466171
	pesos_i(23817) := b"1111111111111111_1111111111111111_1110000001101101_0110001101001100"; -- -0.12333087333168304
	pesos_i(23818) := b"1111111111111111_1111111111111111_1110101110001110_0000001110001100"; -- -0.07986429060213968
	pesos_i(23819) := b"1111111111111111_1111111111111111_1111100000000100_0110011101010001"; -- -0.031182806611311346
	pesos_i(23820) := b"0000000000000000_0000000000000000_0000101011001101_0101101000111110"; -- 0.042195930548721616
	pesos_i(23821) := b"0000000000000000_0000000000000000_0001111000111000_1000001010001011"; -- 0.11804977312881945
	pesos_i(23822) := b"0000000000000000_0000000000000000_0001111000111110_0000010100010110"; -- 0.11813384796503235
	pesos_i(23823) := b"1111111111111111_1111111111111111_1101100110001100_1000110111010111"; -- -0.15019906528272567
	pesos_i(23824) := b"1111111111111111_1111111111111111_1110111110111000_1011010011101100"; -- -0.06358784901069613
	pesos_i(23825) := b"0000000000000000_0000000000000000_0000111100011100_0000000100010001"; -- 0.05902105970641122
	pesos_i(23826) := b"0000000000000000_0000000000000000_0001000010001001_1000001011110100"; -- 0.0645982594956373
	pesos_i(23827) := b"0000000000000000_0000000000000000_0001110111000010_1110101010011101"; -- 0.11625543904122106
	pesos_i(23828) := b"1111111111111111_1111111111111111_1110001001001010_1001010111011100"; -- -0.11604941731539196
	pesos_i(23829) := b"0000000000000000_0000000000000000_0001110010000110_1000010110100110"; -- 0.11142764371095674
	pesos_i(23830) := b"1111111111111111_1111111111111111_1111011011101001_0011000100110011"; -- -0.03550426969611683
	pesos_i(23831) := b"0000000000000000_0000000000000000_0001010101111110_0101001110000101"; -- 0.08395883565356917
	pesos_i(23832) := b"0000000000000000_0000000000000000_0001001001011011_1111100000000111"; -- 0.0717158333588164
	pesos_i(23833) := b"1111111111111111_1111111111111111_1110000110000000_1000101111111011"; -- -0.11913228140718964
	pesos_i(23834) := b"1111111111111111_1111111111111111_1110110111101000_0000000010111010"; -- -0.07067866764285603
	pesos_i(23835) := b"1111111111111111_1111111111111111_1110010111010001_0111001001110000"; -- -0.10227284212871446
	pesos_i(23836) := b"0000000000000000_0000000000000000_0000110110001011_1110110010010010"; -- 0.05291632233726135
	pesos_i(23837) := b"1111111111111111_1111111111111111_1110110100110110_1001001010110011"; -- -0.07338603134291156
	pesos_i(23838) := b"1111111111111111_1111111111111111_1101111101101001_1010101011111101"; -- -0.12729388539455386
	pesos_i(23839) := b"0000000000000000_0000000000000000_0000100000010111_1010010110001011"; -- 0.03161081921725567
	pesos_i(23840) := b"0000000000000000_0000000000000000_0000100111110010_1011100010110111"; -- 0.03885988681349844
	pesos_i(23841) := b"1111111111111111_1111111111111111_1111101011110110_1011001110001101"; -- -0.019673135780952453
	pesos_i(23842) := b"1111111111111111_1111111111111111_1111111000110001_1110011101010010"; -- -0.0070510316686411304
	pesos_i(23843) := b"1111111111111111_1111111111111111_1111101111011111_0000110001100110"; -- -0.016127800994011468
	pesos_i(23844) := b"0000000000000000_0000000000000000_0000001001111111_1000101011111101"; -- 0.009758650569277735
	pesos_i(23845) := b"1111111111111111_1111111111111111_1101101010010100_1100001110011110"; -- -0.14616753955857018
	pesos_i(23846) := b"1111111111111111_1111111111111111_1111101110111000_0010101010001111"; -- -0.01672109621195296
	pesos_i(23847) := b"0000000000000000_0000000000000000_0000010111100111_0111101111001101"; -- 0.023063409448050687
	pesos_i(23848) := b"0000000000000000_0000000000000000_0000111010011101_0110101000011011"; -- 0.05708945428075409
	pesos_i(23849) := b"1111111111111111_1111111111111111_1111011001100001_1100101000100001"; -- -0.03757034970293349
	pesos_i(23850) := b"1111111111111111_1111111111111111_1110010001110111_0010010000000110"; -- -0.10755705701832008
	pesos_i(23851) := b"1111111111111111_1111111111111111_1111111101111001_1100011110100001"; -- -0.00204803776101595
	pesos_i(23852) := b"0000000000000000_0000000000000000_0010000001110010_0110100011001100"; -- 0.12674574834104468
	pesos_i(23853) := b"0000000000000000_0000000000000000_0010010011101011_0001110000001111"; -- 0.14421248780803128
	pesos_i(23854) := b"1111111111111111_1111111111111111_1110101000010000_1101010101011101"; -- -0.0856806419445019
	pesos_i(23855) := b"0000000000000000_0000000000000000_0001001011100110_1011001100001000"; -- 0.07383269246468245
	pesos_i(23856) := b"1111111111111111_1111111111111111_1110100000001000_1000001101001011"; -- -0.0936201041290045
	pesos_i(23857) := b"0000000000000000_0000000000000000_0000001011111100_0111101101111001"; -- 0.011665074388244342
	pesos_i(23858) := b"0000000000000000_0000000000000000_0000101111000011_0011101001010111"; -- 0.0459476912596935
	pesos_i(23859) := b"1111111111111111_1111111111111111_1111010010100101_0000100110001111"; -- -0.044356730130700926
	pesos_i(23860) := b"0000000000000000_0000000000000000_0001100000100111_0000001011101001"; -- 0.09434526613310064
	pesos_i(23861) := b"0000000000000000_0000000000000000_0000100101111010_0111111101101001"; -- 0.037025416584108864
	pesos_i(23862) := b"0000000000000000_0000000000000000_0001000101011110_1100000011101010"; -- 0.06785207482746335
	pesos_i(23863) := b"1111111111111111_1111111111111111_1110000110100100_1111111101001111"; -- -0.11857609098823345
	pesos_i(23864) := b"1111111111111111_1111111111111111_1111000101100111_1110010101000001"; -- -0.05700843016412362
	pesos_i(23865) := b"0000000000000000_0000000000000000_0001010111011100_1100011000000101"; -- 0.08539998639011659
	pesos_i(23866) := b"1111111111111111_1111111111111111_1110011000010011_1011110000110101"; -- -0.10126136504766615
	pesos_i(23867) := b"0000000000000000_0000000000000000_0000101101001000_0000001111001011"; -- 0.04406760892243134
	pesos_i(23868) := b"1111111111111111_1111111111111111_1110101010110101_1110110001100000"; -- -0.08316157011729942
	pesos_i(23869) := b"1111111111111111_1111111111111111_1111000110011110_1111100100000000"; -- -0.05616801986848578
	pesos_i(23870) := b"0000000000000000_0000000000000000_0001010011010001_0010001010110111"; -- 0.0813161561812104
	pesos_i(23871) := b"1111111111111111_1111111111111111_1101111000011100_1000101010100010"; -- -0.13237699068862513
	pesos_i(23872) := b"0000000000000000_0000000000000000_0000000010110111_0101010100010101"; -- 0.002797429592096834
	pesos_i(23873) := b"1111111111111111_1111111111111111_1110011111010110_0110000001101001"; -- -0.09438512255498935
	pesos_i(23874) := b"1111111111111111_1111111111111111_1111110001110101_1011010010010000"; -- -0.013828959400817803
	pesos_i(23875) := b"1111111111111111_1111111111111111_1110111010010111_1011011111000001"; -- -0.06799747015533415
	pesos_i(23876) := b"0000000000000000_0000000000000000_0000000101000001_0011001000000011"; -- 0.004901052141162455
	pesos_i(23877) := b"0000000000000000_0000000000000000_0000110111110011_0111110100011000"; -- 0.05449659192115416
	pesos_i(23878) := b"1111111111111111_1111111111111111_1111100010111101_1011100001111101"; -- -0.02835509243616952
	pesos_i(23879) := b"0000000000000000_0000000000000000_0010010011011010_0001100011111010"; -- 0.14395290472108563
	pesos_i(23880) := b"0000000000000000_0000000000000000_0000100000101011_0101100010001111"; -- 0.031911406360617275
	pesos_i(23881) := b"1111111111111111_1111111111111111_1110100101010100_1111010101111010"; -- -0.08854738022396652
	pesos_i(23882) := b"0000000000000000_0000000000000000_0000101100110010_1100100101100010"; -- 0.0437436927266287
	pesos_i(23883) := b"0000000000000000_0000000000000000_0001100001101001_0010011101101011"; -- 0.09535452238493919
	pesos_i(23884) := b"0000000000000000_0000000000000000_0001110110000100_0001011010000100"; -- 0.11529675211379699
	pesos_i(23885) := b"1111111111111111_1111111111111111_1101100111010110_1100101011110001"; -- -0.1490662729317836
	pesos_i(23886) := b"0000000000000000_0000000000000000_0010010001110101_0001110111010001"; -- 0.14241205559179454
	pesos_i(23887) := b"1111111111111111_1111111111111111_1110011011110010_0110000001010010"; -- -0.09786413184161001
	pesos_i(23888) := b"0000000000000000_0000000000000000_0001001001101110_0010001011010100"; -- 0.07199304260715267
	pesos_i(23889) := b"1111111111111111_1111111111111111_1111110000101110_0101000010011100"; -- -0.014918290912932274
	pesos_i(23890) := b"1111111111111111_1111111111111111_1101101100011011_0110001100100001"; -- -0.14411335410826845
	pesos_i(23891) := b"0000000000000000_0000000000000000_0000001101110000_1011010111001110"; -- 0.013438570709904842
	pesos_i(23892) := b"1111111111111111_1111111111111111_1110101001000101_1101100010011111"; -- -0.0848717319028891
	pesos_i(23893) := b"1111111111111111_1111111111111111_1110011001000010_0010000111110101"; -- -0.10055339598722678
	pesos_i(23894) := b"1111111111111111_1111111111111111_1111011011100111_0111010000100001"; -- -0.03553079781894754
	pesos_i(23895) := b"0000000000000000_0000000000000000_0000110001001010_1001011000010110"; -- 0.04801309629774398
	pesos_i(23896) := b"0000000000000000_0000000000000000_0000011101011111_1010110001111100"; -- 0.028803615853763766
	pesos_i(23897) := b"0000000000000000_0000000000000000_0000101111111000_0010110101111010"; -- 0.046755640297194034
	pesos_i(23898) := b"1111111111111111_1111111111111111_1111111111100011_0000101011010111"; -- -0.00044185873456457854
	pesos_i(23899) := b"0000000000000000_0000000000000000_0001111110110011_1111101111000011"; -- 0.12384007937337219
	pesos_i(23900) := b"0000000000000000_0000000000000000_0000011010010001_1100010001001100"; -- 0.025661724573595997
	pesos_i(23901) := b"0000000000000000_0000000000000000_0001010101100101_1100110111100011"; -- 0.08358465949385967
	pesos_i(23902) := b"1111111111111111_1111111111111111_1110011111100000_0111111000110110"; -- -0.09423075851260673
	pesos_i(23903) := b"1111111111111111_1111111111111111_1111101000000101_0101110100111000"; -- -0.023355649852344312
	pesos_i(23904) := b"1111111111111111_1111111111111111_1110000010000101_0010010110000100"; -- -0.12296834505212963
	pesos_i(23905) := b"1111111111111111_1111111111111111_1110000001011011_1100011100001100"; -- -0.12359958599463615
	pesos_i(23906) := b"1111111111111111_1111111111111111_1111100010010100_0110111001010111"; -- -0.02898512252316025
	pesos_i(23907) := b"0000000000000000_0000000000000000_0001000010101101_0101101110110001"; -- 0.06514523578297388
	pesos_i(23908) := b"0000000000000000_0000000000000000_0000011010100000_0011000000111110"; -- 0.025881781814891768
	pesos_i(23909) := b"0000000000000000_0000000000000000_0010010101110111_0001010101001111"; -- 0.14634831594809594
	pesos_i(23910) := b"1111111111111111_1111111111111111_1101110000110000_0011101101111110"; -- -0.139889032211261
	pesos_i(23911) := b"1111111111111111_1111111111111111_1101111010010000_0000001111110000"; -- -0.13061499965376835
	pesos_i(23912) := b"1111111111111111_1111111111111111_1101110011101000_0000101101010111"; -- -0.13708428514263318
	pesos_i(23913) := b"1111111111111111_1111111111111111_1111100100000011_1100010110000110"; -- -0.027286200215765534
	pesos_i(23914) := b"1111111111111111_1111111111111111_1110110000110100_1101111000010010"; -- -0.07731830644295296
	pesos_i(23915) := b"1111111111111111_1111111111111111_1110010100011101_0100111010011101"; -- -0.10502155946457956
	pesos_i(23916) := b"0000000000000000_0000000000000000_0001010111000000_0000101000110100"; -- 0.08496154565494718
	pesos_i(23917) := b"1111111111111111_1111111111111111_1101101111000101_1100101100101010"; -- -0.14151315899099212
	pesos_i(23918) := b"0000000000000000_0000000000000000_0010001101011000_0101101101000111"; -- 0.13806696388585832
	pesos_i(23919) := b"1111111111111111_1111111111111111_1110111101000011_0101101110000000"; -- -0.06537845739494988
	pesos_i(23920) := b"0000000000000000_0000000000000000_0001000110010001_0111000100011111"; -- 0.06862551693649627
	pesos_i(23921) := b"1111111111111111_1111111111111111_1110011101011000_0100001000000011"; -- -0.0963095420004547
	pesos_i(23922) := b"0000000000000000_0000000000000000_0001111010001100_0011010111011010"; -- 0.11932694023286301
	pesos_i(23923) := b"1111111111111111_1111111111111111_1111111110011110_0111110011000111"; -- -0.001487923967702926
	pesos_i(23924) := b"0000000000000000_0000000000000000_0001101100010000_1111101000101011"; -- 0.10572780179159191
	pesos_i(23925) := b"0000000000000000_0000000000000000_0010000000000110_0110001100001001"; -- 0.12509745560381838
	pesos_i(23926) := b"1111111111111111_1111111111111111_1110011000111001_0110001000010100"; -- -0.10068690311962974
	pesos_i(23927) := b"0000000000000000_0000000000000000_0000001101010001_1001100111011101"; -- 0.01296388293411574
	pesos_i(23928) := b"0000000000000000_0000000000000000_0000010110100001_1100111011101011"; -- 0.022000248421149296
	pesos_i(23929) := b"0000000000000000_0000000000000000_0001011010111011_0011110101010101"; -- 0.08879454932941042
	pesos_i(23930) := b"0000000000000000_0000000000000000_0001100000010000_0010001001100000"; -- 0.09399618957103395
	pesos_i(23931) := b"0000000000000000_0000000000000000_0010001000011001_0000000000001011"; -- 0.13319397219079462
	pesos_i(23932) := b"1111111111111111_1111111111111111_1110110111001001_1000000001011111"; -- -0.0711440819842224
	pesos_i(23933) := b"0000000000000000_0000000000000000_0000110001110111_1010101100000100"; -- 0.048700989249384534
	pesos_i(23934) := b"1111111111111111_1111111111111111_1110011101111001_0101010001101000"; -- -0.09580490559993758
	pesos_i(23935) := b"1111111111111111_1111111111111111_1110000001111010_0001010010011110"; -- -0.12313719885255611
	pesos_i(23936) := b"1111111111111111_1111111111111111_1110011101111010_0101001010001111"; -- -0.0957897568729185
	pesos_i(23937) := b"1111111111111111_1111111111111111_1111100111000001_0111101010000100"; -- -0.02439150114849884
	pesos_i(23938) := b"0000000000000000_0000000000000000_0001101010100101_1101000011010110"; -- 0.10409264782549302
	pesos_i(23939) := b"0000000000000000_0000000000000000_0000001000010111_0110111110100011"; -- 0.008170106130286318
	pesos_i(23940) := b"1111111111111111_1111111111111111_1111001010011010_0011010011001010"; -- -0.0523345000510019
	pesos_i(23941) := b"0000000000000000_0000000000000000_0000010010001010_0100010000001001"; -- 0.017734768057437147
	pesos_i(23942) := b"1111111111111111_1111111111111111_1101111010111101_1110101010011001"; -- -0.12991460585803705
	pesos_i(23943) := b"0000000000000000_0000000000000000_0010010110010010_1001000111010011"; -- 0.14676772489444903
	pesos_i(23944) := b"1111111111111111_1111111111111111_1101101001000000_0000000000101110"; -- -0.1474609267967693
	pesos_i(23945) := b"0000000000000000_0000000000000000_0010001010011111_1010110011010000"; -- 0.13524894783820848
	pesos_i(23946) := b"0000000000000000_0000000000000000_0001000111100100_1110001001001111"; -- 0.06989874296470762
	pesos_i(23947) := b"1111111111111111_1111111111111111_1110011110000001_0011001111000000"; -- -0.09568478158600796
	pesos_i(23948) := b"1111111111111111_1111111111111111_1111111110000011_0100110110010101"; -- -0.001902724492606874
	pesos_i(23949) := b"1111111111111111_1111111111111111_1110011100000011_1011111101100111"; -- -0.0975990650837636
	pesos_i(23950) := b"0000000000000000_0000000000000000_0000101000010000_0011101110010100"; -- 0.03931019182494784
	pesos_i(23951) := b"1111111111111111_1111111111111111_1111010001000100_1110001000110101"; -- -0.0458239194499544
	pesos_i(23952) := b"1111111111111111_1111111111111111_1111001101110110_1000111000100100"; -- -0.04897224061766506
	pesos_i(23953) := b"1111111111111111_1111111111111111_1110110111001110_1110110001110011"; -- -0.07106134596325518
	pesos_i(23954) := b"1111111111111111_1111111111111111_1111001000010111_1001010110000100"; -- -0.05432763603115092
	pesos_i(23955) := b"0000000000000000_0000000000000000_0001111010100101_0100111011100000"; -- 0.11970990160067407
	pesos_i(23956) := b"0000000000000000_0000000000000000_0000000101100101_0011101110010111"; -- 0.005450939484950172
	pesos_i(23957) := b"1111111111111111_1111111111111111_1110101111011011_0011010101000011"; -- -0.07868640051455504
	pesos_i(23958) := b"1111111111111111_1111111111111111_1101110101110000_1001101100011011"; -- -0.1350005206188504
	pesos_i(23959) := b"0000000000000000_0000000000000000_0000100000000110_1100100000010000"; -- 0.03135347729280316
	pesos_i(23960) := b"1111111111111111_1111111111111111_1110110101111011_0100010111001000"; -- -0.07233775967118294
	pesos_i(23961) := b"1111111111111111_1111111111111111_1111000011001000_0010011101111000"; -- -0.05944588966574552
	pesos_i(23962) := b"1111111111111111_1111111111111111_1101101111101011_1011100011100111"; -- -0.14093441351475847
	pesos_i(23963) := b"0000000000000000_0000000000000000_0001100010100111_0101010010101100"; -- 0.09630326455582987
	pesos_i(23964) := b"1111111111111111_1111111111111111_1101110110110111_0011011100000100"; -- -0.13392311231487303
	pesos_i(23965) := b"1111111111111111_1111111111111111_1111001010000101_0000000001111110"; -- -0.05265805178219841
	pesos_i(23966) := b"0000000000000000_0000000000000000_0001100101010110_1011011110011101"; -- 0.09897945005429634
	pesos_i(23967) := b"1111111111111111_1111111111111111_1110001000010101_1101011100100100"; -- -0.11685424214135842
	pesos_i(23968) := b"0000000000000000_0000000000000000_0000011100011011_1010000111110110"; -- 0.027765390924180126
	pesos_i(23969) := b"0000000000000000_0000000000000000_0001001110100101_1101001000101110"; -- 0.07674897782013863
	pesos_i(23970) := b"0000000000000000_0000000000000000_0001110010011111_1010100110110000"; -- 0.111811261509686
	pesos_i(23971) := b"1111111111111111_1111111111111111_1110000111110101_1101011110101110"; -- -0.117342491155734
	pesos_i(23972) := b"1111111111111111_1111111111111111_1110010101010110_0110001000101101"; -- -0.10415064243984459
	pesos_i(23973) := b"1111111111111111_1111111111111111_1110001000001010_0001110011100010"; -- -0.11703319058776362
	pesos_i(23974) := b"0000000000000000_0000000000000000_0000101110010101_0011111101011010"; -- 0.0452460856374116
	pesos_i(23975) := b"1111111111111111_1111111111111111_1101111010010001_0010011011111001"; -- -0.13059765256659156
	pesos_i(23976) := b"0000000000000000_0000000000000000_0001110010011110_0111110100110001"; -- 0.1117933506704223
	pesos_i(23977) := b"1111111111111111_1111111111111111_1101111011111100_1101001001110111"; -- -0.1289547404535756
	pesos_i(23978) := b"0000000000000000_0000000000000000_0001111001101010_0010110101110010"; -- 0.1188076402967638
	pesos_i(23979) := b"1111111111111111_1111111111111111_1110101010110101_0100000111111000"; -- -0.0831717271008018
	pesos_i(23980) := b"0000000000000000_0000000000000000_0001010100010001_0100111100101111"; -- 0.08229536914180742
	pesos_i(23981) := b"0000000000000000_0000000000000000_0000111001011111_0101010011001100"; -- 0.056142139356865774
	pesos_i(23982) := b"0000000000000000_0000000000000000_0001101000000010_1110001110011100"; -- 0.10160658409306397
	pesos_i(23983) := b"1111111111111111_1111111111111111_1110000110010110_0111000101101011"; -- -0.11879817129069266
	pesos_i(23984) := b"0000000000000000_0000000000000000_0001001010000101_1110000101111101"; -- 0.07235535900547808
	pesos_i(23985) := b"1111111111111111_1111111111111111_1101101011111001_1111001111010001"; -- -0.14462352889840496
	pesos_i(23986) := b"1111111111111111_1111111111111111_1110001100011001_1011110101011101"; -- -0.1128884932388369
	pesos_i(23987) := b"1111111111111111_1111111111111111_1110110100001010_1100010001010000"; -- -0.07405446106962332
	pesos_i(23988) := b"1111111111111111_1111111111111111_1110010110010010_0101110111010100"; -- -0.10323537414505725
	pesos_i(23989) := b"0000000000000000_0000000000000000_0001111010100111_0011110101010111"; -- 0.11973937399043685
	pesos_i(23990) := b"0000000000000000_0000000000000000_0010000010011001_1001000000011010"; -- 0.12734318391033497
	pesos_i(23991) := b"1111111111111111_1111111111111111_1110111011110011_0111000001101101"; -- -0.06659791313850727
	pesos_i(23992) := b"1111111111111111_1111111111111111_1110001100101101_1000011011001100"; -- -0.11258657004077642
	pesos_i(23993) := b"0000000000000000_0000000000000000_0000001010100011_1010101100000100"; -- 0.01030987598095114
	pesos_i(23994) := b"1111111111111111_1111111111111111_1111111101110101_1100111011011000"; -- -0.0021086427182921124
	pesos_i(23995) := b"1111111111111111_1111111111111111_1110111111101001_1010001001000110"; -- -0.06284127985650097
	pesos_i(23996) := b"0000000000000000_0000000000000000_0000010000100110_0110001101100011"; -- 0.01621075798731948
	pesos_i(23997) := b"1111111111111111_1111111111111111_1110101001001111_1000010101111000"; -- -0.08472410037166332
	pesos_i(23998) := b"1111111111111111_1111111111111111_1110010101000011_0110000010001100"; -- -0.10444065646966451
	pesos_i(23999) := b"0000000000000000_0000000000000000_0000101110101110_1001111011100101"; -- 0.04563325009960438
	pesos_i(24000) := b"1111111111111111_1111111111111111_1110111110110111_1100000011111110"; -- -0.0636023882824889
	pesos_i(24001) := b"1111111111111111_1111111111111111_1111100010001111_1010110000111010"; -- -0.029057727674656215
	pesos_i(24002) := b"0000000000000000_0000000000000000_0001000011101001_1110001001100001"; -- 0.06606879115576247
	pesos_i(24003) := b"0000000000000000_0000000000000000_0001101110010000_1100100001101110"; -- 0.1076779621117022
	pesos_i(24004) := b"1111111111111111_1111111111111111_1111111100011100_1010000000111100"; -- -0.003469453079204291
	pesos_i(24005) := b"1111111111111111_1111111111111111_1111011011110110_1000000100011100"; -- -0.03530114232251304
	pesos_i(24006) := b"0000000000000000_0000000000000000_0000110010101100_0100000000111001"; -- 0.04950333977536386
	pesos_i(24007) := b"1111111111111111_1111111111111111_1110110111010111_0110011101110011"; -- -0.07093194426182507
	pesos_i(24008) := b"1111111111111111_1111111111111111_1110100000000011_1100000000001011"; -- -0.0936927768691958
	pesos_i(24009) := b"0000000000000000_0000000000000000_0000010111111111_1110111111001101"; -- 0.02343653449881563
	pesos_i(24010) := b"1111111111111111_1111111111111111_1110010111000110_1111110001111110"; -- -0.10243245997926503
	pesos_i(24011) := b"0000000000000000_0000000000000000_0010010000101100_1110101100010001"; -- 0.1413103978335473
	pesos_i(24012) := b"0000000000000000_0000000000000000_0010010101110100_1011111001001011"; -- 0.1463126119141191
	pesos_i(24013) := b"1111111111111111_1111111111111111_1111000100000111_1000001101101101"; -- -0.058479104876188875
	pesos_i(24014) := b"0000000000000000_0000000000000000_0001000101111000_1001010010110001"; -- 0.06824616742324743
	pesos_i(24015) := b"0000000000000000_0000000000000000_0001100100000010_0100101100110101"; -- 0.09769125025115312
	pesos_i(24016) := b"0000000000000000_0000000000000000_0001110010101010_0011011110001101"; -- 0.11197230521345233
	pesos_i(24017) := b"1111111111111111_1111111111111111_1111000110110001_0000000011101101"; -- -0.05589288912216067
	pesos_i(24018) := b"1111111111111111_1111111111111111_1110001101111100_0011011111110010"; -- -0.11138582546428094
	pesos_i(24019) := b"0000000000000000_0000000000000000_0001001110000110_1110001111100111"; -- 0.07627701171056687
	pesos_i(24020) := b"0000000000000000_0000000000000000_0000100110000000_1101011000001000"; -- 0.037122132231028615
	pesos_i(24021) := b"1111111111111111_1111111111111111_1110010000010100_1100010011011011"; -- -0.10905809062742446
	pesos_i(24022) := b"1111111111111111_1111111111111111_1101100011000101_0111100011110000"; -- -0.15323681022556837
	pesos_i(24023) := b"1111111111111111_1111111111111111_1101100110110101_1101010011000110"; -- -0.14956922691388347
	pesos_i(24024) := b"0000000000000000_0000000000000000_0001110111010101_1001001100100101"; -- 0.11654014247555126
	pesos_i(24025) := b"1111111111111111_1111111111111111_1101100000101011_1000100111110110"; -- -0.15558564901805302
	pesos_i(24026) := b"0000000000000000_0000000000000000_0000001101011111_0110011100011101"; -- 0.013174480991780523
	pesos_i(24027) := b"0000000000000000_0000000000000000_0000010001110010_0110010111000101"; -- 0.017370567995289108
	pesos_i(24028) := b"0000000000000000_0000000000000000_0000001010110100_1010101001100010"; -- 0.010569237715065334
	pesos_i(24029) := b"1111111111111111_1111111111111111_1111010011101011_1110010011001110"; -- -0.043275546850325565
	pesos_i(24030) := b"1111111111111111_1111111111111111_1101111011100010_1110010110101100"; -- -0.1293503242652433
	pesos_i(24031) := b"1111111111111111_1111111111111111_1101111110100100_1111011100100101"; -- -0.12638907754474163
	pesos_i(24032) := b"1111111111111111_1111111111111111_1101111100110101_0011010110100000"; -- -0.1280943379526259
	pesos_i(24033) := b"0000000000000000_0000000000000000_0000100011110010_0001001101110100"; -- 0.03494378655953445
	pesos_i(24034) := b"1111111111111111_1111111111111111_1110111010110001_1100001001000110"; -- -0.06760011474981108
	pesos_i(24035) := b"1111111111111111_1111111111111111_1111000111011001_1110101000100010"; -- -0.055268637355860406
	pesos_i(24036) := b"1111111111111111_1111111111111111_1111010111000010_0000101011101010"; -- -0.04000789433689485
	pesos_i(24037) := b"1111111111111111_1111111111111111_1110100000100100_0011000000101000"; -- -0.09319781314292806
	pesos_i(24038) := b"1111111111111111_1111111111111111_1110111000110110_0001100111110011"; -- -0.06948697873392842
	pesos_i(24039) := b"1111111111111111_1111111111111111_1111110011100000_0111000001011110"; -- -0.012200333538081367
	pesos_i(24040) := b"1111111111111111_1111111111111111_1110001000001000_1110101011100000"; -- -0.11705143010049844
	pesos_i(24041) := b"0000000000000000_0000000000000000_0000011001100000_1010011000000011"; -- 0.024912238935513198
	pesos_i(24042) := b"1111111111111111_1111111111111111_1110000100101111_0001111000010110"; -- -0.12037479368684914
	pesos_i(24043) := b"1111111111111111_1111111111111111_1110010111100101_0011100000011001"; -- -0.10197114371853716
	pesos_i(24044) := b"0000000000000000_0000000000000000_0001111001011110_0110011101010101"; -- 0.11862798527852526
	pesos_i(24045) := b"0000000000000000_0000000000000000_0010011001001011_1100110000101011"; -- 0.1495940785846603
	pesos_i(24046) := b"0000000000000000_0000000000000000_0000110100000011_1000000010000001"; -- 0.050834685737484835
	pesos_i(24047) := b"1111111111111111_1111111111111111_1111001010100011_0001010110101011"; -- -0.05219902579643795
	pesos_i(24048) := b"1111111111111111_1111111111111111_1111110010000101_0111000011000001"; -- -0.013588860514474261
	pesos_i(24049) := b"1111111111111111_1111111111111111_1110000100101011_0110000101100101"; -- -0.12043181692659968
	pesos_i(24050) := b"1111111111111111_1111111111111111_1111000001111100_0110011111111100"; -- -0.06060171226221294
	pesos_i(24051) := b"0000000000000000_0000000000000000_0000000011111001_1001101110111011"; -- 0.0038087206583266144
	pesos_i(24052) := b"1111111111111111_1111111111111111_1111011101000100_1101101011000101"; -- -0.03410561257580938
	pesos_i(24053) := b"0000000000000000_0000000000000000_0000010110001110_1010001110001111"; -- 0.021707746785580774
	pesos_i(24054) := b"1111111111111111_1111111111111111_1111100000100101_1111100101001110"; -- -0.030670565024713537
	pesos_i(24055) := b"0000000000000000_0000000000000000_0001101001011101_0011011101010001"; -- 0.10298486453655203
	pesos_i(24056) := b"0000000000000000_0000000000000000_0000011101001001_0111101111110000"; -- 0.028465028863821813
	pesos_i(24057) := b"0000000000000000_0000000000000000_0001000110100010_1100011000100001"; -- 0.06888998330836966
	pesos_i(24058) := b"0000000000000000_0000000000000000_0001110110000111_0101001000011101"; -- 0.11534608094234582
	pesos_i(24059) := b"0000000000000000_0000000000000000_0010000100111100_1000010010010000"; -- 0.12982967868324116
	pesos_i(24060) := b"0000000000000000_0000000000000000_0001110001110010_1001001001101100"; -- 0.11112322947493307
	pesos_i(24061) := b"0000000000000000_0000000000000000_0001011001011000_1011010110000100"; -- 0.08729109251613273
	pesos_i(24062) := b"1111111111111111_1111111111111111_1110100011001111_0101000101000010"; -- -0.09058658731295471
	pesos_i(24063) := b"0000000000000000_0000000000000000_0000110111000010_0010101101111001"; -- 0.053744046321244736
	pesos_i(24064) := b"0000000000000000_0000000000000000_0001000101100101_1010000111111001"; -- 0.06795704207783869
	pesos_i(24065) := b"0000000000000000_0000000000000000_0000111110111101_1011101101110110"; -- 0.06148883471359984
	pesos_i(24066) := b"1111111111111111_1111111111111111_1110010110001101_1000110100000111"; -- -0.10330885492634945
	pesos_i(24067) := b"1111111111111111_1111111111111111_1111001011001011_1001001111100011"; -- -0.05158115108066997
	pesos_i(24068) := b"1111111111111111_1111111111111111_1111111110110100_1001001101000011"; -- -0.0011508905404597936
	pesos_i(24069) := b"0000000000000000_0000000000000000_0001000011101101_0000101000010111"; -- 0.06611693433936881
	pesos_i(24070) := b"1111111111111111_1111111111111111_1110010111000100_0100011110011111"; -- -0.10247375827774159
	pesos_i(24071) := b"0000000000000000_0000000000000000_0001011000111101_1001100110110011"; -- 0.08687744721781569
	pesos_i(24072) := b"1111111111111111_1111111111111111_1111101011110110_0111110010010110"; -- -0.019676411961182926
	pesos_i(24073) := b"1111111111111111_1111111111111111_1110000111101110_1000000011001001"; -- -0.1174544820003627
	pesos_i(24074) := b"0000000000000000_0000000000000000_0000100000111010_0011100101000001"; -- 0.03213842240248128
	pesos_i(24075) := b"0000000000000000_0000000000000000_0001100111011011_0011011001110111"; -- 0.10100117108852938
	pesos_i(24076) := b"0000000000000000_0000000000000000_0010110001010100_0001110101111010"; -- 0.17315849526405833
	pesos_i(24077) := b"1111111111111111_1111111111111111_1111011110101011_1110010001110000"; -- -0.0325333810752951
	pesos_i(24078) := b"0000000000000000_0000000000000000_0000100001000000_1011111111110111"; -- 0.0322380044237784
	pesos_i(24079) := b"1111111111111111_1111111111111111_1111111110100011_1110011011011111"; -- -0.001405306344451125
	pesos_i(24080) := b"1111111111111111_1111111111111111_1110000001010001_0000011100111111"; -- -0.12376360613563178
	pesos_i(24081) := b"0000000000000000_0000000000000000_0001111000000010_1110011110111110"; -- 0.11723183041897285
	pesos_i(24082) := b"0000000000000000_0000000000000000_0000001001110010_1101101111010110"; -- 0.00956510522429474
	pesos_i(24083) := b"1111111111111111_1111111111111111_1101110110001011_1011101000011011"; -- -0.13458668560272125
	pesos_i(24084) := b"1111111111111111_1111111111111111_1110011010000010_0100101001101011"; -- -0.09957442165719732
	pesos_i(24085) := b"1111111111111111_1111111111111111_1101110011011011_1010111011110100"; -- -0.13727289721578967
	pesos_i(24086) := b"1111111111111111_1111111111111111_1110001011010100_0110110101010010"; -- -0.11394612062041459
	pesos_i(24087) := b"1111111111111111_1111111111111111_1110001110011110_0000101001000010"; -- -0.11086974993591239
	pesos_i(24088) := b"1111111111111111_1111111111111111_1111100110100000_0000101111010011"; -- -0.024901639067413897
	pesos_i(24089) := b"0000000000000000_0000000000000000_0000101100011000_0110010011010010"; -- 0.0433409702406361
	pesos_i(24090) := b"1111111111111111_1111111111111111_1110000011111010_0100010000110011"; -- -0.12118123776361962
	pesos_i(24091) := b"1111111111111111_1111111111111111_1110111001101111_1110011010011011"; -- -0.0686050293711696
	pesos_i(24092) := b"1111111111111111_1111111111111111_1111010110110011_0101110010001010"; -- -0.04023191097479183
	pesos_i(24093) := b"1111111111111111_1111111111111111_1110001001011111_1111111010000101"; -- -0.115722744411662
	pesos_i(24094) := b"1111111111111111_1111111111111111_1111101000001110_0001000001010100"; -- -0.023222903612857126
	pesos_i(24095) := b"0000000000000000_0000000000000000_0000111000101000_1011100011110111"; -- 0.05530887633625799
	pesos_i(24096) := b"0000000000000000_0000000000000000_0001011100110111_1101010000100111"; -- 0.09069562865954861
	pesos_i(24097) := b"0000000000000000_0000000000000000_0000110001110010_0001100001111011"; -- 0.04861596120798842
	pesos_i(24098) := b"0000000000000000_0000000000000000_0000101011110100_1111110111010011"; -- 0.042800773650854135
	pesos_i(24099) := b"0000000000000000_0000000000000000_0000111011001001_0000001101000001"; -- 0.05775471050503163
	pesos_i(24100) := b"1111111111111111_1111111111111111_1110111111100111_0111101011110101"; -- -0.062874140874635
	pesos_i(24101) := b"1111111111111111_1111111111111111_1101111111001110_0011111100101111"; -- -0.1257591734272657
	pesos_i(24102) := b"1111111111111111_1111111111111111_1111001000110000_0011010110111001"; -- -0.05395187602043649
	pesos_i(24103) := b"1111111111111111_1111111111111111_1111101000110000_1011000110010001"; -- -0.022694494296137933
	pesos_i(24104) := b"0000000000000000_0000000000000000_0010000011100111_1100010111110100"; -- 0.1285365792436443
	pesos_i(24105) := b"0000000000000000_0000000000000000_0000101111000100_0101011001000111"; -- 0.04596461507341315
	pesos_i(24106) := b"1111111111111111_1111111111111111_1111001001110000_0000111110010010"; -- -0.052977587576182573
	pesos_i(24107) := b"0000000000000000_0000000000000000_0000110000011100_1110110101011001"; -- 0.047316393229666596
	pesos_i(24108) := b"1111111111111111_1111111111111111_1111101100110001_1111101111010111"; -- -0.01876855844630894
	pesos_i(24109) := b"1111111111111111_1111111111111111_1101111100111111_0111010011101110"; -- -0.12793797682149444
	pesos_i(24110) := b"0000000000000000_0000000000000000_0001011110010001_1011110111011011"; -- 0.09206759064254194
	pesos_i(24111) := b"1111111111111111_1111111111111111_1110101100101110_0000110100110111"; -- -0.08132855803977594
	pesos_i(24112) := b"1111111111111111_1111111111111111_1111010110110010_1010110011001110"; -- -0.04024238548395925
	pesos_i(24113) := b"0000000000000000_0000000000000000_0000100101101111_1010101101010100"; -- 0.036860187579772434
	pesos_i(24114) := b"1111111111111111_1111111111111111_1110011011110011_0011110011010001"; -- -0.09785098926039415
	pesos_i(24115) := b"0000000000000000_0000000000000000_0000011111111101_0110100000010010"; -- 0.03121042660701524
	pesos_i(24116) := b"1111111111111111_1111111111111111_1111111101011110_1111101101000001"; -- -0.00245694790282448
	pesos_i(24117) := b"0000000000000000_0000000000000000_0001011011010011_0010101000001100"; -- 0.08915961072039813
	pesos_i(24118) := b"0000000000000000_0000000000000000_0000101011011011_1000111000001110"; -- 0.042412641939284935
	pesos_i(24119) := b"1111111111111111_1111111111111111_1110011101011011_1110110001001001"; -- -0.09625361640636265
	pesos_i(24120) := b"0000000000000000_0000000000000000_0001000110110111_0001011110000101"; -- 0.06920001016948353
	pesos_i(24121) := b"1111111111111111_1111111111111111_1111110100110010_1010001011010101"; -- -0.010946105026243779
	pesos_i(24122) := b"1111111111111111_1111111111111111_1111010111111100_0111100000011100"; -- -0.03911637599751453
	pesos_i(24123) := b"1111111111111111_1111111111111111_1110001010001001_1111001011100100"; -- -0.11508256844708259
	pesos_i(24124) := b"1111111111111111_1111111111111111_1110101100101010_0110011101001110"; -- -0.08138422348178022
	pesos_i(24125) := b"0000000000000000_0000000000000000_0000000010001101_1000111101001000"; -- 0.0021600294998645703
	pesos_i(24126) := b"1111111111111111_1111111111111111_1101101110011110_1111001000111000"; -- -0.14210592398496857
	pesos_i(24127) := b"1111111111111111_1111111111111111_1101100000101100_1101111001101001"; -- -0.15556535653933787
	pesos_i(24128) := b"0000000000000000_0000000000000000_0000010100111010_1110111111111110"; -- 0.02043056435803281
	pesos_i(24129) := b"0000000000000000_0000000000000000_0001110001101001_1000111000000000"; -- 0.11098563678270976
	pesos_i(24130) := b"1111111111111111_1111111111111111_1111100110110111_1101001111000110"; -- -0.024538769008785263
	pesos_i(24131) := b"1111111111111111_1111111111111111_1111001001000110_1010001001100101"; -- -0.053609705357238
	pesos_i(24132) := b"1111111111111111_1111111111111111_1101100000000111_1100000011000110"; -- -0.15613169838282848
	pesos_i(24133) := b"0000000000000000_0000000000000000_0001001010001100_1010000011001111"; -- 0.07245831549514943
	pesos_i(24134) := b"0000000000000000_0000000000000000_0001101001000011_1110101101110110"; -- 0.10259887346367086
	pesos_i(24135) := b"0000000000000000_0000000000000000_0001111010000101_1110100000111100"; -- 0.1192307612930169
	pesos_i(24136) := b"0000000000000000_0000000000000000_0001111010100010_0100011111101001"; -- 0.1196637099426048
	pesos_i(24137) := b"0000000000000000_0000000000000000_0000100011000000_0111101000100001"; -- 0.034186966931161654
	pesos_i(24138) := b"1111111111111111_1111111111111111_1110001011110110_0010011011011000"; -- -0.11343152271801293
	pesos_i(24139) := b"0000000000000000_0000000000000000_0000110010100100_0111011101110011"; -- 0.04938456102727726
	pesos_i(24140) := b"0000000000000000_0000000000000000_0000100011100010_1010011100101111"; -- 0.03470845134776443
	pesos_i(24141) := b"1111111111111111_1111111111111111_1111001000111001_0001101001011101"; -- -0.0538161777039499
	pesos_i(24142) := b"1111111111111111_1111111111111111_1111110001000010_1110000000101100"; -- -0.014604558211886423
	pesos_i(24143) := b"0000000000000000_0000000000000000_0001011000001101_0100111110001111"; -- 0.08614060634414573
	pesos_i(24144) := b"1111111111111111_1111111111111111_1101111100100110_1010000101000010"; -- -0.1283168042985601
	pesos_i(24145) := b"1111111111111111_1111111111111111_1110100010011111_0100010010111101"; -- -0.09131975535949236
	pesos_i(24146) := b"0000000000000000_0000000000000000_0000001101110100_1001010100111101"; -- 0.01349766472611107
	pesos_i(24147) := b"1111111111111111_1111111111111111_1111100001100101_0000100100001001"; -- -0.029708323673941252
	pesos_i(24148) := b"0000000000000000_0000000000000000_0001001110010111_0001011110010000"; -- 0.07652423160258617
	pesos_i(24149) := b"0000000000000000_0000000000000000_0001111011110000_0101000001110111"; -- 0.12085440550578089
	pesos_i(24150) := b"0000000000000000_0000000000000000_0001000111001100_0111110111111011"; -- 0.0695265520060514
	pesos_i(24151) := b"0000000000000000_0000000000000000_0001111011101001_0010001101000110"; -- 0.12074490038153005
	pesos_i(24152) := b"1111111111111111_1111111111111111_1101100011000111_1000111010011010"; -- -0.15320500120860064
	pesos_i(24153) := b"0000000000000000_0000000000000000_0010010110001010_0010101001011101"; -- 0.14663948803294807
	pesos_i(24154) := b"0000000000000000_0000000000000000_0000001100100000_0001001100000101"; -- 0.012208164830946543
	pesos_i(24155) := b"0000000000000000_0000000000000000_0001000011101011_0001101000001100"; -- 0.06608736800019448
	pesos_i(24156) := b"0000000000000000_0000000000000000_0001011011000100_0010010001111001"; -- 0.08893039666772473
	pesos_i(24157) := b"1111111111111111_1111111111111111_1111010101000101_1011110110001110"; -- -0.04190459525860853
	pesos_i(24158) := b"1111111111111111_1111111111111111_1110010011111110_1101100111111011"; -- -0.1054862749354399
	pesos_i(24159) := b"1111111111111111_1111111111111111_1110111001111101_0110110011010010"; -- -0.06839866522181268
	pesos_i(24160) := b"0000000000000000_0000000000000000_0001101100011101_0101000011110000"; -- 0.10591607905083743
	pesos_i(24161) := b"0000000000000000_0000000000000000_0000101011010100_1101101010100110"; -- 0.0423103956850114
	pesos_i(24162) := b"0000000000000000_0000000000000000_0001100111110000_0101010110000000"; -- 0.1013234556691368
	pesos_i(24163) := b"0000000000000000_0000000000000000_0000101010000000_1101100100111001"; -- 0.04102857238171208
	pesos_i(24164) := b"1111111111111111_1111111111111111_1111000111101001_0100111110111000"; -- -0.0550337004306657
	pesos_i(24165) := b"0000000000000000_0000000000000000_0000101000010010_0110111000000001"; -- 0.03934371494773362
	pesos_i(24166) := b"0000000000000000_0000000000000000_0001010100010111_0101000110100010"; -- 0.0823870679525317
	pesos_i(24167) := b"0000000000000000_0000000000000000_0000101001000010_1011100010111010"; -- 0.04008059056996476
	pesos_i(24168) := b"1111111111111111_1111111111111111_1110110011010010_1000000110110101"; -- -0.07491292308345429
	pesos_i(24169) := b"0000000000000000_0000000000000000_0010001010011000_0110000101001000"; -- 0.13513763434474205
	pesos_i(24170) := b"0000000000000000_0000000000000000_0000011100111101_0001010111001101"; -- 0.028275835596595623
	pesos_i(24171) := b"1111111111111111_1111111111111111_1111001111111010_1101011000100000"; -- -0.04695378983963759
	pesos_i(24172) := b"0000000000000000_0000000000000000_0001010011000100_0100010000110010"; -- 0.0811197874645844
	pesos_i(24173) := b"0000000000000000_0000000000000000_0000011111000111_0011010101100100"; -- 0.030383431416184298
	pesos_i(24174) := b"1111111111111111_1111111111111111_1111010000011010_0000111010000000"; -- -0.0464774071143413
	pesos_i(24175) := b"1111111111111111_1111111111111111_1110100100100110_1100101001011010"; -- -0.0892518550324978
	pesos_i(24176) := b"0000000000000000_0000000000000000_0001110000101011_0111000010100000"; -- 0.11003784078729115
	pesos_i(24177) := b"1111111111111111_1111111111111111_1110011111011101_1000011100001111"; -- -0.09427600740630601
	pesos_i(24178) := b"1111111111111111_1111111111111111_1101010111001110_1101000010100000"; -- -0.16481300433566776
	pesos_i(24179) := b"1111111111111111_1111111111111111_1110011101110110_0111011101000011"; -- -0.09584860441312665
	pesos_i(24180) := b"0000000000000000_0000000000000000_0000001101101101_0110000100011100"; -- 0.013387746179800819
	pesos_i(24181) := b"1111111111111111_1111111111111111_1110011000100101_0011111001101011"; -- -0.1009942045174645
	pesos_i(24182) := b"1111111111111111_1111111111111111_1101101010100110_0110010101001111"; -- -0.14589850261660067
	pesos_i(24183) := b"1111111111111111_1111111111111111_1111001111001010_0100101100100100"; -- -0.047694495781344104
	pesos_i(24184) := b"0000000000000000_0000000000000000_0010001110111101_1011110001010011"; -- 0.13961388617791354
	pesos_i(24185) := b"1111111111111111_1111111111111111_1111001111001001_0010000111011010"; -- -0.047712215691874595
	pesos_i(24186) := b"1111111111111111_1111111111111111_1101101011100001_0111001010101101"; -- -0.14499743722091804
	pesos_i(24187) := b"0000000000000000_0000000000000000_0010001001101111_1010001101001110"; -- 0.13451595929320254
	pesos_i(24188) := b"1111111111111111_1111111111111111_1110001000000101_1011111100101010"; -- -0.11709981185433777
	pesos_i(24189) := b"0000000000000000_0000000000000000_0010011000011010_0110000110010001"; -- 0.14884004391721145
	pesos_i(24190) := b"1111111111111111_1111111111111111_1101101011010110_1010010011110001"; -- -0.14516228784160026
	pesos_i(24191) := b"1111111111111111_1111111111111111_1110100111001100_1110111111011111"; -- -0.08671665948715937
	pesos_i(24192) := b"0000000000000000_0000000000000000_0001000100101111_0000110000111100"; -- 0.06712414236753786
	pesos_i(24193) := b"1111111111111111_1111111111111111_1110100011101110_1110111100111010"; -- -0.09010414930154584
	pesos_i(24194) := b"0000000000000000_0000000000000000_0000101101111000_0000100010000111"; -- 0.044800312851549576
	pesos_i(24195) := b"1111111111111111_1111111111111111_1101110111111010_0010111001000011"; -- -0.13290129531782544
	pesos_i(24196) := b"1111111111111111_1111111111111111_1110011101011101_1110110000001011"; -- -0.09622311344015641
	pesos_i(24197) := b"0000000000000000_0000000000000000_0000000011101010_0000000000110011"; -- 0.0035705684958015917
	pesos_i(24198) := b"1111111111111111_1111111111111111_1101111101001011_0001100001001100"; -- -0.1277603926467656
	pesos_i(24199) := b"0000000000000000_0000000000000000_0001101101110110_0100101101101101"; -- 0.10727378291371416
	pesos_i(24200) := b"1111111111111111_1111111111111111_1101111011111010_1010010001110010"; -- -0.1289880010925865
	pesos_i(24201) := b"0000000000000000_0000000000000000_0001010100110010_1011110101100101"; -- 0.08280547823406806
	pesos_i(24202) := b"1111111111111111_1111111111111111_1111111010010101_1110001001010001"; -- -0.005525450944750744
	pesos_i(24203) := b"0000000000000000_0000000000000000_0000000111011000_0011110010110001"; -- 0.007205765861862082
	pesos_i(24204) := b"1111111111111111_1111111111111111_1110001100000010_0001000110100100"; -- -0.11324968107217653
	pesos_i(24205) := b"1111111111111111_1111111111111111_1110110111011001_0011011110000101"; -- -0.0709042834963045
	pesos_i(24206) := b"0000000000000000_0000000000000000_0010000000010011_1101110010101000"; -- 0.12530306920622084
	pesos_i(24207) := b"1111111111111111_1111111111111111_1110111110100101_1111001000010111"; -- -0.06387412018327658
	pesos_i(24208) := b"1111111111111111_1111111111111111_1111000111001000_0110001000011001"; -- -0.05553614502924441
	pesos_i(24209) := b"1111111111111111_1111111111111111_1111100000000101_0000111110100010"; -- -0.03117277420714402
	pesos_i(24210) := b"1111111111111111_1111111111111111_1101100010101011_0001001110100110"; -- -0.15363957604455306
	pesos_i(24211) := b"1111111111111111_1111111111111111_1101110101000100_0110101000011110"; -- -0.1356748273435717
	pesos_i(24212) := b"1111111111111111_1111111111111111_1101110001111101_1011110100011011"; -- -0.1387063798273471
	pesos_i(24213) := b"0000000000000000_0000000000000000_0010010100101101_1110001101111111"; -- 0.14523145529766882
	pesos_i(24214) := b"1111111111111111_1111111111111111_1110010100011010_1010010101100100"; -- -0.10506216349834584
	pesos_i(24215) := b"0000000000000000_0000000000000000_0000101100100011_0011001100111100"; -- 0.043505861355085954
	pesos_i(24216) := b"1111111111111111_1111111111111111_1110011000111111_0010011000110100"; -- -0.1005989192305312
	pesos_i(24217) := b"1111111111111111_1111111111111111_1111000000110100_1100010100010110"; -- -0.06169479565551434
	pesos_i(24218) := b"1111111111111111_1111111111111111_1110110011010010_1001100011010111"; -- -0.07491154433498572
	pesos_i(24219) := b"1111111111111111_1111111111111111_1110010110110011_0001010010001111"; -- -0.1027362013263379
	pesos_i(24220) := b"0000000000000000_0000000000000000_0001100000110111_1101111110111010"; -- 0.09460256860850075
	pesos_i(24221) := b"0000000000000000_0000000000000000_0001001111101110_1011100100111100"; -- 0.07786138274117521
	pesos_i(24222) := b"0000000000000000_0000000000000000_0010000011110111_0011001110101000"; -- 0.1287719998185305
	pesos_i(24223) := b"1111111111111111_1111111111111111_1110110100110110_0010100001110101"; -- -0.07339236386145653
	pesos_i(24224) := b"1111111111111111_1111111111111111_1111101100011100_0001001001011000"; -- -0.01910291058286852
	pesos_i(24225) := b"0000000000000000_0000000000000000_0000000011100111_1001010110101001"; -- 0.0035337008219869194
	pesos_i(24226) := b"1111111111111111_1111111111111111_1111011111001101_1000000100110111"; -- -0.032020496443297096
	pesos_i(24227) := b"1111111111111111_1111111111111111_1111011101011110_0110011110001010"; -- -0.0337157523944782
	pesos_i(24228) := b"0000000000000000_0000000000000000_0000111001001100_0010110100110001"; -- 0.055849861509506035
	pesos_i(24229) := b"0000000000000000_0000000000000000_0000110101010111_1010011110100100"; -- 0.052118756851012915
	pesos_i(24230) := b"1111111111111111_1111111111111111_1110101100101010_1010100001110101"; -- -0.08138034003312249
	pesos_i(24231) := b"0000000000000000_0000000000000000_0001100101101011_1011110100100110"; -- 0.09930021448939204
	pesos_i(24232) := b"0000000000000000_0000000000000000_0010000111101111_1000101101101101"; -- 0.13256141100015995
	pesos_i(24233) := b"0000000000000000_0000000000000000_0001011110011111_1011000011001010"; -- 0.09228043489577875
	pesos_i(24234) := b"1111111111111111_1111111111111111_1101100101101010_1011111111000010"; -- -0.15071488880316475
	pesos_i(24235) := b"1111111111111111_1111111111111111_1110010101010111_0011000100001110"; -- -0.10413831144924372
	pesos_i(24236) := b"1111111111111111_1111111111111111_1101110001011100_1000011000001100"; -- -0.13921320162908546
	pesos_i(24237) := b"1111111111111111_1111111111111111_1111011010111101_0000010011100111"; -- -0.0361782965863323
	pesos_i(24238) := b"0000000000000000_0000000000000000_0001101110011010_0111010100010010"; -- 0.10782558144543947
	pesos_i(24239) := b"0000000000000000_0000000000000000_0001001000001010_1100011110000111"; -- 0.07047698058188043
	pesos_i(24240) := b"1111111111111111_1111111111111111_1111110010010100_1001001100011001"; -- -0.013357931589555177
	pesos_i(24241) := b"0000000000000000_0000000000000000_0001001111010110_0011001111110111"; -- 0.07748722817776373
	pesos_i(24242) := b"1111111111111111_1111111111111111_1110101000101111_0110010011000100"; -- -0.085214330754129
	pesos_i(24243) := b"1111111111111111_1111111111111111_1111110010011011_0010000101110000"; -- -0.013257894587302078
	pesos_i(24244) := b"0000000000000000_0000000000000000_0000000111100110_0111110010110000"; -- 0.007423203323865223
	pesos_i(24245) := b"0000000000000000_0000000000000000_0010001010100010_0111101010100100"; -- 0.13529173371415815
	pesos_i(24246) := b"1111111111111111_1111111111111111_1111010101011101_0010100100101001"; -- -0.04154722932070723
	pesos_i(24247) := b"0000000000000000_0000000000000000_0010000101111111_0101001010111011"; -- 0.130849047235908
	pesos_i(24248) := b"1111111111111111_1111111111111111_1101111111000110_0001010101000101"; -- -0.12588374193033028
	pesos_i(24249) := b"0000000000000000_0000000000000000_0000100100010101_1110001011100101"; -- 0.035490208447456234
	pesos_i(24250) := b"1111111111111111_1111111111111111_1111011000111110_0111101100011001"; -- -0.03810911798254673
	pesos_i(24251) := b"1111111111111111_1111111111111111_1101101001100111_0010101111001100"; -- -0.1468632342785824
	pesos_i(24252) := b"0000000000000000_0000000000000000_0000110110011101_1000111111110111"; -- 0.053185460884908456
	pesos_i(24253) := b"1111111111111111_1111111111111111_1111001001001011_1110101110100101"; -- -0.05352904527659353
	pesos_i(24254) := b"1111111111111111_1111111111111111_1111100111011111_0011010101000011"; -- -0.023937865392791656
	pesos_i(24255) := b"1111111111111111_1111111111111111_1111111100001100_0111011000000010"; -- -0.003716110632926431
	pesos_i(24256) := b"1111111111111111_1111111111111111_1111101011010001_1010010101010000"; -- -0.020238559807025353
	pesos_i(24257) := b"1111111111111111_1111111111111111_1111101011011110_1111010110101010"; -- -0.020035406210348803
	pesos_i(24258) := b"1111111111111111_1111111111111111_1101100110000100_0011111111000000"; -- -0.15032579015046726
	pesos_i(24259) := b"1111111111111111_1111111111111111_1111010110111011_1110001110100111"; -- -0.04010178720547836
	pesos_i(24260) := b"1111111111111111_1111111111111111_1110110001100100_0100111001001100"; -- -0.07659445425002169
	pesos_i(24261) := b"0000000000000000_0000000000000000_0000111100010011_0000100010000001"; -- 0.058884173818409206
	pesos_i(24262) := b"1111111111111111_1111111111111111_1101100100001010_0100111001011101"; -- -0.15218649132761
	pesos_i(24263) := b"1111111111111111_1111111111111111_1110010010000100_1011011011001100"; -- -0.10734994441118073
	pesos_i(24264) := b"0000000000000000_0000000000000000_0001100010110001_1110010001011101"; -- 0.09646441713848197
	pesos_i(24265) := b"0000000000000000_0000000000000000_0001100111101001_0001101110011001"; -- 0.1012131926891
	pesos_i(24266) := b"1111111111111111_1111111111111111_1110110010000111_0010101100011100"; -- -0.07606249398529819
	pesos_i(24267) := b"0000000000000000_0000000000000000_0001001100000011_1000100000000001"; -- 0.07427263290443072
	pesos_i(24268) := b"0000000000000000_0000000000000000_0000011010101010_1111111111001101"; -- 0.026046741108107126
	pesos_i(24269) := b"1111111111111111_1111111111111111_1101101011110010_0100011010011110"; -- -0.14474066392856907
	pesos_i(24270) := b"0000000000000000_0000000000000000_0000110011101001_0101010001000000"; -- 0.05043531961503209
	pesos_i(24271) := b"1111111111111111_1111111111111111_1111011101100011_1110101110111001"; -- -0.03363157976665367
	pesos_i(24272) := b"0000000000000000_0000000000000000_0010100100111110_0101111001011000"; -- 0.16110791831770718
	pesos_i(24273) := b"1111111111111111_1111111111111111_1111000100111101_0101111010001111"; -- -0.05765732772778297
	pesos_i(24274) := b"0000000000000000_0000000000000000_0001111110001110_0010110100010111"; -- 0.12326318550893244
	pesos_i(24275) := b"0000000000000000_0000000000000000_0001011001010110_1100000001110110"; -- 0.08726122732444005
	pesos_i(24276) := b"1111111111111111_1111111111111111_1111111111011101_1111100101011110"; -- -0.0005191941934811756
	pesos_i(24277) := b"0000000000000000_0000000000000000_0001001111111011_0110101011011110"; -- 0.07805507580247942
	pesos_i(24278) := b"0000000000000000_0000000000000000_0001111001011101_0101001011100101"; -- 0.11861150838097319
	pesos_i(24279) := b"0000000000000000_0000000000000000_0001111011110101_1100111111110000"; -- 0.12093829736609839
	pesos_i(24280) := b"0000000000000000_0000000000000000_0001011001111001_1101111001001110"; -- 0.08779706385195436
	pesos_i(24281) := b"1111111111111111_1111111111111111_1110001011110001_1011100111000001"; -- -0.11349906009771936
	pesos_i(24282) := b"0000000000000000_0000000000000000_0010011111111010_0110111011011011"; -- 0.15616505470093878
	pesos_i(24283) := b"0000000000000000_0000000000000000_0000011011011010_1111110001101100"; -- 0.02677896156303486
	pesos_i(24284) := b"1111111111111111_1111111111111111_1111000110000011_0111011101111011"; -- -0.05658772694374015
	pesos_i(24285) := b"0000000000000000_0000000000000000_0001100110001110_1011100010111101"; -- 0.09983400919496062
	pesos_i(24286) := b"1111111111111111_1111111111111111_1101011111110010_0100000010010111"; -- -0.1564597730992922
	pesos_i(24287) := b"0000000000000000_0000000000000000_0001000100100101_0000111010010101"; -- 0.06697169438247218
	pesos_i(24288) := b"0000000000000000_0000000000000000_0010001101001001_1111111111101000"; -- 0.13784789469934486
	pesos_i(24289) := b"0000000000000000_0000000000000000_0000111000001110_0000011010111010"; -- 0.05490152388313969
	pesos_i(24290) := b"1111111111111111_1111111111111111_1101111100101011_0010100100100001"; -- -0.12824767054071143
	pesos_i(24291) := b"0000000000000000_0000000000000000_0001011011101001_1011011010010010"; -- 0.08950367994380672
	pesos_i(24292) := b"0000000000000000_0000000000000000_0000110010101101_1001011010100110"; -- 0.04952374978275154
	pesos_i(24293) := b"1111111111111111_1111111111111111_1110010111111011_0010001100111011"; -- -0.10163669413486277
	pesos_i(24294) := b"1111111111111111_1111111111111111_1101101100100111_0101110000110111"; -- -0.1439306608606437
	pesos_i(24295) := b"1111111111111111_1111111111111111_1110101111010011_1101000101110101"; -- -0.07879916100920992
	pesos_i(24296) := b"1111111111111111_1111111111111111_1111111011111011_1001101110100101"; -- -0.0039732668951226865
	pesos_i(24297) := b"0000000000000000_0000000000000000_0010000011011001_1001110001100010"; -- 0.12832047825390125
	pesos_i(24298) := b"0000000000000000_0000000000000000_0000000111010000_0000011100010111"; -- 0.007080500805321777
	pesos_i(24299) := b"1111111111111111_1111111111111111_1111111100000110_1111110100100001"; -- -0.0037996094908003776
	pesos_i(24300) := b"1111111111111111_1111111111111111_1110100000101001_0110000011000110"; -- -0.0931186215424848
	pesos_i(24301) := b"1111111111111111_1111111111111111_1111101111010010_1011000100100000"; -- -0.01631634677407169
	pesos_i(24302) := b"0000000000000000_0000000000000000_0010001010011111_0101010101100101"; -- 0.13524373739567258
	pesos_i(24303) := b"0000000000000000_0000000000000000_0001101001010011_1101011100000110"; -- 0.10284179586554243
	pesos_i(24304) := b"0000000000000000_0000000000000000_0000011111100111_0011000010111101"; -- 0.030871435196840283
	pesos_i(24305) := b"0000000000000000_0000000000000000_0001001101101011_1011000110101010"; -- 0.07586202999850007
	pesos_i(24306) := b"1111111111111111_1111111111111111_1110001101000100_0111011111010010"; -- -0.112236510489053
	pesos_i(24307) := b"0000000000000000_0000000000000000_0001110111000100_0111001001011001"; -- 0.11627878822519762
	pesos_i(24308) := b"1111111111111111_1111111111111111_1110110111111011_1101010100001100"; -- -0.07037609541418967
	pesos_i(24309) := b"0000000000000000_0000000000000000_0001010001110110_0101000001010001"; -- 0.07993032440210053
	pesos_i(24310) := b"0000000000000000_0000000000000000_0001011010111011_1111010100010101"; -- 0.08880550169334364
	pesos_i(24311) := b"1111111111111111_1111111111111111_1101110110100110_1010001001010110"; -- -0.13417611504703372
	pesos_i(24312) := b"1111111111111111_1111111111111111_1101110101100001_1111101101001001"; -- -0.1352236697514477
	pesos_i(24313) := b"0000000000000000_0000000000000000_0000000000011111_1111000011011110"; -- 0.0004873793572438779
	pesos_i(24314) := b"1111111111111111_1111111111111111_1111101101110010_0101100010001101"; -- -0.01778647001927936
	pesos_i(24315) := b"1111111111111111_1111111111111111_1101101000001001_0011100101100001"; -- -0.14829675087320124
	pesos_i(24316) := b"1111111111111111_1111111111111111_1111101111100111_1111011011100001"; -- -0.01599175451012368
	pesos_i(24317) := b"1111111111111111_1111111111111111_1110011001011001_1110011101110100"; -- -0.10019067206681019
	pesos_i(24318) := b"0000000000000000_0000000000000000_0000011101110101_1111110010010101"; -- 0.02914408339789896
	pesos_i(24319) := b"1111111111111111_1111111111111111_1111110011011110_0001100101000001"; -- -0.01223604365064234
	pesos_i(24320) := b"0000000000000000_0000000000000000_0000101011001001_1111011000110111"; -- 0.04214419211599412
	pesos_i(24321) := b"0000000000000000_0000000000000000_0000011110101111_0011110110000101"; -- 0.03001770502669405
	pesos_i(24322) := b"0000000000000000_0000000000000000_0001101101011001_0010100010011000"; -- 0.10682920176815712
	pesos_i(24323) := b"1111111111111111_1111111111111111_1110001010001111_1100011010110001"; -- -0.11499365018007035
	pesos_i(24324) := b"0000000000000000_0000000000000000_0001100010011101_1011000101110011"; -- 0.09615620670832908
	pesos_i(24325) := b"1111111111111111_1111111111111111_1111101010011110_1110001110000111"; -- -0.021013049671991614
	pesos_i(24326) := b"0000000000000000_0000000000000000_0001100101110101_1000001001001001"; -- 0.09944929401758687
	pesos_i(24327) := b"0000000000000000_0000000000000000_0000100101000110_0001010001000110"; -- 0.036225573733853114
	pesos_i(24328) := b"0000000000000000_0000000000000000_0010000111010000_0110000100010000"; -- 0.13208586346713744
	pesos_i(24329) := b"0000000000000000_0000000000000000_0010100000110101_1000111000101110"; -- 0.15706719034308472
	pesos_i(24330) := b"0000000000000000_0000000000000000_0000001000010110_1110001110101111"; -- 0.008161764399224456
	pesos_i(24331) := b"0000000000000000_0000000000000000_0000100001001101_1111110010101101"; -- 0.032439987408662115
	pesos_i(24332) := b"1111111111111111_1111111111111111_1110010001011100_1001110010110111"; -- -0.10796185038364604
	pesos_i(24333) := b"1111111111111111_1111111111111111_1110010111110010_0000101100011100"; -- -0.1017754607972559
	pesos_i(24334) := b"0000000000000000_0000000000000000_0000111111011101_0010001000111101"; -- 0.06196798304275742
	pesos_i(24335) := b"1111111111111111_1111111111111111_1110101110111100_1001101101000100"; -- -0.07915334301672798
	pesos_i(24336) := b"1111111111111111_1111111111111111_1101100101010110_1111101010110110"; -- -0.15101655060643931
	pesos_i(24337) := b"1111111111111111_1111111111111111_1111010010110010_1000000001111100"; -- -0.04415127720172011
	pesos_i(24338) := b"0000000000000000_0000000000000000_0000001000001100_0101111011101101"; -- 0.00800126353349315
	pesos_i(24339) := b"0000000000000000_0000000000000000_0010001001000000_1100110100100010"; -- 0.13380128944521286
	pesos_i(24340) := b"0000000000000000_0000000000000000_0000110100100101_1111000101001000"; -- 0.05136020664392841
	pesos_i(24341) := b"1111111111111111_1111111111111111_1110111011000110_1100001010111011"; -- -0.06727965288233304
	pesos_i(24342) := b"0000000000000000_0000000000000000_0001000100001001_0011110011010100"; -- 0.06654720476692037
	pesos_i(24343) := b"1111111111111111_1111111111111111_1110001111010010_1101111100111001"; -- -0.11006359909757803
	pesos_i(24344) := b"1111111111111111_1111111111111111_1111101110110110_0111001010000000"; -- -0.016747325684704006
	pesos_i(24345) := b"1111111111111111_1111111111111111_1110010111000001_0001001010111001"; -- -0.10252268775500778
	pesos_i(24346) := b"1111111111111111_1111111111111111_1111001011111010_1101111010010100"; -- -0.05085953599898444
	pesos_i(24347) := b"0000000000000000_0000000000000000_0001111100111010_1000111110110001"; -- 0.12198732455374
	pesos_i(24348) := b"0000000000000000_0000000000000000_0000011010101110_0111101000000011"; -- 0.026099801857194432
	pesos_i(24349) := b"0000000000000000_0000000000000000_0001001011001101_0011001011101100"; -- 0.07344358699725542
	pesos_i(24350) := b"0000000000000000_0000000000000000_0001010111011110_1000111110110100"; -- 0.08542726666157312
	pesos_i(24351) := b"0000000000000000_0000000000000000_0000011101001111_1011001000010000"; -- 0.028559807777003027
	pesos_i(24352) := b"1111111111111111_1111111111111111_1111110101110101_1001010010101101"; -- -0.009924609888631078
	pesos_i(24353) := b"0000000000000000_0000000000000000_0001010100101110_1000101001011010"; -- 0.08274140074486516
	pesos_i(24354) := b"0000000000000000_0000000000000000_0001100011100100_0100010010011110"; -- 0.09723309383658044
	pesos_i(24355) := b"0000000000000000_0000000000000000_0000001100011111_0000000011100000"; -- 0.012191824586749077
	pesos_i(24356) := b"1111111111111111_1111111111111111_1110100111001101_1100100000100011"; -- -0.08670376919088434
	pesos_i(24357) := b"1111111111111111_1111111111111111_1101101001011101_1001000100111010"; -- -0.1470097765266031
	pesos_i(24358) := b"0000000000000000_0000000000000000_0001100101110101_1111000001011001"; -- 0.09945585407462744
	pesos_i(24359) := b"1111111111111111_1111111111111111_1111100111011100_0011111011100100"; -- -0.023983067797210808
	pesos_i(24360) := b"1111111111111111_1111111111111111_1110001101110000_0101000100111010"; -- -0.11156742410845773
	pesos_i(24361) := b"1111111111111111_1111111111111111_1111001001110110_1011010110111000"; -- -0.052876131694448436
	pesos_i(24362) := b"1111111111111111_1111111111111111_1110100110110101_1110001010110001"; -- -0.0870683973895013
	pesos_i(24363) := b"1111111111111111_1111111111111111_1110111111111101_1001101101001010"; -- -0.06253652042336923
	pesos_i(24364) := b"0000000000000000_0000000000000000_0000000011001111_0010001010100001"; -- 0.0031606333599272845
	pesos_i(24365) := b"0000000000000000_0000000000000000_0001011101111011_1010000111010001"; -- 0.09173022605059816
	pesos_i(24366) := b"1111111111111111_1111111111111111_1110100111100101_1110001101111111"; -- -0.08633592758553332
	pesos_i(24367) := b"0000000000000000_0000000000000000_0000101000110110_0011000011110010"; -- 0.03988939187192623
	pesos_i(24368) := b"1111111111111111_1111111111111111_1110110110110101_0011111110101011"; -- -0.07145311431915687
	pesos_i(24369) := b"0000000000000000_0000000000000000_0001100100100111_1011110000000010"; -- 0.09826254901577205
	pesos_i(24370) := b"0000000000000000_0000000000000000_0010000000010110_1000101010011001"; -- 0.1253439543101487
	pesos_i(24371) := b"1111111111111111_1111111111111111_1110100101110000_0110000100111001"; -- -0.08812897081684458
	pesos_i(24372) := b"0000000000000000_0000000000000000_0000110100010011_1100100011011010"; -- 0.05108313859201881
	pesos_i(24373) := b"1111111111111111_1111111111111111_1111111011100111_1010110100111100"; -- -0.0042773941064300994
	pesos_i(24374) := b"0000000000000000_0000000000000000_0000000111110010_0010100000001101"; -- 0.0076012642515606845
	pesos_i(24375) := b"1111111111111111_1111111111111111_1111100011100101_1110001100100111"; -- -0.02774219787607793
	pesos_i(24376) := b"0000000000000000_0000000000000000_0001111110000010_1000010001101100"; -- 0.1230852855529202
	pesos_i(24377) := b"1111111111111111_1111111111111111_1110001000110100_1010000110010001"; -- -0.11638441278269661
	pesos_i(24378) := b"1111111111111111_1111111111111111_1110010010100110_1110101100011101"; -- -0.10682802714097499
	pesos_i(24379) := b"0000000000000000_0000000000000000_0001000101110000_0011011101000111"; -- 0.06811852920068281
	pesos_i(24380) := b"1111111111111111_1111111111111111_1110101111000011_1111101100101101"; -- -0.07904081494451165
	pesos_i(24381) := b"1111111111111111_1111111111111111_1110000011100110_1000010000010010"; -- -0.12148260657350926
	pesos_i(24382) := b"0000000000000000_0000000000000000_0000111101111100_0100000100100111"; -- 0.060489723326842555
	pesos_i(24383) := b"1111111111111111_1111111111111111_1110000111101111_0110010010111101"; -- -0.11744089486598407
	pesos_i(24384) := b"1111111111111111_1111111111111111_1110010001001111_1010111100111000"; -- -0.10815911181877866
	pesos_i(24385) := b"1111111111111111_1111111111111111_1111110101111110_0010001010111000"; -- -0.009794073092505224
	pesos_i(24386) := b"0000000000000000_0000000000000000_0000110110011101_0101100100101000"; -- 0.05318219399887978
	pesos_i(24387) := b"0000000000000000_0000000000000000_0001101000001001_0101011001110101"; -- 0.1017049822537959
	pesos_i(24388) := b"0000000000000000_0000000000000000_0001101111001001_1011101100101101"; -- 0.10854692311950977
	pesos_i(24389) := b"0000000000000000_0000000000000000_0001101110100010_0000101011011110"; -- 0.10794132159178647
	pesos_i(24390) := b"1111111111111111_1111111111111111_1111110101111001_1010010010001110"; -- -0.009862628395760157
	pesos_i(24391) := b"1111111111111111_1111111111111111_1111010010101100_1011111000100110"; -- -0.044239154531024144
	pesos_i(24392) := b"0000000000000000_0000000000000000_0000100111011010_1100110010001000"; -- 0.038494857083051434
	pesos_i(24393) := b"0000000000000000_0000000000000000_0001011101001011_0111100100010101"; -- 0.0909953761248858
	pesos_i(24394) := b"1111111111111111_1111111111111111_1110000111011010_1100101110110010"; -- -0.11775519273743441
	pesos_i(24395) := b"1111111111111111_1111111111111111_1110010101101011_0100010111100101"; -- -0.10383189360433319
	pesos_i(24396) := b"1111111111111111_1111111111111111_1110100100011001_0111111101100001"; -- -0.08945468797149538
	pesos_i(24397) := b"1111111111111111_1111111111111111_1111011111011000_0110001111010001"; -- -0.0318544019882233
	pesos_i(24398) := b"1111111111111111_1111111111111111_1111111010011111_0001010111011000"; -- -0.00538505062290478
	pesos_i(24399) := b"0000000000000000_0000000000000000_0000010111010101_1110101111100101"; -- 0.02279543242658861
	pesos_i(24400) := b"0000000000000000_0000000000000000_0001010101101010_0000110101010010"; -- 0.08364947548123985
	pesos_i(24401) := b"0000000000000000_0000000000000000_0010010000011101_1010010101000000"; -- 0.1410773545656239
	pesos_i(24402) := b"1111111111111111_1111111111111111_1101110001100101_0001001010101101"; -- -0.1390827491873663
	pesos_i(24403) := b"1111111111111111_1111111111111111_1110011001100111_1001110101101101"; -- -0.09998146131871605
	pesos_i(24404) := b"0000000000000000_0000000000000000_0001001011100000_1000101100001110"; -- 0.0737387570479447
	pesos_i(24405) := b"1111111111111111_1111111111111111_1111100101110111_1111000001111011"; -- -0.025513620297662555
	pesos_i(24406) := b"1111111111111111_1111111111111111_1110001100010001_1011011111101110"; -- -0.11301088763771108
	pesos_i(24407) := b"1111111111111111_1111111111111111_1101110001100101_1010111000001000"; -- -0.13907348923187499
	pesos_i(24408) := b"1111111111111111_1111111111111111_1101010010110110_1110100001101010"; -- -0.16908404747440112
	pesos_i(24409) := b"0000000000000000_0000000000000000_0000111010101000_1001111010101000"; -- 0.05726043310740936
	pesos_i(24410) := b"1111111111111111_1111111111111111_1111000110001010_0011101101010111"; -- -0.05648450015536675
	pesos_i(24411) := b"0000000000000000_0000000000000000_0010000001100010_0000011111100111"; -- 0.12649583245207693
	pesos_i(24412) := b"1111111111111111_1111111111111111_1110110111011101_1110010011001101"; -- -0.0708329200271457
	pesos_i(24413) := b"1111111111111111_1111111111111111_1110111001010001_1001010110111001"; -- -0.06906761394784114
	pesos_i(24414) := b"1111111111111111_1111111111111111_1110011010010100_1001001010111110"; -- -0.09929545260105045
	pesos_i(24415) := b"1111111111111111_1111111111111111_1110000111111100_1101000110010011"; -- -0.11723604355809697
	pesos_i(24416) := b"0000000000000000_0000000000000000_0001111001111000_0110110010000110"; -- 0.11902502311910329
	pesos_i(24417) := b"0000000000000000_0000000000000000_0000110010101100_1011001011101001"; -- 0.04951017562775822
	pesos_i(24418) := b"0000000000000000_0000000000000000_0000011011001001_0100011000000010"; -- 0.026508689340342458
	pesos_i(24419) := b"1111111111111111_1111111111111111_1110100011000110_0011101111100010"; -- -0.09072519051133796
	pesos_i(24420) := b"0000000000000000_0000000000000000_0001011010110110_0111001101011110"; -- 0.08872147609852205
	pesos_i(24421) := b"0000000000000000_0000000000000000_0000000000110100_1111110111000100"; -- 0.0008085827078681559
	pesos_i(24422) := b"1111111111111111_1111111111111111_1111001100001011_0101010000011101"; -- -0.0506083896753327
	pesos_i(24423) := b"1111111111111111_1111111111111111_1110111101101000_1101001101110101"; -- -0.06480673202731149
	pesos_i(24424) := b"1111111111111111_1111111111111111_1110111100011110_0010101100101000"; -- -0.06594591405338827
	pesos_i(24425) := b"0000000000000000_0000000000000000_0010001101000011_0110111100101001"; -- 0.1377477144573152
	pesos_i(24426) := b"0000000000000000_0000000000000000_0001011011111111_1000000101010010"; -- 0.08983619931137994
	pesos_i(24427) := b"0000000000000000_0000000000000000_0010010010011010_0100111110011100"; -- 0.1429795985896644
	pesos_i(24428) := b"1111111111111111_1111111111111111_1110100000001110_1001100001011001"; -- -0.09352729626976088
	pesos_i(24429) := b"0000000000000000_0000000000000000_0000101110010010_0101100001100010"; -- 0.04520180125372176
	pesos_i(24430) := b"0000000000000000_0000000000000000_0001011001001001_0110011000110001"; -- 0.08705748265787268
	pesos_i(24431) := b"1111111111111111_1111111111111111_1111110100110010_0010100001101110"; -- -0.010953400775081603
	pesos_i(24432) := b"1111111111111111_1111111111111111_1110011100011110_1111001100010000"; -- -0.09718399877542769
	pesos_i(24433) := b"1111111111111111_1111111111111111_1110010100001111_0101000111010100"; -- -0.10523499087292275
	pesos_i(24434) := b"1111111111111111_1111111111111111_1110100001111001_0110000111001001"; -- -0.09189785815912993
	pesos_i(24435) := b"0000000000000000_0000000000000000_0000101100011110_0110001000111100"; -- 0.04343236896653291
	pesos_i(24436) := b"1111111111111111_1111111111111111_1101111110110110_1000000000010000"; -- -0.12612151727656745
	pesos_i(24437) := b"0000000000000000_0000000000000000_0001111100111111_1110110000111010"; -- 0.12206913397968165
	pesos_i(24438) := b"1111111111111111_1111111111111111_1111110011100110_1111001001001010"; -- -0.012101037060743421
	pesos_i(24439) := b"1111111111111111_1111111111111111_1110101101010010_0001011000000000"; -- -0.08077871788722368
	pesos_i(24440) := b"0000000000000000_0000000000000000_0000101000101010_0101111101100001"; -- 0.039709054238911856
	pesos_i(24441) := b"0000000000000000_0000000000000000_0010011100111001_0001110110010101"; -- 0.15321526426518178
	pesos_i(24442) := b"0000000000000000_0000000000000000_0000001110111110_1101110100011100"; -- 0.014631099099093615
	pesos_i(24443) := b"1111111111111111_1111111111111111_1101110110011100_1010110010101100"; -- -0.13432808684132622
	pesos_i(24444) := b"0000000000000000_0000000000000000_0001100111111001_1111110001001111"; -- 0.10147072729701419
	pesos_i(24445) := b"1111111111111111_1111111111111111_1110011001001000_0111111010111000"; -- -0.10045631414177221
	pesos_i(24446) := b"1111111111111111_1111111111111111_1111000000110100_1101011001100010"; -- -0.06169376466435937
	pesos_i(24447) := b"0000000000000000_0000000000000000_0000110001010010_0110001000111001"; -- 0.048132075171582904
	pesos_i(24448) := b"0000000000000000_0000000000000000_0000001101111000_0100001001001000"; -- 0.013553755251828729
	pesos_i(24449) := b"1111111111111111_1111111111111111_1110111111011000_1011100001100000"; -- -0.06309936190857193
	pesos_i(24450) := b"0000000000000000_0000000000000000_0001101110100000_0100001001001100"; -- 0.107914107808535
	pesos_i(24451) := b"1111111111111111_1111111111111111_1111001000010111_0110100001001101"; -- -0.05433033111867421
	pesos_i(24452) := b"0000000000000000_0000000000000000_0001110001010111_1111111111001001"; -- 0.1107177605377447
	pesos_i(24453) := b"0000000000000000_0000000000000000_0000101001011110_0001011110110000"; -- 0.04049823802675907
	pesos_i(24454) := b"0000000000000000_0000000000000000_0010001111101000_1000011010101110"; -- 0.14026681666507237
	pesos_i(24455) := b"1111111111111111_1111111111111111_1101111100100010_1101010010001011"; -- -0.12837478257776783
	pesos_i(24456) := b"0000000000000000_0000000000000000_0001100100101000_1010011101011101"; -- 0.09827657712749133
	pesos_i(24457) := b"1111111111111111_1111111111111111_1111110011100110_1110101100111101"; -- -0.012101457162752655
	pesos_i(24458) := b"1111111111111111_1111111111111111_1111111100101001_1001001100100010"; -- -0.0032718699478893006
	pesos_i(24459) := b"1111111111111111_1111111111111111_1101111010010001_0111000110010001"; -- -0.13059320658391244
	pesos_i(24460) := b"1111111111111111_1111111111111111_1110111010010011_1101100100000010"; -- -0.0680565233489432
	pesos_i(24461) := b"1111111111111111_1111111111111111_1110010101100111_0111111101011000"; -- -0.10388950440641616
	pesos_i(24462) := b"1111111111111111_1111111111111111_1111110110010111_0011010101000100"; -- -0.009411497880103292
	pesos_i(24463) := b"0000000000000000_0000000000000000_0010000000110100_1011001110000010"; -- 0.12580415648218543
	pesos_i(24464) := b"0000000000000000_0000000000000000_0000001111110100_1000101101100110"; -- 0.015450203245551951
	pesos_i(24465) := b"1111111111111111_1111111111111111_1110100011001010_0001110010000111"; -- -0.0906660242120994
	pesos_i(24466) := b"0000000000000000_0000000000000000_0000100111000000_0110110000111111"; -- 0.038092389510329824
	pesos_i(24467) := b"0000000000000000_0000000000000000_0000100010111001_1011011101001001"; -- 0.034083800509033334
	pesos_i(24468) := b"0000000000000000_0000000000000000_0000111111000000_0110000111111100"; -- 0.06152927792823688
	pesos_i(24469) := b"0000000000000000_0000000000000000_0000011111100000_0101000101111101"; -- 0.030766575917832127
	pesos_i(24470) := b"1111111111111111_1111111111111111_1110101110101011_0011000110100111"; -- -0.07941903749801242
	pesos_i(24471) := b"0000000000000000_0000000000000000_0001010100001101_1000000000101101"; -- 0.08223725413990028
	pesos_i(24472) := b"1111111111111111_1111111111111111_1111010010000111_0010101001100101"; -- -0.04481253665795874
	pesos_i(24473) := b"1111111111111111_1111111111111111_1110110111110011_0010000001101111"; -- -0.07050893102680801
	pesos_i(24474) := b"0000000000000000_0000000000000000_0010010010010110_0000010000010011"; -- 0.14291406111116964
	pesos_i(24475) := b"1111111111111111_1111111111111111_1111011001110010_1111001110000100"; -- -0.03730848332697774
	pesos_i(24476) := b"0000000000000000_0000000000000000_0000011110101010_1011111100100101"; -- 0.029949137141473597
	pesos_i(24477) := b"0000000000000000_0000000000000000_0010001001100100_0011001010000011"; -- 0.13434138967032472
	pesos_i(24478) := b"0000000000000000_0000000000000000_0000010000001101_1011011001011101"; -- 0.015834233894530633
	pesos_i(24479) := b"1111111111111111_1111111111111111_1111100101011010_0101101110100111"; -- -0.025964995980164305
	pesos_i(24480) := b"1111111111111111_1111111111111111_1110000111110100_0100110100110111"; -- -0.11736600315460596
	pesos_i(24481) := b"1111111111111111_1111111111111111_1110101110100101_0101010100101011"; -- -0.07950847333613177
	pesos_i(24482) := b"0000000000000000_0000000000000000_0001001100011001_0010000101001111"; -- 0.0746022051411857
	pesos_i(24483) := b"1111111111111111_1111111111111111_1111000010010001_1110011101111110"; -- -0.060273677522273444
	pesos_i(24484) := b"1111111111111111_1111111111111111_1110110110010011_0110011111111000"; -- -0.07196951092567513
	pesos_i(24485) := b"0000000000000000_0000000000000000_0000000110100010_1000000010001010"; -- 0.006385835444218181
	pesos_i(24486) := b"0000000000000000_0000000000000000_0001001100000100_0010001001010000"; -- 0.07428183029938853
	pesos_i(24487) := b"0000000000000000_0000000000000000_0001100101001010_0010100000011101"; -- 0.09878779139911349
	pesos_i(24488) := b"1111111111111111_1111111111111111_1110010110000101_1100001001010110"; -- -0.1034277477002392
	pesos_i(24489) := b"0000000000000000_0000000000000000_0001010010010001_0000001011110100"; -- 0.08033770034011778
	pesos_i(24490) := b"0000000000000000_0000000000000000_0000010011111001_1010001101111000"; -- 0.01943418197210515
	pesos_i(24491) := b"1111111111111111_1111111111111111_1111111101110001_1111110110000011"; -- -0.0021668963536467965
	pesos_i(24492) := b"1111111111111111_1111111111111111_1110010001110100_0001010000100111"; -- -0.10760377938410669
	pesos_i(24493) := b"0000000000000000_0000000000000000_0010001000100111_0001001110001010"; -- 0.13340875738880878
	pesos_i(24494) := b"0000000000000000_0000000000000000_0001101101101010_1100010111100101"; -- 0.10709797718487452
	pesos_i(24495) := b"1111111111111111_1111111111111111_1101011011101101_0001011100100011"; -- -0.1604447878970459
	pesos_i(24496) := b"1111111111111111_1111111111111111_1101110100110101_1101011001101000"; -- -0.1358972545013412
	pesos_i(24497) := b"0000000000000000_0000000000000000_0000111100100001_1000000110110001"; -- 0.059105020276965486
	pesos_i(24498) := b"1111111111111111_1111111111111111_1110100100111001_0111111101101101"; -- -0.08896640375127533
	pesos_i(24499) := b"1111111111111111_1111111111111111_1111001110101100_1111000010110000"; -- -0.04814239210357577
	pesos_i(24500) := b"0000000000000000_0000000000000000_0001101100110100_1001110010001011"; -- 0.1062715377832624
	pesos_i(24501) := b"1111111111111111_1111111111111111_1111111000101000_1111100101100101"; -- -0.007187283383477914
	pesos_i(24502) := b"1111111111111111_1111111111111111_1111010011000110_1101010111101100"; -- -0.04384100897920543
	pesos_i(24503) := b"1111111111111111_1111111111111111_1110110010111001_1001101100101001"; -- -0.0752928757608975
	pesos_i(24504) := b"0000000000000000_0000000000000000_0000010011010101_0011101010011101"; -- 0.018878615683351523
	pesos_i(24505) := b"1111111111111111_1111111111111111_1110111010000100_1110010001111111"; -- -0.06828472049978979
	pesos_i(24506) := b"1111111111111111_1111111111111111_1111000101111001_1110001010010100"; -- -0.0567339315277004
	pesos_i(24507) := b"0000000000000000_0000000000000000_0000001000000011_1010110001101011"; -- 0.007868553348699967
	pesos_i(24508) := b"0000000000000000_0000000000000000_0001100000001100_1000001100111001"; -- 0.09394092701297557
	pesos_i(24509) := b"0000000000000000_0000000000000000_0000110011100010_1110000011111001"; -- 0.05033689577764147
	pesos_i(24510) := b"0000000000000000_0000000000000000_0000000110100010_0100000001001001"; -- 0.0063820056209444075
	pesos_i(24511) := b"1111111111111111_1111111111111111_1111111010010011_1001011111010001"; -- -0.005560409103377199
	pesos_i(24512) := b"0000000000000000_0000000000000000_0000101100100111_0101100001000110"; -- 0.04356910432023769
	pesos_i(24513) := b"1111111111111111_1111111111111111_1101110000111011_0000111100101011"; -- -0.13972382727739388
	pesos_i(24514) := b"1111111111111111_1111111111111111_1110001111101101_0000101111101111"; -- -0.1096642056888351
	pesos_i(24515) := b"0000000000000000_0000000000000000_0000000001100100_0010100010101010"; -- 0.0015283025810445558
	pesos_i(24516) := b"1111111111111111_1111111111111111_1110110010000010_0111010001010100"; -- -0.0761344237469292
	pesos_i(24517) := b"1111111111111111_1111111111111111_1111011111111001_0100110111010001"; -- -0.03135217325246126
	pesos_i(24518) := b"0000000000000000_0000000000000000_0000010101010000_1110111010000000"; -- 0.02076616894458604
	pesos_i(24519) := b"0000000000000000_0000000000000000_0000010111001011_0000000111011001"; -- 0.022628894240832125
	pesos_i(24520) := b"1111111111111111_1111111111111111_1110110100101011_0101000100010001"; -- -0.07355779021699013
	pesos_i(24521) := b"1111111111111111_1111111111111111_1110001010000100_0011110101000100"; -- -0.11516968806854198
	pesos_i(24522) := b"0000000000000000_0000000000000000_0001011101001010_0101100111111011"; -- 0.09097826363721669
	pesos_i(24523) := b"1111111111111111_1111111111111111_1110111100110111_1100000011010101"; -- -0.06555552298091406
	pesos_i(24524) := b"1111111111111111_1111111111111111_1101111011001001_0100011111101111"; -- -0.12974119592526978
	pesos_i(24525) := b"1111111111111111_1111111111111111_1110010010011101_0100000110000001"; -- -0.10697546582880282
	pesos_i(24526) := b"0000000000000000_0000000000000000_0000101111011011_1101011010001001"; -- 0.04632321204323401
	pesos_i(24527) := b"0000000000000000_0000000000000000_0010001101001111_0100000001010100"; -- 0.1379280286167651
	pesos_i(24528) := b"1111111111111111_1111111111111111_1110010101101001_1010001000101010"; -- -0.10385691135584957
	pesos_i(24529) := b"0000000000000000_0000000000000000_0001100110111110_0010000101100111"; -- 0.1005574108858329
	pesos_i(24530) := b"1111111111111111_1111111111111111_1111101100001010_0110001110010110"; -- -0.019372726270535812
	pesos_i(24531) := b"0000000000000000_0000000000000000_0001110101101110_1001100011110011"; -- 0.11496883323159676
	pesos_i(24532) := b"1111111111111111_1111111111111111_1101110001101010_0001011110010111"; -- -0.13900616222837625
	pesos_i(24533) := b"0000000000000000_0000000000000000_0001010011001110_0110001001010100"; -- 0.08127417146014272
	pesos_i(24534) := b"1111111111111111_1111111111111111_1110100100000101_1000101010110101"; -- -0.08975918836723218
	pesos_i(24535) := b"0000000000000000_0000000000000000_0001100101011011_1101101100001111"; -- 0.09905785660596562
	pesos_i(24536) := b"0000000000000000_0000000000000000_0001101100101110_0111111011100100"; -- 0.10617821759707616
	pesos_i(24537) := b"1111111111111111_1111111111111111_1111111011000010_1110111100010111"; -- -0.004838044080892591
	pesos_i(24538) := b"1111111111111111_1111111111111111_1110101111000000_1111010101011111"; -- -0.07908693713287766
	pesos_i(24539) := b"1111111111111111_1111111111111111_1111111000101011_1000011101101101"; -- -0.007148299964047154
	pesos_i(24540) := b"1111111111111111_1111111111111111_1111001101010000_0001110111111100"; -- -0.049558759708194906
	pesos_i(24541) := b"1111111111111111_1111111111111111_1111011011101001_0100101111010000"; -- -0.03550268328114637
	pesos_i(24542) := b"0000000000000000_0000000000000000_0000011001010100_1111010111000010"; -- 0.024733886511353356
	pesos_i(24543) := b"0000000000000000_0000000000000000_0001101011101010_1001011111100011"; -- 0.10514210975335368
	pesos_i(24544) := b"1111111111111111_1111111111111111_1110101001110010_0100110011100000"; -- -0.08419341586815633
	pesos_i(24545) := b"0000000000000000_0000000000000000_0000011010000101_1100101000101101"; -- 0.025478969561006808
	pesos_i(24546) := b"0000000000000000_0000000000000000_0000100000100101_1110100011110000"; -- 0.03182845939854437
	pesos_i(24547) := b"0000000000000000_0000000000000000_0000110111011001_0111000110000110"; -- 0.05409917385044165
	pesos_i(24548) := b"0000000000000000_0000000000000000_0010000001010000_0111000000010000"; -- 0.12622738267395933
	pesos_i(24549) := b"1111111111111111_1111111111111111_1111011001110011_1111000101000100"; -- -0.037293358625787636
	pesos_i(24550) := b"0000000000000000_0000000000000000_0001010000010000_1011100110011001"; -- 0.07838020318893764
	pesos_i(24551) := b"0000000000000000_0000000000000000_0011001110000000_1000011101101101"; -- 0.2011799469809753
	pesos_i(24552) := b"0000000000000000_0000000000000000_0001100101100010_1100100110010011"; -- 0.09916362619902866
	pesos_i(24553) := b"1111111111111111_1111111111111111_1101101010011101_1010110010100001"; -- -0.14603158062544228
	pesos_i(24554) := b"1111111111111111_1111111111111111_1110110111001101_1111111011010111"; -- -0.07107550869821587
	pesos_i(24555) := b"0000000000000000_0000000000000000_0001010110101110_1101000100110110"; -- 0.08469874920451856
	pesos_i(24556) := b"1111111111111111_1111111111111111_1111101100010001_0100100001011111"; -- -0.019267537008016866
	pesos_i(24557) := b"0000000000000000_0000000000000000_0001110100001110_1001110110111101"; -- 0.11350427488555596
	pesos_i(24558) := b"0000000000000000_0000000000000000_0001010101111010_0001010100001011"; -- 0.0838940764258058
	pesos_i(24559) := b"1111111111111111_1111111111111111_1110111000010101_1010010110001001"; -- -0.06998219886797899
	pesos_i(24560) := b"0000000000000000_0000000000000000_0010000101011001_0110011000110011"; -- 0.13027037384223883
	pesos_i(24561) := b"0000000000000000_0000000000000000_0010001100001111_0100110111011000"; -- 0.13695227172129862
	pesos_i(24562) := b"0000000000000000_0000000000000000_0000101111001100_1100111111111110"; -- 0.04609394032535134
	pesos_i(24563) := b"1111111111111111_1111111111111111_1111001010011110_0000111111010110"; -- -0.052275667473921
	pesos_i(24564) := b"1111111111111111_1111111111111111_1110101100000001_0011111000000101"; -- -0.08201229460032265
	pesos_i(24565) := b"1111111111111111_1111111111111111_1111110010001110_1111110000001100"; -- -0.013443228738315091
	pesos_i(24566) := b"1111111111111111_1111111111111111_1101111111011000_0010010100110100"; -- -0.12560813403643256
	pesos_i(24567) := b"1111111111111111_1111111111111111_1110100000000111_0001011101011101"; -- -0.09364179589500489
	pesos_i(24568) := b"0000000000000000_0000000000000000_0001011110100011_0100101100110010"; -- 0.09233541468611235
	pesos_i(24569) := b"1111111111111111_1111111111111111_1110000001000101_0110101010101100"; -- -0.12394078551301281
	pesos_i(24570) := b"0000000000000000_0000000000000000_0000000100101110_0010110100011100"; -- 0.004610842976404561
	pesos_i(24571) := b"1111111111111111_1111111111111111_1110101010011100_0001001100000100"; -- -0.08355599545248169
	pesos_i(24572) := b"1111111111111111_1111111111111111_1111000101101001_0100011101100010"; -- -0.05698732233062228
	pesos_i(24573) := b"1111111111111111_1111111111111111_1110000110101110_1110100110011001"; -- -0.11842479709947573
	pesos_i(24574) := b"1111111111111111_1111111111111111_1110100010111111_0001101011101110"; -- -0.09083396610730467
	pesos_i(24575) := b"1111111111111111_1111111111111111_1101101011001111_1110010011100000"; -- -0.1452652886010199
	pesos_i(24576) := b"1111111111111111_1111111111111111_1101001001011111_0011110010000111"; -- -0.1782343074206376
	pesos_i(24577) := b"0000000000000000_0000000000000000_0011001010010010_1101101110111111"; -- 0.19755338108846893
	pesos_i(24578) := b"1111111111111111_1111111111111111_1110010010010000_1000011001111011"; -- -0.10716971877682592
	pesos_i(24579) := b"0000000000000000_0000000000000000_0000101110111111_0111110000110011"; -- 0.045890581526175936
	pesos_i(24580) := b"1111111111111111_1111111111111111_1111101111010011_0011101011000100"; -- -0.016308142793445897
	pesos_i(24581) := b"0000000000000000_0000000000000000_0010000110100011_1000100010001011"; -- 0.1314015712885445
	pesos_i(24582) := b"0000000000000000_0000000000000000_0010000100111111_0100001100011100"; -- 0.12987155372877454
	pesos_i(24583) := b"0000000000000000_0000000000000000_0010110010100010_1111111011011100"; -- 0.17436211453656172
	pesos_i(24584) := b"1111111111111111_1111111111111111_1110010101010010_1010110110011100"; -- -0.10420718140390824
	pesos_i(24585) := b"1111111111111111_1111111111111111_1111011101110001_1011111101011101"; -- -0.03342060065144326
	pesos_i(24586) := b"0000000000000000_0000000000000000_0001101100100011_1110001110010111"; -- 0.10601637300326584
	pesos_i(24587) := b"0000000000000000_0000000000000000_0010110110101100_0010110011010100"; -- 0.17840843357032085
	pesos_i(24588) := b"1111111111111111_1111111111111111_1110010101100011_1111001110110100"; -- -0.10394360398496996
	pesos_i(24589) := b"0000000000000000_0000000000000000_0010111001111010_1001100001010111"; -- 0.18155815248390528
	pesos_i(24590) := b"1111111111111111_1111111111111111_1111100001001000_1010111100100101"; -- -0.030140927859181255
	pesos_i(24591) := b"1111111111111111_1111111111111111_1110001110011111_0010010100010001"; -- -0.1108528933144811
	pesos_i(24592) := b"1111111111111111_1111111111111111_1111011001011111_0010101111000011"; -- -0.03761030653702906
	pesos_i(24593) := b"1111111111111111_1111111111111111_1110100110110011_0011101101000100"; -- -0.08710889435581824
	pesos_i(24594) := b"0000000000000000_0000000000000000_0010000110010101_0010100001100110"; -- 0.13118221755294576
	pesos_i(24595) := b"1111111111111111_1111111111111111_1110010100110010_1110011000101110"; -- -0.10469209073797997
	pesos_i(24596) := b"1111111111111111_1111111111111111_1101010100000001_0100101001111100"; -- -0.16794905164340118
	pesos_i(24597) := b"0000000000000000_0000000000000000_0001001011011000_1100101010011010"; -- 0.07362047438165291
	pesos_i(24598) := b"0000000000000000_0000000000000000_0001110011010001_0100011001110010"; -- 0.11256828586779263
	pesos_i(24599) := b"0000000000000000_0000000000000000_0001110111010001_0111101001111100"; -- 0.11647763746657953
	pesos_i(24600) := b"0000000000000000_0000000000000000_0011000101101110_0000011010110111"; -- 0.1930851169264048
	pesos_i(24601) := b"0000000000000000_0000000000000000_0010010010111110_0110111100110010"; -- 0.14353079766002466
	pesos_i(24602) := b"0000000000000000_0000000000000000_0011000000001101_1110110110110010"; -- 0.18771253201602908
	pesos_i(24603) := b"0000000000000000_0000000000000000_0010110111000100_0101011111000000"; -- 0.17877720287486024
	pesos_i(24604) := b"1111111111111111_1111111111111111_1101110011110001_1001001011000011"; -- -0.13693888412833863
	pesos_i(24605) := b"0000000000000000_0000000000000000_0001101011111001_1101110010110011"; -- 0.1053750932207588
	pesos_i(24606) := b"0000000000000000_0000000000000000_0001100001101001_0111000110110111"; -- 0.09535895088139688
	pesos_i(24607) := b"1111111111111111_1111111111111111_1110110101100000_1001101101011011"; -- -0.07274464622873276
	pesos_i(24608) := b"0000000000000000_0000000000000000_0001101001101010_1101110001100111"; -- 0.10319306856200011
	pesos_i(24609) := b"1111111111111111_1111111111111111_1111011000110110_0110111000001000"; -- -0.03823196696423825
	pesos_i(24610) := b"0000000000000000_0000000000000000_0001011110001011_0000011110000000"; -- 0.09196516861743353
	pesos_i(24611) := b"0000000000000000_0000000000000000_0001101010111101_1100001110110011"; -- 0.10445807570348652
	pesos_i(24612) := b"0000000000000000_0000000000000000_0001111011111010_0110001110100111"; -- 0.12100813699389595
	pesos_i(24613) := b"0000000000000000_0000000000000000_0011000001010010_0101001011111011"; -- 0.18875616678968735
	pesos_i(24614) := b"1111111111111111_1111111111111111_1100111011011100_0101000111110100"; -- -0.19195068161868578
	pesos_i(24615) := b"0000000000000000_0000000000000000_0001100101100110_1010000101000101"; -- 0.0992222588581211
	pesos_i(24616) := b"1111111111111111_1111111111111111_1110000011110011_0111000110001000"; -- -0.12128534715157036
	pesos_i(24617) := b"1111111111111111_1111111111111111_1101000011110001_0001001010010001"; -- -0.18382152508545763
	pesos_i(24618) := b"1111111111111111_1111111111111111_1101011000111011_1101010010000000"; -- -0.1631495654761716
	pesos_i(24619) := b"1111111111111111_1111111111111111_1111011101010110_1110101000110111"; -- -0.03383003385028968
	pesos_i(24620) := b"0000000000000000_0000000000000000_0000000000000101_1001000110001001"; -- 8.49685002907991e-05
	pesos_i(24621) := b"0000000000000000_0000000000000000_0000001110111010_1100011010111110"; -- 0.014568730801480655
	pesos_i(24622) := b"1111111111111111_1111111111111111_1101110101011001_0001011101011100"; -- -0.1353593255491378
	pesos_i(24623) := b"0000000000000000_0000000000000000_0000100000100110_1111001110110010"; -- 0.031844359264434324
	pesos_i(24624) := b"0000000000000000_0000000000000000_0010001001011011_1010100000101101"; -- 0.1342110738008562
	pesos_i(24625) := b"0000000000000000_0000000000000000_0000011110101100_0110001011111101"; -- 0.029974161981285836
	pesos_i(24626) := b"0000000000000000_0000000000000000_0000101011000101_1100100111101101"; -- 0.042080517223528874
	pesos_i(24627) := b"1111111111111111_1111111111111111_1110100111001000_0101110011100011"; -- -0.08678645567346394
	pesos_i(24628) := b"0000000000000000_0000000000000000_0000001110110110_1001000111100001"; -- 0.014504544730285552
	pesos_i(24629) := b"0000000000000000_0000000000000000_0001110000110011_0111111101000001"; -- 0.11016078315123057
	pesos_i(24630) := b"1111111111111111_1111111111111111_1101111110101111_0110110010000001"; -- -0.12622949449898338
	pesos_i(24631) := b"0000000000000000_0000000000000000_0000011110101111_0101011000001111"; -- 0.030019167611399604
	pesos_i(24632) := b"0000000000000000_0000000000000000_0010011000110010_0011100000101010"; -- 0.14920378710878202
	pesos_i(24633) := b"0000000000000000_0000000000000000_0000101010111000_1101010000100000"; -- 0.04188276081533072
	pesos_i(24634) := b"1111111111111111_1111111111111111_1111011001010100_0101100111010111"; -- -0.0377754068033376
	pesos_i(24635) := b"0000000000000000_0000000000000000_0001101101110010_1111100111011000"; -- 0.10722314380991627
	pesos_i(24636) := b"0000000000000000_0000000000000000_0000011110100110_0101100110100011"; -- 0.029882051732079088
	pesos_i(24637) := b"1111111111111111_1111111111111111_1101001101110101_1110111011011010"; -- -0.17398173493611446
	pesos_i(24638) := b"0000000000000000_0000000000000000_0010110100011111_0110110001011100"; -- 0.1762607310734346
	pesos_i(24639) := b"0000000000000000_0000000000000000_0010110011110000_0010000010111111"; -- 0.17553906122382204
	pesos_i(24640) := b"1111111111111111_1111111111111111_1111110000101011_0101101110001001"; -- -0.014963416137724787
	pesos_i(24641) := b"1111111111111111_1111111111111111_1100110111001101_0011110110000000"; -- -0.19608703245954848
	pesos_i(24642) := b"0000000000000000_0000000000000000_0010011001001001_1111110100101011"; -- 0.14956648158076602
	pesos_i(24643) := b"0000000000000000_0000000000000000_0001111000101000_1000000101001001"; -- 0.11780555756261675
	pesos_i(24644) := b"0000000000000000_0000000000000000_0001101100010011_1110000001000000"; -- 0.10577203336021511
	pesos_i(24645) := b"0000000000000000_0000000000000000_0011010001001100_0010000011100111"; -- 0.20428662909338854
	pesos_i(24646) := b"0000000000000000_0000000000000000_0010111000011101_0110001001011011"; -- 0.18013586721844044
	pesos_i(24647) := b"1111111111111111_1111111111111111_1110001001000011_1010010001010111"; -- -0.11615536573233463
	pesos_i(24648) := b"0000000000000000_0000000000000000_0000000101001110_0000011101011011"; -- 0.005096873946882984
	pesos_i(24649) := b"1111111111111111_1111111111111111_1101101010011001_0011100001011100"; -- -0.14609954604120584
	pesos_i(24650) := b"1111111111111111_1111111111111111_1101100110010110_0111000101101111"; -- -0.15004817051699326
	pesos_i(24651) := b"1111111111111111_1111111111111111_1110101000010001_1000001111101000"; -- -0.0856702383455553
	pesos_i(24652) := b"0000000000000000_0000000000000000_0000010100101001_0000001000101000"; -- 0.020156988947829274
	pesos_i(24653) := b"0000000000000000_0000000000000000_0001101010111010_1101100110110110"; -- 0.10441361143771202
	pesos_i(24654) := b"0000000000000000_0000000000000000_0001111101101001_0110011000011100"; -- 0.12270200895924849
	pesos_i(24655) := b"1111111111111111_1111111111111111_1110100001101000_0111010100000100"; -- -0.09215611118274843
	pesos_i(24656) := b"0000000000000000_0000000000000000_0000101111000011_0100000110001110"; -- 0.045948121238536956
	pesos_i(24657) := b"0000000000000000_0000000000000000_0001101000111001_0001101101100101"; -- 0.10243388377647508
	pesos_i(24658) := b"0000000000000000_0000000000000000_0010110001011101_0100110001110111"; -- 0.17329862506890245
	pesos_i(24659) := b"0000000000000000_0000000000000000_0000101110000111_0001011101011100"; -- 0.04503007874326521
	pesos_i(24660) := b"0000000000000000_0000000000000000_0001101000010011_0101000000110100"; -- 0.1018571975667943
	pesos_i(24661) := b"0000000000000000_0000000000000000_0000001000110101_0011001011101010"; -- 0.008624250436111564
	pesos_i(24662) := b"1111111111111111_1111111111111111_1110110001011011_0001110110101111"; -- -0.0767346809564535
	pesos_i(24663) := b"0000000000000000_0000000000000000_0000101011100101_1000000001110001"; -- 0.04256441840006209
	pesos_i(24664) := b"1111111111111111_1111111111111111_1111011000101100_0100101110010001"; -- -0.03838660928166795
	pesos_i(24665) := b"0000000000000000_0000000000000000_0010101110010011_1001001101100010"; -- 0.1702205766831502
	pesos_i(24666) := b"1111111111111111_1111111111111111_1111000100110100_1100000100011111"; -- -0.057788782078959405
	pesos_i(24667) := b"1111111111111111_1111111111111111_1101101010111001_0111011011101001"; -- -0.1456075364606538
	pesos_i(24668) := b"0000000000000000_0000000000000000_0010111100011100_0111100100111101"; -- 0.18402822248837286
	pesos_i(24669) := b"1111111111111111_1111111111111111_1111110001000000_1100001110000010"; -- -0.014636784300035148
	pesos_i(24670) := b"1111111111111111_1111111111111111_1111100011111101_0011111000011110"; -- -0.027385823929853254
	pesos_i(24671) := b"1111111111111111_1111111111111111_1101010111011010_0011101010011011"; -- -0.16463884093784537
	pesos_i(24672) := b"1111111111111111_1111111111111111_1110001001110110_0100101011001011"; -- -0.11538250492380356
	pesos_i(24673) := b"0000000000000000_0000000000000000_0010100110101010_0101010010010110"; -- 0.16275528581558707
	pesos_i(24674) := b"0000000000000000_0000000000000000_0010000011001000_0010000010000110"; -- 0.12805369625240215
	pesos_i(24675) := b"1111111111111111_1111111111111111_1110110101110000_1100000000010111"; -- -0.0724983161414091
	pesos_i(24676) := b"1111111111111111_1111111111111111_1110001101101010_0000010100001100"; -- -0.11166351754080449
	pesos_i(24677) := b"1111111111111111_1111111111111111_1110111110000100_1110000011010101"; -- -0.0643786888989466
	pesos_i(24678) := b"1111111111111111_1111111111111111_1111111110011110_0000011010101010"; -- -0.001494964201540822
	pesos_i(24679) := b"0000000000000000_0000000000000000_0001111111111100_0101000110110011"; -- 0.1249438345991597
	pesos_i(24680) := b"0000000000000000_0000000000000000_0001000000011010_1010110011010000"; -- 0.06290702898703766
	pesos_i(24681) := b"0000000000000000_0000000000000000_0000010010010001_1100001111101110"; -- 0.01784920281386909
	pesos_i(24682) := b"1111111111111111_1111111111111111_1101101011001101_1011000110111011"; -- -0.145298854570955
	pesos_i(24683) := b"0000000000000000_0000000000000000_0000001001111111_0100100100101011"; -- 0.00975472742305259
	pesos_i(24684) := b"0000000000000000_0000000000000000_0000110000110010_0111010000101011"; -- 0.04764486371030421
	pesos_i(24685) := b"1111111111111111_1111111111111111_1110101111001101_1011001010110110"; -- -0.07889254625246939
	pesos_i(24686) := b"0000000000000000_0000000000000000_0010111010000100_1111000010000000"; -- 0.18171599516203285
	pesos_i(24687) := b"1111111111111111_1111111111111111_1101101101001100_1001100110001101"; -- -0.1433624297260185
	pesos_i(24688) := b"0000000000000000_0000000000000000_0001000111011101_0110101001001000"; -- 0.06978477726269657
	pesos_i(24689) := b"1111111111111111_1111111111111111_1111100001000111_0010100100100100"; -- -0.030164173848953316
	pesos_i(24690) := b"0000000000000000_0000000000000000_0000101110101011_1001101101101010"; -- 0.045587266313183286
	pesos_i(24691) := b"1111111111111111_1111111111111111_1101111001110011_0011001000111111"; -- -0.1310547443631768
	pesos_i(24692) := b"0000000000000000_0000000000000000_0010001010010110_0001110011000111"; -- 0.13510303360327422
	pesos_i(24693) := b"0000000000000000_0000000000000000_0010000101011111_0011000111110011"; -- 0.13035881206715771
	pesos_i(24694) := b"1111111111111111_1111111111111111_1111100101001110_0110001001101111"; -- -0.026147697365816316
	pesos_i(24695) := b"1111111111111111_1111111111111111_1111011000100110_1110110101100010"; -- -0.038468516923557405
	pesos_i(24696) := b"1111111111111111_1111111111111111_1101100111010000_1000100110101101"; -- -0.1491617157179435
	pesos_i(24697) := b"0000000000000000_0000000000000000_0001000111010100_1101111111001001"; -- 0.06965445200435301
	pesos_i(24698) := b"0000000000000000_0000000000000000_0001001011100111_1011001101000111"; -- 0.07384796597207816
	pesos_i(24699) := b"1111111111111111_1111111111111111_1101101111010001_1110111001111100"; -- -0.14132794837271934
	pesos_i(24700) := b"1111111111111111_1111111111111111_1111111101001100_0110101100111000"; -- -0.002740191259077865
	pesos_i(24701) := b"1111111111111111_1111111111111111_1111101010111101_1011000011000100"; -- -0.02054305289528728
	pesos_i(24702) := b"0000000000000000_0000000000000000_0001100010111100_0100110110111000"; -- 0.09662328467729994
	pesos_i(24703) := b"1111111111111111_1111111111111111_1110011110100110_1110001001100111"; -- -0.0951097963801716
	pesos_i(24704) := b"1111111111111111_1111111111111111_1111001011110000_1111101110110101"; -- -0.05101038763821493
	pesos_i(24705) := b"1111111111111111_1111111111111111_1111111111100001_1000110001111001"; -- -0.0004646497536465038
	pesos_i(24706) := b"0000000000000000_0000000000000000_0000100011000010_0100101100100100"; -- 0.034214683811761605
	pesos_i(24707) := b"0000000000000000_0000000000000000_0010100010111111_1100101001010101"; -- 0.1591764886774045
	pesos_i(24708) := b"1111111111111111_1111111111111111_1100111011101000_0100001001101010"; -- -0.19176850228263068
	pesos_i(24709) := b"1111111111111111_1111111111111111_1101100100010010_1000000100101101"; -- -0.15206139239871846
	pesos_i(24710) := b"0000000000000000_0000000000000000_0001110001010100_1011110110011011"; -- 0.11066803954032771
	pesos_i(24711) := b"0000000000000000_0000000000000000_0001011111100011_1011110101110111"; -- 0.09331878805823043
	pesos_i(24712) := b"1111111111111111_1111111111111111_1101100011001000_1101101100101100"; -- -0.15318517853320676
	pesos_i(24713) := b"0000000000000000_0000000000000000_0010111010110101_1001110111000000"; -- 0.18245874335506032
	pesos_i(24714) := b"0000000000000000_0000000000000000_0010101101111111_1010001011110001"; -- 0.16991632837335557
	pesos_i(24715) := b"0000000000000000_0000000000000000_0000101111010010_0001001101000100"; -- 0.046174243965042494
	pesos_i(24716) := b"0000000000000000_0000000000000000_0001111000110000_0011100110010001"; -- 0.11792335300811174
	pesos_i(24717) := b"0000000000000000_0000000000000000_0001011011001100_0010011010000111"; -- 0.08905258932802285
	pesos_i(24718) := b"1111111111111111_1111111111111111_1101000000001001_1001001100011000"; -- -0.18735390348177394
	pesos_i(24719) := b"0000000000000000_0000000000000000_0010001011000001_1001100001010110"; -- 0.1357665262562839
	pesos_i(24720) := b"0000000000000000_0000000000000000_0000001111001100_1011110010001101"; -- 0.014842781555094236
	pesos_i(24721) := b"1111111111111111_1111111111111111_1111101000010010_1000111101011110"; -- -0.023154296331555132
	pesos_i(24722) := b"1111111111111111_1111111111111111_1110110011001111_1011001010000100"; -- -0.07495579023122115
	pesos_i(24723) := b"1111111111111111_1111111111111111_1111111110011001_1011010011111110"; -- -0.0015608672583136644
	pesos_i(24724) := b"0000000000000000_0000000000000000_0000100111000010_1111110101011000"; -- 0.03813155557865102
	pesos_i(24725) := b"0000000000000000_0000000000000000_0000101110000000_0101111000110100"; -- 0.04492748999697143
	pesos_i(24726) := b"1111111111111111_1111111111111111_1110001100000111_0010111110100001"; -- -0.11317159967857444
	pesos_i(24727) := b"1111111111111111_1111111111111111_1111011101111111_0100000010010011"; -- -0.03321453476080884
	pesos_i(24728) := b"1111111111111111_1111111111111111_1101100011110101_0101010010110010"; -- -0.15250654855000803
	pesos_i(24729) := b"0000000000000000_0000000000000000_0000010110010101_1000110010111011"; -- 0.02181319772630854
	pesos_i(24730) := b"1111111111111111_1111111111111111_1110001100010111_0111110000101100"; -- -0.11292289652334085
	pesos_i(24731) := b"1111111111111111_1111111111111111_1110011011000000_0100010110011001"; -- -0.09862866419267609
	pesos_i(24732) := b"1111111111111111_1111111111111111_1100110001001011_0101010000010011"; -- -0.2019755796745154
	pesos_i(24733) := b"1111111111111111_1111111111111111_1111010000100000_1001000010011010"; -- -0.04637809990654517
	pesos_i(24734) := b"1111111111111111_1111111111111111_1111010001001101_1000001110000001"; -- -0.045692234959367105
	pesos_i(24735) := b"0000000000000000_0000000000000000_0001010011111110_1110101101101001"; -- 0.08201476386750242
	pesos_i(24736) := b"1111111111111111_1111111111111111_1111101111001110_0100001001110011"; -- -0.01638397886595918
	pesos_i(24737) := b"0000000000000000_0000000000000000_0000001010100010_0111011000001001"; -- 0.010291459381026725
	pesos_i(24738) := b"1111111111111111_1111111111111111_1110011010101001_0101111010000001"; -- -0.09897813175898605
	pesos_i(24739) := b"1111111111111111_1111111111111111_1111010100100110_0011001000000111"; -- -0.04238593416629706
	pesos_i(24740) := b"0000000000000000_0000000000000000_0000010010110001_1100100110010100"; -- 0.018337820712020385
	pesos_i(24741) := b"1111111111111111_1111111111111111_1100101110000001_1001001010010001"; -- -0.20505413024162525
	pesos_i(24742) := b"1111111111111111_1111111111111111_1100110011011011_0001000001100001"; -- -0.1997823489053117
	pesos_i(24743) := b"0000000000000000_0000000000000000_0000110110001000_0101100010101101"; -- 0.05286173078904515
	pesos_i(24744) := b"0000000000000000_0000000000000000_0000001100100110_0101010001100001"; -- 0.012303613425963101
	pesos_i(24745) := b"1111111111111111_1111111111111111_1111001101111100_0011101011010000"; -- -0.04888565457028399
	pesos_i(24746) := b"1111111111111111_1111111111111111_1101011011010110_1100111000101010"; -- -0.16078483077624622
	pesos_i(24747) := b"1111111111111111_1111111111111111_1110001010101000_1100001000111110"; -- -0.11461244565586677
	pesos_i(24748) := b"0000000000000000_0000000000000000_0000110011101110_0010001100110010"; -- 0.050508689674954525
	pesos_i(24749) := b"0000000000000000_0000000000000000_0010111011011011_0000111110110110"; -- 0.18303011133595973
	pesos_i(24750) := b"1111111111111111_1111111111111111_1110100110111010_0011101011000110"; -- -0.08700211195874867
	pesos_i(24751) := b"0000000000000000_0000000000000000_0000111110011001_1110010100101101"; -- 0.06094200463736432
	pesos_i(24752) := b"0000000000000000_0000000000000000_0001100101110011_0010010101010111"; -- 0.09941323632610106
	pesos_i(24753) := b"1111111111111111_1111111111111111_1101010001111111_1100111101000111"; -- -0.1699247790238764
	pesos_i(24754) := b"0000000000000000_0000000000000000_0001110000101010_0100110010011111"; -- 0.11002043605149096
	pesos_i(24755) := b"1111111111111111_1111111111111111_1110111100100100_0100111010101111"; -- -0.06585224379108673
	pesos_i(24756) := b"1111111111111111_1111111111111111_1110110000110000_0110011100010011"; -- -0.0773864345372392
	pesos_i(24757) := b"0000000000000000_0000000000000000_0001000001010111_1101100000001110"; -- 0.06384039242040772
	pesos_i(24758) := b"0000000000000000_0000000000000000_0010101101011000_1010101000011010"; -- 0.16932166219856304
	pesos_i(24759) := b"0000000000000000_0000000000000000_0010010000100010_1011101110001100"; -- 0.14115497748311967
	pesos_i(24760) := b"0000000000000000_0000000000000000_0010101000100111_1111111110001111"; -- 0.1646728251672855
	pesos_i(24761) := b"1111111111111111_1111111111111111_1101001000111100_1100010110100101"; -- -0.17876019220096376
	pesos_i(24762) := b"1111111111111111_1111111111111111_1111011000000000_0001001001000100"; -- -0.03906141129667683
	pesos_i(24763) := b"1111111111111111_1111111111111111_1111010000000001_1100000111001011"; -- -0.046848190176456916
	pesos_i(24764) := b"1111111111111111_1111111111111111_1110011110101101_0000110110111101"; -- -0.09501566073130861
	pesos_i(24765) := b"1111111111111111_1111111111111111_1110101101010110_0000100011101101"; -- -0.08071846202884274
	pesos_i(24766) := b"0000000000000000_0000000000000000_0010101001110100_1011110001011100"; -- 0.16584374667750543
	pesos_i(24767) := b"1111111111111111_1111111111111111_1110110000111111_1100001110111100"; -- -0.07715202962415665
	pesos_i(24768) := b"0000000000000000_0000000000000000_0000110110101010_0110111010001000"; -- 0.05338183227073204
	pesos_i(24769) := b"1111111111111111_1111111111111111_1101011100001100_0100010010100001"; -- -0.15996905385834756
	pesos_i(24770) := b"1111111111111111_1111111111111111_1111000001100101_0111101010010100"; -- -0.0609515561466954
	pesos_i(24771) := b"1111111111111111_1111111111111111_1101001000011101_1010111111111110"; -- -0.17923450511140226
	pesos_i(24772) := b"0000000000000000_0000000000000000_0011010010001000_0011001101010011"; -- 0.20520325444597592
	pesos_i(24773) := b"1111111111111111_1111111111111111_1110111100111111_0100100110000110"; -- -0.06544056397724725
	pesos_i(24774) := b"1111111111111111_1111111111111111_1111000011000110_0001000111110010"; -- -0.05947769008135035
	pesos_i(24775) := b"1111111111111111_1111111111111111_1101000100111010_0001110000100001"; -- -0.1827070635173484
	pesos_i(24776) := b"0000000000000000_0000000000000000_0001000000010111_1110100101100101"; -- 0.06286486343537068
	pesos_i(24777) := b"0000000000000000_0000000000000000_0010000101101001_0011110111011001"; -- 0.13051210937209487
	pesos_i(24778) := b"0000000000000000_0000000000000000_0010011100100101_0010100101111110"; -- 0.1529107983790919
	pesos_i(24779) := b"0000000000000000_0000000000000000_0000100111111110_1010111001111100"; -- 0.039042382393745856
	pesos_i(24780) := b"0000000000000000_0000000000000000_0010000001001000_1110111100100110"; -- 0.12611288721426306
	pesos_i(24781) := b"0000000000000000_0000000000000000_0000101011010110_0010011101101110"; -- 0.04233023095384254
	pesos_i(24782) := b"0000000000000000_0000000000000000_0001111110110110_0011101001010100"; -- 0.12387432633204817
	pesos_i(24783) := b"1111111111111111_1111111111111111_1101000110010001_0110000010010000"; -- -0.18137547007415628
	pesos_i(24784) := b"1111111111111111_1111111111111111_1111111101001111_1100101110001010"; -- -0.0026886737320508574
	pesos_i(24785) := b"0000000000000000_0000000000000000_0010010000101011_0100111111110001"; -- 0.14128589278595288
	pesos_i(24786) := b"1111111111111111_1111111111111111_1111001110011111_1111001100010110"; -- -0.04834061349118296
	pesos_i(24787) := b"1111111111111111_1111111111111111_1101111100111000_0001001010011010"; -- -0.12805064908496336
	pesos_i(24788) := b"1111111111111111_1111111111111111_1101110001010111_1101001100101110"; -- -0.1392848980253439
	pesos_i(24789) := b"1111111111111111_1111111111111111_1110000010010000_1110111100101011"; -- -0.12278847893308928
	pesos_i(24790) := b"0000000000000000_0000000000000000_0011000000110010_1100110100011110"; -- 0.1882751653558355
	pesos_i(24791) := b"0000000000000000_0000000000000000_0010001101101000_0111100100100110"; -- 0.13831288499632133
	pesos_i(24792) := b"0000000000000000_0000000000000000_0010101011101111_1010101010101000"; -- 0.16771952254864897
	pesos_i(24793) := b"0000000000000000_0000000000000000_0001010000011000_0111001011010111"; -- 0.07849805581520344
	pesos_i(24794) := b"1111111111111111_1111111111111111_1101101011001101_0100110101110010"; -- -0.14530483213859466
	pesos_i(24795) := b"1111111111111111_1111111111111111_1111000001001011_1000100100010001"; -- -0.06134742095840421
	pesos_i(24796) := b"1111111111111111_1111111111111111_1101000011011101_0010101001010010"; -- -0.18412528513340742
	pesos_i(24797) := b"1111111111111111_1111111111111111_1110101010101110_0011010110001101"; -- -0.08327927886560167
	pesos_i(24798) := b"1111111111111111_1111111111111111_1111001011010110_0011100001011011"; -- -0.05141875997843197
	pesos_i(24799) := b"0000000000000000_0000000000000000_0000001101110001_0010100010101010"; -- 0.013445416990435333
	pesos_i(24800) := b"0000000000000000_0000000000000000_0010110110010100_0100000011100001"; -- 0.17804341782454258
	pesos_i(24801) := b"1111111111111111_1111111111111111_1101101010100011_1100001111010110"; -- -0.14593864462233996
	pesos_i(24802) := b"1111111111111111_1111111111111111_1101101000001111_1100000100100101"; -- -0.14819710577997683
	pesos_i(24803) := b"0000000000000000_0000000000000000_0001110011001101_0000100110111000"; -- 0.11250363106852977
	pesos_i(24804) := b"0000000000000000_0000000000000000_0010110101100101_0011011001010100"; -- 0.17732562594002987
	pesos_i(24805) := b"0000000000000000_0000000000000000_0000101110000101_1111110101001110"; -- 0.04501326713939818
	pesos_i(24806) := b"0000000000000000_0000000000000000_0000001001111110_1101100110100010"; -- 0.009748079340773935
	pesos_i(24807) := b"1111111111111111_1111111111111111_1111101100111110_1110100001010101"; -- -0.01857135711494412
	pesos_i(24808) := b"1111111111111111_1111111111111111_1111101000010101_1111000000001100"; -- -0.023102757492144372
	pesos_i(24809) := b"0000000000000000_0000000000000000_0000110011111011_0011101101010110"; -- 0.050708492636359674
	pesos_i(24810) := b"1111111111111111_1111111111111111_1111011101111011_0011011000011110"; -- -0.03327619326707418
	pesos_i(24811) := b"0000000000000000_0000000000000000_0011000111001010_0001011001001000"; -- 0.19448985340197958
	pesos_i(24812) := b"1111111111111111_1111111111111111_1101110010010000_1100100010011100"; -- -0.13841577716656187
	pesos_i(24813) := b"1111111111111111_1111111111111111_1111111100000100_0110010000001101"; -- -0.0038392513060402232
	pesos_i(24814) := b"0000000000000000_0000000000000000_0010010111000000_1110101110111011"; -- 0.14747498819327867
	pesos_i(24815) := b"0000000000000000_0000000000000000_0000111000110010_0000011011100111"; -- 0.05545085088916098
	pesos_i(24816) := b"1111111111111111_1111111111111111_1110101100111101_0001101010110011"; -- -0.08109887242152511
	pesos_i(24817) := b"1111111111111111_1111111111111111_1101001100000101_0011010111000010"; -- -0.17570175192821025
	pesos_i(24818) := b"0000000000000000_0000000000000000_0001010100001011_0011010110100111"; -- 0.08220229455449476
	pesos_i(24819) := b"0000000000000000_0000000000000000_0000001001111001_0110111001100011"; -- 0.009665393118604516
	pesos_i(24820) := b"0000000000000000_0000000000000000_0001011010100110_0011101000010101"; -- 0.0884739208910951
	pesos_i(24821) := b"1111111111111111_1111111111111111_1110101111010001_1000010000001111"; -- -0.07883429187192278
	pesos_i(24822) := b"1111111111111111_1111111111111111_1111111010011100_0000011111110110"; -- -0.005431654463720993
	pesos_i(24823) := b"1111111111111111_1111111111111111_1101010000101101_0010110101001011"; -- -0.17118565482541312
	pesos_i(24824) := b"0000000000000000_0000000000000000_0001111010111110_1001101110001100"; -- 0.12009594131028507
	pesos_i(24825) := b"1111111111111111_1111111111111111_1101010010011001_1110011001011011"; -- -0.16952667495375556
	pesos_i(24826) := b"0000000000000000_0000000000000000_0000000001101110_1010111101000110"; -- 0.0016889138212785326
	pesos_i(24827) := b"0000000000000000_0000000000000000_0001001001110010_1001111001010110"; -- 0.07206143949887862
	pesos_i(24828) := b"1111111111111111_1111111111111111_1110000010100101_1110101101011001"; -- -0.12246827190021074
	pesos_i(24829) := b"0000000000000000_0000000000000000_0010001001111000_1101001011001111"; -- 0.13465611995420615
	pesos_i(24830) := b"1111111111111111_1111111111111111_1101101111111011_1001000111000110"; -- -0.1406926051786012
	pesos_i(24831) := b"1111111111111111_1111111111111111_1101000011011010_1010001110101010"; -- -0.18416382873743095
	pesos_i(24832) := b"1111111111111111_1111111111111111_1110010100001101_0101011011100100"; -- -0.10526520677015139
	pesos_i(24833) := b"1111111111111111_1111111111111111_1110001011010101_1000111011000110"; -- -0.11392886791937605
	pesos_i(24834) := b"1111111111111111_1111111111111111_1101111011100001_1110011000010001"; -- -0.1293655594569032
	pesos_i(24835) := b"0000000000000000_0000000000000000_0001011110100010_1100111001010110"; -- 0.09232797235442398
	pesos_i(24836) := b"0000000000000000_0000000000000000_0000010000111111_0001001111010001"; -- 0.016587484972621244
	pesos_i(24837) := b"1111111111111111_1111111111111111_1101000111110101_1010100101101011"; -- -0.1798452486972005
	pesos_i(24838) := b"0000000000000000_0000000000000000_0000010010101001_0000011100001110"; -- 0.01820415591277564
	pesos_i(24839) := b"0000000000000000_0000000000000000_0010110011010011_0100000000110000"; -- 0.17509843045103857
	pesos_i(24840) := b"0000000000000000_0000000000000000_0001110110101010_0011011100000011"; -- 0.11587852311640369
	pesos_i(24841) := b"1111111111111111_1111111111111111_1111001000001110_1101110010011100"; -- -0.054460727664585214
	pesos_i(24842) := b"1111111111111111_1111111111111111_1111110001101100_1101001101110111"; -- -0.013964446453826034
	pesos_i(24843) := b"1111111111111111_1111111111111111_1111011000010001_1000111010110010"; -- -0.03879459520620363
	pesos_i(24844) := b"0000000000000000_0000000000000000_0011010010101111_0100001001110001"; -- 0.20579924838625688
	pesos_i(24845) := b"0000000000000000_0000000000000000_0000010011111110_1100100101111001"; -- 0.019512741086069776
	pesos_i(24846) := b"1111111111111111_1111111111111111_1111111101101100_0110011001110000"; -- -0.0022521951190540798
	pesos_i(24847) := b"1111111111111111_1111111111111111_1101101100101111_1100011000100010"; -- -0.14380227729851583
	pesos_i(24848) := b"0000000000000000_0000000000000000_0001001100001000_0110011100101010"; -- 0.07434696933508676
	pesos_i(24849) := b"0000000000000000_0000000000000000_0001000011011011_0010111010001010"; -- 0.06584444868813324
	pesos_i(24850) := b"1111111111111111_1111111111111111_1101100010011000_1100011101001110"; -- -0.15391878453267807
	pesos_i(24851) := b"0000000000000000_0000000000000000_0000011000000100_0011101010010111"; -- 0.023502027383538224
	pesos_i(24852) := b"0000000000000000_0000000000000000_0001100110100101_1111000110001101"; -- 0.1001883477669217
	pesos_i(24853) := b"0000000000000000_0000000000000000_0000110110000100_0000100000101000"; -- 0.052795896355506584
	pesos_i(24854) := b"0000000000000000_0000000000000000_0001000011010001_0110000011010010"; -- 0.06569485780837263
	pesos_i(24855) := b"1111111111111111_1111111111111111_1101000101110111_1000110001110110"; -- -0.1817695819018521
	pesos_i(24856) := b"0000000000000000_0000000000000000_0000011010010011_0000100011001001"; -- 0.02568106569787201
	pesos_i(24857) := b"0000000000000000_0000000000000000_0010101110010100_0011100111100100"; -- 0.17023050128370623
	pesos_i(24858) := b"0000000000000000_0000000000000000_0001110000000110_1100110111111010"; -- 0.10947882992383073
	pesos_i(24859) := b"0000000000000000_0000000000000000_0001111111010111_1001100010111111"; -- 0.12438349407382708
	pesos_i(24860) := b"1111111111111111_1111111111111111_1100111011000001_1001100001111001"; -- -0.19235846565531683
	pesos_i(24861) := b"1111111111111111_1111111111111111_1100110010000010_0011100000000011"; -- -0.20113801886575544
	pesos_i(24862) := b"0000000000000000_0000000000000000_0010101011001011_0101100100101001"; -- 0.16716534860670829
	pesos_i(24863) := b"1111111111111111_1111111111111111_1110100100100101_1101100110100111"; -- -0.08926620178315568
	pesos_i(24864) := b"0000000000000000_0000000000000000_0000010101001111_0110100111111111"; -- 0.020743012241809054
	pesos_i(24865) := b"1111111111111111_1111111111111111_1110100101011100_1111011010101000"; -- -0.08842523956714857
	pesos_i(24866) := b"1111111111111111_1111111111111111_1110011010011100_0111101111001111"; -- -0.09917474942032116
	pesos_i(24867) := b"1111111111111111_1111111111111111_1110010110110010_1100010101000110"; -- -0.10274092723588568
	pesos_i(24868) := b"1111111111111111_1111111111111111_1101110111110100_0111101010010010"; -- -0.13298829973156867
	pesos_i(24869) := b"1111111111111111_1111111111111111_1101110101110010_0111010100110011"; -- -0.13497226240338703
	pesos_i(24870) := b"1111111111111111_1111111111111111_1101010100111110_0110001101010100"; -- -0.16701678459336178
	pesos_i(24871) := b"0000000000000000_0000000000000000_0000011000110001_0111110111110110"; -- 0.0241926885855768
	pesos_i(24872) := b"0000000000000000_0000000000000000_0010111100000111_1000101111001010"; -- 0.18370889363751866
	pesos_i(24873) := b"1111111111111111_1111111111111111_1111111001010111_1110110100100111"; -- -0.006470850068731455
	pesos_i(24874) := b"1111111111111111_1111111111111111_1110011101000110_1101110110101101"; -- -0.0965749218875541
	pesos_i(24875) := b"0000000000000000_0000000000000000_0010100000100101_1100001011011101"; -- 0.15682618994929579
	pesos_i(24876) := b"0000000000000000_0000000000000000_0000011011111011_1111011011100001"; -- 0.02728217129569234
	pesos_i(24877) := b"1111111111111111_1111111111111111_1110110101101111_0011110010100111"; -- -0.07252140932631757
	pesos_i(24878) := b"1111111111111111_1111111111111111_1101110110011100_0100111011010000"; -- -0.13433368120475112
	pesos_i(24879) := b"1111111111111111_1111111111111111_1111110111111110_0001001111100000"; -- -0.007841832909675493
	pesos_i(24880) := b"1111111111111111_1111111111111111_1110110100010001_1011100110011010"; -- -0.0739482878025995
	pesos_i(24881) := b"1111111111111111_1111111111111111_1101001111000011_0101111010111010"; -- -0.17280013991631238
	pesos_i(24882) := b"1111111111111111_1111111111111111_1111000110001110_0010101010011000"; -- -0.05642446315440202
	pesos_i(24883) := b"0000000000000000_0000000000000000_0000011110001101_0010000011010101"; -- 0.02949719628604836
	pesos_i(24884) := b"0000000000000000_0000000000000000_0000010111101011_0001111010110010"; -- 0.02311889512510387
	pesos_i(24885) := b"1111111111111111_1111111111111111_1101000100001101_0100100000011000"; -- -0.18339108860776673
	pesos_i(24886) := b"1111111111111111_1111111111111111_1101011000100010_1010001100010111"; -- -0.16353398027016405
	pesos_i(24887) := b"0000000000000000_0000000000000000_0010101110001001_0100100000010010"; -- 0.17006349991617606
	pesos_i(24888) := b"1111111111111111_1111111111111111_1101011011000001_1101110100100000"; -- -0.16110437367042107
	pesos_i(24889) := b"1111111111111111_1111111111111111_1111000010100111_1110000001001001"; -- -0.05993841367748748
	pesos_i(24890) := b"0000000000000000_0000000000000000_0000100100110000_0111001011111101"; -- 0.03589552565557325
	pesos_i(24891) := b"0000000000000000_0000000000000000_0001000101111110_1000001000101110"; -- 0.06833661663179007
	pesos_i(24892) := b"0000000000000000_0000000000000000_0001000101101100_0010101111100010"; -- 0.06805681488501131
	pesos_i(24893) := b"0000000000000000_0000000000000000_0000011011001101_0010101110011010"; -- 0.02656815064031757
	pesos_i(24894) := b"0000000000000000_0000000000000000_0001011001110110_1001111001111010"; -- 0.08774748313362894
	pesos_i(24895) := b"0000000000000000_0000000000000000_0000100100000100_1011100010001010"; -- 0.035228284599477196
	pesos_i(24896) := b"1111111111111111_1111111111111111_1101111111110001_0010100011101101"; -- -0.12522644255322674
	pesos_i(24897) := b"1111111111111111_1111111111111111_1101110110100110_1101001101110101"; -- -0.13417318721875784
	pesos_i(24898) := b"1111111111111111_1111111111111111_1111101011101011_1100001010101011"; -- -0.01984008137227393
	pesos_i(24899) := b"1111111111111111_1111111111111111_1110000110010010_1111011100101011"; -- -0.1188512344163662
	pesos_i(24900) := b"0000000000000000_0000000000000000_0000011011001111_1010011100011110"; -- 0.026606030261696084
	pesos_i(24901) := b"0000000000000000_0000000000000000_0000011011100000_0011000000111011"; -- 0.02685834345424156
	pesos_i(24902) := b"0000000000000000_0000000000000000_0000110001110100_0110011001011010"; -- 0.04865112027177745
	pesos_i(24903) := b"1111111111111111_1111111111111111_1101011111011011_1011101001000001"; -- -0.1568034736777797
	pesos_i(24904) := b"1111111111111111_1111111111111111_1111010110000001_0110011010110110"; -- -0.040994244128169224
	pesos_i(24905) := b"0000000000000000_0000000000000000_0000110011100100_1001011110010000"; -- 0.05036303783523884
	pesos_i(24906) := b"0000000000000000_0000000000000000_0010111110000001_0101010101111100"; -- 0.18556722904574904
	pesos_i(24907) := b"0000000000000000_0000000000000000_0001101001011010_0010011110100100"; -- 0.10293815377347675
	pesos_i(24908) := b"1111111111111111_1111111111111111_1101001100101100_0001111000110001"; -- -0.17510806377027818
	pesos_i(24909) := b"0000000000000000_0000000000000000_0010000000010110_1101101011100110"; -- 0.1253487407593362
	pesos_i(24910) := b"1111111111111111_1111111111111111_1110100010110101_1110001000100000"; -- -0.09097468102641716
	pesos_i(24911) := b"0000000000000000_0000000000000000_0001011110110110_1101011010110111"; -- 0.09263364767005891
	pesos_i(24912) := b"0000000000000000_0000000000000000_0000101100110001_0111101000100111"; -- 0.04372371151536362
	pesos_i(24913) := b"0000000000000000_0000000000000000_0010110011100110_1101100100110101"; -- 0.1753974680050891
	pesos_i(24914) := b"0000000000000000_0000000000000000_0000000010110010_0110000011110111"; -- 0.0027218440278144285
	pesos_i(24915) := b"1111111111111111_1111111111111111_1111100101110001_1100111010010100"; -- -0.02560719380078829
	pesos_i(24916) := b"1111111111111111_1111111111111111_1111110001100111_0000010010011010"; -- -0.01405307051074831
	pesos_i(24917) := b"1111111111111111_1111111111111111_1110011010100000_0011110001110011"; -- -0.09911749078544901
	pesos_i(24918) := b"0000000000000000_0000000000000000_0000101011101111_1101111011000101"; -- 0.042722628667041775
	pesos_i(24919) := b"1111111111111111_1111111111111111_1101010101101000_0010011011000010"; -- -0.16637952579282414
	pesos_i(24920) := b"0000000000000000_0000000000000000_0000010011110011_0011101000111110"; -- 0.019336357295831358
	pesos_i(24921) := b"0000000000000000_0000000000000000_0001111101110001_1010001011100101"; -- 0.12282770239929003
	pesos_i(24922) := b"0000000000000000_0000000000000000_0010001000100000_1000011100000011"; -- 0.13330882851320155
	pesos_i(24923) := b"1111111111111111_1111111111111111_1110010101000000_0000101100010110"; -- -0.1044915268085401
	pesos_i(24924) := b"0000000000000000_0000000000000000_0000000011100001_0001010011000011"; -- 0.0034344650300622984
	pesos_i(24925) := b"0000000000000000_0000000000000000_0001011001001111_1001111110010000"; -- 0.08715245503309496
	pesos_i(24926) := b"1111111111111111_1111111111111111_1110110011101000_1000010001101010"; -- -0.07457706842183796
	pesos_i(24927) := b"1111111111111111_1111111111111111_1111111100000111_0000000011110011"; -- -0.0037993818220623727
	pesos_i(24928) := b"0000000000000000_0000000000000000_0010010001101000_1000100001010110"; -- 0.1422200403020276
	pesos_i(24929) := b"0000000000000000_0000000000000000_0001100010111010_0101001000010101"; -- 0.09659302717322946
	pesos_i(24930) := b"1111111111111111_1111111111111111_1101011001010001_1101100011100000"; -- -0.16281361138608705
	pesos_i(24931) := b"1111111111111111_1111111111111111_1110100100011100_1001001101101011"; -- -0.08940771713991139
	pesos_i(24932) := b"0000000000000000_0000000000000000_0000000010011000_1011011110111001"; -- 0.002330286580720972
	pesos_i(24933) := b"0000000000000000_0000000000000000_0010101101110110_1101100111010111"; -- 0.16978227144929423
	pesos_i(24934) := b"1111111111111111_1111111111111111_1110111110111101_1110100001010101"; -- -0.06350849082501539
	pesos_i(24935) := b"1111111111111111_1111111111111111_1111011000100011_1101011000100101"; -- -0.03851567837406105
	pesos_i(24936) := b"1111111111111111_1111111111111111_1110110001100010_0101110100111010"; -- -0.07662408184571713
	pesos_i(24937) := b"1111111111111111_1111111111111111_1111101010011111_0110010010101011"; -- -0.021005352262335592
	pesos_i(24938) := b"1111111111111111_1111111111111111_1101000110011110_1100100000001110"; -- -0.18117093725010688
	pesos_i(24939) := b"1111111111111111_1111111111111111_1101011100100100_0101011101111010"; -- -0.15960171958880884
	pesos_i(24940) := b"0000000000000000_0000000000000000_0000101000000001_0001010010100000"; -- 0.03907898802381923
	pesos_i(24941) := b"1111111111111111_1111111111111111_1110011101001011_1110000000011111"; -- -0.0964984821596994
	pesos_i(24942) := b"1111111111111111_1111111111111111_1110111101100011_1111110000011000"; -- -0.06488060392404929
	pesos_i(24943) := b"0000000000000000_0000000000000000_0011010011111101_1111110011010100"; -- 0.20700054330040113
	pesos_i(24944) := b"0000000000000000_0000000000000000_0000011111000100_1110110111011101"; -- 0.03034865033742872
	pesos_i(24945) := b"1111111111111111_1111111111111111_1101001010011110_0111111110010000"; -- -0.17726900799174955
	pesos_i(24946) := b"1111111111111111_1111111111111111_1101010011100110_0010111100110110"; -- -0.16836266452812054
	pesos_i(24947) := b"1111111111111111_1111111111111111_1101000010000011_1110101010110110"; -- -0.18548710887281808
	pesos_i(24948) := b"1111111111111111_1111111111111111_1110101111111100_1011000011001000"; -- -0.07817549808926894
	pesos_i(24949) := b"0000000000000000_0000000000000000_0001110101010001_1111010011100110"; -- 0.11453180888874616
	pesos_i(24950) := b"0000000000000000_0000000000000000_0010110110011110_1000010000100011"; -- 0.17820001452238635
	pesos_i(24951) := b"0000000000000000_0000000000000000_0000000101100100_0110010000111101"; -- 0.005438103564091025
	pesos_i(24952) := b"1111111111111111_1111111111111111_1110001101100001_1010110011101101"; -- -0.11179084025541237
	pesos_i(24953) := b"0000000000000000_0000000000000000_0001100010101110_1001000110011101"; -- 0.09641370863816755
	pesos_i(24954) := b"0000000000000000_0000000000000000_0001111110110111_1100001010110101"; -- 0.12389771393213528
	pesos_i(24955) := b"0000000000000000_0000000000000000_0010111000101110_1011111100011000"; -- 0.1804007943206277
	pesos_i(24956) := b"1111111111111111_1111111111111111_1101111000110001_1110000011111001"; -- -0.1320514099645429
	pesos_i(24957) := b"0000000000000000_0000000000000000_0000101100111010_0111111000111101"; -- 0.043861284227930994
	pesos_i(24958) := b"1111111111111111_1111111111111111_1100111010010001_0011101000010001"; -- -0.1930965144675867
	pesos_i(24959) := b"1111111111111111_1111111111111111_1111010000110110_0110011001110111"; -- -0.04604491795635022
	pesos_i(24960) := b"1111111111111111_1111111111111111_1110101000101100_1001000001100110"; -- -0.08525750649998064
	pesos_i(24961) := b"0000000000000000_0000000000000000_0000110100100001_0001000110000000"; -- 0.05128583316868481
	pesos_i(24962) := b"0000000000000000_0000000000000000_0001010111011110_0001110000110100"; -- 0.0854203822409074
	pesos_i(24963) := b"0000000000000000_0000000000000000_0001111111101011_1111011001010101"; -- 0.12469424793934564
	pesos_i(24964) := b"0000000000000000_0000000000000000_0011010100100000_0100010110110101"; -- 0.20752368611688415
	pesos_i(24965) := b"1111111111111111_1111111111111111_1111110000111101_0011001011000000"; -- -0.01469118902412443
	pesos_i(24966) := b"1111111111111111_1111111111111111_1101110110010111_0110001010100011"; -- -0.13440879364890004
	pesos_i(24967) := b"1111111111111111_1111111111111111_1110011011100111_1100101100111001"; -- -0.09802560676471049
	pesos_i(24968) := b"1111111111111111_1111111111111111_1111010000101101_1110001000001011"; -- -0.0461748813253599
	pesos_i(24969) := b"1111111111111111_1111111111111111_1101001010111111_0110111101100111"; -- -0.1767664312759494
	pesos_i(24970) := b"0000000000000000_0000000000000000_0010100101110101_1110000001111011"; -- 0.16195490840236224
	pesos_i(24971) := b"0000000000000000_0000000000000000_0001100000001000_0111111001000001"; -- 0.09387959565746513
	pesos_i(24972) := b"0000000000000000_0000000000000000_0010000010011101_1011000001000001"; -- 0.12740613536594805
	pesos_i(24973) := b"1111111111111111_1111111111111111_1111011011010111_1100101000011100"; -- -0.035769813603677904
	pesos_i(24974) := b"0000000000000000_0000000000000000_0000100000111001_1011101001010100"; -- 0.03213085696646421
	pesos_i(24975) := b"0000000000000000_0000000000000000_0010111111001101_0000011110000110"; -- 0.1867222502146092
	pesos_i(24976) := b"0000000000000000_0000000000000000_0001010000111010_0011001100101111"; -- 0.07901306059922625
	pesos_i(24977) := b"0000000000000000_0000000000000000_0001011111101101_0001011110011110"; -- 0.0934614905865533
	pesos_i(24978) := b"0000000000000000_0000000000000000_0010011000101010_1101100001000010"; -- 0.14909125921096267
	pesos_i(24979) := b"1111111111111111_1111111111111111_1101011000010010_0010000111011001"; -- -0.16378582440621053
	pesos_i(24980) := b"0000000000000000_0000000000000000_0001001000110111_0001101011101001"; -- 0.0711533372695393
	pesos_i(24981) := b"1111111111111111_1111111111111111_1100111110000011_0010011101111001"; -- -0.18940499580520087
	pesos_i(24982) := b"1111111111111111_1111111111111111_1101101110110001_0101011011111010"; -- -0.14182526014676614
	pesos_i(24983) := b"1111111111111111_1111111111111111_1111101101010111_0101111111110101"; -- -0.018198015771199016
	pesos_i(24984) := b"1111111111111111_1111111111111111_1110101011101100_0000011111110011"; -- -0.0823359520871665
	pesos_i(24985) := b"1111111111111111_1111111111111111_1101010011000100_0001001011111010"; -- -0.16888314628819986
	pesos_i(24986) := b"0000000000000000_0000000000000000_0000110000111111_0100110001010011"; -- 0.04784085297027006
	pesos_i(24987) := b"0000000000000000_0000000000000000_0000100011001111_0001100101000110"; -- 0.034410075818119897
	pesos_i(24988) := b"0000000000000000_0000000000000000_0001001111011100_0000001111001101"; -- 0.07757591004102596
	pesos_i(24989) := b"0000000000000000_0000000000000000_0010000110110110_0111000000010010"; -- 0.13169002944472
	pesos_i(24990) := b"1111111111111111_1111111111111111_1110001110110110_0000001111010010"; -- -0.11050392269244257
	pesos_i(24991) := b"0000000000000000_0000000000000000_0001000111011111_1010110011111001"; -- 0.06981927002428313
	pesos_i(24992) := b"0000000000000000_0000000000000000_0000000010010101_0011111111001010"; -- 0.0022773615800243028
	pesos_i(24993) := b"1111111111111111_1111111111111111_1101110001010011_0000010101001110"; -- -0.1393582042882058
	pesos_i(24994) := b"1111111111111111_1111111111111111_1110100000101100_1010001110000110"; -- -0.09306886649606692
	pesos_i(24995) := b"0000000000000000_0000000000000000_0001010110000100_0111100010010011"; -- 0.08405259700555602
	pesos_i(24996) := b"1111111111111111_1111111111111111_1110011101100110_0011111101000010"; -- -0.09609608305509233
	pesos_i(24997) := b"0000000000000000_0000000000000000_0000100010110101_1011101101010100"; -- 0.03402300646474498
	pesos_i(24998) := b"0000000000000000_0000000000000000_0000000001111110_0100101010111001"; -- 0.0019270611539875476
	pesos_i(24999) := b"1111111111111111_1111111111111111_1100111100111111_1000100111101011"; -- -0.19043672568404268
	pesos_i(25000) := b"1111111111111111_1111111111111111_1101010011111011_0001111100110101"; -- -0.16804318396483217
	pesos_i(25001) := b"1111111111111111_1111111111111111_1111100100010011_1111010001101100"; -- -0.02703926437354106
	pesos_i(25002) := b"0000000000000000_0000000000000000_0010110111101011_0001001111011010"; -- 0.17936824865203554
	pesos_i(25003) := b"1111111111111111_1111111111111111_1110100001100110_0011011001010100"; -- -0.09219036530965649
	pesos_i(25004) := b"1111111111111111_1111111111111111_1101010101011110_1010001111110110"; -- -0.1665246511088812
	pesos_i(25005) := b"0000000000000000_0000000000000000_0001000001011000_0110101110001101"; -- 0.06384918391190163
	pesos_i(25006) := b"0000000000000000_0000000000000000_0000111100011110_0001111100001100"; -- 0.05905336420633972
	pesos_i(25007) := b"1111111111111111_1111111111111111_1111110010010001_0011110110100110"; -- -0.013408801164968842
	pesos_i(25008) := b"1111111111111111_1111111111111111_1111001000100000_1100010111000010"; -- -0.05418743145745317
	pesos_i(25009) := b"0000000000000000_0000000000000000_0001111011111010_0001110011001001"; -- 0.12100391300483353
	pesos_i(25010) := b"0000000000000000_0000000000000000_0001110110100001_0010111100000001"; -- 0.11574071667649155
	pesos_i(25011) := b"1111111111111111_1111111111111111_1110000001110011_1001011101101001"; -- -0.12323621452400352
	pesos_i(25012) := b"1111111111111111_1111111111111111_1101000101101110_1001110111011100"; -- -0.1819058739723932
	pesos_i(25013) := b"0000000000000000_0000000000000000_0000101011000001_1100111011000111"; -- 0.042019771261387416
	pesos_i(25014) := b"0000000000000000_0000000000000000_0001011000110111_1010111011101000"; -- 0.08678715864288282
	pesos_i(25015) := b"0000000000000000_0000000000000000_0000100000001101_0101001010000100"; -- 0.0314532824845297
	pesos_i(25016) := b"1111111111111111_1111111111111111_1101010000101100_1011000000001000"; -- -0.17119312095157085
	pesos_i(25017) := b"1111111111111111_1111111111111111_1110101000110011_1000101000010010"; -- -0.08515107215866208
	pesos_i(25018) := b"0000000000000000_0000000000000000_0000110110110010_1000000100000011"; -- 0.05350500418931971
	pesos_i(25019) := b"1111111111111111_1111111111111111_1111101001110011_1010000010010101"; -- -0.02167316770740672
	pesos_i(25020) := b"0000000000000000_0000000000000000_0010101110101101_1011111101110011"; -- 0.1706199317290058
	pesos_i(25021) := b"0000000000000000_0000000000000000_0000110011101011_1100001010110100"; -- 0.05047242064563364
	pesos_i(25022) := b"0000000000000000_0000000000000000_0000000101100100_0100001001100010"; -- 0.005436085627984894
	pesos_i(25023) := b"0000000000000000_0000000000000000_0001001001001100_1110011100000011"; -- 0.07148593731541027
	pesos_i(25024) := b"1111111111111111_1111111111111111_1110110000000110_0110001101101011"; -- -0.07802752151285615
	pesos_i(25025) := b"0000000000000000_0000000000000000_0010110100110111_0000001001101011"; -- 0.17662062748779891
	pesos_i(25026) := b"0000000000000000_0000000000000000_0000111111110010_0100011011011111"; -- 0.06229060129892991
	pesos_i(25027) := b"0000000000000000_0000000000000000_0001101101100111_1011101001100100"; -- 0.10705151504324681
	pesos_i(25028) := b"0000000000000000_0000000000000000_0001000100110110_0111101011011101"; -- 0.06723754773400308
	pesos_i(25029) := b"1111111111111111_1111111111111111_1100110011001000_1010010000010010"; -- -0.20006346283482213
	pesos_i(25030) := b"1111111111111111_1111111111111111_1110011001000101_1101000010100011"; -- -0.10049720788062144
	pesos_i(25031) := b"1111111111111111_1111111111111111_1110111110010101_0100010101100110"; -- -0.0641285540677553
	pesos_i(25032) := b"1111111111111111_1111111111111111_1111100010010000_0001000010010111"; -- -0.029051745641975033
	pesos_i(25033) := b"0000000000000000_0000000000000000_0001001101010001_1011100001000111"; -- 0.07546569567041904
	pesos_i(25034) := b"0000000000000000_0000000000000000_0000110110010100_1110010111000110"; -- 0.05305324629736169
	pesos_i(25035) := b"0000000000000000_0000000000000000_0010100101100000_0001100111110101"; -- 0.16162264087845987
	pesos_i(25036) := b"0000000000000000_0000000000000000_0010111111001011_1111011010001110"; -- 0.1867059800377046
	pesos_i(25037) := b"0000000000000000_0000000000000000_0010010011100010_1100110101111100"; -- 0.14408573411688214
	pesos_i(25038) := b"1111111111111111_1111111111111111_1110010101010000_1000100110110110"; -- -0.10423983857940353
	pesos_i(25039) := b"0000000000000000_0000000000000000_0001100100010100_0100011110111111"; -- 0.09796570209368306
	pesos_i(25040) := b"1111111111111111_1111111111111111_1101001100001000_0100110000111111"; -- -0.1756546350785741
	pesos_i(25041) := b"0000000000000000_0000000000000000_0000111101110001_0000111000111011"; -- 0.06031884137847621
	pesos_i(25042) := b"0000000000000000_0000000000000000_0001011001101100_0101011011001000"; -- 0.08759062184485991
	pesos_i(25043) := b"0000000000000000_0000000000000000_0000101110110000_1101100110100010"; -- 0.045667268770307176
	pesos_i(25044) := b"0000000000000000_0000000000000000_0001011100010101_1001000110011001"; -- 0.0901728629685392
	pesos_i(25045) := b"1111111111111111_1111111111111111_1111111101110110_0011110100100100"; -- -0.002102068725775122
	pesos_i(25046) := b"1111111111111111_1111111111111111_1100100001100110_0100000000110100"; -- -0.21718977674685924
	pesos_i(25047) := b"1111111111111111_1111111111111111_1110001101110110_1001101101111011"; -- -0.11147144545392025
	pesos_i(25048) := b"0000000000000000_0000000000000000_0010101010100001_0101100101111010"; -- 0.1665244981871073
	pesos_i(25049) := b"1111111111111111_1111111111111111_1111100110000011_1111010101010000"; -- -0.025330226827650047
	pesos_i(25050) := b"1111111111111111_1111111111111111_1111000110101001_1000000001111000"; -- -0.05600735727098558
	pesos_i(25051) := b"1111111111111111_1111111111111111_1111110000110001_1000110111011011"; -- -0.014868864016146142
	pesos_i(25052) := b"0000000000000000_0000000000000000_0010101010100110_0011110101110111"; -- 0.1665991226186076
	pesos_i(25053) := b"1111111111111111_1111111111111111_1110101110110011_0001110000111101"; -- -0.07929824370539162
	pesos_i(25054) := b"1111111111111111_1111111111111111_1110110101010010_0011000011111111"; -- -0.07296460884468685
	pesos_i(25055) := b"0000000000000000_0000000000000000_0010010100001010_1110100000101101"; -- 0.1446976765914795
	pesos_i(25056) := b"0000000000000000_0000000000000000_0001011010101111_1101110010110101"; -- 0.08862094329831399
	pesos_i(25057) := b"1111111111111111_1111111111111111_1100110111111000_0010010100100110"; -- -0.19543235619378874
	pesos_i(25058) := b"0000000000000000_0000000000000000_0010010000100011_1110101000110011"; -- 0.14117301698265802
	pesos_i(25059) := b"0000000000000000_0000000000000000_0000110000100111_1011110110010100"; -- 0.04748139260176896
	pesos_i(25060) := b"0000000000000000_0000000000000000_0001001000001110_0110111100110011"; -- 0.07053275104463388
	pesos_i(25061) := b"0000000000000000_0000000000000000_0011001111000011_0000110101100101"; -- 0.20219501215371796
	pesos_i(25062) := b"1111111111111111_1111111111111111_1110100100110101_1010000100000100"; -- -0.08902543678602644
	pesos_i(25063) := b"0000000000000000_0000000000000000_0000111011100101_1101001010111011"; -- 0.05819432323793825
	pesos_i(25064) := b"1111111111111111_1111111111111111_1110010000101000_1110111011110000"; -- -0.10875040653808982
	pesos_i(25065) := b"0000000000000000_0000000000000000_0000111011010010_1101101111110111"; -- 0.05790495665997399
	pesos_i(25066) := b"1111111111111111_1111111111111111_1100101111010001_1101010111001110"; -- -0.20382941928551265
	pesos_i(25067) := b"1111111111111111_1111111111111111_1101110010000111_1010111110101111"; -- -0.13855459193182473
	pesos_i(25068) := b"0000000000000000_0000000000000000_0001001001011111_0110001110110100"; -- 0.07176802779161043
	pesos_i(25069) := b"0000000000000000_0000000000000000_0000111001001111_0011010110111011"; -- 0.055896146907801786
	pesos_i(25070) := b"0000000000000000_0000000000000000_0001010011001010_1010011011101110"; -- 0.08121722517538113
	pesos_i(25071) := b"1111111111111111_1111111111111111_1111001001100111_1100111010011011"; -- -0.05310353018274249
	pesos_i(25072) := b"0000000000000000_0000000000000000_0000100000110010_1101000100011100"; -- 0.032025403418370055
	pesos_i(25073) := b"0000000000000000_0000000000000000_0010000010111011_0110001111010101"; -- 0.12785934411746136
	pesos_i(25074) := b"0000000000000000_0000000000000000_0001000011111100_1010111001001001"; -- 0.06635560315623869
	pesos_i(25075) := b"0000000000000000_0000000000000000_0010000010000011_0000001000000110"; -- 0.1269990220173844
	pesos_i(25076) := b"0000000000000000_0000000000000000_0010010111001110_1101101110011010"; -- 0.1476876497395095
	pesos_i(25077) := b"0000000000000000_0000000000000000_0011001001010110_0110101111101011"; -- 0.19663118819340125
	pesos_i(25078) := b"1111111111111111_1111111111111111_1110111001000100_1010110101111011"; -- -0.06926456202372536
	pesos_i(25079) := b"0000000000000000_0000000000000000_0001111101000010_0000010110010100"; -- 0.1221011625967133
	pesos_i(25080) := b"1111111111111111_1111111111111111_1110010000110101_0100100000100011"; -- -0.10856198446513447
	pesos_i(25081) := b"0000000000000000_0000000000000000_0010001101001111_0011011001011001"; -- 0.13792743380676029
	pesos_i(25082) := b"1111111111111111_1111111111111111_1101100000000000_0000000110110110"; -- -0.15624989803288536
	pesos_i(25083) := b"0000000000000000_0000000000000000_0000000110010111_1100011111000000"; -- 0.006222233233577035
	pesos_i(25084) := b"1111111111111111_1111111111111111_1101111010011010_1101001111111011"; -- -0.13045001154558494
	pesos_i(25085) := b"0000000000000000_0000000000000000_0000110101110010_1100111110110011"; -- 0.05253313182699146
	pesos_i(25086) := b"1111111111111111_1111111111111111_1110000010010000_0011110110111101"; -- -0.12279905452239742
	pesos_i(25087) := b"0000000000000000_0000000000000000_0000000000100010_0000111101000101"; -- 0.0005197089876763063
	pesos_i(25088) := b"0000000000000000_0000000000000000_0001100101101011_1001001111010111"; -- 0.09929775225679813
	pesos_i(25089) := b"0000000000000000_0000000000000000_0010100011110111_1010110000110001"; -- 0.1600291843764145
	pesos_i(25090) := b"1111111111111111_1111111111111111_1110100010010001_1110001101011011"; -- -0.09152392413999812
	pesos_i(25091) := b"0000000000000000_0000000000000000_0001101000101010_1010111010101101"; -- 0.10221378064115774
	pesos_i(25092) := b"1111111111111111_1111111111111111_1110101111010100_1110100110001000"; -- -0.0787824670677973
	pesos_i(25093) := b"1111111111111111_1111111111111111_1101010101010000_1101011110101100"; -- -0.16673519188591449
	pesos_i(25094) := b"1111111111111111_1111111111111111_1110001111001100_0001000111000110"; -- -0.11016739760352953
	pesos_i(25095) := b"0000000000000000_0000000000000000_0010010101001001_1000111110010111"; -- 0.14565370025678093
	pesos_i(25096) := b"0000000000000000_0000000000000000_0010111010101101_1011111111100101"; -- 0.18233870841979907
	pesos_i(25097) := b"1111111111111111_1111111111111111_1101001101011010_0011011011001011"; -- -0.1744046931013217
	pesos_i(25098) := b"1111111111111111_1111111111111111_1110101010101101_1100001001001111"; -- -0.08328614787165535
	pesos_i(25099) := b"1111111111111111_1111111111111111_1110011110100111_0000110011100100"; -- -0.09510726388591507
	pesos_i(25100) := b"0000000000000000_0000000000000000_0000001001100111_0110101000100101"; -- 0.00939048191206394
	pesos_i(25101) := b"1111111111111111_1111111111111111_1101000010001110_0010011011010110"; -- -0.1853309372081655
	pesos_i(25102) := b"0000000000000000_0000000000000000_0010010000000011_0000101001010110"; -- 0.14067139251992203
	pesos_i(25103) := b"1111111111111111_1111111111111111_1110111000111100_0100111100011101"; -- -0.06939225712455097
	pesos_i(25104) := b"0000000000000000_0000000000000000_0001111111011110_1011010110110110"; -- 0.12449203193223624
	pesos_i(25105) := b"0000000000000000_0000000000000000_0000000101001100_0011110100000000"; -- 0.005069553889720377
	pesos_i(25106) := b"0000000000000000_0000000000000000_0000100001101100_1101111000000110"; -- 0.03291118295626492
	pesos_i(25107) := b"0000000000000000_0000000000000000_0010111111110010_0000110001110101"; -- 0.18728711940891637
	pesos_i(25108) := b"0000000000000000_0000000000000000_0010110010000011_0001110110011001"; -- 0.17387566559761583
	pesos_i(25109) := b"0000000000000000_0000000000000000_0010100101101001_0000001011001011"; -- 0.16175858931604944
	pesos_i(25110) := b"0000000000000000_0000000000000000_0000000110011000_0111011100100110"; -- 0.006232687656921861
	pesos_i(25111) := b"1111111111111111_1111111111111111_1110010110011011_0111001000110000"; -- -0.10309683163085627
	pesos_i(25112) := b"1111111111111111_1111111111111111_1100110111110000_1010011001110110"; -- -0.1955467187237049
	pesos_i(25113) := b"1111111111111111_1111111111111111_1100111000111010_0010101101111000"; -- -0.1944248993501507
	pesos_i(25114) := b"0000000000000000_0000000000000000_0000001110101000_1111011001011110"; -- 0.014296911135328159
	pesos_i(25115) := b"0000000000000000_0000000000000000_0001100100111101_0000001100001111"; -- 0.09858721846600917
	pesos_i(25116) := b"0000000000000000_0000000000000000_0000110110110101_1000111010011101"; -- 0.05355159134859417
	pesos_i(25117) := b"1111111111111111_1111111111111111_1101000011000000_1001011100000011"; -- -0.1845613116034117
	pesos_i(25118) := b"1111111111111111_1111111111111111_1111110011101010_1111101010000011"; -- -0.012039511772071899
	pesos_i(25119) := b"1111111111111111_1111111111111111_1110111101111001_0001011010011100"; -- -0.06455858890841132
	pesos_i(25120) := b"0000000000000000_0000000000000000_0000010001011000_0010010010111000"; -- 0.016969962027003953
	pesos_i(25121) := b"1111111111111111_1111111111111111_1111011000000101_0111010010010100"; -- -0.03897925743223004
	pesos_i(25122) := b"1111111111111111_1111111111111111_1110100111010110_0010100110111100"; -- -0.0865758816452094
	pesos_i(25123) := b"0000000000000000_0000000000000000_0001001010011100_1011010010000100"; -- 0.0727036306122636
	pesos_i(25124) := b"1111111111111111_1111111111111111_1110101100111111_1111100100101111"; -- -0.08105509378292355
	pesos_i(25125) := b"0000000000000000_0000000000000000_0000110010110010_1101010111010100"; -- 0.04960380967003202
	pesos_i(25126) := b"1111111111111111_1111111111111111_1110011001010001_1101101111000011"; -- -0.1003134392550312
	pesos_i(25127) := b"0000000000000000_0000000000000000_0010000100001010_1101001011011110"; -- 0.12907140647589316
	pesos_i(25128) := b"0000000000000000_0000000000000000_0001010001101100_1100000111000100"; -- 0.07978449845239385
	pesos_i(25129) := b"0000000000000000_0000000000000000_0010000011011100_1011001100111001"; -- 0.12836761606807442
	pesos_i(25130) := b"1111111111111111_1111111111111111_1111101001011011_0110101111011111"; -- -0.022042520467674503
	pesos_i(25131) := b"1111111111111111_1111111111111111_1100101011000000_0000010001100000"; -- -0.20800755166829937
	pesos_i(25132) := b"0000000000000000_0000000000000000_0000001100011101_0010110111001001"; -- 0.012163983973171802
	pesos_i(25133) := b"1111111111111111_1111111111111111_1110010010100000_1011100100111001"; -- -0.10692255366300804
	pesos_i(25134) := b"0000000000000000_0000000000000000_0010000001101000_1001101010110100"; -- 0.12659613505389442
	pesos_i(25135) := b"1111111111111111_1111111111111111_1110101011101101_0010101001000111"; -- -0.0823186471395388
	pesos_i(25136) := b"0000000000000000_0000000000000000_0010111111010110_0101010000010111"; -- 0.1868641429956626
	pesos_i(25137) := b"0000000000000000_0000000000000000_0001111110000100_0011010111110011"; -- 0.12311112585943698
	pesos_i(25138) := b"0000000000000000_0000000000000000_0000001010110010_0110010101101010"; -- 0.010534609296858611
	pesos_i(25139) := b"1111111111111111_1111111111111111_1101010100010111_0101110011011100"; -- -0.16761226296388587
	pesos_i(25140) := b"0000000000000000_0000000000000000_0001001111001000_0000101100000000"; -- 0.07727116354987279
	pesos_i(25141) := b"0000000000000000_0000000000000000_0010101101011100_0000011101000010"; -- 0.16937299112546672
	pesos_i(25142) := b"0000000000000000_0000000000000000_0001011001111111_1011101101101001"; -- 0.08788653679173931
	pesos_i(25143) := b"1111111111111111_1111111111111111_1100110010000011_0111100111011111"; -- -0.20111883466110922
	pesos_i(25144) := b"0000000000000000_0000000000000000_0000000111001100_0011100110000100"; -- 0.0070224712259780156
	pesos_i(25145) := b"0000000000000000_0000000000000000_0001011011011100_1000101001000011"; -- 0.08930267464940646
	pesos_i(25146) := b"0000000000000000_0000000000000000_0000111111000100_1010011110111111"; -- 0.061594471019909496
	pesos_i(25147) := b"1111111111111111_1111111111111111_1111010101100001_1010100010011110"; -- -0.04147859700303206
	pesos_i(25148) := b"1111111111111111_1111111111111111_1111001111100100_0010101101001001"; -- -0.04729966618488665
	pesos_i(25149) := b"1111111111111111_1111111111111111_1110010110111111_0110111100110010"; -- -0.10254769354957227
	pesos_i(25150) := b"0000000000000000_0000000000000000_0010011111110011_0011101011100011"; -- 0.15605514564882175
	pesos_i(25151) := b"0000000000000000_0000000000000000_0010101011100001_1101110100011001"; -- 0.1675089059929911
	pesos_i(25152) := b"1111111111111111_1111111111111111_1111101110101011_1011101111110100"; -- -0.01691079416783616
	pesos_i(25153) := b"0000000000000000_0000000000000000_0000011111000110_1110110011000100"; -- 0.030379102623572105
	pesos_i(25154) := b"1111111111111111_1111111111111111_1111101000011100_0000100010010101"; -- -0.0230097424134539
	pesos_i(25155) := b"0000000000000000_0000000000000000_0001110000000110_1110010100000110"; -- 0.10948020353697585
	pesos_i(25156) := b"0000000000000000_0000000000000000_0011000010111001_0100011101011001"; -- 0.19032712872826849
	pesos_i(25157) := b"0000000000000000_0000000000000000_0000001101011110_0010110011010011"; -- 0.013155747970271116
	pesos_i(25158) := b"1111111111111111_1111111111111111_1111111100101001_1000111000001001"; -- -0.0032721735774358532
	pesos_i(25159) := b"0000000000000000_0000000000000000_0001101100000000_1100100000111001"; -- 0.10548068421408327
	pesos_i(25160) := b"1111111111111111_1111111111111111_1110010110011000_0111111111001010"; -- -0.10314179721079791
	pesos_i(25161) := b"1111111111111111_1111111111111111_1110101110110111_0011011101100010"; -- -0.07923559052930372
	pesos_i(25162) := b"0000000000000000_0000000000000000_0000001111001011_0010101001011100"; -- 0.014818809040917308
	pesos_i(25163) := b"1111111111111111_1111111111111111_1111101011011111_1000011000000110"; -- -0.020026801628445782
	pesos_i(25164) := b"0000000000000000_0000000000000000_0001001001100011_1000101100111010"; -- 0.07183141861134601
	pesos_i(25165) := b"0000000000000000_0000000000000000_0010000000010100_1001010011000111"; -- 0.12531404354086503
	pesos_i(25166) := b"1111111111111111_1111111111111111_1110001100000000_0001001101100101"; -- -0.11328009401149954
	pesos_i(25167) := b"1111111111111111_1111111111111111_1111010100111001_0011010010000000"; -- -0.04209586980041161
	pesos_i(25168) := b"0000000000000000_0000000000000000_0000000010000101_1000011010110010"; -- 0.002037447331871093
	pesos_i(25169) := b"0000000000000000_0000000000000000_0010001000010100_0011000100000001"; -- 0.13312059663152812
	pesos_i(25170) := b"1111111111111111_1111111111111111_1101010010101001_0000011000011001"; -- -0.16929590111399573
	pesos_i(25171) := b"0000000000000000_0000000000000000_0001000000000101_1010101110110010"; -- 0.06258652777791955
	pesos_i(25172) := b"0000000000000000_0000000000000000_0001010110111001_1100001010010101"; -- 0.08486572388031867
	pesos_i(25173) := b"1111111111111111_1111111111111111_1101000101001101_1001000000100001"; -- -0.18241023243535212
	pesos_i(25174) := b"1111111111111111_1111111111111111_1110010110000000_0110001001011101"; -- -0.10350976201544221
	pesos_i(25175) := b"0000000000000000_0000000000000000_0000001011110001_0101011100110110"; -- 0.011495066330203944
	pesos_i(25176) := b"0000000000000000_0000000000000000_0001010001011011_1011000100010001"; -- 0.07952410387591821
	pesos_i(25177) := b"0000000000000000_0000000000000000_0000010110110100_0111010110111100"; -- 0.022284849512155223
	pesos_i(25178) := b"0000000000000000_0000000000000000_0001110001101001_1010011010111100"; -- 0.11098711094066954
	pesos_i(25179) := b"1111111111111111_1111111111111111_1111000110100010_0100001000100011"; -- -0.0561178840825369
	pesos_i(25180) := b"0000000000000000_0000000000000000_0001101111100101_1101111100001000"; -- 0.10897630650823995
	pesos_i(25181) := b"0000000000000000_0000000000000000_0001100100001100_0011000001000000"; -- 0.09784223127747126
	pesos_i(25182) := b"1111111111111111_1111111111111111_1100110000110101_1001111110110001"; -- -0.20230676586808843
	pesos_i(25183) := b"1111111111111111_1111111111111111_1111101101110101_1000100011001010"; -- -0.017737818476146732
	pesos_i(25184) := b"0000000000000000_0000000000000000_0000001111010010_0000000001010100"; -- 0.014923115279700565
	pesos_i(25185) := b"0000000000000000_0000000000000000_0010100010000011_0010110111101100"; -- 0.15825163854920632
	pesos_i(25186) := b"1111111111111111_1111111111111111_1111011101001101_0010100011111111"; -- -0.03397887968882801
	pesos_i(25187) := b"0000000000000000_0000000000000000_0010001010100000_1011111101011000"; -- 0.1352653112591501
	pesos_i(25188) := b"1111111111111111_1111111111111111_1111111110111001_0000110100111010"; -- -0.0010825856449231917
	pesos_i(25189) := b"0000000000000000_0000000000000000_0011010000000101_0011011110101101"; -- 0.2032046125911541
	pesos_i(25190) := b"0000000000000000_0000000000000000_0000001011001101_0011110100000110"; -- 0.010944188994916506
	pesos_i(25191) := b"1111111111111111_1111111111111111_1110001101111110_0100011000001001"; -- -0.111354468215931
	pesos_i(25192) := b"1111111111111111_1111111111111111_1110000101101010_1001000010101011"; -- -0.11946769536459768
	pesos_i(25193) := b"0000000000000000_0000000000000000_0001001001001110_1111000100010101"; -- 0.07151705509952735
	pesos_i(25194) := b"1111111111111111_1111111111111111_1111001100110011_0000110101011000"; -- -0.05000225647493399
	pesos_i(25195) := b"0000000000000000_0000000000000000_0000010101110011_1011111011011010"; -- 0.021297386290565955
	pesos_i(25196) := b"0000000000000000_0000000000000000_0001001010000010_0011111011101001"; -- 0.07229989234297535
	pesos_i(25197) := b"1111111111111111_1111111111111111_1110000011011011_0000101100011111"; -- -0.12165766232930317
	pesos_i(25198) := b"1111111111111111_1111111111111111_1110011010010111_0001101111000111"; -- -0.09925676726531049
	pesos_i(25199) := b"1111111111111111_1111111111111111_1110011010001011_0000011111010101"; -- -0.09944106144867296
	pesos_i(25200) := b"1111111111111111_1111111111111111_1110000011011110_1011011100001000"; -- -0.1216016392620216
	pesos_i(25201) := b"0000000000000000_0000000000000000_0001001111010000_0011111111110110"; -- 0.07739639041152661
	pesos_i(25202) := b"1111111111111111_1111111111111111_1101000110100000_1011000100111011"; -- -0.18114177994805655
	pesos_i(25203) := b"0000000000000000_0000000000000000_0010101011011100_0010000000000110"; -- 0.16742134228526975
	pesos_i(25204) := b"1111111111111111_1111111111111111_1101100010101010_0110010001000010"; -- -0.15365003002452626
	pesos_i(25205) := b"0000000000000000_0000000000000000_0001110010000100_0001000011010110"; -- 0.11139016368246063
	pesos_i(25206) := b"0000000000000000_0000000000000000_0010100000001110_1011010011001101"; -- 0.1564743997035564
	pesos_i(25207) := b"0000000000000000_0000000000000000_0001110100010101_0010011100101111"; -- 0.11360402017316917
	pesos_i(25208) := b"0000000000000000_0000000000000000_0010100001101011_0110110000001110"; -- 0.15788913093615375
	pesos_i(25209) := b"0000000000000000_0000000000000000_0000110001111000_0111111001111111"; -- 0.04871359449551662
	pesos_i(25210) := b"1111111111111111_1111111111111111_1111011010101101_1011111000001001"; -- -0.036411402600037474
	pesos_i(25211) := b"1111111111111111_1111111111111111_1100111111100100_0101011011001000"; -- -0.18792207358198942
	pesos_i(25212) := b"0000000000000000_0000000000000000_0000000011011010_1010111101110100"; -- 0.003336873772706614
	pesos_i(25213) := b"0000000000000000_0000000000000000_0011000101101110_0101001011111001"; -- 0.1930896622799049
	pesos_i(25214) := b"1111111111111111_1111111111111111_1101000111100100_1101001100100100"; -- -0.18010216124563447
	pesos_i(25215) := b"1111111111111111_1111111111111111_1110000001101100_1001110110010111"; -- -0.12334265777552121
	pesos_i(25216) := b"0000000000000000_0000000000000000_0010011101010100_0001011011000110"; -- 0.15362684578617883
	pesos_i(25217) := b"0000000000000000_0000000000000000_0001011110000111_0000001100111111"; -- 0.09190388002895972
	pesos_i(25218) := b"0000000000000000_0000000000000000_0010101011110110_0110000110010011"; -- 0.16782197800130355
	pesos_i(25219) := b"0000000000000000_0000000000000000_0001000101001000_1110111000111001"; -- 0.06751908202072884
	pesos_i(25220) := b"1111111111111111_1111111111111111_1111111010010001_0100011101010111"; -- -0.005595723290426736
	pesos_i(25221) := b"1111111111111111_1111111111111111_1101101101100110_1010011111111100"; -- -0.1429648407790556
	pesos_i(25222) := b"1111111111111111_1111111111111111_1101100001001101_0111100111001011"; -- -0.1550678137900152
	pesos_i(25223) := b"1111111111111111_1111111111111111_1101011100110101_1100001100100110"; -- -0.1593359024650088
	pesos_i(25224) := b"0000000000000000_0000000000000000_0001111101101011_1111101111000010"; -- 0.12274144644082315
	pesos_i(25225) := b"0000000000000000_0000000000000000_0001100101101000_1110001001000101"; -- 0.09925665088161255
	pesos_i(25226) := b"0000000000000000_0000000000000000_0010111001001100_1100011101110111"; -- 0.18085905703657926
	pesos_i(25227) := b"0000000000000000_0000000000000000_0000011000100110_0010010010100101"; -- 0.024019518155764592
	pesos_i(25228) := b"1111111111111111_1111111111111111_1111111011100000_1011110011011100"; -- -0.004383274417610669
	pesos_i(25229) := b"1111111111111111_1111111111111111_1101001101010011_0111110010011011"; -- -0.1745073434783149
	pesos_i(25230) := b"1111111111111111_1111111111111111_1100101111000001_0100101110011111"; -- -0.20408179631617882
	pesos_i(25231) := b"1111111111111111_1111111111111111_1111011000100011_1000010111101000"; -- -0.038520460988687846
	pesos_i(25232) := b"0000000000000000_0000000000000000_0011001000101101_1000100010011100"; -- 0.19600728807149911
	pesos_i(25233) := b"0000000000000000_0000000000000000_0010101010010010_0101000100001001"; -- 0.16629511325431104
	pesos_i(25234) := b"1111111111111111_1111111111111111_1101010000110110_1110110110111111"; -- -0.17103685460475498
	pesos_i(25235) := b"0000000000000000_0000000000000000_0001001001001010_1100110110110100"; -- 0.07145391125375299
	pesos_i(25236) := b"0000000000000000_0000000000000000_0000111010011001_0000000010110110"; -- 0.05702213699183533
	pesos_i(25237) := b"0000000000000000_0000000000000000_0000100110000110_1100110100100001"; -- 0.037213154336588665
	pesos_i(25238) := b"1111111111111111_1111111111111111_1101000101000011_1010111000111100"; -- -0.18256102602024085
	pesos_i(25239) := b"1111111111111111_1111111111111111_1111010101010100_1101010100110111"; -- -0.04167430307023667
	pesos_i(25240) := b"1111111111111111_1111111111111111_1111101111001101_0011100011010110"; -- -0.016399810667225668
	pesos_i(25241) := b"0000000000000000_0000000000000000_0001100100101110_0101001010110110"; -- 0.09836308427134706
	pesos_i(25242) := b"0000000000000000_0000000000000000_0000110010100110_1110110001011010"; -- 0.04942204673794894
	pesos_i(25243) := b"0000000000000000_0000000000000000_0010001010111011_1111100110111111"; -- 0.13568077948381368
	pesos_i(25244) := b"1111111111111111_1111111111111111_1111101111011011_1000111110110110"; -- -0.01618100946393174
	pesos_i(25245) := b"1111111111111111_1111111111111111_1101110000001010_1010000100100110"; -- -0.14046280693108576
	pesos_i(25246) := b"1111111111111111_1111111111111111_1111010101001101_0010011000101000"; -- -0.04179154896411341
	pesos_i(25247) := b"1111111111111111_1111111111111111_1111010110001111_0100001110000100"; -- -0.04078271891993334
	pesos_i(25248) := b"1111111111111111_1111111111111111_1110010010011011_0010011101011110"; -- -0.10700754123606857
	pesos_i(25249) := b"0000000000000000_0000000000000000_0010000100111101_0111000010000000"; -- 0.12984374158528264
	pesos_i(25250) := b"1111111111111111_1111111111111111_1110011011101100_0011101100111111"; -- -0.09795789453398178
	pesos_i(25251) := b"1111111111111111_1111111111111111_1110101101101000_0000001110000100"; -- -0.08044412627431982
	pesos_i(25252) := b"1111111111111111_1111111111111111_1111111100010010_1011100100100100"; -- -0.0036205565441247865
	pesos_i(25253) := b"0000000000000000_0000000000000000_0001111000100111_0011110101010110"; -- 0.11778624866706087
	pesos_i(25254) := b"1111111111111111_1111111111111111_1111011000110010_1111011010001001"; -- -0.03828486583290944
	pesos_i(25255) := b"1111111111111111_1111111111111111_1101110001101000_0101000000100101"; -- -0.13903330894989244
	pesos_i(25256) := b"1111111111111111_1111111111111111_1101110011001111_1000001000000011"; -- -0.1374586813959994
	pesos_i(25257) := b"0000000000000000_0000000000000000_0001000000000011_1000001010110010"; -- 0.06255356642999262
	pesos_i(25258) := b"0000000000000000_0000000000000000_0001001011011101_1100100000101000"; -- 0.07369662263181888
	pesos_i(25259) := b"1111111111111111_1111111111111111_1110011101000001_0110011000101000"; -- -0.09665833979203199
	pesos_i(25260) := b"0000000000000000_0000000000000000_0000010101011000_0011010101011010"; -- 0.020877203470330567
	pesos_i(25261) := b"0000000000000000_0000000000000000_0000010010010111_1001010000010110"; -- 0.017937903653946482
	pesos_i(25262) := b"1111111111111111_1111111111111111_1111001001000010_0011100110010011"; -- -0.05367698817639524
	pesos_i(25263) := b"1111111111111111_1111111111111111_1111001011001000_1101011111011101"; -- -0.05162287581672719
	pesos_i(25264) := b"0000000000000000_0000000000000000_0000011111000110_1010100001001110"; -- 0.03037502194604423
	pesos_i(25265) := b"1111111111111111_1111111111111111_1110011010101100_1110101110010101"; -- -0.09892394644644402
	pesos_i(25266) := b"1111111111111111_1111111111111111_1101011110001000_0110110011001111"; -- -0.15807456923547356
	pesos_i(25267) := b"0000000000000000_0000000000000000_0000000011111001_0010001011110001"; -- 0.0038015212202957257
	pesos_i(25268) := b"1111111111111111_1111111111111111_1110001101100011_1111111010010111"; -- -0.11175545505044543
	pesos_i(25269) := b"0000000000000000_0000000000000000_0001010010100111_0010011101010011"; -- 0.08067556168972226
	pesos_i(25270) := b"1111111111111111_1111111111111111_1110100110111010_1000111101010011"; -- -0.0869970723726729
	pesos_i(25271) := b"0000000000000000_0000000000000000_0010010110011111_0101010101111110"; -- 0.14696249321764418
	pesos_i(25272) := b"0000000000000000_0000000000000000_0001100010001100_1100110001000001"; -- 0.09589840487517456
	pesos_i(25273) := b"1111111111111111_1111111111111111_1101110100100110_0101110000101010"; -- -0.1361334225550954
	pesos_i(25274) := b"1111111111111111_1111111111111111_1111111010110011_1000011111110010"; -- -0.005073073869300655
	pesos_i(25275) := b"0000000000000000_0000000000000000_0001011011101101_0011101011011100"; -- 0.08955734123038642
	pesos_i(25276) := b"1111111111111111_1111111111111111_1101001111011011_1111011110010011"; -- -0.1724248186317637
	pesos_i(25277) := b"0000000000000000_0000000000000000_0000000001100101_1000100001001000"; -- 0.0015492605906281536
	pesos_i(25278) := b"0000000000000000_0000000000000000_0000100010011111_0011001010100001"; -- 0.03367916513483672
	pesos_i(25279) := b"1111111111111111_1111111111111111_1101001011110001_1101001010101001"; -- -0.17599757557123732
	pesos_i(25280) := b"1111111111111111_1111111111111111_1101101101110010_0011100011011011"; -- -0.1427883591685529
	pesos_i(25281) := b"1111111111111111_1111111111111111_1101010111100110_1011011100110111"; -- -0.16444830814562383
	pesos_i(25282) := b"1111111111111111_1111111111111111_1110011001101111_0110010001110011"; -- -0.0998627871052333
	pesos_i(25283) := b"0000000000000000_0000000000000000_0010111000110010_0010011001100001"; -- 0.1804527269196661
	pesos_i(25284) := b"0000000000000000_0000000000000000_0010111000100010_0101001100111100"; -- 0.1802112600961637
	pesos_i(25285) := b"0000000000000000_0000000000000000_0010100100110101_0100011001101111"; -- 0.16096916397462277
	pesos_i(25286) := b"0000000000000000_0000000000000000_0000101101011011_0111010111101101"; -- 0.04436432884275381
	pesos_i(25287) := b"0000000000000000_0000000000000000_0001010100110100_1010011001001011"; -- 0.08283461890556806
	pesos_i(25288) := b"0000000000000000_0000000000000000_0000000100100011_0101110111101011"; -- 0.004445905477971886
	pesos_i(25289) := b"0000000000000000_0000000000000000_0000011001001111_1111001010000011"; -- 0.024657399109123602
	pesos_i(25290) := b"0000000000000000_0000000000000000_0010101110011010_0100100011111001"; -- 0.17032295296532915
	pesos_i(25291) := b"0000000000000000_0000000000000000_0010100000110010_0011010111111010"; -- 0.15701615675479277
	pesos_i(25292) := b"0000000000000000_0000000000000000_0001001011111110_0011000011011001"; -- 0.07419114406877624
	pesos_i(25293) := b"0000000000000000_0000000000000000_0001011100101110_0101011010100111"; -- 0.09055081913248016
	pesos_i(25294) := b"0000000000000000_0000000000000000_0011011011001011_0111111100000010"; -- 0.2140426044904447
	pesos_i(25295) := b"0000000000000000_0000000000000000_0010101000011110_1011111010111110"; -- 0.164531632888009
	pesos_i(25296) := b"0000000000000000_0000000000000000_0001001100100110_1011001111101110"; -- 0.0748093086379275
	pesos_i(25297) := b"1111111111111111_1111111111111111_1101010101001100_0101000000001111"; -- -0.1668043102509256
	pesos_i(25298) := b"1111111111111111_1111111111111111_1111101110000001_0100111101011010"; -- -0.017558136591397915
	pesos_i(25299) := b"1111111111111111_1111111111111111_1110111111001001_0001110110001110"; -- -0.0633374718690114
	pesos_i(25300) := b"1111111111111111_1111111111111111_1111111010011000_0001000011010001"; -- -0.005492161754833638
	pesos_i(25301) := b"0000000000000000_0000000000000000_0001111011111110_0110110000101011"; -- 0.12106967966829935
	pesos_i(25302) := b"0000000000000000_0000000000000000_0001001011111011_1001100100100011"; -- 0.07415158380038464
	pesos_i(25303) := b"0000000000000000_0000000000000000_0010111101000001_0100111001001110"; -- 0.18459023856302786
	pesos_i(25304) := b"0000000000000000_0000000000000000_0000110011110111_1010101001011010"; -- 0.0506540747389466
	pesos_i(25305) := b"1111111111111111_1111111111111111_1110001110001000_0001011100111001"; -- -0.11120467057619168
	pesos_i(25306) := b"0000000000000000_0000000000000000_0010010001100111_1110110100011101"; -- 0.14221078822868205
	pesos_i(25307) := b"1111111111111111_1111111111111111_1101101111111101_1111110101110110"; -- -0.1406556689587131
	pesos_i(25308) := b"0000000000000000_0000000000000000_0010000011001001_1001111101000110"; -- 0.12807651001457165
	pesos_i(25309) := b"0000000000000000_0000000000000000_0001111010111111_1101110110001010"; -- 0.12011513351625365
	pesos_i(25310) := b"0000000000000000_0000000000000000_0000010110100011_0101000111000000"; -- 0.022023305186490323
	pesos_i(25311) := b"1111111111111111_1111111111111111_1111111110001111_1001010110111100"; -- -0.0017153183483613612
	pesos_i(25312) := b"1111111111111111_1111111111111111_1101111101010000_1101110011010100"; -- -0.1276723845536904
	pesos_i(25313) := b"0000000000000000_0000000000000000_0001110100101110_1101101110001111"; -- 0.11399624097520203
	pesos_i(25314) := b"0000000000000000_0000000000000000_0010001011011101_1011001010100001"; -- 0.13619533939448986
	pesos_i(25315) := b"0000000000000000_0000000000000000_0000001111010011_0010001011101011"; -- 0.014940435840827507
	pesos_i(25316) := b"0000000000000000_0000000000000000_0001001010110011_1010100100010011"; -- 0.07305390078453514
	pesos_i(25317) := b"1111111111111111_1111111111111111_1100110110010101_0111101000001000"; -- -0.1969379167691498
	pesos_i(25318) := b"1111111111111111_1111111111111111_1110110010001001_1010101010101011"; -- -0.07602437318528715
	pesos_i(25319) := b"0000000000000000_0000000000000000_0010000010110000_1100010101001101"; -- 0.127697307027743
	pesos_i(25320) := b"0000000000000000_0000000000000000_0000110011111110_0101110001101000"; -- 0.05075624019890915
	pesos_i(25321) := b"0000000000000000_0000000000000000_0001011011110000_1111111000010001"; -- 0.08961475302250947
	pesos_i(25322) := b"1111111111111111_1111111111111111_1101011101010011_1001101111111010"; -- -0.15888047358135654
	pesos_i(25323) := b"1111111111111111_1111111111111111_1110110111011111_0100110100010101"; -- -0.07081144569424637
	pesos_i(25324) := b"1111111111111111_1111111111111111_1101010011100011_1011011101000101"; -- -0.16840033105975963
	pesos_i(25325) := b"0000000000000000_0000000000000000_0001110000000100_0100101001110000"; -- 0.10944047193183079
	pesos_i(25326) := b"1111111111111111_1111111111111111_1110100010110111_0001100110111010"; -- -0.09095610813135568
	pesos_i(25327) := b"0000000000000000_0000000000000000_0001011101000000_0010100110001010"; -- 0.09082278850920714
	pesos_i(25328) := b"0000000000000000_0000000000000000_0011001011100101_1000010001100011"; -- 0.19881465349161015
	pesos_i(25329) := b"1111111111111111_1111111111111111_1101010001110010_0110001001101001"; -- -0.17012963224717698
	pesos_i(25330) := b"0000000000000000_0000000000000000_0001111001111110_1101111101101011"; -- 0.11912342422851158
	pesos_i(25331) := b"0000000000000000_0000000000000000_0000011111000110_0001010100010101"; -- 0.030366246887330167
	pesos_i(25332) := b"1111111111111111_1111111111111111_1101000101101010_1100001100000000"; -- -0.18196469556611847
	pesos_i(25333) := b"1111111111111111_1111111111111111_1111111110010100_1011100011010001"; -- -0.0016369332782573483
	pesos_i(25334) := b"0000000000000000_0000000000000000_0010100101000000_0010011101111101"; -- 0.1611351661126095
	pesos_i(25335) := b"0000000000000000_0000000000000000_0010100101011000_0101010111001101"; -- 0.16150413764729388
	pesos_i(25336) := b"0000000000000000_0000000000000000_0000101000110010_0111010111111110"; -- 0.03983247238693948
	pesos_i(25337) := b"0000000000000000_0000000000000000_0001010001001001_0100101011010110"; -- 0.07924335217442952
	pesos_i(25338) := b"1111111111111111_1111111111111111_1111000001110110_1101100111111000"; -- -0.06068647102775075
	pesos_i(25339) := b"1111111111111111_1111111111111111_1101110000000110_1100010010110111"; -- -0.14052172221714695
	pesos_i(25340) := b"0000000000000000_0000000000000000_0001100001010110_0100001010111110"; -- 0.09506623393108882
	pesos_i(25341) := b"0000000000000000_0000000000000000_0001110110011110_0010100001110001"; -- 0.11569454919616161
	pesos_i(25342) := b"1111111111111111_1111111111111111_1101000100010101_1111011111101110"; -- -0.18325853765360356
	pesos_i(25343) := b"0000000000000000_0000000000000000_0000010011111111_1010010101111111"; -- 0.019525855645352377
	pesos_i(25344) := b"1111111111111111_1111111111111111_1111000001001101_1010000001001000"; -- -0.06131551977925069
	pesos_i(25345) := b"1111111111111111_1111111111111111_1111000010110010_0111110100000110"; -- -0.059776483674841945
	pesos_i(25346) := b"0000000000000000_0000000000000000_0001111100100110_1110110101001100"; -- 0.12168772807255426
	pesos_i(25347) := b"0000000000000000_0000000000000000_0001101110011000_0101101110100010"; -- 0.10779354765941285
	pesos_i(25348) := b"1111111111111111_1111111111111111_1101010100100110_1100011101010110"; -- -0.16737703463395892
	pesos_i(25349) := b"1111111111111111_1111111111111111_1110000101100011_0000011001110101"; -- -0.1195827448998972
	pesos_i(25350) := b"1111111111111111_1111111111111111_1101001010101010_0101100101101101"; -- -0.1770881757304456
	pesos_i(25351) := b"1111111111111111_1111111111111111_1101010011101001_1000010110000110"; -- -0.16831174354692813
	pesos_i(25352) := b"1111111111111111_1111111111111111_1100110011101111_0011100010111001"; -- -0.19947476848928114
	pesos_i(25353) := b"1111111111111111_1111111111111111_1111011010100101_1000011110100011"; -- -0.03653671528674293
	pesos_i(25354) := b"0000000000000000_0000000000000000_0000011101110000_0100111111001001"; -- 0.029057490045503186
	pesos_i(25355) := b"0000000000000000_0000000000000000_0010011111001100_0010000101100100"; -- 0.15545853327452613
	pesos_i(25356) := b"1111111111111111_1111111111111111_1111100101110100_1110111011001000"; -- -0.025559498026032048
	pesos_i(25357) := b"1111111111111111_1111111111111111_1111100010110101_1101100110100011"; -- -0.028475186959659456
	pesos_i(25358) := b"1111111111111111_1111111111111111_1110001110100010_0010101001100011"; -- -0.11080679962436447
	pesos_i(25359) := b"0000000000000000_0000000000000000_0001011010111110_1111100000100101"; -- 0.08885146037438864
	pesos_i(25360) := b"0000000000000000_0000000000000000_0010000111011011_1100110101101001"; -- 0.13226016817103842
	pesos_i(25361) := b"0000000000000000_0000000000000000_0000001010010011_0110101101101001"; -- 0.010061944071665985
	pesos_i(25362) := b"1111111111111111_1111111111111111_1101100001111111_1011000010101000"; -- -0.15430160435450027
	pesos_i(25363) := b"0000000000000000_0000000000000000_0001111011111011_0101111111001110"; -- 0.12102316645838083
	pesos_i(25364) := b"0000000000000000_0000000000000000_0000001011001010_1001110111110011"; -- 0.010904189868966463
	pesos_i(25365) := b"0000000000000000_0000000000000000_0001000110111111_0101110000111100"; -- 0.06932617638714762
	pesos_i(25366) := b"1111111111111111_1111111111111111_1111010011010001_1000011000011110"; -- -0.043677919028978336
	pesos_i(25367) := b"1111111111111111_1111111111111111_1111101001101110_1110010111010111"; -- -0.021745333586858845
	pesos_i(25368) := b"0000000000000000_0000000000000000_0000100111100101_1100011101001110"; -- 0.03866239223033087
	pesos_i(25369) := b"1111111111111111_1111111111111111_1101011101110110_0001110110100110"; -- -0.15835394559460644
	pesos_i(25370) := b"1111111111111111_1111111111111111_1110100011111001_1010110101111100"; -- -0.08994022113182913
	pesos_i(25371) := b"0000000000000000_0000000000000000_0010000001101000_1111001010001110"; -- 0.12660137139349664
	pesos_i(25372) := b"0000000000000000_0000000000000000_0001001001111110_0111001010111001"; -- 0.07224194553820965
	pesos_i(25373) := b"1111111111111111_1111111111111111_1101010011010111_1001101001110110"; -- -0.16858515385326256
	pesos_i(25374) := b"0000000000000000_0000000000000000_0001010010101100_1101110010001011"; -- 0.0807626571898736
	pesos_i(25375) := b"0000000000000000_0000000000000000_0000010010011100_0001111000011000"; -- 0.01800716483422227
	pesos_i(25376) := b"1111111111111111_1111111111111111_1101001010000000_0011111110111001"; -- -0.17773057689244914
	pesos_i(25377) := b"0000000000000000_0000000000000000_0000000111101011_0010110001011000"; -- 0.007494708592377812
	pesos_i(25378) := b"1111111111111111_1111111111111111_1111010010100111_1111111110110000"; -- -0.04431154199706433
	pesos_i(25379) := b"0000000000000000_0000000000000000_0010000011110001_0100101011001110"; -- 0.12868182690317434
	pesos_i(25380) := b"0000000000000000_0000000000000000_0001110111000100_0001010110010010"; -- 0.1162732584278949
	pesos_i(25381) := b"1111111111111111_1111111111111111_1111110110011001_0011011001001111"; -- -0.00938091825402239
	pesos_i(25382) := b"1111111111111111_1111111111111111_1110011100101001_0010111010000001"; -- -0.09702786779320369
	pesos_i(25383) := b"0000000000000000_0000000000000000_0001110011101001_1010011110100011"; -- 0.11294028973538885
	pesos_i(25384) := b"1111111111111111_1111111111111111_1101101111111011_0010101100100100"; -- -0.14069872251870422
	pesos_i(25385) := b"1111111111111111_1111111111111111_1110110000010111_0010000010110111"; -- -0.07777209781234344
	pesos_i(25386) := b"1111111111111111_1111111111111111_1110101000010101_1010011101110110"; -- -0.08560708405399702
	pesos_i(25387) := b"1111111111111111_1111111111111111_1111000000000101_1010010010111010"; -- -0.06241388752579891
	pesos_i(25388) := b"1111111111111111_1111111111111111_1101010111100110_1011100100110010"; -- -0.16444818997788335
	pesos_i(25389) := b"1111111111111111_1111111111111111_1110001101100110_0000010001101011"; -- -0.11172459020051441
	pesos_i(25390) := b"1111111111111111_1111111111111111_1101111110111010_1101010001111011"; -- -0.12605545042689417
	pesos_i(25391) := b"0000000000000000_0000000000000000_0010000010111010_0100011011001111"; -- 0.12784235528633936
	pesos_i(25392) := b"1111111111111111_1111111111111111_1101001100011011_1010100110111010"; -- -0.17535914611844855
	pesos_i(25393) := b"1111111111111111_1111111111111111_1101011011000101_1110010101110111"; -- -0.16104284143064276
	pesos_i(25394) := b"0000000000000000_0000000000000000_0010000100001010_0001011110010001"; -- 0.12906024257498558
	pesos_i(25395) := b"1111111111111111_1111111111111111_1101010001101001_0101100111111101"; -- -0.17026746343621377
	pesos_i(25396) := b"0000000000000000_0000000000000000_0010010010010011_1000001010000011"; -- 0.14287582105056326
	pesos_i(25397) := b"1111111111111111_1111111111111111_1101111001000111_1011001100000100"; -- -0.13171845575726981
	pesos_i(25398) := b"0000000000000000_0000000000000000_0000011011111010_1110110011100111"; -- 0.027266317727472487
	pesos_i(25399) := b"1111111111111111_1111111111111111_1110010001010111_0010000000010110"; -- -0.10804557296011787
	pesos_i(25400) := b"1111111111111111_1111111111111111_1100110111100111_1000011101101100"; -- -0.19568589784471807
	pesos_i(25401) := b"0000000000000000_0000000000000000_0010100011010111_0111011010010011"; -- 0.15953770720249333
	pesos_i(25402) := b"1111111111111111_1111111111111111_1101010100100001_1010110000010100"; -- -0.16745495325247892
	pesos_i(25403) := b"1111111111111111_1111111111111111_1101011110110001_1011000111000110"; -- -0.15744484816636897
	pesos_i(25404) := b"0000000000000000_0000000000000000_0000100011111010_1001111111011100"; -- 0.03507422559184939
	pesos_i(25405) := b"1111111111111111_1111111111111111_1111100000110101_1001101001010111"; -- -0.03043208487435876
	pesos_i(25406) := b"1111111111111111_1111111111111111_1111110001011101_0101000111001011"; -- -0.0142010572750281
	pesos_i(25407) := b"1111111111111111_1111111111111111_1111000000101000_1100111111100010"; -- -0.06187725760539911
	pesos_i(25408) := b"0000000000000000_0000000000000000_0000101000010110_0110101010010101"; -- 0.039404546041387996
	pesos_i(25409) := b"1111111111111111_1111111111111111_1111010001011111_0111111101111001"; -- -0.045417817045269
	pesos_i(25410) := b"0000000000000000_0000000000000000_0000110010101110_1110001000011010"; -- 0.0495435059983336
	pesos_i(25411) := b"0000000000000000_0000000000000000_0010100000111100_0010011110110001"; -- 0.157167893081648
	pesos_i(25412) := b"1111111111111111_1111111111111111_1111001010100100_0111010011011001"; -- -0.0521780940113727
	pesos_i(25413) := b"0000000000000000_0000000000000000_0000110110010001_1110110011101100"; -- 0.05300789598120194
	pesos_i(25414) := b"0000000000000000_0000000000000000_0001111100001100_0110001101110110"; -- 0.12128278373588909
	pesos_i(25415) := b"1111111111111111_1111111111111111_1101011010110010_0001101001111111"; -- -0.16134485620960826
	pesos_i(25416) := b"1111111111111111_1111111111111111_1110010011010111_1001111010010100"; -- -0.10608490846657108
	pesos_i(25417) := b"0000000000000000_0000000000000000_0001010110001101_0001110000001111"; -- 0.0841844117191823
	pesos_i(25418) := b"1111111111111111_1111111111111111_1101101111100010_1100001110111111"; -- -0.1410710963017408
	pesos_i(25419) := b"1111111111111111_1111111111111111_1101100011101000_0011111001111110"; -- -0.15270623616076262
	pesos_i(25420) := b"1111111111111111_1111111111111111_1100101110101000_1011011100001110"; -- -0.20445686262631085
	pesos_i(25421) := b"0000000000000000_0000000000000000_0000010001011000_0000000011010101"; -- 0.016967823019923146
	pesos_i(25422) := b"1111111111111111_1111111111111111_1111000110001101_0001000100001110"; -- -0.05644124409590297
	pesos_i(25423) := b"0000000000000000_0000000000000000_0000100111001010_1110001100100011"; -- 0.038252063788023684
	pesos_i(25424) := b"0000000000000000_0000000000000000_0000001100000010_1111100101101111"; -- 0.011764134910018695
	pesos_i(25425) := b"0000000000000000_0000000000000000_0001010111101010_1111101110110010"; -- 0.08561680889586164
	pesos_i(25426) := b"0000000000000000_0000000000000000_0000100000001111_0101000111101111"; -- 0.031483765490178096
	pesos_i(25427) := b"1111111111111111_1111111111111111_1100111100010101_1110001101010001"; -- -0.19107226638493882
	pesos_i(25428) := b"1111111111111111_1111111111111111_1111100001001011_0101010111110100"; -- -0.03010046759351635
	pesos_i(25429) := b"1111111111111111_1111111111111111_1111110001011111_0110010011000010"; -- -0.014169409516022606
	pesos_i(25430) := b"0000000000000000_0000000000000000_0010101010010001_1011100100111001"; -- 0.16628606464372322
	pesos_i(25431) := b"1111111111111111_1111111111111111_1111110001000000_1101011110000011"; -- -0.014635591918023343
	pesos_i(25432) := b"1111111111111111_1111111111111111_1111110010101001_1110111000110001"; -- -0.013032067303145123
	pesos_i(25433) := b"1111111111111111_1111111111111111_1110001100101000_1001100110110010"; -- -0.11266173743181442
	pesos_i(25434) := b"1111111111111111_1111111111111111_1110101011011100_0000000001001011"; -- -0.08258054886807346
	pesos_i(25435) := b"1111111111111111_1111111111111111_1110111000000010_0111000011001000"; -- -0.07027526019050918
	pesos_i(25436) := b"1111111111111111_1111111111111111_1110011011100010_0011101011101011"; -- -0.09811050180507411
	pesos_i(25437) := b"1111111111111111_1111111111111111_1101000010001001_1011101110111001"; -- -0.1853983568392694
	pesos_i(25438) := b"0000000000000000_0000000000000000_0000011100011100_1101011101101110"; -- 0.027783836755554358
	pesos_i(25439) := b"0000000000000000_0000000000000000_0000100010101010_1101100000001100"; -- 0.033856871615157325
	pesos_i(25440) := b"1111111111111111_1111111111111111_1111000111011111_0101101011101011"; -- -0.05518562093731261
	pesos_i(25441) := b"0000000000000000_0000000000000000_0000110101100110_0000011001000100"; -- 0.05233802004624778
	pesos_i(25442) := b"1111111111111111_1111111111111111_1111010010011100_0011110011111110"; -- -0.044490993392802526
	pesos_i(25443) := b"1111111111111111_1111111111111111_1111011000010011_0001100110010100"; -- -0.03877105836770012
	pesos_i(25444) := b"1111111111111111_1111111111111111_1101000001110001_0000000011101011"; -- -0.18577570214186245
	pesos_i(25445) := b"1111111111111111_1111111111111111_1110001011111100_1111111000110100"; -- -0.11332713343588074
	pesos_i(25446) := b"1111111111111111_1111111111111111_1101000110100110_0101000110100010"; -- -0.18105592522057565
	pesos_i(25447) := b"0000000000000000_0000000000000000_0010101011101010_1100000010010011"; -- 0.16764453502854818
	pesos_i(25448) := b"1111111111111111_1111111111111111_1111011110111111_0001110101100101"; -- -0.032240069289118864
	pesos_i(25449) := b"0000000000000000_0000000000000000_0010001011000101_1000000001011000"; -- 0.13582613131777002
	pesos_i(25450) := b"1111111111111111_1111111111111111_1111111110010100_0101111111010000"; -- -0.0016422384438015572
	pesos_i(25451) := b"0000000000000000_0000000000000000_0010110011100000_1100100000001011"; -- 0.17530489235555347
	pesos_i(25452) := b"1111111111111111_1111111111111111_1100111100110011_0000011010110111"; -- -0.19062765144343496
	pesos_i(25453) := b"1111111111111111_1111111111111111_1101001010010001_1101100000101000"; -- -0.1774620916360202
	pesos_i(25454) := b"0000000000000000_0000000000000000_0010001001000010_0000000101010101"; -- 0.13381965936133752
	pesos_i(25455) := b"1111111111111111_1111111111111111_1111011111011010_1110101011010111"; -- -0.031815836482488626
	pesos_i(25456) := b"1111111111111111_1111111111111111_1111001011101101_0100000011111111"; -- -0.05106729282600311
	pesos_i(25457) := b"1111111111111111_1111111111111111_1110000111101110_0100011000100010"; -- -0.11745797784852954
	pesos_i(25458) := b"0000000000000000_0000000000000000_0010111011101101_1110010001111101"; -- 0.18331745189973453
	pesos_i(25459) := b"0000000000000000_0000000000000000_0010011001011010_1010011001100011"; -- 0.14982070836531514
	pesos_i(25460) := b"0000000000000000_0000000000000000_0010100100000001_1010110100100011"; -- 0.16018182846566095
	pesos_i(25461) := b"1111111111111111_1111111111111111_1111000001101001_0100111011001001"; -- -0.06089313117369017
	pesos_i(25462) := b"1111111111111111_1111111111111111_1110000111010111_0110100111001111"; -- -0.11780680362855853
	pesos_i(25463) := b"1111111111111111_1111111111111111_1110110110001111_1010000101011000"; -- -0.07202712635747262
	pesos_i(25464) := b"0000000000000000_0000000000000000_0001010011100011_0110110110111110"; -- 0.08159528628041457
	pesos_i(25465) := b"0000000000000000_0000000000000000_0010001101101100_1000000100101010"; -- 0.13837439809693053
	pesos_i(25466) := b"0000000000000000_0000000000000000_0000011001010010_0010000110101000"; -- 0.024690726799530535
	pesos_i(25467) := b"1111111111111111_1111111111111111_1110001111101111_0001101010110001"; -- -0.10963280842577132
	pesos_i(25468) := b"0000000000000000_0000000000000000_0011000111011110_0010100101100110"; -- 0.19479616861176116
	pesos_i(25469) := b"0000000000000000_0000000000000000_0001101101010010_0110100111000010"; -- 0.10672627438723838
	pesos_i(25470) := b"0000000000000000_0000000000000000_0010011011011000_0011101000000101"; -- 0.15173685664465575
	pesos_i(25471) := b"1111111111111111_1111111111111111_1111010100000101_0111111101011001"; -- -0.04288486559827768
	pesos_i(25472) := b"1111111111111111_1111111111111111_1111001000001111_0010100010101000"; -- -0.054456194938660635
	pesos_i(25473) := b"1111111111111111_1111111111111111_1111011101001100_1000001010110110"; -- -0.03398879094696768
	pesos_i(25474) := b"0000000000000000_0000000000000000_0001000100111010_1010000010101101"; -- 0.067300836882869
	pesos_i(25475) := b"1111111111111111_1111111111111111_1111001010111110_1000110110000111"; -- -0.05177989444155719
	pesos_i(25476) := b"0000000000000000_0000000000000000_0010100000100110_0000011000111111"; -- 0.1568302062106541
	pesos_i(25477) := b"1111111111111111_1111111111111111_1111010011111000_0000000010010100"; -- -0.04309078576598729
	pesos_i(25478) := b"1111111111111111_1111111111111111_1111111111001000_1101011000001111"; -- -0.0008417331914205119
	pesos_i(25479) := b"0000000000000000_0000000000000000_0000001101111101_1011000000111010"; -- 0.013636602670176084
	pesos_i(25480) := b"0000000000000000_0000000000000000_0000100010101010_1110011110101001"; -- 0.03385780224844478
	pesos_i(25481) := b"1111111111111111_1111111111111111_1101100111000000_0100001111010000"; -- -0.14941002053236968
	pesos_i(25482) := b"0000000000000000_0000000000000000_0010101110001001_0111000011000100"; -- 0.17006592556151282
	pesos_i(25483) := b"0000000000000000_0000000000000000_0000010101110110_0111111000000001"; -- 0.02133929762026265
	pesos_i(25484) := b"0000000000000000_0000000000000000_0011000001100001_0111001101001100"; -- 0.18898697485826993
	pesos_i(25485) := b"1111111111111111_1111111111111111_1111111101111110_0101011100011100"; -- -0.001978450413147884
	pesos_i(25486) := b"0000000000000000_0000000000000000_0010100110010110_1100111111010000"; -- 0.16245745489920752
	pesos_i(25487) := b"0000000000000000_0000000000000000_0001111101011110_1011111111110010"; -- 0.1225395170360307
	pesos_i(25488) := b"1111111111111111_1111111111111111_1110000001001011_0110110000110111"; -- -0.12384914077218849
	pesos_i(25489) := b"1111111111111111_1111111111111111_1111110101101001_0010110100110011"; -- -0.010113883150520652
	pesos_i(25490) := b"1111111111111111_1111111111111111_1110010101001110_1111010010000111"; -- -0.10426398943827332
	pesos_i(25491) := b"0000000000000000_0000000000000000_0010110101010110_0000000011100101"; -- 0.17709355914973468
	pesos_i(25492) := b"0000000000000000_0000000000000000_0001010001110010_1110010000100101"; -- 0.07987810050362541
	pesos_i(25493) := b"1111111111111111_1111111111111111_1111111101000010_0111110101011101"; -- -0.002891697640105018
	pesos_i(25494) := b"0000000000000000_0000000000000000_0010011000100111_1011011000011000"; -- 0.14904344648191808
	pesos_i(25495) := b"1111111111111111_1111111111111111_1101101101110010_0111001011010000"; -- -0.14278490463917304
	pesos_i(25496) := b"1111111111111111_1111111111111111_1100101111001111_0111111010101101"; -- -0.2038651301690852
	pesos_i(25497) := b"1111111111111111_1111111111111111_1111101000011010_0110110000001110"; -- -0.023034330897713968
	pesos_i(25498) := b"0000000000000000_0000000000000000_0010000101111000_0011010000000011"; -- 0.1307404048175471
	pesos_i(25499) := b"1111111111111111_1111111111111111_1111001001010101_1111000110110111"; -- -0.05337609568891744
	pesos_i(25500) := b"1111111111111111_1111111111111111_1101101101011011_1011010000110111"; -- -0.14313195860213623
	pesos_i(25501) := b"0000000000000000_0000000000000000_0000010100111001_0111101010000100"; -- 0.020408303410064638
	pesos_i(25502) := b"1111111111111111_1111111111111111_1111101000101000_0110001000011100"; -- -0.02282130066930556
	pesos_i(25503) := b"0000000000000000_0000000000000000_0000110011000000_1111110010110010"; -- 0.04981974920423905
	pesos_i(25504) := b"1111111111111111_1111111111111111_1111100100111101_0110100001110111"; -- -0.026406737329895465
	pesos_i(25505) := b"0000000000000000_0000000000000000_0010100111111000_1110010110100111"; -- 0.16395411799285362
	pesos_i(25506) := b"1111111111111111_1111111111111111_1101001111100011_1001010110100101"; -- -0.17230858546200864
	pesos_i(25507) := b"0000000000000000_0000000000000000_0000010101000001_0011011100101000"; -- 0.02052635885852125
	pesos_i(25508) := b"0000000000000000_0000000000000000_0010100100110101_0000110001101111"; -- 0.1609657070302562
	pesos_i(25509) := b"0000000000000000_0000000000000000_0001100010101011_0110100100000111"; -- 0.09636551294780063
	pesos_i(25510) := b"1111111111111111_1111111111111111_1111110000100011_0111001001000100"; -- -0.015084131680570602
	pesos_i(25511) := b"1111111111111111_1111111111111111_1100101010001111_1011010111000110"; -- -0.20874465870762027
	pesos_i(25512) := b"1111111111111111_1111111111111111_1110101011010110_0110010111001101"; -- -0.0826660512337903
	pesos_i(25513) := b"0000000000000000_0000000000000000_0001010011001100_0011000110101111"; -- 0.08124075432917607
	pesos_i(25514) := b"0000000000000000_0000000000000000_0010110101011001_1100001100101011"; -- 0.17715091512797487
	pesos_i(25515) := b"0000000000000000_0000000000000000_0000101011001000_0011101000110011"; -- 0.04211772683306586
	pesos_i(25516) := b"1111111111111111_1111111111111111_1110111000010010_0010110101010111"; -- -0.0700351393084586
	pesos_i(25517) := b"0000000000000000_0000000000000000_0010111000110101_1110000010000011"; -- 0.1805095978107646
	pesos_i(25518) := b"0000000000000000_0000000000000000_0001010101101100_1000100100111000"; -- 0.08368737820859876
	pesos_i(25519) := b"0000000000000000_0000000000000000_0011001010101100_1100101110011111"; -- 0.19794914839847605
	pesos_i(25520) := b"1111111111111111_1111111111111111_1110011011100000_0110010001100100"; -- -0.09813854749943486
	pesos_i(25521) := b"1111111111111111_1111111111111111_1111111100001000_0110001100101101"; -- -0.003778268331698433
	pesos_i(25522) := b"0000000000000000_0000000000000000_0000000000101011_1010010010000100"; -- 0.0006659337242110231
	pesos_i(25523) := b"0000000000000000_0000000000000000_0001010000101010_1111010001000001"; -- 0.07878042779908143
	pesos_i(25524) := b"1111111111111111_1111111111111111_1111001010110011_1111101010111101"; -- -0.05194123159357902
	pesos_i(25525) := b"0000000000000000_0000000000000000_0000110101100111_1011010110010100"; -- 0.05236372819824886
	pesos_i(25526) := b"0000000000000000_0000000000000000_0010110011000000_1100011101111010"; -- 0.174816577132248
	pesos_i(25527) := b"0000000000000000_0000000000000000_0001111100100110_0000101001100111"; -- 0.1216742040085136
	pesos_i(25528) := b"0000000000000000_0000000000000000_0011010001110100_1100010011010101"; -- 0.2049067516064925
	pesos_i(25529) := b"0000000000000000_0000000000000000_0001010010000101_1010011111011010"; -- 0.08016442361771613
	pesos_i(25530) := b"0000000000000000_0000000000000000_0001001001000101_0111111111100110"; -- 0.0713729797279132
	pesos_i(25531) := b"1111111111111111_1111111111111111_1101000111000101_1100100101111011"; -- -0.18057575932867204
	pesos_i(25532) := b"0000000000000000_0000000000000000_0010000110010101_1110111010100001"; -- 0.1311940329719194
	pesos_i(25533) := b"0000000000000000_0000000000000000_0000110001101011_0100101110001111"; -- 0.04851219399620127
	pesos_i(25534) := b"1111111111111111_1111111111111111_1100101110100001_0000100100001000"; -- -0.20457404655371772
	pesos_i(25535) := b"0000000000000000_0000000000000000_0010111001001010_0001110111010100"; -- 0.18081842833245745
	pesos_i(25536) := b"1111111111111111_1111111111111111_1101100001001100_1001010110010010"; -- -0.15508141684991011
	pesos_i(25537) := b"0000000000000000_0000000000000000_0001101001001010_0010101101101100"; -- 0.10269423847049312
	pesos_i(25538) := b"0000000000000000_0000000000000000_0000101000101011_0101111011111001"; -- 0.0397242888273587
	pesos_i(25539) := b"0000000000000000_0000000000000000_0010010111011000_1100011101000001"; -- 0.14783902480902159
	pesos_i(25540) := b"0000000000000000_0000000000000000_0001000101101100_1010010010000010"; -- 0.06806400463714268
	pesos_i(25541) := b"1111111111111111_1111111111111111_1111000100100110_1000100010111011"; -- -0.05800576624182874
	pesos_i(25542) := b"0000000000000000_0000000000000000_0000101111011000_1001001110010111"; -- 0.0462734454688286
	pesos_i(25543) := b"1111111111111111_1111111111111111_1101101100101000_0000101011110011"; -- -0.14392024579405052
	pesos_i(25544) := b"1111111111111111_1111111111111111_1110101010011000_0111010001010100"; -- -0.0836112303875636
	pesos_i(25545) := b"1111111111111111_1111111111111111_1101100000001100_1010001011010011"; -- -0.15605718952441733
	pesos_i(25546) := b"0000000000000000_0000000000000000_0001101100001101_1000111001000001"; -- 0.10567559323968471
	pesos_i(25547) := b"1111111111111111_1111111111111111_1101100000110101_0110101100001001"; -- -0.15543490435545892
	pesos_i(25548) := b"0000000000000000_0000000000000000_0001110111101010_0110000101000111"; -- 0.11685760491061287
	pesos_i(25549) := b"0000000000000000_0000000000000000_0001010110110011_1111000001000011"; -- 0.08477689401089011
	pesos_i(25550) := b"1111111111111111_1111111111111111_1101001010100001_0111110011111000"; -- -0.1772233861832565
	pesos_i(25551) := b"1111111111111111_1111111111111111_1111000011110011_1100100010100000"; -- -0.05878015599927115
	pesos_i(25552) := b"0000000000000000_0000000000000000_0000101111110111_0010110111010100"; -- 0.04674040237463764
	pesos_i(25553) := b"1111111111111111_1111111111111111_1101110011110101_0111000110101101"; -- -0.13687982114876415
	pesos_i(25554) := b"1111111111111111_1111111111111111_1111110000101011_0100101010001110"; -- -0.01496442822476483
	pesos_i(25555) := b"0000000000000000_0000000000000000_0000001110000011_0000001011010000"; -- 0.013717819012860382
	pesos_i(25556) := b"0000000000000000_0000000000000000_0001111101001001_0010100100010011"; -- 0.12221008983283588
	pesos_i(25557) := b"0000000000000000_0000000000000000_0001100001011110_0010000100000001"; -- 0.0951862933206741
	pesos_i(25558) := b"1111111111111111_1111111111111111_1101011110000010_1000000101001100"; -- -0.15816490070000955
	pesos_i(25559) := b"0000000000000000_0000000000000000_0010101010011111_1001011001011000"; -- 0.16649760865619329
	pesos_i(25560) := b"0000000000000000_0000000000000000_0001001011101001_1011101110110001"; -- 0.07387898512440502
	pesos_i(25561) := b"0000000000000000_0000000000000000_0001100000111100_0011011000000010"; -- 0.0946687463884821
	pesos_i(25562) := b"0000000000000000_0000000000000000_0001000100100100_1110111001011111"; -- 0.06696977453229831
	pesos_i(25563) := b"1111111111111111_1111111111111111_1101111101100100_1100010000111111"; -- -0.12736867384664202
	pesos_i(25564) := b"1111111111111111_1111111111111111_1101001000011111_0001001011111001"; -- -0.17921334678523593
	pesos_i(25565) := b"0000000000000000_0000000000000000_0000001011111010_0000100110111111"; -- 0.011627778265524033
	pesos_i(25566) := b"1111111111111111_1111111111111111_1111111011111100_1110010001100010"; -- -0.003953672419022305
	pesos_i(25567) := b"0000000000000000_0000000000000000_0001111010111000_0101111101001011"; -- 0.12000079712514398
	pesos_i(25568) := b"0000000000000000_0000000000000000_0000011110111001_0000001010100101"; -- 0.030166783532063177
	pesos_i(25569) := b"1111111111111111_1111111111111111_1110111111000110_0010101001101000"; -- -0.0633824822661035
	pesos_i(25570) := b"1111111111111111_1111111111111111_1111011000110011_1101000110000111"; -- -0.03827181299881824
	pesos_i(25571) := b"1111111111111111_1111111111111111_1110101011001111_1111110110001100"; -- -0.08276381804911176
	pesos_i(25572) := b"0000000000000000_0000000000000000_0010001010000101_0110000011011001"; -- 0.13484769161840396
	pesos_i(25573) := b"0000000000000000_0000000000000000_0000100011101100_0100010100000100"; -- 0.03485518794526007
	pesos_i(25574) := b"1111111111111111_1111111111111111_1110101111100000_0110010011001011"; -- -0.07860727341630755
	pesos_i(25575) := b"1111111111111111_1111111111111111_1111010110001110_1010011000111110"; -- -0.04079209313422888
	pesos_i(25576) := b"1111111111111111_1111111111111111_1111100010111001_0010001000100110"; -- -0.028425088546907007
	pesos_i(25577) := b"1111111111111111_1111111111111111_1110011011101110_0011101011111101"; -- -0.09792739222714321
	pesos_i(25578) := b"0000000000000000_0000000000000000_0000000000101010_0011100100100101"; -- 0.0006442752222747971
	pesos_i(25579) := b"1111111111111111_1111111111111111_1101110100111011_1000010001110001"; -- -0.13581058736346233
	pesos_i(25580) := b"1111111111111111_1111111111111111_1111000100010010_0000010000101010"; -- -0.05831884360522011
	pesos_i(25581) := b"0000000000000000_0000000000000000_0010000100101001_0110010101000101"; -- 0.12953789652822428
	pesos_i(25582) := b"0000000000000000_0000000000000000_0001110101110101_1100011001111000"; -- 0.11507835806342949
	pesos_i(25583) := b"0000000000000000_0000000000000000_0001110101101010_0111000001010111"; -- 0.1149053775527065
	pesos_i(25584) := b"1111111111111111_1111111111111111_1101111110100011_0111011100101010"; -- -0.12641196476293584
	pesos_i(25585) := b"0000000000000000_0000000000000000_0010111011011001_0100111001010000"; -- 0.1830033250555644
	pesos_i(25586) := b"0000000000000000_0000000000000000_0010111110111011_1101000100110100"; -- 0.18645961292740176
	pesos_i(25587) := b"1111111111111111_1111111111111111_1100110100100100_0100101000011001"; -- -0.1986650170778974
	pesos_i(25588) := b"0000000000000000_0000000000000000_0010100100000100_1111100101100001"; -- 0.16023214923680087
	pesos_i(25589) := b"1111111111111111_1111111111111111_1110100011110001_1000100101011110"; -- -0.0900644441365153
	pesos_i(25590) := b"1111111111111111_1111111111111111_1111100010110001_1000111001001000"; -- -0.028540713804959986
	pesos_i(25591) := b"0000000000000000_0000000000000000_0011000001010010_1111011100101111"; -- 0.18876595397205537
	pesos_i(25592) := b"0000000000000000_0000000000000000_0010100010000110_1011000111001000"; -- 0.1583052744381729
	pesos_i(25593) := b"0000000000000000_0000000000000000_0001000000110111_1110110011000010"; -- 0.06335334528770178
	pesos_i(25594) := b"1111111111111111_1111111111111111_1111010101011001_0000111110000111"; -- -0.04160979228099449
	pesos_i(25595) := b"0000000000000000_0000000000000000_0010011011100111_0110001010110011"; -- 0.15196816327433482
	pesos_i(25596) := b"1111111111111111_1111111111111111_1111101100110010_1001110000010011"; -- -0.018759007875751514
	pesos_i(25597) := b"0000000000000000_0000000000000000_0000001100010111_1001110100011011"; -- 0.012079066271309356
	pesos_i(25598) := b"1111111111111111_1111111111111111_1110000010000000_1111100111100011"; -- -0.1230319806936993
	pesos_i(25599) := b"1111111111111111_1111111111111111_1111110110110011_1010101100100101"; -- -0.00897722571800373
	pesos_i(25600) := b"0000000000000000_0000000000000000_0011000010110000_1111100001010010"; -- 0.1902003480092257
	pesos_i(25601) := b"0000000000000000_0000000000000000_0000110100110000_1001010011111010"; -- 0.05152255166669732
	pesos_i(25602) := b"0000000000000000_0000000000000000_0001110000001001_1100011001000111"; -- 0.10952414736321028
	pesos_i(25603) := b"0000000000000000_0000000000000000_0000110100011011_1010000111000011"; -- 0.05120287912450139
	pesos_i(25604) := b"0000000000000000_0000000000000000_0010000101011010_1000000001110101"; -- 0.13028719756521118
	pesos_i(25605) := b"0000000000000000_0000000000000000_0001000000110110_1010101010111010"; -- 0.06333415071159934
	pesos_i(25606) := b"1111111111111111_1111111111111111_1111010011111100_1110101101000111"; -- -0.043015761644376524
	pesos_i(25607) := b"1111111111111111_1111111111111111_1101111100001110_1011101111000011"; -- -0.12868143543113347
	pesos_i(25608) := b"0000000000000000_0000000000000000_0001001101001111_0101111001111110"; -- 0.07542982641169217
	pesos_i(25609) := b"0000000000000000_0000000000000000_0000001001000111_1111010101010111"; -- 0.008910497365142982
	pesos_i(25610) := b"0000000000000000_0000000000000000_0010110110011110_0110101000001000"; -- 0.17819845862947467
	pesos_i(25611) := b"1111111111111111_1111111111111111_1111000010110101_0000001111011000"; -- -0.05973793018233761
	pesos_i(25612) := b"1111111111111111_1111111111111111_1111111001000001_0001011110101011"; -- -0.006819268052944852
	pesos_i(25613) := b"0000000000000000_0000000000000000_0001110100001100_1100100111100101"; -- 0.11347638922891318
	pesos_i(25614) := b"1111111111111111_1111111111111111_1110101000111000_1101110001101001"; -- -0.08506987034094884
	pesos_i(25615) := b"0000000000000000_0000000000000000_0011000000010000_1110001001101111"; -- 0.18775763700518563
	pesos_i(25616) := b"0000000000000000_0000000000000000_0001011010000011_1101100100111001"; -- 0.08794934889064833
	pesos_i(25617) := b"0000000000000000_0000000000000000_0001010100001000_0001110011101001"; -- 0.08215504356739027
	pesos_i(25618) := b"0000000000000000_0000000000000000_0010101100001011_0001011110010010"; -- 0.16813800163188508
	pesos_i(25619) := b"1111111111111111_1111111111111111_1101001010100110_1011101000001101"; -- -0.1771434515153562
	pesos_i(25620) := b"0000000000000000_0000000000000000_0000111001110010_0111110010111100"; -- 0.056434436660187354
	pesos_i(25621) := b"0000000000000000_0000000000000000_0010100111110111_1100111010011100"; -- 0.1639374858567894
	pesos_i(25622) := b"0000000000000000_0000000000000000_0000011101010101_0001100101101010"; -- 0.028642261910427392
	pesos_i(25623) := b"1111111111111111_1111111111111111_1110000000110010_1101100111011101"; -- -0.12422407486910901
	pesos_i(25624) := b"0000000000000000_0000000000000000_0001010001110100_1100011000000100"; -- 0.07990682214563918
	pesos_i(25625) := b"0000000000000000_0000000000000000_0001000100100100_1000011101001100"; -- 0.06696363078415592
	pesos_i(25626) := b"0000000000000000_0000000000000000_0000011110001110_1000011111111111"; -- 0.02951860394329227
	pesos_i(25627) := b"1111111111111111_1111111111111111_1111010001011101_1001101010010011"; -- -0.04544671916555025
	pesos_i(25628) := b"1111111111111111_1111111111111111_1100110100000110_1100101011001100"; -- -0.1991151096544606
	pesos_i(25629) := b"0000000000000000_0000000000000000_0010000001110011_1100010010110111"; -- 0.12676648575720342
	pesos_i(25630) := b"1111111111111111_1111111111111111_1110111000000011_0000000101001000"; -- -0.07026664733245533
	pesos_i(25631) := b"1111111111111111_1111111111111111_1101001101010000_1010101000010001"; -- -0.17455041002383573
	pesos_i(25632) := b"0000000000000000_0000000000000000_0001001101111000_1111101111110111"; -- 0.0760648228713086
	pesos_i(25633) := b"1111111111111111_1111111111111111_1110001000010111_1111110011100111"; -- -0.11682147373422597
	pesos_i(25634) := b"1111111111111111_1111111111111111_1111101010001110_0110010100101011"; -- -0.021264721985494336
	pesos_i(25635) := b"1111111111111111_1111111111111111_1110100000000111_0111011000001100"; -- -0.09363615223359324
	pesos_i(25636) := b"1111111111111111_1111111111111111_1110101110000111_1011011101011110"; -- -0.07996038395441621
	pesos_i(25637) := b"0000000000000000_0000000000000000_0001001101110000_1101111010011010"; -- 0.07594100243420081
	pesos_i(25638) := b"1111111111111111_1111111111111111_1101100001010000_0000100001001010"; -- -0.155028802884143
	pesos_i(25639) := b"1111111111111111_1111111111111111_1110010101010100_0110011100000111"; -- -0.10418087089110224
	pesos_i(25640) := b"0000000000000000_0000000000000000_0000011101000010_0001000000000110"; -- 0.028351785115094886
	pesos_i(25641) := b"0000000000000000_0000000000000000_0001000000101011_0001000010110100"; -- 0.06315712345953825
	pesos_i(25642) := b"1111111111111111_1111111111111111_1110011010001100_0100001000011111"; -- -0.09942232847532766
	pesos_i(25643) := b"1111111111111111_1111111111111111_1110011000100101_1011001000011110"; -- -0.10098730813599835
	pesos_i(25644) := b"1111111111111111_1111111111111111_1100111000000000_0111100011011000"; -- -0.19530529714964365
	pesos_i(25645) := b"0000000000000000_0000000000000000_0000011101101000_1010001111000011"; -- 0.02894042495166807
	pesos_i(25646) := b"1111111111111111_1111111111111111_1111101111010101_0011000110000010"; -- -0.016278177066333877
	pesos_i(25647) := b"0000000000000000_0000000000000000_0001100110011110_1011000111010100"; -- 0.10007773809659248
	pesos_i(25648) := b"1111111111111111_1111111111111111_1101101011000111_1010100000010001"; -- -0.1453909833900256
	pesos_i(25649) := b"1111111111111111_1111111111111111_1111101110001100_0101001001001001"; -- -0.017390115034828943
	pesos_i(25650) := b"1111111111111111_1111111111111111_1101100101010110_1101100010001110"; -- -0.151018586462837
	pesos_i(25651) := b"0000000000000000_0000000000000000_0001100111001011_0000100111000001"; -- 0.10075436557548768
	pesos_i(25652) := b"0000000000000000_0000000000000000_0000010110000101_0000010011101000"; -- 0.021560961323645336
	pesos_i(25653) := b"1111111111111111_1111111111111111_1110010000010010_1011101101011010"; -- -0.109089174751911
	pesos_i(25654) := b"1111111111111111_1111111111111111_1110111010100101_1111110001010001"; -- -0.0677797605900122
	pesos_i(25655) := b"0000000000000000_0000000000000000_0000100000101111_0010111100010010"; -- 0.03196996864016078
	pesos_i(25656) := b"0000000000000000_0000000000000000_0000011011010101_1111111111111010"; -- 0.026702879515089938
	pesos_i(25657) := b"1111111111111111_1111111111111111_1110110111001101_0001111011110110"; -- -0.07108885278749211
	pesos_i(25658) := b"0000000000000000_0000000000000000_0000101101011011_1001101110011011"; -- 0.044366574696994315
	pesos_i(25659) := b"0000000000000000_0000000000000000_0010001000101101_1010001110010101"; -- 0.13350889581074887
	pesos_i(25660) := b"1111111111111111_1111111111111111_1111001101011001_1111010100010011"; -- -0.049408610133806964
	pesos_i(25661) := b"0000000000000000_0000000000000000_0010111111100101_0101000010101111"; -- 0.18709282170695088
	pesos_i(25662) := b"1111111111111111_1111111111111111_1111001000001001_1011001111000001"; -- -0.0545394567044499
	pesos_i(25663) := b"0000000000000000_0000000000000000_0011000110011100_0001111001100011"; -- 0.19378843235375587
	pesos_i(25664) := b"0000000000000000_0000000000000000_0010011110011010_0101000000010101"; -- 0.1546983768152166
	pesos_i(25665) := b"1111111111111111_1111111111111111_1111001010010010_1111000000100100"; -- -0.05244540325027749
	pesos_i(25666) := b"0000000000000000_0000000000000000_0010011101110110_0001010111101111"; -- 0.1541455944947944
	pesos_i(25667) := b"1111111111111111_1111111111111111_1110100111101000_1010100100010001"; -- -0.086293633751508
	pesos_i(25668) := b"1111111111111111_1111111111111111_1111111000010100_1000011011100100"; -- -0.007499284152084496
	pesos_i(25669) := b"0000000000000000_0000000000000000_0000000100001110_0001001011100100"; -- 0.004120999075460576
	pesos_i(25670) := b"0000000000000000_0000000000000000_0010010011001010_0000111111011111"; -- 0.14370822136055866
	pesos_i(25671) := b"0000000000000000_0000000000000000_0011000001001110_1101111101011011"; -- 0.18870349855706595
	pesos_i(25672) := b"0000000000000000_0000000000000000_0000000101001111_0001101000100100"; -- 0.005113252409327359
	pesos_i(25673) := b"0000000000000000_0000000000000000_0010111111001111_1100001111111100"; -- 0.18676400090150963
	pesos_i(25674) := b"1111111111111111_1111111111111111_1101010000100110_1101011011110001"; -- -0.17128235455045657
	pesos_i(25675) := b"0000000000000000_0000000000000000_0010001010101110_1111000010111100"; -- 0.13548187811983514
	pesos_i(25676) := b"0000000000000000_0000000000000000_0000010010011111_1100101101111101"; -- 0.018063276366424606
	pesos_i(25677) := b"1111111111111111_1111111111111111_1101011011101111_1011111001101000"; -- -0.16040430038628184
	pesos_i(25678) := b"0000000000000000_0000000000000000_0001110011010011_1100100011101000"; -- 0.11260657934050071
	pesos_i(25679) := b"0000000000000000_0000000000000000_0000011111111100_1011010010001110"; -- 0.031199726844140123
	pesos_i(25680) := b"0000000000000000_0000000000000000_0000001111110110_1111111100101101"; -- 0.015487621701055023
	pesos_i(25681) := b"1111111111111111_1111111111111111_1100111111010101_0010111101011011"; -- -0.18815330521380813
	pesos_i(25682) := b"0000000000000000_0000000000000000_0001010000110110_0010001011011110"; -- 0.07895105280349571
	pesos_i(25683) := b"0000000000000000_0000000000000000_0000011001011011_0010110010001011"; -- 0.02482870470364122
	pesos_i(25684) := b"1111111111111111_1111111111111111_1101111000111010_0111101011001001"; -- -0.13192017176214416
	pesos_i(25685) := b"1111111111111111_1111111111111111_1111010101101001_1110010001101101"; -- -0.04135296201363954
	pesos_i(25686) := b"1111111111111111_1111111111111111_1111011111000100_1000110110110110"; -- -0.03215708060770982
	pesos_i(25687) := b"0000000000000000_0000000000000000_0000001001010111_1000110000010101"; -- 0.00914836417468843
	pesos_i(25688) := b"1111111111111111_1111111111111111_1110010000001111_1000101000110011"; -- -0.10913788075102668
	pesos_i(25689) := b"1111111111111111_1111111111111111_1111011011001111_1100100011011100"; -- -0.0358919585222567
	pesos_i(25690) := b"0000000000000000_0000000000000000_0010000001101011_1000110100111011"; -- 0.1266411083314096
	pesos_i(25691) := b"0000000000000000_0000000000000000_0000011100010000_0100111111000100"; -- 0.02759264512021267
	pesos_i(25692) := b"0000000000000000_0000000000000000_0000100100011011_1010000010011010"; -- 0.03557781000104336
	pesos_i(25693) := b"0000000000000000_0000000000000000_0011011001010011_0001101011011011"; -- 0.21220558022065034
	pesos_i(25694) := b"0000000000000000_0000000000000000_0001000010001000_1010001000011111"; -- 0.06458485844402048
	pesos_i(25695) := b"0000000000000000_0000000000000000_0001111001111100_0011101111001010"; -- 0.1190831534350647
	pesos_i(25696) := b"1111111111111111_1111111111111111_1101101111100001_0011111001011011"; -- -0.14109430588174904
	pesos_i(25697) := b"1111111111111111_1111111111111111_1110010000101110_0010101001100111"; -- -0.10867056837023405
	pesos_i(25698) := b"0000000000000000_0000000000000000_0010010101111000_1101011011000110"; -- 0.14637510609472063
	pesos_i(25699) := b"0000000000000000_0000000000000000_0011000111110000_0000000111000000"; -- 0.19506846372882056
	pesos_i(25700) := b"0000000000000000_0000000000000000_0000010100010001_1011111101100010"; -- 0.019802056789096075
	pesos_i(25701) := b"0000000000000000_0000000000000000_0000000100110100_1111000100100010"; -- 0.004714079609180652
	pesos_i(25702) := b"0000000000000000_0000000000000000_0000001111000110_1100100000000101"; -- 0.01475191237944639
	pesos_i(25703) := b"1111111111111111_1111111111111111_1110101111011000_0101001001111010"; -- -0.07873043552156408
	pesos_i(25704) := b"1111111111111111_1111111111111111_1100110101011010_1001111111101100"; -- -0.19783592691814678
	pesos_i(25705) := b"0000000000000000_0000000000000000_0000011111010100_0100101101001001"; -- 0.030583100533772858
	pesos_i(25706) := b"0000000000000000_0000000000000000_0001100001100101_1101110010010010"; -- 0.09530428472288677
	pesos_i(25707) := b"1111111111111111_1111111111111111_1100110110010101_0000000110110001"; -- -0.19694508956729473
	pesos_i(25708) := b"0000000000000000_0000000000000000_0001001100100001_1110011001100110"; -- 0.0747360227516715
	pesos_i(25709) := b"0000000000000000_0000000000000000_0000001010100100_1001111101001011"; -- 0.01032443598850636
	pesos_i(25710) := b"1111111111111111_1111111111111111_1110100101000001_0101001011100100"; -- -0.08884698797796588
	pesos_i(25711) := b"1111111111111111_1111111111111111_1111110111100000_0001111011000001"; -- -0.008298948289896945
	pesos_i(25712) := b"0000000000000000_0000000000000000_0010111011100100_0001011011011100"; -- 0.18316786653500342
	pesos_i(25713) := b"0000000000000000_0000000000000000_0000011100000011_1011011001011100"; -- 0.027400395752230484
	pesos_i(25714) := b"0000000000000000_0000000000000000_0000100101101001_1111010111000101"; -- 0.03677307187487813
	pesos_i(25715) := b"0000000000000000_0000000000000000_0001110100010101_0001010100011110"; -- 0.11360294331146072
	pesos_i(25716) := b"0000000000000000_0000000000000000_0000000000000100_1001000000110010"; -- 6.962975473387282e-05
	pesos_i(25717) := b"1111111111111111_1111111111111111_1111111010010010_1111001101010001"; -- -0.005570213983359863
	pesos_i(25718) := b"1111111111111111_1111111111111111_1110100010111100_1001110011111111"; -- -0.09087199005088081
	pesos_i(25719) := b"1111111111111111_1111111111111111_1101100001100110_0111000111110110"; -- -0.15468681087307273
	pesos_i(25720) := b"1111111111111111_1111111111111111_1110111100011000_0100100001000100"; -- -0.06603573179273478
	pesos_i(25721) := b"0000000000000000_0000000000000000_0010111010001111_0110001110010011"; -- 0.18187544194662883
	pesos_i(25722) := b"1111111111111111_1111111111111111_1111010000011100_1100011111001110"; -- -0.046435844561348937
	pesos_i(25723) := b"0000000000000000_0000000000000000_0000001110010011_1101001110100001"; -- 0.013974405970908144
	pesos_i(25724) := b"0000000000000000_0000000000000000_0011001110101101_0111111110111010"; -- 0.20186613350414667
	pesos_i(25725) := b"1111111111111111_1111111111111111_1110101101101101_1101011101010101"; -- -0.08035520719516429
	pesos_i(25726) := b"0000000000000000_0000000000000000_0010110001100101_0100010110000110"; -- 0.17342028161211473
	pesos_i(25727) := b"1111111111111111_1111111111111111_1111101011101101_1011010001100110"; -- -0.019810414404403513
	pesos_i(25728) := b"0000000000000000_0000000000000000_0000010111010000_0001011100100100"; -- 0.022706457461564036
	pesos_i(25729) := b"0000000000000000_0000000000000000_0001011100100010_0110010110110110"; -- 0.09036861134276068
	pesos_i(25730) := b"0000000000000000_0000000000000000_0010101001010001_1101001010000101"; -- 0.165311009740836
	pesos_i(25731) := b"0000000000000000_0000000000000000_0001001011111111_1110011110100010"; -- 0.07421729748935982
	pesos_i(25732) := b"0000000000000000_0000000000000000_0001110100010000_1100101001100010"; -- 0.11353745353331177
	pesos_i(25733) := b"1111111111111111_1111111111111111_1111100101110010_1110010010011111"; -- -0.025590621188077606
	pesos_i(25734) := b"1111111111111111_1111111111111111_1111111001111001_0011000011100010"; -- -0.005963272933909682
	pesos_i(25735) := b"1111111111111111_1111111111111111_1111110100010001_0011110110101011"; -- -0.01145567481922739
	pesos_i(25736) := b"1111111111111111_1111111111111111_1111111100101110_0100110010010010"; -- -0.0031997818423674515
	pesos_i(25737) := b"1111111111111111_1111111111111111_1111101000110011_0100011011001101"; -- -0.022655081748891165
	pesos_i(25738) := b"0000000000000000_0000000000000000_0010010101010001_0110110011010101"; -- 0.14577369870257517
	pesos_i(25739) := b"0000000000000000_0000000000000000_0000001100010100_0101011011101100"; -- 0.012029106842594775
	pesos_i(25740) := b"0000000000000000_0000000000000000_0001000110000100_0001101100011010"; -- 0.06842202557325489
	pesos_i(25741) := b"1111111111111111_1111111111111111_1110101100000001_1010101110000000"; -- -0.08200576910405172
	pesos_i(25742) := b"1111111111111111_1111111111111111_1101101011010110_1001110000010010"; -- -0.14516281669560704
	pesos_i(25743) := b"0000000000000000_0000000000000000_0011010001101110_0110011010111110"; -- 0.2048095907829541
	pesos_i(25744) := b"0000000000000000_0000000000000000_0000100011100011_1111111001010110"; -- 0.03472890463139662
	pesos_i(25745) := b"1111111111111111_1111111111111111_1111111110000101_0000111111101100"; -- -0.0018758819310856541
	pesos_i(25746) := b"1111111111111111_1111111111111111_1111101100010011_0100010111010010"; -- -0.019237171321923065
	pesos_i(25747) := b"0000000000000000_0000000000000000_0000101011001001_0111010010100100"; -- 0.04213646901520693
	pesos_i(25748) := b"0000000000000000_0000000000000000_0001001000001101_0011100110111101"; -- 0.07051430575049587
	pesos_i(25749) := b"1111111111111111_1111111111111111_1101011011110010_0111101010001101"; -- -0.1603625684080163
	pesos_i(25750) := b"1111111111111111_1111111111111111_1110111000000100_0110100011111010"; -- -0.07024520782536535
	pesos_i(25751) := b"1111111111111111_1111111111111111_1101100101101101_1001011110001110"; -- -0.1506715086654288
	pesos_i(25752) := b"1111111111111111_1111111111111111_1111110110011101_1101001011001100"; -- -0.009310555646548287
	pesos_i(25753) := b"0000000000000000_0000000000000000_0010001001011110_0000101010001111"; -- 0.13424745540576466
	pesos_i(25754) := b"1111111111111111_1111111111111111_1110101001010001_0010001011000001"; -- -0.08469946656309253
	pesos_i(25755) := b"1111111111111111_1111111111111111_1110111111101011_1001101001000000"; -- -0.06281124045943325
	pesos_i(25756) := b"1111111111111111_1111111111111111_1110000000111010_1111011011001011"; -- -0.12410028031855916
	pesos_i(25757) := b"0000000000000000_0000000000000000_0000100111110110_1011111010010011"; -- 0.0389212713136787
	pesos_i(25758) := b"1111111111111111_1111111111111111_1111111011110001_1111110100110011"; -- -0.004120039945618226
	pesos_i(25759) := b"1111111111111111_1111111111111111_1101101111001011_1001010001010010"; -- -0.14142487524356445
	pesos_i(25760) := b"0000000000000000_0000000000000000_0000001101000111_0100010000010110"; -- 0.012806182155605889
	pesos_i(25761) := b"1111111111111111_1111111111111111_1110010011001011_0010010010101110"; -- -0.10627527964817435
	pesos_i(25762) := b"0000000000000000_0000000000000000_0010000011100110_0010111011100011"; -- 0.12851231617733705
	pesos_i(25763) := b"1111111111111111_1111111111111111_1111100100011011_0010001001110101"; -- -0.02692970883964338
	pesos_i(25764) := b"1111111111111111_1111111111111111_1111110010001010_1101000100100001"; -- -0.013506822063949772
	pesos_i(25765) := b"1111111111111111_1111111111111111_1101101000001110_1110001011010110"; -- -0.1482103564922077
	pesos_i(25766) := b"1111111111111111_1111111111111111_1101111101000000_1011001001010111"; -- -0.12791905762916175
	pesos_i(25767) := b"1111111111111111_1111111111111111_1110000011111110_0010001100111111"; -- -0.12112216674863878
	pesos_i(25768) := b"0000000000000000_0000000000000000_0010000000000110_0010000010100111"; -- 0.1250934990497302
	pesos_i(25769) := b"1111111111111111_1111111111111111_1111001011000110_1011011010000011"; -- -0.051655381232141834
	pesos_i(25770) := b"1111111111111111_1111111111111111_1111101110101010_0001010110111101"; -- -0.016935960168540595
	pesos_i(25771) := b"1111111111111111_1111111111111111_1111111001011011_0111011010110011"; -- -0.006416875228768609
	pesos_i(25772) := b"1111111111111111_1111111111111111_1101100100000100_0001100011000101"; -- -0.15228123852486364
	pesos_i(25773) := b"1111111111111111_1111111111111111_1110101001000001_1010100001110110"; -- -0.08493563759494906
	pesos_i(25774) := b"0000000000000000_0000000000000000_0001010010000100_1100011011011110"; -- 0.08015101361862247
	pesos_i(25775) := b"1111111111111111_1111111111111111_1110010101011101_0001111000111100"; -- -0.10404788056181176
	pesos_i(25776) := b"1111111111111111_1111111111111111_1110100100111100_0011000101110101"; -- -0.08892527484736465
	pesos_i(25777) := b"0000000000000000_0000000000000000_0000011011101000_1010000010000100"; -- 0.02698710643107919
	pesos_i(25778) := b"0000000000000000_0000000000000000_0001001101100010_1001010011110101"; -- 0.0757229898705111
	pesos_i(25779) := b"1111111111111111_1111111111111111_1100111111010001_1111000111100111"; -- -0.18820274460430486
	pesos_i(25780) := b"1111111111111111_1111111111111111_1110101001010000_0100011001110011"; -- -0.0847125978637343
	pesos_i(25781) := b"1111111111111111_1111111111111111_1101001100000001_1010110100010010"; -- -0.1757556754992708
	pesos_i(25782) := b"0000000000000000_0000000000000000_0001011111010001_1111011101111100"; -- 0.0930475881140048
	pesos_i(25783) := b"0000000000000000_0000000000000000_0001000011111110_1010001001001011"; -- 0.0663854057754903
	pesos_i(25784) := b"1111111111111111_1111111111111111_1101101111100111_1111000011101001"; -- -0.1409921103006195
	pesos_i(25785) := b"0000000000000000_0000000000000000_0010011011101010_0010110110100011"; -- 0.15201077682768482
	pesos_i(25786) := b"1111111111111111_1111111111111111_1100111000101110_0010101010111011"; -- -0.19460804865610848
	pesos_i(25787) := b"1111111111111111_1111111111111111_1110010000111010_1010111111001111"; -- -0.10847951133327002
	pesos_i(25788) := b"0000000000000000_0000000000000000_0001010000111101_0111000100101110"; -- 0.07906253209187307
	pesos_i(25789) := b"1111111111111111_1111111111111111_1111111110001011_1000000011101100"; -- -0.0017775940673060888
	pesos_i(25790) := b"1111111111111111_1111111111111111_1111011111000100_0001010110000010"; -- -0.032164245424267913
	pesos_i(25791) := b"0000000000000000_0000000000000000_0010001010100101_1100011000101100"; -- 0.13534201227371523
	pesos_i(25792) := b"1111111111111111_1111111111111111_1110010000101000_1000001111100010"; -- -0.10875678760517514
	pesos_i(25793) := b"1111111111111111_1111111111111111_1111111010000100_0010010111001000"; -- -0.005796087859085729
	pesos_i(25794) := b"1111111111111111_1111111111111111_1111111010101111_1001010100000100"; -- -0.0051333298098369265
	pesos_i(25795) := b"0000000000000000_0000000000000000_0001011000000101_0111101111101100"; -- 0.086021180215525
	pesos_i(25796) := b"0000000000000000_0000000000000000_0001100110110000_0010010000100101"; -- 0.10034395125466904
	pesos_i(25797) := b"0000000000000000_0000000000000000_0001110100001100_0110000001000100"; -- 0.11347009342415194
	pesos_i(25798) := b"0000000000000000_0000000000000000_0000001101011100_1010011001111110"; -- 0.013132482234423015
	pesos_i(25799) := b"0000000000000000_0000000000000000_0000001000011111_0011011011101100"; -- 0.008288796024529995
	pesos_i(25800) := b"0000000000000000_0000000000000000_0001001011100010_0111000011110000"; -- 0.07376771793692057
	pesos_i(25801) := b"1111111111111111_1111111111111111_1110010011000000_1000000101011000"; -- -0.10643760306189999
	pesos_i(25802) := b"0000000000000000_0000000000000000_0000000110101001_1001110010100010"; -- 0.006494321469073733
	pesos_i(25803) := b"0000000000000000_0000000000000000_0010000111100001_1011001110001010"; -- 0.13235017891946008
	pesos_i(25804) := b"0000000000000000_0000000000000000_0001111111100000_1110011010010000"; -- 0.12452546124636685
	pesos_i(25805) := b"1111111111111111_1111111111111111_1100111100000111_1011001001100101"; -- -0.19128880544459947
	pesos_i(25806) := b"1111111111111111_1111111111111111_1101011010001110_1101111100100110"; -- -0.16188245121474004
	pesos_i(25807) := b"0000000000000000_0000000000000000_0010011011000011_0110000010110100"; -- 0.15141872773268716
	pesos_i(25808) := b"1111111111111111_1111111111111111_1111010001001111_1101000011011001"; -- -0.04565710732760757
	pesos_i(25809) := b"0000000000000000_0000000000000000_0010000101100001_1111101101100111"; -- 0.13040133721661987
	pesos_i(25810) := b"1111111111111111_1111111111111111_1101110001011101_1010110000011011"; -- -0.139195674418455
	pesos_i(25811) := b"1111111111111111_1111111111111111_1101010101001101_0010110100001100"; -- -0.16679113825471878
	pesos_i(25812) := b"0000000000000000_0000000000000000_0000001101101000_1110010100001110"; -- 0.013319316735267813
	pesos_i(25813) := b"0000000000000000_0000000000000000_0000000110100001_0000011101001111"; -- 0.006363350563428759
	pesos_i(25814) := b"0000000000000000_0000000000000000_0000111101010101_0111111001000011"; -- 0.05989827280764813
	pesos_i(25815) := b"0000000000000000_0000000000000000_0001010011001011_1001011001000000"; -- 0.08123148985820335
	pesos_i(25816) := b"1111111111111111_1111111111111111_1101000100011100_1000100110010000"; -- -0.18315830445878162
	pesos_i(25817) := b"1111111111111111_1111111111111111_1101111101000001_0010001101011101"; -- -0.12791232090499066
	pesos_i(25818) := b"0000000000000000_0000000000000000_0001001110101101_1001011001100111"; -- 0.07686748528256787
	pesos_i(25819) := b"1111111111111111_1111111111111111_1110101101111001_1011010100101011"; -- -0.08017413810363298
	pesos_i(25820) := b"1111111111111111_1111111111111111_1111100110110011_0011101110110010"; -- -0.02460886855007048
	pesos_i(25821) := b"0000000000000000_0000000000000000_0010010001101110_1000010110010101"; -- 0.14231142894951274
	pesos_i(25822) := b"1111111111111111_1111111111111111_1111110001000101_0010110011111000"; -- -0.014569463111125027
	pesos_i(25823) := b"0000000000000000_0000000000000000_0001100111000100_1010111000101011"; -- 0.1006573538746318
	pesos_i(25824) := b"0000000000000000_0000000000000000_0010101110111001_0001011011100011"; -- 0.1707929901399053
	pesos_i(25825) := b"1111111111111111_1111111111111111_1100111000110111_0011110110101111"; -- -0.19446959003584455
	pesos_i(25826) := b"0000000000000000_0000000000000000_0001110110101011_1111100001011110"; -- 0.11590530680219394
	pesos_i(25827) := b"0000000000000000_0000000000000000_0000110101010110_1000110111000101"; -- 0.05210195597620202
	pesos_i(25828) := b"0000000000000000_0000000000000000_0010001100110000_1001010010000100"; -- 0.1374600241595097
	pesos_i(25829) := b"0000000000000000_0000000000000000_0000100000010000_1111111010100001"; -- 0.03150931777026796
	pesos_i(25830) := b"1111111111111111_1111111111111111_1101010000110110_1000110000100010"; -- -0.17104267293947123
	pesos_i(25831) := b"0000000000000000_0000000000000000_0000001011110000_0110101011011001"; -- 0.011480978094146593
	pesos_i(25832) := b"1111111111111111_1111111111111111_1101111111000010_0101000100001010"; -- -0.12594121465048144
	pesos_i(25833) := b"1111111111111111_1111111111111111_1100110000110111_0100011001010001"; -- -0.20228157531624408
	pesos_i(25834) := b"0000000000000000_0000000000000000_0010010100100011_1101001010011100"; -- 0.14507786093041883
	pesos_i(25835) := b"0000000000000000_0000000000000000_0010000001100101_1100010100011010"; -- 0.12655288585036395
	pesos_i(25836) := b"1111111111111111_1111111111111111_1111001001111000_1111011011001111"; -- -0.05284173441506054
	pesos_i(25837) := b"1111111111111111_1111111111111111_1111001010110001_1100101011110101"; -- -0.051974597123881874
	pesos_i(25838) := b"0000000000000000_0000000000000000_0011001011111110_0011110001011001"; -- 0.19919182945667088
	pesos_i(25839) := b"0000000000000000_0000000000000000_0010101001110100_1111100011000111"; -- 0.165847347897833
	pesos_i(25840) := b"1111111111111111_1111111111111111_1111011101101100_0101110010110000"; -- -0.03350277622320291
	pesos_i(25841) := b"0000000000000000_0000000000000000_0001011010001110_0111010111110000"; -- 0.08811127758731158
	pesos_i(25842) := b"0000000000000000_0000000000000000_0001111010101000_0011010110010011"; -- 0.11975416993554287
	pesos_i(25843) := b"1111111111111111_1111111111111111_1110110001010011_0101000000110101"; -- -0.0768537398199284
	pesos_i(25844) := b"0000000000000000_0000000000000000_0011001100101010_0111101100101000"; -- 0.1998669597119907
	pesos_i(25845) := b"1111111111111111_1111111111111111_1111111110110110_1011110110101001"; -- -0.0011178458677121932
	pesos_i(25846) := b"1111111111111111_1111111111111111_1101101000000100_1011000010111001"; -- -0.14836593128248135
	pesos_i(25847) := b"1111111111111111_1111111111111111_1110000011100001_1100110001101000"; -- -0.12155458890162374
	pesos_i(25848) := b"0000000000000000_0000000000000000_0001111110010111_0101011111101101"; -- 0.12340306803749247
	pesos_i(25849) := b"1111111111111111_1111111111111111_1111001110000100_0111000010010001"; -- -0.048760380332869974
	pesos_i(25850) := b"0000000000000000_0000000000000000_0010110110111100_1101001111111101"; -- 0.17866253775310248
	pesos_i(25851) := b"1111111111111111_1111111111111111_1101101100100000_1110100010101101"; -- -0.14402910016503825
	pesos_i(25852) := b"0000000000000000_0000000000000000_0011010000100110_1010111100110001"; -- 0.2037152763012653
	pesos_i(25853) := b"0000000000000000_0000000000000000_0001001011001111_0010000100101011"; -- 0.07347304627757707
	pesos_i(25854) := b"0000000000000000_0000000000000000_0001000000111100_1001001010010011"; -- 0.06342426374467741
	pesos_i(25855) := b"0000000000000000_0000000000000000_0000100111111001_0001011010110111"; -- 0.03895704234680931
    return pesos_i;
    end function;
end package body mnist_weights;
    