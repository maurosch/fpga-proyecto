
-- ARCHIVO AUTOGENERADO CON ../../generate_weights_package.py

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.perceptron_package.perceptron_input;

package mnist_inputs_1 is
    function GetInputs1(Dummy: natural)
    return perceptron_input;
end package mnist_inputs_1;

package body mnist_inputs_1 is
    function GetInputs1(Dummy: natural) return perceptron_input is
        variable pesos_i : perceptron_input(63 downto 0);
    begin
	pesos_i(0) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(1) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(2) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(3) := b"0000000000000000_0000000000001100_0000000000000000_0000000000000000"; -- 12.0
	pesos_i(4) := b"0000000000000000_0000000000001101_0000000000000000_0000000000000000"; -- 13.0
	pesos_i(5) := b"0000000000000000_0000000000000101_0000000000000000_0000000000000000"; -- 5.0
	pesos_i(6) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(7) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(8) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(9) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(10) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(11) := b"0000000000000000_0000000000001011_0000000000000000_0000000000000000"; -- 11.0
	pesos_i(12) := b"0000000000000000_0000000000010000_0000000000000000_0000000000000000"; -- 16.0
	pesos_i(13) := b"0000000000000000_0000000000001001_0000000000000000_0000000000000000"; -- 9.0
	pesos_i(14) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(15) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(16) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(17) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(18) := b"0000000000000000_0000000000000011_0000000000000000_0000000000000000"; -- 3.0
	pesos_i(19) := b"0000000000000000_0000000000001111_0000000000000000_0000000000000000"; -- 15.0
	pesos_i(20) := b"0000000000000000_0000000000010000_0000000000000000_0000000000000000"; -- 16.0
	pesos_i(21) := b"0000000000000000_0000000000000110_0000000000000000_0000000000000000"; -- 6.0
	pesos_i(22) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(23) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(24) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(25) := b"0000000000000000_0000000000000111_0000000000000000_0000000000000000"; -- 7.0
	pesos_i(26) := b"0000000000000000_0000000000001111_0000000000000000_0000000000000000"; -- 15.0
	pesos_i(27) := b"0000000000000000_0000000000010000_0000000000000000_0000000000000000"; -- 16.0
	pesos_i(28) := b"0000000000000000_0000000000010000_0000000000000000_0000000000000000"; -- 16.0
	pesos_i(29) := b"0000000000000000_0000000000000010_0000000000000000_0000000000000000"; -- 2.0
	pesos_i(30) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(31) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(32) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(33) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(34) := b"0000000000000000_0000000000000001_0000000000000000_0000000000000000"; -- 1.0
	pesos_i(35) := b"0000000000000000_0000000000010000_0000000000000000_0000000000000000"; -- 16.0
	pesos_i(36) := b"0000000000000000_0000000000010000_0000000000000000_0000000000000000"; -- 16.0
	pesos_i(37) := b"0000000000000000_0000000000000011_0000000000000000_0000000000000000"; -- 3.0
	pesos_i(38) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(39) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(40) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(41) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(42) := b"0000000000000000_0000000000000001_0000000000000000_0000000000000000"; -- 1.0
	pesos_i(43) := b"0000000000000000_0000000000010000_0000000000000000_0000000000000000"; -- 16.0
	pesos_i(44) := b"0000000000000000_0000000000010000_0000000000000000_0000000000000000"; -- 16.0
	pesos_i(45) := b"0000000000000000_0000000000000110_0000000000000000_0000000000000000"; -- 6.0
	pesos_i(46) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(47) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(48) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(49) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(50) := b"0000000000000000_0000000000000001_0000000000000000_0000000000000000"; -- 1.0
	pesos_i(51) := b"0000000000000000_0000000000010000_0000000000000000_0000000000000000"; -- 16.0
	pesos_i(52) := b"0000000000000000_0000000000010000_0000000000000000_0000000000000000"; -- 16.0
	pesos_i(53) := b"0000000000000000_0000000000000110_0000000000000000_0000000000000000"; -- 6.0
	pesos_i(54) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(55) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(56) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(57) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(58) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(59) := b"0000000000000000_0000000000001011_0000000000000000_0000000000000000"; -- 11.0
	pesos_i(60) := b"0000000000000000_0000000000010000_0000000000000000_0000000000000000"; -- 16.0
	pesos_i(61) := b"0000000000000000_0000000000001010_0000000000000000_0000000000000000"; -- 10.0
	pesos_i(62) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(63) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
    return pesos_i;
    end function;
end package body mnist_inputs_1;
    