
-- ARCHIVO AUTOGENERADO CON generate_weights_package.py

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.perceptron_package.perceptron_input;

package mnist_biases is
    function GetBiases(Dummy: natural)
    return perceptron_input;
end package mnist_biases;

package body mnist_biases is
    function GetBiases(Dummy: natural) return perceptron_input is
        variable pesos_i : perceptron_input(265 downto 0);
    begin
	pesos_i(0) := b"1111111111111111_1111111111111111_1101110101101110_0100100010100100"; -- -0.1350359535341312
	pesos_i(1) := b"1111111111111111_1111111111111111_1111110011110100_1001101100001010"; -- -0.011892614424570399
	pesos_i(2) := b"0000000000000000_0000000000000000_0010100011110011_1100100011100011"; -- 0.1599698595987859
	pesos_i(3) := b"0000000000000000_0000000000000000_0010010011011110_1111111111111011"; -- 0.14402770875317616
	pesos_i(4) := b"0000000000000000_0000000000000000_0000010000000010_1000001010001110"; -- 0.015663299341968032
	pesos_i(5) := b"1111111111111111_1111111111111111_1110001100010111_0011100111101011"; -- -0.11292684574775753
	pesos_i(6) := b"0000000000000000_0000000000000000_0000001001110110_0000100010001100"; -- 0.009613546515039149
	pesos_i(7) := b"1111111111111111_1111111111111111_1110001111000100_0100000010100110"; -- -0.11028667398704388
	pesos_i(8) := b"1111111111111111_1111111111111111_1110101101111001_1011011000111001"; -- -0.08017407532108937
	pesos_i(9) := b"0000000000000000_0000000000000000_0000010010110100_1011011011001001"; -- 0.018382476827610125
	pesos_i(10) := b"0000000000000000_0000000000000000_0001001011010010_0010111101100010"; -- 0.07351966990199012
	pesos_i(11) := b"1111111111111111_1111111111111111_1111111000001000_0011001010010001"; -- -0.007687415799496988
	pesos_i(12) := b"0000000000000000_0000000000000000_0000101010010111_1110001011001011"; -- 0.04138009510588794
	pesos_i(13) := b"0000000000000000_0000000000000000_0001000101100011_0101000110000101"; -- 0.06792172912707425
	pesos_i(14) := b"0000000000000000_0000000000000000_0001000000101010_1101101010000010"; -- 0.06315389323539393
	pesos_i(15) := b"0000000000000000_0000000000000000_0010001101001111_0111101010011000"; -- 0.13793150155842407
	pesos_i(16) := b"0000000000000000_0000000000000000_0010100110010011_0101000100011000"; -- 0.16240412560525244
	pesos_i(17) := b"1111111111111111_1111111111111111_1101101000110010_1101100100101000"; -- -0.1476616171309888
	pesos_i(18) := b"0000000000000000_0000000000000000_0000011110001111_1000011101000011"; -- 0.029533818987653757
	pesos_i(19) := b"1111111111111111_1111111111111111_1111010000010001_0100100001110000"; -- -0.04661128292240073
	pesos_i(20) := b"1111111111111111_1111111111111111_1101101010010001_1100111001110101"; -- -0.14621266990189902
	pesos_i(21) := b"1111111111111111_1111111111111111_1111000101000101_0010010011100111"; -- -0.05753869393698238
	pesos_i(22) := b"1111111111111111_1111111111111111_1110010001100010_0001110110000101"; -- -0.10787787919214277
	pesos_i(23) := b"0000000000000000_0000000000000000_0001011101110011_0011011100010110"; -- 0.09160179410418168
	pesos_i(24) := b"1111111111111111_1111111111111111_1101111000100100_1110101101000101"; -- -0.13224916044338064
	pesos_i(25) := b"0000000000000000_0000000000000000_0000110111011100_1101010010010111"; -- 0.05415085489259466
	pesos_i(26) := b"0000000000000000_0000000000000000_0010011111001011_0000001010001110"; -- 0.1554414364825157
	pesos_i(27) := b"1111111111111111_1111111111111111_1101110110111111_0011100011111000"; -- -0.13380092557889273
	pesos_i(28) := b"0000000000000000_0000000000000000_0001111001011101_0100001101001001"; -- 0.11861057783218962
	pesos_i(29) := b"1111111111111111_1111111111111111_1111101010101000_0100101011111100"; -- -0.02086955408093424
	pesos_i(30) := b"1111111111111111_1111111111111111_1110001101111111_0101100111111010"; -- -0.11133802081955016
	pesos_i(31) := b"0000000000000000_0000000000000000_0010010010000010_1011111111100111"; -- 0.1426200809542133
	pesos_i(32) := b"0000000000000000_0000000000000000_0010001100100010_1110101000101110"; -- 0.13725150693794216
	pesos_i(33) := b"0000000000000000_0000000000000000_0010111001000100_0011000111101011"; -- 0.18072807308270522
	pesos_i(34) := b"0000000000000000_0000000000000000_0001110011000011_0111000011110110"; -- 0.11235719693057421
	pesos_i(35) := b"1111111111111111_1111111111111111_1110100100101001_1011001101000101"; -- -0.08920745434471457
	pesos_i(36) := b"0000000000000000_0000000000000000_0000100100100001_1100100001010110"; -- 0.035671731030766846
	pesos_i(37) := b"0000000000000000_0000000000000000_0010011111010111_0011010010101110"; -- 0.1556275296746553
	pesos_i(38) := b"0000000000000000_0000000000000000_0010000001100000_1011011011000011"; -- 0.12647573709336324
	pesos_i(39) := b"1111111111111111_1111111111111111_1111101101111101_0010010010001100"; -- -0.01762172309811969
	pesos_i(40) := b"1111111111111111_1111111111111111_1111100101100000_0000011011010011"; -- -0.025878499436476975
	pesos_i(41) := b"0000000000000000_0000000000000000_0010001100001001_0110011111100110"; -- 0.13686227181954008
	pesos_i(42) := b"1111111111111111_1111111111111111_1111011011000100_0000111100001010"; -- -0.03607088102313171
	pesos_i(43) := b"0000000000000000_0000000000000000_0010101010110010_1101011101111011"; -- 0.16679140819386692
	pesos_i(44) := b"0000000000000000_0000000000000000_0000100110001001_0100110111010000"; -- 0.03725134219453724
	pesos_i(45) := b"1111111111111111_1111111111111111_1110110000011100_1111010001010101"; -- -0.07768319052939009
	pesos_i(46) := b"1111111111111111_1111111111111111_1111011010100011_1110001111101010"; -- -0.036561732738629255
	pesos_i(47) := b"1111111111111111_1111111111111111_1110111100100100_1101110110101010"; -- -0.06584372133122388
	pesos_i(48) := b"0000000000000000_0000000000000000_0001110010011011_0101100000011011"; -- 0.11174536383016505
	pesos_i(49) := b"1111111111111111_1111111111111111_1110001100001011_1111111111100111"; -- -0.1130981503834217
	pesos_i(50) := b"1111111111111111_1111111111111111_1111000001101011_0111110111000001"; -- -0.06085981399138467
	pesos_i(51) := b"0000000000000000_0000000000000000_0001010111010001_0110000110000101"; -- 0.08522614954333929
	pesos_i(52) := b"0000000000000000_0000000000000000_0000100100110100_0010100110001000"; -- 0.0359521824628369
	pesos_i(53) := b"0000000000000000_0000000000000000_0010001111100101_0001011000011010"; -- 0.14021433015007423
	pesos_i(54) := b"0000000000000000_0000000000000000_0010010000110011_0111101000001001"; -- 0.14141047220411737
	pesos_i(55) := b"0000000000000000_0000000000000000_0010100101100010_0110101110001011"; -- 0.16165802138172317
	pesos_i(56) := b"1111111111111111_1111111111111111_1110100110110011_0110111111101010"; -- -0.08710575613000787
	pesos_i(57) := b"1111111111111111_1111111111111111_1111010100100001_0110011001000010"; -- -0.04245911502001535
	pesos_i(58) := b"1111111111111111_1111111111111111_1111011001101000_0011001111110000"; -- -0.0374724902991876
	pesos_i(59) := b"1111111111111111_1111111111111111_1111000110110101_0011000111010110"; -- -0.05582893871646137
	pesos_i(60) := b"0000000000000000_0000000000000000_0000001110000000_0000001011110010"; -- 0.013672050653750436
	pesos_i(61) := b"0000000000000000_0000000000000000_0010001111101001_1100111000000001"; -- 0.1402863265358549
	pesos_i(62) := b"0000000000000000_0000000000000000_0010101000101001_0001010110101111"; -- 0.1646894027146692
	pesos_i(63) := b"1111111111111111_1111111111111111_1110010011000100_0100010011001000"; -- -0.10638017759325118
	pesos_i(64) := b"0000000000000000_0000000000000000_0001110100001010_0000100011001111"; -- 0.11343436292908465
	pesos_i(65) := b"0000000000000000_0000000000000000_0010100000100011_1101101110010001"; -- 0.15679714471039666
	pesos_i(66) := b"0000000000000000_0000000000000000_0000000010111100_1001110010101101"; -- 0.002877990933952552
	pesos_i(67) := b"0000000000000000_0000000000000000_0000101100101110_1100011111011100"; -- 0.04368256673112424
	pesos_i(68) := b"0000000000000000_0000000000000000_0000110111111101_1100011001010100"; -- 0.054653544953798996
	pesos_i(69) := b"1111111111111111_1111111111111111_1111011110100000_1101100000011010"; -- -0.03270196318001552
	pesos_i(70) := b"0000000000000000_0000000000000000_0010000110101010_1101110001110101"; -- 0.13151338449077016
	pesos_i(71) := b"1111111111111111_1111111111111111_1110010011100001_1111001100100011"; -- -0.10592728044341615
	pesos_i(72) := b"0000000000000000_0000000000000000_0001101000000001_0001111100110000"; -- 0.10157961780889246
	pesos_i(73) := b"1111111111111111_1111111111111111_1111111100011010_1101011101010010"; -- -0.003496687369832857
	pesos_i(74) := b"1111111111111111_1111111111111111_1111110001001000_0111010100001111"; -- -0.014519389999365813
	pesos_i(75) := b"0000000000000000_0000000000000000_0010010011100110_0000000010111001"; -- 0.14413456447909348
	pesos_i(76) := b"0000000000000000_0000000000000000_0000100101101100_1011101110001110"; -- 0.03681537838282905
	pesos_i(77) := b"0000000000000000_0000000000000000_0000101111000001_1100010110010111"; -- 0.045925473677544196
	pesos_i(78) := b"0000000000000000_0000000000000000_0010010111010010_1010110001110000"; -- 0.14774587386477786
	pesos_i(79) := b"0000000000000000_0000000000000000_0010011111011001_1010001001000110"; -- 0.15566457957751764
	pesos_i(80) := b"0000000000000000_0000000000000000_0001100010001001_1010010111010101"; -- 0.0958503384975496
	pesos_i(81) := b"1111111111111111_1111111111111111_1110100101110100_0010001011011011"; -- -0.0880716528600765
	pesos_i(82) := b"1111111111111111_1111111111111111_1110110110000000_1000100101100011"; -- -0.07225743602508936
	pesos_i(83) := b"0000000000000000_0000000000000000_0010010100101001_0101100100000010"; -- 0.14516216555496986
	pesos_i(84) := b"1111111111111111_1111111111111111_1110001111011011_1000000001011101"; -- -0.10993192406329003
	pesos_i(85) := b"1111111111111111_1111111111111111_1110100010000110_0011001110001010"; -- -0.09170225027533188
	pesos_i(86) := b"0000000000000000_0000000000000000_0010000100111001_1110110111010110"; -- 0.12979017706918097
	pesos_i(87) := b"1111111111111111_1111111111111111_1111001101001011_1111111000001010"; -- -0.04962169885101447
	pesos_i(88) := b"1111111111111111_1111111111111111_1101101111011100_0111000101011110"; -- -0.14116755925834099
	pesos_i(89) := b"1111111111111111_1111111111111111_1110110110110010_0011111001010110"; -- -0.07149897004167402
	pesos_i(90) := b"0000000000000000_0000000000000000_0010001011010000_0001011111111001"; -- 0.13598775707591496
	pesos_i(91) := b"0000000000000000_0000000000000000_0010001111100001_0010101110111101"; -- 0.1401545844301488
	pesos_i(92) := b"1111111111111111_1111111111111111_1111100100110010_1011011011010011"; -- -0.02656991336785594
	pesos_i(93) := b"0000000000000000_0000000000000000_0010011001111000_1111010011101011"; -- 0.15028315299529843
	pesos_i(94) := b"0000000000000000_0000000000000000_0001101010111010_1010100110011001"; -- 0.10441074359051081
	pesos_i(95) := b"1111111111111111_1111111111111111_1111000110001100_1001000100110101"; -- -0.05644886454116038
	pesos_i(96) := b"0000000000000000_0000000000000000_0010000111111011_0001010011011010"; -- 0.13273744883718622
	pesos_i(97) := b"0000000000000000_0000000000000000_0010100110101101_1011101011100101"; -- 0.1628071602159637
	pesos_i(98) := b"0000000000000000_0000000000000000_0001111001000100_0110011011110110"; -- 0.11823123458205649
	pesos_i(99) := b"1111111111111111_1111111111111111_1101110001100111_1010000011110000"; -- -0.1390437521331466
	pesos_i(100) := b"0000000000000000_0000000000000000_0001010011100100_0111110111100110"; -- 0.08161150793322527
	pesos_i(101) := b"1111111111111111_1111111111111111_1110110101011100_0101111110001000"; -- -0.0728092473276585
	pesos_i(102) := b"0000000000000000_0000000000000000_0000010111010111_0111011010000001"; -- 0.02281895305405156
	pesos_i(103) := b"1111111111111111_1111111111111111_1110101001100010_1101101010110110"; -- -0.0844291024536489
	pesos_i(104) := b"1111111111111111_1111111111111111_1110011111111110_1101011011010000"; -- -0.09376771378175552
	pesos_i(105) := b"0000000000000000_0000000000000000_0001111010010110_1100000111011101"; -- 0.11948787360499687
	pesos_i(106) := b"1111111111111111_1111111111111111_1101111101010001_1001111001100011"; -- -0.12766084746736114
	pesos_i(107) := b"0000000000000000_0000000000000000_0001010111100111_1011010100101111"; -- 0.08556682966968368
	pesos_i(108) := b"1111111111111111_1111111111111111_1101101111110100_1111001110001001"; -- -0.14079358960257762
	pesos_i(109) := b"0000000000000000_0000000000000000_0000000100000000_0000000100100000"; -- 0.003906317168295407
	pesos_i(110) := b"1111111111111111_1111111111111111_1111011011000010_1001000101001100"; -- -0.03609363465638104
	pesos_i(111) := b"1111111111111111_1111111111111111_1111000010110100_0010000110000101"; -- -0.059751419977000585
	pesos_i(112) := b"1111111111111111_1111111111111111_1101001111100001_1111101100011101"; -- -0.17233305491429984
	pesos_i(113) := b"0000000000000000_0000000000000000_0000110111100011_1010101010011111"; -- 0.05425516486741021
	pesos_i(114) := b"1111111111111111_1111111111111111_1110001011110110_0100000001110010"; -- -0.11342999659600124
	pesos_i(115) := b"0000000000000000_0000000000000000_0000111011101111_0001000011011000"; -- 0.05833535450802444
	pesos_i(116) := b"1111111111111111_1111111111111111_1110011000101000_1001100001100011"; -- -0.10094306542213745
	pesos_i(117) := b"0000000000000000_0000000000000000_0001101011111110_1010111010101101"; -- 0.10544864387848876
	pesos_i(118) := b"0000000000000000_0000000000000000_0001000101101001_1011010000110110"; -- 0.06801916421480662
	pesos_i(119) := b"0000000000000000_0000000000000000_0001010010111101_0110100011000110"; -- 0.08101515609867492
	pesos_i(120) := b"1111111111111111_1111111111111111_1110000111000110_0110001110110000"; -- -0.1180665679815449
	pesos_i(121) := b"1111111111111111_1111111111111111_1111101110001000_1010000101010011"; -- -0.017446439107842784
	pesos_i(122) := b"0000000000000000_0000000000000000_0000111000100011_1011101100010101"; -- 0.05523270855206253
	pesos_i(123) := b"0000000000000000_0000000000000000_0000100101001001_1101111110111111"; -- 0.03628347795609252
	pesos_i(124) := b"0000000000000000_0000000000000000_0001011110101001_0111100100100011"; -- 0.09242970566919921
	pesos_i(125) := b"0000000000000000_0000000000000000_0001110000101000_1001101010111000"; -- 0.10999457343327712
	pesos_i(126) := b"0000000000000000_0000000000000000_0000010101110111_0001000010011001"; -- 0.021348035241444224
	pesos_i(127) := b"0000000000000000_0000000000000000_0001010010101000_1110100000101011"; -- 0.08070231493563812
	pesos_i(128) := b"0000000000000000_0000000000000000_0001110101101101_1010001000101111"; -- 0.11495412496365982
	pesos_i(129) := b"0000000000000000_0000000000000000_0000110001010010_0001100111001011"; -- 0.048127758117575754
	pesos_i(130) := b"0000000000000000_0000000000000000_0001000111000111_1010011111111100"; -- 0.06945276166521293
	pesos_i(131) := b"1111111111111111_1111111111111111_1110111001001101_0011101001001111"; -- -0.06913409781589396
	pesos_i(132) := b"1111111111111111_1111111111111111_1110100100001111_0101110010010111"; -- -0.08960934941355624
	pesos_i(133) := b"1111111111111111_1111111111111111_1110011100110010_0110001010100111"; -- -0.09688743036616648
	pesos_i(134) := b"0000000000000000_0000000000000000_0000101111011111_0011100000011000"; -- 0.046374803297339465
	pesos_i(135) := b"0000000000000000_0000000000000000_0000011001101000_1010011000011100"; -- 0.025034314837915485
	pesos_i(136) := b"1111111111111111_1111111111111111_1110101101110011_0000011111101111"; -- -0.08027601646056177
	pesos_i(137) := b"1111111111111111_1111111111111111_1110011101011011_0011111000110001"; -- -0.0962639932910737
	pesos_i(138) := b"1111111111111111_1111111111111111_1111101010111011_1000100001001001"; -- -0.02057598331514297
	pesos_i(139) := b"0000000000000000_0000000000000000_0010011011101100_0100000000010110"; -- 0.15204239410951959
	pesos_i(140) := b"0000000000000000_0000000000000000_0010000101011111_0111101100001000"; -- 0.1303631682276769
	pesos_i(141) := b"0000000000000000_0000000000000000_0000010100110111_1010110000010001"; -- 0.02038073935682177
	pesos_i(142) := b"1111111111111111_1111111111111111_1111110110111110_1100000010111010"; -- -0.008808092658016398
	pesos_i(143) := b"0000000000000000_0000000000000000_0001011000100110_1101111111001011"; -- 0.08653067307325048
	pesos_i(144) := b"1111111111111111_1111111111111111_1110111100100001_1010100001101110"; -- -0.06589267082304083
	pesos_i(145) := b"1111111111111111_1111111111111111_1111100110111110_0001101000001100"; -- -0.024443027539960832
	pesos_i(146) := b"0000000000000000_0000000000000000_0000100010011011_1010010000111001"; -- 0.0336249007327132
	pesos_i(147) := b"0000000000000000_0000000000000000_0000010011001000_1100110001010111"; -- 0.01868893736264226
	pesos_i(148) := b"1111111111111111_1111111111111111_1110011001010100_0110000000101101"; -- -0.10027502931161117
	pesos_i(149) := b"0000000000000000_0000000000000000_0001001101101011_0101000111000110"; -- 0.07585631456169734
	pesos_i(150) := b"1111111111111111_1111111111111111_1111101000101011_0100101111011000"; -- -0.022776851423374628
	pesos_i(151) := b"0000000000000000_0000000000000000_0001101100100010_0011001011101100"; -- 0.1059905839532164
	pesos_i(152) := b"0000000000000000_0000000000000000_0000001110001100_0010010111011000"; -- 0.013857236159396658
	pesos_i(153) := b"1111111111111111_1111111111111111_1111100111111101_1100111110111011"; -- -0.02347089459307635
	pesos_i(154) := b"0000000000000000_0000000000000000_0000100100111111_0010010100100001"; -- 0.03611976684133228
	pesos_i(155) := b"1111111111111111_1111111111111111_1111000110110111_1000001001100100"; -- -0.0557936198039341
	pesos_i(156) := b"0000000000000000_0000000000000000_0001101111110001_0011100011111000"; -- 0.10914951375639251
	pesos_i(157) := b"0000000000000000_0000000000000000_0001100111110000_1001011001100100"; -- 0.10132732343902692
	pesos_i(158) := b"1111111111111111_1111111111111111_1111101111010010_0000001101010111"; -- -0.01632670528842127
	pesos_i(159) := b"1111111111111111_1111111111111111_1101111111110010_0111000111011001"; -- -0.12520683724122825
	pesos_i(160) := b"0000000000000000_0000000000000000_0010011010010100_1010111000001101"; -- 0.15070617495517424
	pesos_i(161) := b"0000000000000000_0000000000000000_0000011111110000_1011010000001000"; -- 0.031016590092876682
	pesos_i(162) := b"1111111111111111_1111111111111111_1101110000010000_1111011010000110"; -- -0.1403661654563001
	pesos_i(163) := b"1111111111111111_1111111111111111_1110100101001011_0101011010000110"; -- -0.0886941836649579
	pesos_i(164) := b"0000000000000000_0000000000000000_0001010111111110_0011000110001110"; -- 0.08590993616196733
	pesos_i(165) := b"1111111111111111_1111111111111111_1110000011001110_1100101001100111"; -- -0.12184462541758677
	pesos_i(166) := b"0000000000000000_0000000000000000_0000000111000001_0100011100101010"; -- 0.006855437933019849
	pesos_i(167) := b"0000000000000000_0000000000000000_0010000010101110_1101001000100011"; -- 0.12766755450900763
	pesos_i(168) := b"0000000000000000_0000000000000000_0001111101110010_0010101110110011"; -- 0.12283585654890164
	pesos_i(169) := b"1111111111111111_1111111111111111_1110100100000100_0001010011010010"; -- -0.08978147380773062
	pesos_i(170) := b"0000000000000000_0000000000000000_0000010110001100_0000001101010011"; -- 0.02166767851129414
	pesos_i(171) := b"0000000000000000_0000000000000000_0000111000111010_0000010111100000"; -- 0.05557285992326075
	pesos_i(172) := b"1111111111111111_1111111111111111_1111111110111000_1010110001010001"; -- -0.0010883620359936003
	pesos_i(173) := b"1111111111111111_1111111111111111_1111011001111011_0001001111110010"; -- -0.037184480100054325
	pesos_i(174) := b"1111111111111111_1111111111111111_1101101101100011_0110111100110101"; -- -0.14301400144311732
	pesos_i(175) := b"0000000000000000_0000000000000000_0010010000001101_1000110101101011"; -- 0.14083179333892068
	pesos_i(176) := b"1111111111111111_1111111111111111_1110001111001001_1011011110001111"; -- -0.11020329245775144
	pesos_i(177) := b"1111111111111111_1111111111111111_1110000111011001_1111100101010010"; -- -0.11776773212059136
	pesos_i(178) := b"1111111111111111_1111111111111111_1101111001110000_0111011101000001"; -- -0.13109640757630686
	pesos_i(179) := b"0000000000000000_0000000000000000_0010011100101001_1001111001000101"; -- 0.15297879391635186
	pesos_i(180) := b"1111111111111111_1111111111111111_1110011101101101_1101110110010001"; -- -0.09597983550547415
	pesos_i(181) := b"0000000000000000_0000000000000000_0010010011111101_1011101011101010"; -- 0.14449661453231963
	pesos_i(182) := b"0000000000000000_0000000000000000_0001011010001001_1101111110101001"; -- 0.08804128534113569
	pesos_i(183) := b"0000000000000000_0000000000000000_0000111100000011_0000011110011101"; -- 0.058639980075212414
	pesos_i(184) := b"0000000000000000_0000000000000000_0001101011011111_0100011001111111"; -- 0.10496941190140935
	pesos_i(185) := b"0000000000000000_0000000000000000_0010001110001111_1111110001110011"; -- 0.1389158040171386
	pesos_i(186) := b"1111111111111111_1111111111111111_1110110001010101_0001010001011111"; -- -0.07682678881052461
	pesos_i(187) := b"1111111111111111_1111111111111111_1111011111111111_0100011100111101"; -- -0.03126101255974925
	pesos_i(188) := b"1111111111111111_1111111111111111_1111000010110010_1001000100011000"; -- -0.059775287327868507
	pesos_i(189) := b"1111111111111111_1111111111111111_1111100110111110_1111011010010101"; -- -0.02442988272073828
	pesos_i(190) := b"1111111111111111_1111111111111111_1111101001101000_1111111111011111"; -- -0.021835334872490737
	pesos_i(191) := b"1111111111111111_1111111111111111_1111000100011000_0100111000111010"; -- -0.058222876473798035
	pesos_i(192) := b"1111111111111111_1111111111111111_1110110111010110_1100011001111101"; -- -0.07094153832016406
	pesos_i(193) := b"0000000000000000_0000000000000000_0000101110001000_1110000010100000"; -- 0.0450573340425211
	pesos_i(194) := b"0000000000000000_0000000000000000_0010011011110010_0010010011110101"; -- 0.15213232976151467
	pesos_i(195) := b"0000000000000000_0000000000000000_0000110110000111_1000101110001010"; -- 0.052849503739421023
	pesos_i(196) := b"0000000000000000_0000000000000000_0001010000000001_0111100100111010"; -- 0.07814748434558377
	pesos_i(197) := b"0000000000000000_0000000000000000_0001001010110001_1101100111011011"; -- 0.07302629086453037
	pesos_i(198) := b"1111111111111111_1111111111111111_1111000101011110_0101000011001101"; -- -0.05715460778579488
	pesos_i(199) := b"0000000000000000_0000000000000000_0000000110010100_0110111111110010"; -- 0.006171223188607941
	pesos_i(200) := b"0000000000000000_0000000000000000_0001011111001111_1100100001111011"; -- 0.09301426887935134
	pesos_i(201) := b"1111111111111111_1111111111111111_1110101101100011_1110000000100101"; -- -0.08050726979543063
	pesos_i(202) := b"0000000000000000_0000000000000000_0000010000001110_0000111011111001"; -- 0.01583951556310679
	pesos_i(203) := b"0000000000000000_0000000000000000_0001011111001011_1001110110001011"; -- 0.09295067436126966
	pesos_i(204) := b"1111111111111111_1111111111111111_1101101110101011_0101000110000000"; -- -0.14191713929515704
	pesos_i(205) := b"1111111111111111_1111111111111111_1111111100001110_1001100001001100"; -- -0.003683549239850729
	pesos_i(206) := b"1111111111111111_1111111111111111_1111100000010011_1000010000111111"; -- -0.03095220061745052
	pesos_i(207) := b"1111111111111111_1111111111111111_1110011000011100_1111001001101101"; -- -0.10112080410196223
	pesos_i(208) := b"1111111111111111_1111111111111111_1101111000011010_0001011000001101"; -- -0.13241445721643738
	pesos_i(209) := b"1111111111111111_1111111111111111_1110110000110100_0011011011100101"; -- -0.0773282710864104
	pesos_i(210) := b"1111111111111111_1111111111111111_1111101001011100_0000010000010110"; -- -0.02203344794430074
	pesos_i(211) := b"1111111111111111_1111111111111111_1111011111111100_0110101010111010"; -- -0.03130467386306667
	pesos_i(212) := b"0000000000000000_0000000000000000_0000000010011000_1010010111100110"; -- 0.0023292241690095116
	pesos_i(213) := b"1111111111111111_1111111111111111_1110001111000111_1010100010001101"; -- -0.11023470458018496
	pesos_i(214) := b"1111111111111111_1111111111111111_1110111111011010_1001111100000111"; -- -0.06307035530317191
	pesos_i(215) := b"0000000000000000_0000000000000000_0000010011110000_1011001011011000"; -- 0.019297769301954225
	pesos_i(216) := b"0000000000000000_0000000000000000_0001001000011111_0110101011100110"; -- 0.07079189419479777
	pesos_i(217) := b"1111111111111111_1111111111111111_1111100111111010_1001000100101100"; -- -0.023520399816128666
	pesos_i(218) := b"1111111111111111_1111111111111111_1111000010001100_0100011010111001"; -- -0.06035955420507093
	pesos_i(219) := b"1111111111111111_1111111111111111_1101111100111000_0001110000110001"; -- -0.12805007739337587
	pesos_i(220) := b"0000000000000000_0000000000000000_0001000001111001_0001001100110110"; -- 0.06434745846368282
	pesos_i(221) := b"1111111111111111_1111111111111111_1110001111010010_0100111101100000"; -- -0.1100721732705777
	pesos_i(222) := b"0000000000000000_0000000000000000_0000000000010011_0100001110000000"; -- 0.0002939403977093312
	pesos_i(223) := b"0000000000000000_0000000000000000_0001011011101010_1001010010101001"; -- 0.08951691742719659
	pesos_i(224) := b"1111111111111111_1111111111111111_1101111000111111_1101110101001001"; -- -0.13183800668050422
	pesos_i(225) := b"0000000000000000_0000000000000000_0000100100001101_0010101010001110"; -- 0.03535715079943706
	pesos_i(226) := b"1111111111111111_1111111111111111_1111001010101101_0101000001111010"; -- -0.05204293264860037
	pesos_i(227) := b"1111111111111111_1111111111111111_1111111111000101_0110110110011001"; -- -0.0008937360145663192
	pesos_i(228) := b"1111111111111111_1111111111111111_1110101100001110_1110010100001010"; -- -0.08180397518232378
	pesos_i(229) := b"1111111111111111_1111111111111111_1110001100110101_1010010100111011"; -- -0.11246268565163928
	pesos_i(230) := b"1111111111111111_1111111111111111_1110010000010000_0011100100111111"; -- -0.10912744725282665
	pesos_i(231) := b"0000000000000000_0000000000000000_0000010001111011_0011100101100101"; -- 0.017505251993836905
	pesos_i(232) := b"1111111111111111_1111111111111111_1110000011100000_0011110101100010"; -- -0.12157837252606266
	pesos_i(233) := b"0000000000000000_0000000000000000_0001101001110001_1101011110100110"; -- 0.10329959683246884
	pesos_i(234) := b"0000000000000000_0000000000000000_0010001010001010_0011111111000011"; -- 0.13492201328917394
	pesos_i(235) := b"0000000000000000_0000000000000000_0000101001111011_1100001010111011"; -- 0.040950937863221994
	pesos_i(236) := b"1111111111111111_1111111111111111_1111010101010110_1100010011100000"; -- -0.041644759475358055
	pesos_i(237) := b"1111111111111111_1111111111111111_1110001110101001_0000000101111011"; -- -0.11070242637599169
	pesos_i(238) := b"1111111111111111_1111111111111111_1111000010111100_0010000101011001"; -- -0.05962935991704599
	pesos_i(239) := b"0000000000000000_0000000000000000_0010010011011110_1110000000111010"; -- 0.14402581612690168
	pesos_i(240) := b"0000000000000000_0000000000000000_0001101110111100_0000011001001011"; -- 0.10833777740296915
	pesos_i(241) := b"1111111111111111_1111111111111111_1111111010010010_0101000001010111"; -- -0.0055799282376694315
	pesos_i(242) := b"0000000000000000_0000000000000000_0000100101110110_1000110110101110"; -- 0.03696523197751435
	pesos_i(243) := b"0000000000000000_0000000000000000_0001010111000001_1001101001001101"; -- 0.08498539336728475
	pesos_i(244) := b"1111111111111111_1111111111111111_1110010001110101_1011011100101010"; -- -0.10757880418597636
	pesos_i(245) := b"1111111111111111_1111111111111111_1110100010111011_1101011111011010"; -- -0.09088374077882376
	pesos_i(246) := b"1111111111111111_1111111111111111_1110010100011100_0001001010111000"; -- -0.10504038821295054
	pesos_i(247) := b"1111111111111111_1111111111111111_1111000000001010_0111000100100001"; -- -0.062340669043731756
	pesos_i(248) := b"1111111111111111_1111111111111111_1110000111011011_1000100001010011"; -- -0.11774394960499106
	pesos_i(249) := b"0000000000000000_0000000000000000_0000101011101011_1011110001101100"; -- 0.042659546230206534
	pesos_i(250) := b"0000000000000000_0000000000000000_0000110111010000_0010010100001001"; -- 0.05395728567261878
	pesos_i(251) := b"0000000000000000_0000000000000000_0000111110111010_1011101011000000"; -- 0.061443016005332106
	pesos_i(252) := b"1111111111111111_1111111111111111_1110000000011010_1001100111111001"; -- -0.12459409403998953
	pesos_i(253) := b"0000000000000000_0000000000000000_0000101001110100_1010111110001001"; -- 0.040842982179166
	pesos_i(254) := b"0000000000000000_0000000000000000_0010001001001100_0010101001111011"; -- 0.13397470008074094
	pesos_i(255) := b"0000000000000000_0000000000000000_0001010011011100_1011011101101100"; -- 0.0814928662792012
	pesos_i(256) := b"0000000000000000_0000000000000000_0001101100111010_0100111110011010"; -- 0.10635850432886756
	pesos_i(257) := b"1111111111111111_1111111111111111_1101011101110101_1001110111100101"; -- -0.15836156041279864
	pesos_i(258) := b"1111111111111111_1111111111111111_1101101010001110_0111000111110010"; -- -0.14626396037404404
	pesos_i(259) := b"1111111111111111_1111111111111111_1111010011010010_1000111011001000"; -- -0.043662143892466136
	pesos_i(260) := b"1111111111111111_1111111111111111_1101001000000011_1011011101110100"; -- -0.17963078903636343
	pesos_i(261) := b"0000000000000000_0000000000000000_0000110000000101_0010111011101101"; -- 0.046954091013566436
	pesos_i(262) := b"1111111111111111_1111111111111111_1110000101010101_0111110010100001"; -- -0.11978932436406942
	pesos_i(263) := b"0000000000000000_0000000000000000_0010001111010011_1101111011011101"; -- 0.13995163825199627
	pesos_i(264) := b"0000000000000000_0000000000000000_0001010011010100_1110100100101010"; -- 0.0813737608359553
	pesos_i(265) := b"1111111111111111_1111111111111111_1110001001110110_1111000101100110"; -- -0.11537257431688128
    return pesos_i;
    end function;
end package body mnist_biases;
    