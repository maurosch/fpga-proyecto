
-- ARCHIVO AUTOGENERADO CON generate_weights_package.py

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.perceptron_package.perceptron_input;

package mnist_biases is
    function GetBiases(Dummy: natural)
    return perceptron_input;
end package mnist_biases;

package body mnist_biases is
    function GetBiases(Dummy: natural) return perceptron_input is
        variable pesos_i : perceptron_input(265 downto 0);
    begin
	pesos_i(0) := b"1111111111111111_1111111111111111_1111110110011001_0001000000010011"; -- -0.009383197153153382
	pesos_i(1) := b"0000000000000000_0000000000000000_0010110111110101_1110100010010101"; -- 0.17953351637376913
	pesos_i(2) := b"0000000000000000_0000000000000000_0010011000000100_0000111010001010"; -- 0.14849940177163448
	pesos_i(3) := b"1111111111111111_1111111111111111_1110101010001111_1111110111100111"; -- -0.08374035931118998
	pesos_i(4) := b"1111111111111111_1111111111111111_1111000101001000_1011101001001000"; -- -0.057484013982823934
	pesos_i(5) := b"1111111111111111_1111111111111111_1110000011011000_0111110101000100"; -- -0.12169663518285156
	pesos_i(6) := b"0000000000000000_0000000000000000_0010000101101000_0000101000100000"; -- 0.13049376747325298
	pesos_i(7) := b"0000000000000000_0000000000000000_0010010011111110_0010101100111001"; -- 0.1445033088001187
	pesos_i(8) := b"0000000000000000_0000000000000000_0000011111011110_0111001001100100"; -- 0.030738019342439336
	pesos_i(9) := b"0000000000000000_0000000000000000_0001010011110111_0000001111000000"; -- 0.08189414444745871
	pesos_i(10) := b"0000000000000000_0000000000000000_0001111010100001_0100001011001100"; -- 0.11964814639462142
	pesos_i(11) := b"0000000000000000_0000000000000000_0000011010101011_0111101110111101"; -- 0.026054128305457516
	pesos_i(12) := b"1111111111111111_1111111111111111_1101111110010100_0010000110011010"; -- -0.12664594640442747
	pesos_i(13) := b"0000000000000000_0000000000000000_0000010001011010_1110010010111001"; -- 0.017011923871158907
	pesos_i(14) := b"1111111111111111_1111111111111111_1110111111000101_0011100110100111"; -- -0.0633968321659488
	pesos_i(15) := b"0000000000000000_0000000000000000_0001101101100100_0001110111101001"; -- 0.10699641167711407
	pesos_i(16) := b"0000000000000000_0000000000000000_0001010000101101_1100011010001011"; -- 0.07882347951092596
	pesos_i(17) := b"1111111111111111_1111111111111111_1111001111100011_0000011011110111"; -- -0.04731708973081464
	pesos_i(18) := b"0000000000000000_0000000000000000_0001110010000110_0011011110011110"; -- 0.11142299276253821
	pesos_i(19) := b"1111111111111111_1111111111111111_1110000011000011_1000010001010101"; -- -0.12201664841526794
	pesos_i(20) := b"0000000000000000_0000000000000000_0001000011001001_1010101100101011"; -- 0.06557721911756575
	pesos_i(21) := b"1111111111111111_1111111111111111_1111001001101110_0000101001001001"; -- -0.053008420115651225
	pesos_i(22) := b"0000000000000000_0000000000000000_0001001111101101_0011110010000111"; -- 0.07783869081543911
	pesos_i(23) := b"1111111111111111_1111111111111111_1110111010101011_0110110111011011"; -- -0.06769669906302725
	pesos_i(24) := b"0000000000000000_0000000000000000_0000110110011100_0001010111000110"; -- 0.05316291890654342
	pesos_i(25) := b"0000000000000000_0000000000000000_0000011100110010_0100000010000001"; -- 0.028110534278575888
	pesos_i(26) := b"0000000000000000_0000000000000000_0001000110111010_1011011110110010"; -- 0.06925533381124425
	pesos_i(27) := b"1111111111111111_1111111111111111_1111110001101101_1001110001010000"; -- -0.013952474934220532
	pesos_i(28) := b"1111111111111111_1111111111111111_1111110110110110_1110011110101110"; -- -0.008927841093504123
	pesos_i(29) := b"1111111111111111_1111111111111111_1101100110000101_0100111001011111"; -- -0.15030965977145058
	pesos_i(30) := b"0000000000000000_0000000000000000_0001111100100101_0101100100110011"; -- 0.12166364186108153
	pesos_i(31) := b"1111111111111111_1111111111111111_1110011001101100_0110000111011100"; -- -0.09990871786128065
	pesos_i(32) := b"1111111111111111_1111111111111111_1101101000010011_1110110010011001"; -- -0.14813348061900153
	pesos_i(33) := b"0000000000000000_0000000000000000_0000010010111101_1101011010000011"; -- 0.018521697117166072
	pesos_i(34) := b"0000000000000000_0000000000000000_0000010001001001_0010010000000010"; -- 0.016741037847119982
	pesos_i(35) := b"0000000000000000_0000000000000000_0001011100111011_1101010001101101"; -- 0.09075668015438212
	pesos_i(36) := b"1111111111111111_1111111111111111_1110011111110101_0101111010110101"; -- -0.09391220158847748
	pesos_i(37) := b"0000000000000000_0000000000000000_0001111000010111_0101001000111000"; -- 0.11754335267975556
	pesos_i(38) := b"1111111111111111_1111111111111111_1101011011010110_1011011011011011"; -- -0.16078622005910048
	pesos_i(39) := b"0000000000000000_0000000000000000_0001101011011101_1111111011000100"; -- 0.1049498776108671
	pesos_i(40) := b"1111111111111111_1111111111111111_1111011100010000_0000100011001010"; -- -0.03491158546631003
	pesos_i(41) := b"0000000000000000_0000000000000000_0000101110101111_0001011001011110"; -- 0.04564037131183811
	pesos_i(42) := b"1111111111111111_1111111111111111_1111111101111101_1101000010101011"; -- -0.0019864637757097503
	pesos_i(43) := b"1111111111111111_1111111111111111_1101111110111011_1011010011000100"; -- -0.12604208205321943
	pesos_i(44) := b"1111111111111111_1111111111111111_1110010100110011_0110101011101001"; -- -0.10468417950568205
	pesos_i(45) := b"0000000000000000_0000000000000000_0001110110110101_0100000110101101"; -- 0.11604700551712811
	pesos_i(46) := b"0000000000000000_0000000000000000_0001001010001000_0011110110111000"; -- 0.07239137394050617
	pesos_i(47) := b"1111111111111111_1111111111111111_1110001010101010_0101101110001000"; -- -0.11458805018445842
	pesos_i(48) := b"0000000000000000_0000000000000000_0010100011111111_1001000010101111"; -- 0.16014961496777866
	pesos_i(49) := b"0000000000000000_0000000000000000_0010010010101111_1100000000110000"; -- 0.1433067434549253
	pesos_i(50) := b"1111111111111111_1111111111111111_1110011001010010_0111001011101001"; -- -0.10030443012269587
	pesos_i(51) := b"1111111111111111_1111111111111111_1111110100111010_0011000001110100"; -- -0.01083085226330652
	pesos_i(52) := b"0000000000000000_0000000000000000_0000111001010000_0011111100110111"; -- 0.055911971076233434
	pesos_i(53) := b"1111111111111111_1111111111111111_1110101100100000_0111000010100011"; -- -0.0815362550206136
	pesos_i(54) := b"0000000000000000_0000000000000000_0001100011001001_1011110111100011"; -- 0.09682833461752295
	pesos_i(55) := b"1111111111111111_1111111111111111_1111111000010111_0110101010100110"; -- -0.007455191062507179
	pesos_i(56) := b"1111111111111111_1111111111111111_1110100001011000_0110100101011100"; -- -0.09240094666658212
	pesos_i(57) := b"1111111111111111_1111111111111111_1111111000100110_0011101010011011"; -- -0.0072291729377653244
	pesos_i(58) := b"0000000000000000_0000000000000000_0010010011000011_1100100011011001"; -- 0.1436124353696695
	pesos_i(59) := b"1111111111111111_1111111111111111_1111110011110111_0000001001110011"; -- -0.011855933020428436
	pesos_i(60) := b"0000000000000000_0000000000000000_0000111101110110_0010001001000110"; -- 0.06039632984939652
	pesos_i(61) := b"1111111111111111_1111111111111111_1101010111111010_0001011000010110"; -- -0.16415273624012933
	pesos_i(62) := b"0000000000000000_0000000000000000_0010111011100101_1111000010101010"; -- 0.18319610741955014
	pesos_i(63) := b"1111111111111111_1111111111111111_1111111010000101_1011010011110011"; -- -0.00577229556577803
	pesos_i(64) := b"1111111111111111_1111111111111111_1111101010011100_0011111010111000"; -- -0.021053390528404266
	pesos_i(65) := b"1111111111111111_1111111111111111_1110101101001110_1110101100000011"; -- -0.08082705660746922
	pesos_i(66) := b"1111111111111111_1111111111111111_1110010011111000_1101111110010011"; -- -0.10557749435420125
	pesos_i(67) := b"1111111111111111_1111111111111111_1101111010101100_0110110001010100"; -- -0.13018153138444202
	pesos_i(68) := b"0000000000000000_0000000000000000_0001111111000011_0101111001011011"; -- 0.12407483788333767
	pesos_i(69) := b"0000000000000000_0000000000000000_0000001011011111_1001000101011100"; -- 0.01122387394937672
	pesos_i(70) := b"0000000000000000_0000000000000000_0001010100110100_0111100110110100"; -- 0.08283196119017351
	pesos_i(71) := b"0000000000000000_0000000000000000_0000101110001011_0011100111111000"; -- 0.04509317687835767
	pesos_i(72) := b"0000000000000000_0000000000000000_0001000101101001_0001101010100011"; -- 0.06801001053311878
	pesos_i(73) := b"1111111111111111_1111111111111111_1111010010111100_0011111110101111"; -- -0.04400255187087084
	pesos_i(74) := b"0000000000000000_0000000000000000_0010001000111100_0011011010110101"; -- 0.13373128802387166
	pesos_i(75) := b"1111111111111111_1111111111111111_1110001011111011_0110010100101100"; -- -0.11335151352312782
	pesos_i(76) := b"0000000000000000_0000000000000000_0001110010001000_0000000111111001"; -- 0.11145031295691685
	pesos_i(77) := b"0000000000000000_0000000000000000_0000100110101000_1110011111011000"; -- 0.03773354556676659
	pesos_i(78) := b"1111111111111111_1111111111111111_1111000011100101_1001001110001000"; -- -0.05899694370787892
	pesos_i(79) := b"1111111111111111_1111111111111111_1110010101011000_0001100111111001"; -- -0.1041244285527508
	pesos_i(80) := b"1111111111111111_1111111111111111_1110110111000011_1101001111110001"; -- -0.07123065333200711
	pesos_i(81) := b"1111111111111111_1111111111111111_1111110001011110_0101010101110010"; -- -0.014185580989679555
	pesos_i(82) := b"0000000000000000_0000000000000000_0000001100101110_0100000101100111"; -- 0.012424552637081438
	pesos_i(83) := b"0000000000000000_0000000000000000_0001110010011001_1000100110011001"; -- 0.11171779616470662
	pesos_i(84) := b"0000000000000000_0000000000000000_0000101101010101_0011011101010110"; -- 0.04426904528022765
	pesos_i(85) := b"1111111111111111_1111111111111111_1110100101010011_1100110010101010"; -- -0.08856507149007453
	pesos_i(86) := b"1111111111111111_1111111111111111_1110000010001100_0100010100111011"; -- -0.12285964314213457
	pesos_i(87) := b"0000000000000000_0000000000000000_0000010111010100_0111011100001001"; -- 0.022773208314691564
	pesos_i(88) := b"0000000000000000_0000000000000000_0010001001001011_0111111111010111"; -- 0.13396452893475622
	pesos_i(89) := b"0000000000000000_0000000000000000_0001100000011100_0001010110111100"; -- 0.09417854144971233
	pesos_i(90) := b"0000000000000000_0000000000000000_0000000110111011_1001101001101000"; -- 0.006768846891552505
	pesos_i(91) := b"1111111111111111_1111111111111111_1101110001010100_1101111111001101"; -- -0.1393299221284637
	pesos_i(92) := b"0000000000000000_0000000000000000_0010100111101011_0001001101001100"; -- 0.1637432156919677
	pesos_i(93) := b"1111111111111111_1111111111111111_1101100000011111_1011001000000100"; -- -0.15576636705408006
	pesos_i(94) := b"1111111111111111_1111111111111111_1110010010011100_1101111101100101"; -- -0.10698131362597077
	pesos_i(95) := b"1111111111111111_1111111111111111_1110101100111110_0110110010000000"; -- -0.08107873794652617
	pesos_i(96) := b"1111111111111111_1111111111111111_1111000111010111_1100100010011111"; -- -0.05530115232767677
	pesos_i(97) := b"0000000000000000_0000000000000000_0001101110011101_0001110110111011"; -- 0.10786615196139575
	pesos_i(98) := b"1111111111111111_1111111111111111_1101011001010111_0111110100011000"; -- -0.16272752913826746
	pesos_i(99) := b"1111111111111111_1111111111111111_1111100111101110_1111100000000011"; -- -0.023697375517604855
	pesos_i(100) := b"0000000000000000_0000000000000000_0000100100000111_0001111010100000"; -- 0.03526488680392551
	pesos_i(101) := b"0000000000000000_0000000000000000_0010010000111000_1010110111100010"; -- 0.14148985630282288
	pesos_i(102) := b"0000000000000000_0000000000000000_0000100100000011_1001011111101111"; -- 0.03521108229574548
	pesos_i(103) := b"0000000000000000_0000000000000000_0010011000101001_0100011001010111"; -- 0.1490673028271701
	pesos_i(104) := b"1111111111111111_1111111111111111_1111010010111011_1000111110101001"; -- -0.04401304357170771
	pesos_i(105) := b"0000000000000000_0000000000000000_0000111100010011_0010001101010010"; -- 0.058885772154054286
	pesos_i(106) := b"1111111111111111_1111111111111111_1110001111000110_1000010100011001"; -- -0.1102520765737921
	pesos_i(107) := b"1111111111111111_1111111111111111_1110011000111100_0100110010000001"; -- -0.10064241269286492
	pesos_i(108) := b"0000000000000000_0000000000000000_0000000100101100_0010101001011110"; -- 0.004580162048822645
	pesos_i(109) := b"1111111111111111_1111111111111111_1111000100101000_0000101011110111"; -- -0.0579827449088674
	pesos_i(110) := b"0000000000000000_0000000000000000_0001100000000110_0001111100000111"; -- 0.09384340216367135
	pesos_i(111) := b"0000000000000000_0000000000000000_0001100101011101_1101010111000000"; -- 0.09908805786348665
	pesos_i(112) := b"0000000000000000_0000000000000000_0000101100010011_1010100110101000"; -- 0.04326877924408718
	pesos_i(113) := b"0000000000000000_0000000000000000_0001001000010101_0010101011110001"; -- 0.07063549415852804
	pesos_i(114) := b"0000000000000000_0000000000000000_0000011011011111_1011101100111001"; -- 0.026851369365889815
	pesos_i(115) := b"0000000000000000_0000000000000000_0010001111100100_1111101000000000"; -- 0.14021265518145734
	pesos_i(116) := b"0000000000000000_0000000000000000_0010010010010100_0001101011111010"; -- 0.14288490871771306
	pesos_i(117) := b"1111111111111111_1111111111111111_1110100001110101_1110111100101010"; -- -0.09195046644523293
	pesos_i(118) := b"1111111111111111_1111111111111111_1111110000100110_1101010011010000"; -- -0.015032481321834018
	pesos_i(119) := b"1111111111111111_1111111111111111_1111010111010000_1000011011101011"; -- -0.03978688023020434
	pesos_i(120) := b"1111111111111111_1111111111111111_1101101100000011_1101010000101110"; -- -0.1444728267188174
	pesos_i(121) := b"1111111111111111_1111111111111111_1110111001000001_1100101001111101"; -- -0.06930860951759182
	pesos_i(122) := b"0000000000000000_0000000000000000_0000111111110011_1111101100011101"; -- 0.062316603340217755
	pesos_i(123) := b"0000000000000000_0000000000000000_0000110011100110_0011111010101101"; -- 0.05038825733794477
	pesos_i(124) := b"0000000000000000_0000000000000000_0010000000101010_1100001111011100"; -- 0.12565254326495592
	pesos_i(125) := b"0000000000000000_0000000000000000_0001011010100001_0101010011000011"; -- 0.08839921717022552
	pesos_i(126) := b"0000000000000000_0000000000000000_0001000001010110_1011010100010111"; -- 0.06382304967952772
	pesos_i(127) := b"1111111111111111_1111111111111111_1101110101000001_0011000011111001"; -- -0.13572400968500523
	pesos_i(128) := b"1111111111111111_1111111111111111_1111111000100111_0000001100110000"; -- -0.007217217265337623
	pesos_i(129) := b"1111111111111111_1111111111111111_1111011000111010_0111111001101111"; -- -0.03816995422779551
	pesos_i(130) := b"0000000000000000_0000000000000000_0001100011100000_0010011011111101"; -- 0.09717029253995196
	pesos_i(131) := b"1111111111111111_1111111111111111_1111001101111000_1110100111001000"; -- -0.04893626074857809
	pesos_i(132) := b"0000000000000000_0000000000000000_0010010111000001_0011111100100100"; -- 0.1474799596743777
	pesos_i(133) := b"1111111111111111_1111111111111111_1111110101111111_0110111101010000"; -- -0.009774249085931604
	pesos_i(134) := b"0000000000000000_0000000000000000_0000101000010011_0010101001010101"; -- 0.03935494024450136
	pesos_i(135) := b"0000000000000000_0000000000000000_0000110001010111_0100100000001010"; -- 0.04820680841476364
	pesos_i(136) := b"0000000000000000_0000000000000000_0000011100010000_1111010000111011"; -- 0.027602447892004098
	pesos_i(137) := b"0000000000000000_0000000000000000_0010000111000010_0011001101110101"; -- 0.13186952215188585
	pesos_i(138) := b"1111111111111111_1111111111111111_1110101000101011_0001101011001001"; -- -0.08527977554441901
	pesos_i(139) := b"1111111111111111_1111111111111111_1101101100101011_1101110001111101"; -- -0.14386197998998837
	pesos_i(140) := b"1111111111111111_1111111111111111_1110111000101101_1000111010110111"; -- -0.0696173481312193
	pesos_i(141) := b"1111111111111111_1111111111111111_1111011101110001_1100110000000100"; -- -0.03341984666989403
	pesos_i(142) := b"1111111111111111_1111111111111111_1101110001001010_1010000101101101"; -- -0.13948622793635893
	pesos_i(143) := b"0000000000000000_0000000000000000_0001011100110110_0011010011110110"; -- 0.09067088144090196
	pesos_i(144) := b"0000000000000000_0000000000000000_0001000111100000_1001110101100100"; -- 0.06983359997695168
	pesos_i(145) := b"0000000000000000_0000000000000000_0000011111100110_0001000001101001"; -- 0.030854249662322333
	pesos_i(146) := b"0000000000000000_0000000000000000_0001100110100011_1010000100100110"; -- 0.10015303778517352
	pesos_i(147) := b"0000000000000000_0000000000000000_0001101111011010_1111110110101000"; -- 0.10881028500251862
	pesos_i(148) := b"0000000000000000_0000000000000000_0000010100111001_0100111001100100"; -- 0.020405673428939255
	pesos_i(149) := b"1111111111111111_1111111111111111_1110110101101001_1011010110001000"; -- -0.07260575708441612
	pesos_i(150) := b"1111111111111111_1111111111111111_1110101111000101_1000010111011011"; -- -0.07901729012227478
	pesos_i(151) := b"0000000000000000_0000000000000000_0000111011100110_0101011101010011"; -- 0.05820222636570341
	pesos_i(152) := b"0000000000000000_0000000000000000_0000011100001101_1110000000011101"; -- 0.02755547238460168
	pesos_i(153) := b"1111111111111111_1111111111111111_1111011001101001_1001101100000101"; -- -0.037451087375909714
	pesos_i(154) := b"1111111111111111_1111111111111111_1111101111011000_1100110010010110"; -- -0.01622315740401783
	pesos_i(155) := b"0000000000000000_0000000000000000_0000111001110000_0111101000011100"; -- 0.056403762576719134
	pesos_i(156) := b"1111111111111111_1111111111111111_1110000111000001_1100010101110100"; -- -0.11813703450497912
	pesos_i(157) := b"1111111111111111_1111111111111111_1111100101000101_1010011010101100"; -- -0.026280959091116426
	pesos_i(158) := b"1111111111111111_1111111111111111_1101100100000010_0010110000110101"; -- -0.15231059736503816
	pesos_i(159) := b"1111111111111111_1111111111111111_1111100000000110_1001011001011110"; -- -0.031149484705643635
	pesos_i(160) := b"1111111111111111_1111111111111111_1110011001011101_1100110010010110"; -- -0.10013123834703848
	pesos_i(161) := b"1111111111111111_1111111111111111_1110001010000010_0001001101100010"; -- -0.11520270211538414
	pesos_i(162) := b"1111111111111111_1111111111111111_1111110010110100_0110111000011111"; -- -0.012871854288006931
	pesos_i(163) := b"1111111111111111_1111111111111111_1111111110010000_0001011100011000"; -- -0.001707607853097499
	pesos_i(164) := b"1111111111111111_1111111111111111_1111101011011011_1010000101101011"; -- -0.020086203914859484
	pesos_i(165) := b"1111111111111111_1111111111111111_1111101011111000_1101101011011110"; -- -0.019640274926724294
	pesos_i(166) := b"1111111111111111_1111111111111111_1101111110111011_0011101000010100"; -- -0.12604939465467968
	pesos_i(167) := b"1111111111111111_1111111111111111_1101110001010111_0110101010000100"; -- -0.1392911366403112
	pesos_i(168) := b"1111111111111111_1111111111111111_1111010001111100_1010011011000100"; -- -0.044972970135872405
	pesos_i(169) := b"0000000000000000_0000000000000000_0000001000111101_0001111110000111"; -- 0.008745165423098951
	pesos_i(170) := b"0000000000000000_0000000000000000_0000000011101100_1100101110101101"; -- 0.0036132143391202536
	pesos_i(171) := b"0000000000000000_0000000000000000_0001111011101000_1001010111001001"; -- 0.1207364669492226
	pesos_i(172) := b"1111111111111111_1111111111111111_1110101111000001_1111110010111011"; -- -0.07907123974643727
	pesos_i(173) := b"1111111111111111_1111111111111111_1101110011000001_1001000011110010"; -- -0.13767141440580177
	pesos_i(174) := b"1111111111111111_1111111111111111_1111011101011111_1111011010010011"; -- -0.033691968179382026
	pesos_i(175) := b"0000000000000000_0000000000000000_0010000110101100_0001101100010000"; -- 0.13153237472959908
	pesos_i(176) := b"1111111111111111_1111111111111111_1111110111111101_0100111100010010"; -- -0.007853563317847817
	pesos_i(177) := b"0000000000000000_0000000000000000_0001110001100011_1110100000000010"; -- 0.11089944891526958
	pesos_i(178) := b"1111111111111111_1111111111111111_1110101111001010_0110011011010010"; -- -0.07894284593755921
	pesos_i(179) := b"1111111111111111_1111111111111111_1110110000010101_1110100010101110"; -- -0.07779069669660003
	pesos_i(180) := b"1111111111111111_1111111111111111_1111011100000001_1001101001000001"; -- -0.03513179702188162
	pesos_i(181) := b"1111111111111111_1111111111111111_1110110110100010_0100111011001011"; -- -0.07174212964991489
	pesos_i(182) := b"1111111111111111_1111111111111111_1101110011101110_0000000100110011"; -- -0.13699333678227224
	pesos_i(183) := b"0000000000000000_0000000000000000_0000101110111011_0001001010010011"; -- 0.04582325073124378
	pesos_i(184) := b"0000000000000000_0000000000000000_0001000010011010_1011011101010110"; -- 0.06486078127444965
	pesos_i(185) := b"0000000000000000_0000000000000000_0001111001100011_1001001101111101"; -- 0.11870691109021407
	pesos_i(186) := b"0000000000000000_0000000000000000_0010011001011101_1110010000110010"; -- 0.1498701688050842
	pesos_i(187) := b"0000000000000000_0000000000000000_0000100100010111_1101011011001100"; -- 0.035520005007665716
	pesos_i(188) := b"1111111111111111_1111111111111111_1101101010101111_1111101100001001"; -- -0.14575224911527157
	pesos_i(189) := b"1111111111111111_1111111111111111_1111110010001011_1100001111110000"; -- -0.01349234945419928
	pesos_i(190) := b"1111111111111111_1111111111111111_1111011010001110_0010111100110010"; -- -0.03689293887187958
	pesos_i(191) := b"1111111111111111_1111111111111111_1101110110110010_1010010000010000"; -- -0.13399290674118997
	pesos_i(192) := b"0000000000000000_0000000000000000_0000010101010011_1101100000010100"; -- 0.020810608640535334
	pesos_i(193) := b"0000000000000000_0000000000000000_0000000011010111_1000011011000011"; -- 0.0032886721212512064
	pesos_i(194) := b"0000000000000000_0000000000000000_0001100101011101_1100001000010101"; -- 0.09908688560756154
	pesos_i(195) := b"1111111111111111_1111111111111111_1111010110100011_1111010101001111"; -- -0.0404669459399445
	pesos_i(196) := b"0000000000000000_0000000000000000_0010000010000111_1000011100010111"; -- 0.12706798858219862
	pesos_i(197) := b"1111111111111111_1111111111111111_1110010001101110_0000111101100110"; -- -0.10769561545063763
	pesos_i(198) := b"1111111111111111_1111111111111111_1110110101000000_0111111101001011"; -- -0.07323460013666985
	pesos_i(199) := b"0000000000000000_0000000000000000_0010000110100111_0100011000111110"; -- 0.13145865453359967
	pesos_i(200) := b"1111111111111111_1111111111111111_1111100010100101_1010111111110110"; -- -0.028721811765427215
	pesos_i(201) := b"0000000000000000_0000000000000000_0000010101000011_0000111010100001"; -- 0.020554460812969216
	pesos_i(202) := b"1111111111111111_1111111111111111_1110111111001110_1011011011110110"; -- -0.06325203423803849
	pesos_i(203) := b"1111111111111111_1111111111111111_1110100101011101_0001011011000000"; -- -0.08842332654176449
	pesos_i(204) := b"1111111111111111_1111111111111111_1111100110000001_0011110010011111"; -- -0.02537175280770027
	pesos_i(205) := b"1111111111111111_1111111111111111_1111010001001110_0001010111000000"; -- -0.045683518141267025
	pesos_i(206) := b"0000000000000000_0000000000000000_0000100110000000_1100001101111011"; -- 0.03712102661750307
	pesos_i(207) := b"0000000000000000_0000000000000000_0000000100010101_1101100110111111"; -- 0.0042396632468996035
	pesos_i(208) := b"1111111111111111_1111111111111111_1110111011001011_0101001101001001"; -- -0.06721000154510999
	pesos_i(209) := b"0000000000000000_0000000000000000_0010001110010000_1001011111000011"; -- 0.13892506143947939
	pesos_i(210) := b"0000000000000000_0000000000000000_0010001111011001_1101100011001100"; -- 0.14004282931612572
	pesos_i(211) := b"0000000000000000_0000000000000000_0000011111011110_1110101110100110"; -- 0.03074524679837155
	pesos_i(212) := b"0000000000000000_0000000000000000_0010000011000011_1100110001111010"; -- 0.1279876515164792
	pesos_i(213) := b"1111111111111111_1111111111111111_1111101111011001_0111011000110010"; -- -0.016213047785996748
	pesos_i(214) := b"0000000000000000_0000000000000000_0001100101111001_0100100111110010"; -- 0.09950697103545007
	pesos_i(215) := b"1111111111111111_1111111111111111_1111111000101110_1110110001010101"; -- -0.007096509179970749
	pesos_i(216) := b"0000000000000000_0000000000000000_0001010010110100_1001010110010010"; -- 0.08088049719403453
	pesos_i(217) := b"0000000000000000_0000000000000000_0000011100110101_1110111111111111"; -- 0.02816677077326505
	pesos_i(218) := b"0000000000000000_0000000000000000_0001011111001111_0110010111010101"; -- 0.0930083889401501
	pesos_i(219) := b"1111111111111111_1111111111111111_1110111100110000_0000001111010010"; -- -0.06567360032745974
	pesos_i(220) := b"1111111111111111_1111111111111111_1110011100100000_1100110010001100"; -- -0.09715577690617645
	pesos_i(221) := b"1111111111111111_1111111111111111_1111111001110000_0010101110111100"; -- -0.006100908852936932
	pesos_i(222) := b"0000000000000000_0000000000000000_0001111001011100_0100110010110101"; -- 0.11859588068325294
	pesos_i(223) := b"0000000000000000_0000000000000000_0000011101001101_1110000001101111"; -- 0.028532054027379922
	pesos_i(224) := b"1111111111111111_1111111111111111_1111011001011101_0110101010100101"; -- -0.03763707600514111
	pesos_i(225) := b"0000000000000000_0000000000000000_0010001000011111_1000111001101011"; -- 0.13329401119482906
	pesos_i(226) := b"0000000000000000_0000000000000000_0000100100011111_0000000100100101"; -- 0.03562934074029467
	pesos_i(227) := b"0000000000000000_0000000000000000_0001111100101001_0000101010000101"; -- 0.12171998734637526
	pesos_i(228) := b"1111111111111111_1111111111111111_1110101111000011_0000010010111001"; -- -0.07905550461984645
	pesos_i(229) := b"1111111111111111_1111111111111111_1111010010110111_0111101010111110"; -- -0.044075325513627604
	pesos_i(230) := b"0000000000000000_0000000000000000_0000000101110111_1001011111001100"; -- 0.005731093806210861
	pesos_i(231) := b"0000000000000000_0000000000000000_0001000000111101_1111010111010101"; -- 0.06344543877882733
	pesos_i(232) := b"0000000000000000_0000000000000000_0001111000110110_0001001111001101"; -- 0.11801265494355206
	pesos_i(233) := b"1111111111111111_1111111111111111_1110111101010011_1000011011100011"; -- -0.0651317306307242
	pesos_i(234) := b"0000000000000000_0000000000000000_0010010110011011_0001001100000101"; -- 0.14689749590354295
	pesos_i(235) := b"0000000000000000_0000000000000000_0001100011110100_0010001000110100"; -- 0.09747518328383485
	pesos_i(236) := b"0000000000000000_0000000000000000_0000110010001111_1100101000101110"; -- 0.04906905776610572
	pesos_i(237) := b"0000000000000000_0000000000000000_0001100010101000_1101010010110000"; -- 0.09632615363944809
	pesos_i(238) := b"1111111111111111_1111111111111111_1110111110111011_1001000000100110"; -- -0.06354426445277486
	pesos_i(239) := b"1111111111111111_1111111111111111_1111001101111110_1100001000000101"; -- -0.048847078206796894
	pesos_i(240) := b"0000000000000000_0000000000000000_0001111101100011_1110111000101100"; -- 0.12261856637914481
	pesos_i(241) := b"1111111111111111_1111111111111111_1111010010000101_1010011011000010"; -- -0.04483564143814308
	pesos_i(242) := b"0000000000000000_0000000000000000_0000111110100001_0010010010111100"; -- 0.06105260464759899
	pesos_i(243) := b"1111111111111111_1111111111111111_1101110111100111_0100000101100001"; -- -0.13319007278375747
	pesos_i(244) := b"1111111111111111_1111111111111111_1111000110100101_1010111111100001"; -- -0.05606556656824531
	pesos_i(245) := b"0000000000000000_0000000000000000_0000110101011000_1011001101100111"; -- 0.05213471669665903
	pesos_i(246) := b"1111111111111111_1111111111111111_1110001000010010_1001100101100000"; -- -0.11690369993853204
	pesos_i(247) := b"0000000000000000_0000000000000000_0001011001100011_0100101100010100"; -- 0.08745259503099942
	pesos_i(248) := b"1111111111111111_1111111111111111_1111100100001010_0100000011000011"; -- -0.027187302104085466
	pesos_i(249) := b"1111111111111111_1111111111111111_1111001100011111_1111011001000000"; -- -0.0502935498548852
	pesos_i(250) := b"0000000000000000_0000000000000000_0010010010111111_0010000110101110"; -- 0.14354143622018298
	pesos_i(251) := b"0000000000000000_0000000000000000_0001010111011100_0000100011110001"; -- 0.08538871657369546
	pesos_i(252) := b"0000000000000000_0000000000000000_0010011011000110_0101100000011010"; -- 0.15146399149590603
	pesos_i(253) := b"0000000000000000_0000000000000000_0000100101010010_0000101001010111"; -- 0.03640808692206069
	pesos_i(254) := b"1111111111111111_1111111111111111_1111111100000100_0100000011010001"; -- -0.003841351370584754
	pesos_i(255) := b"1111111111111111_1111111111111111_1101101100011101_1100100101010000"; -- -0.14407674606916476
	pesos_i(256) := b"0000000000000000_0000000000000000_0000111101110110_1001001011001010"; -- 0.06040303649641018
	pesos_i(257) := b"1111111111111111_1111111111111111_1110110010100101_1110011111111111"; -- -0.07559347165252632
	pesos_i(258) := b"1111111111111111_1111111111111111_1111010111001011_1000101111111110"; -- -0.03986287160164401
	pesos_i(259) := b"1111111111111111_1111111111111111_1101111001010101_1110111001111010"; -- -0.1315012885467465
	pesos_i(260) := b"0000000000000000_0000000000000000_0011000101011111_0010000100110100"; -- 0.19285781392007292
	pesos_i(261) := b"0000000000000000_0000000000000000_0011001111011001_0000101001111101"; -- 0.20253053227958367
	pesos_i(262) := b"1111111111111111_1111111111111111_1110001110010100_0000100101101010"; -- -0.11102238818034395
	pesos_i(263) := b"0000000000000000_0000000000000000_0001111101010110_0111111110010101"; -- 0.12241361025715332
	pesos_i(264) := b"0000000000000000_0000000000000000_0000110101100000_0010010010111011"; -- 0.05224828307379944
	pesos_i(265) := b"1111111111111111_1111111111111111_1101010010001011_1110100100010111"; -- -0.16974013507228983
    return pesos_i;
    end function;
end package body mnist_biases;
    