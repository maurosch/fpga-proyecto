
-- ARCHIVO AUTOGENERADO CON generate_weights_package.py

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.perceptron_package.perceptron_input;

package mnist_weights is
    function GetWeights(Dummy: natural)
    return perceptron_input;
end package mnist_weights;

package body mnist_weights is
    function GetWeights(Dummy: natural) return perceptron_input is
        variable pesos_i : perceptron_input(7399 downto 0);
    begin
	pesos_i(0) := b"0000000000000000_0000000000000000_0010100101100100_0111011000010100"; -- 0.16168916695520524
	pesos_i(1) := b"1111111111111111_1111111111111111_1101010111101011_1000011001111001"; -- -0.16437491946130176
	pesos_i(2) := b"1111111111111111_1111111111111111_1111010011111100_0100111001110101"; -- -0.04302510872444143
	pesos_i(3) := b"1111111111111111_1111111111111111_1110111101010110_1110010111010101"; -- -0.06508029514611458
	pesos_i(4) := b"1111111111111111_1111111111111111_1110111010010101_1110000110110010"; -- -0.0680254880454667
	pesos_i(5) := b"1111111111111111_1111111111111111_1111001110110100_1101001111000101"; -- -0.0480220454926166
	pesos_i(6) := b"0000000000000000_0000000000000000_0011000000100011_0011011110000010"; -- 0.1880373660907228
	pesos_i(7) := b"1111111111111111_1111111111111111_1111000000101100_1010100000101100"; -- -0.061818589459907425
	pesos_i(8) := b"0000000000000000_0000000000000000_0001010011101100_1010110100100111"; -- 0.08173639483657602
	pesos_i(9) := b"1111111111111111_1111111111111111_1101111101101101_0100000111000001"; -- -0.12723912286435302
	pesos_i(10) := b"0000000000000000_0000000000000000_0010000110101011_1100100010111011"; -- 0.13152746737022608
	pesos_i(11) := b"1111111111111111_1111111111111111_1111000010111001_1000001110100100"; -- -0.05966927751518403
	pesos_i(12) := b"0000000000000000_0000000000000000_0010011100101100_0111101100011000"; -- 0.1530224736070871
	pesos_i(13) := b"1111111111111111_1111111111111111_1101101001111110_0110000000000101"; -- -0.14650916931145053
	pesos_i(14) := b"0000000000000000_0000000000000000_0001001110010011_0011001101111010"; -- 0.07646486033335059
	pesos_i(15) := b"1111111111111111_1111111111111111_1101010111010000_0101000011001101"; -- -0.1647901058347812
	pesos_i(16) := b"0000000000000000_0000000000000000_0001110001001101_1011101110100000"; -- 0.11056111014598546
	pesos_i(17) := b"1111111111111111_1111111111111111_1110000010110011_0100011010000111"; -- -0.12226447310613246
	pesos_i(18) := b"1111111111111111_1111111111111111_1101011011001001_0010110110100100"; -- -0.16099276302933554
	pesos_i(19) := b"1111111111111111_1111111111111111_1101100001010000_1100101011111100"; -- -0.15501719812333434
	pesos_i(20) := b"0000000000000000_0000000000000000_0001110100100011_0000010100010010"; -- 0.11381560984387501
	pesos_i(21) := b"0000000000000000_0000000000000000_0000111111001111_1011001001111100"; -- 0.06176295782888641
	pesos_i(22) := b"1111111111111111_1111111111111111_1101000101111101_0001011010101000"; -- -0.18168505095978982
	pesos_i(23) := b"0000000000000000_0000000000000000_0000110010011101_1010001110110110"; -- 0.049280387893639394
	pesos_i(24) := b"1111111111111111_1111111111111111_1111011101000011_0111000111011101"; -- -0.034127124240091705
	pesos_i(25) := b"1111111111111111_1111111111111111_1110000101110100_0000000111110111"; -- -0.11932361343632147
	pesos_i(26) := b"0000000000000000_0000000000000000_0001001000000011_0011001100110001"; -- 0.07036132764086905
	pesos_i(27) := b"1111111111111111_1111111111111111_1110000011001011_1101100011111011"; -- -0.12188953278908743
	pesos_i(28) := b"0000000000000000_0000000000000000_0010100110110010_0011001111000101"; -- 0.16287540005880996
	pesos_i(29) := b"0000000000000000_0000000000000000_0010101100000011_1111101000101011"; -- 0.16802943747837096
	pesos_i(30) := b"1111111111111111_1111111111111111_1101100110000101_0001101101000100"; -- -0.1503127059395032
	pesos_i(31) := b"0000000000000000_0000000000000000_0000001110010101_0010111101000100"; -- 0.01399512676443862
	pesos_i(32) := b"0000000000000000_0000000000000000_0001000101011101_0011111111010001"; -- 0.06782912122402635
	pesos_i(33) := b"0000000000000000_0000000000000000_0001100111010010_0110010111011110"; -- 0.10086666736552818
	pesos_i(34) := b"0000000000000000_0000000000000000_0000101110110110_1100001000010000"; -- 0.04575741665085242
	pesos_i(35) := b"0000000000000000_0000000000000000_0010001111010101_0101011000111101"; -- 0.13997401229316325
	pesos_i(36) := b"1111111111111111_1111111111111111_1110000111000101_1101100000010010"; -- -0.11807488987503206
	pesos_i(37) := b"0000000000000000_0000000000000000_0001100110110110_0100110010110010"; -- 0.10043792094292986
	pesos_i(38) := b"0000000000000000_0000000000000000_0000011110011000_1110000110011011"; -- 0.029676533116245712
	pesos_i(39) := b"1111111111111111_1111111111111111_1111110110111001_0100100011101111"; -- -0.008891526793067955
	pesos_i(40) := b"0000000000000000_0000000000000000_0010001101001010_0011011010011001"; -- 0.13785115467176112
	pesos_i(41) := b"1111111111111111_1111111111111111_1101010010111000_0101111001111110"; -- -0.16906175068475626
	pesos_i(42) := b"0000000000000000_0000000000000000_0010101011010001_0101000001100100"; -- 0.16725637861243858
	pesos_i(43) := b"0000000000000000_0000000000000000_0000101100010000_0010101010000110"; -- 0.04321542519750912
	pesos_i(44) := b"1111111111111111_1111111111111111_1101110001110011_0011110000100111"; -- -0.13886665386498687
	pesos_i(45) := b"0000000000000000_0000000000000000_0010101001111001_1100100011001100"; -- 0.16592078183303205
	pesos_i(46) := b"1111111111111111_1111111111111111_1111000111100111_0001010111101001"; -- -0.055067663793373633
	pesos_i(47) := b"0000000000000000_0000000000000000_0000010000010001_1110000010000000"; -- 0.015897780686757845
	pesos_i(48) := b"0000000000000000_0000000000000000_0001110101010011_0000101000010111"; -- 0.11454833088586641
	pesos_i(49) := b"0000000000000000_0000000000000000_0000100011101001_0100111111011110"; -- 0.03481005826906314
	pesos_i(50) := b"1111111111111111_1111111111111111_1101001101111010_1101001100001011"; -- -0.17390709855683886
	pesos_i(51) := b"1111111111111111_1111111111111111_1101010111010001_0100010101001010"; -- -0.16477553310425003
	pesos_i(52) := b"0000000000000000_0000000000000000_0001101010100010_0000001111000000"; -- 0.10403464736574625
	pesos_i(53) := b"0000000000000000_0000000000000000_0010001100101000_0001000111111000"; -- 0.13733017262521513
	pesos_i(54) := b"1111111111111111_1111111111111111_1110000000101000_0111111011111111"; -- -0.12438207876577743
	pesos_i(55) := b"0000000000000000_0000000000000000_0010011111011101_1111110001001101"; -- 0.15573098062017704
	pesos_i(56) := b"1111111111111111_1111111111111111_1100111111101001_1010110000100001"; -- -0.1878406924999155
	pesos_i(57) := b"1111111111111111_1111111111111111_1110111101001010_1001100011011110"; -- -0.06526798795987351
	pesos_i(58) := b"1111111111111111_1111111111111111_1101111101000110_1101011011010110"; -- -0.12782532957934217
	pesos_i(59) := b"1111111111111111_1111111111111111_1110111010101111_1011010010101100"; -- -0.06763144302596782
	pesos_i(60) := b"0000000000000000_0000000000000000_0010111011110101_1011101101001111"; -- 0.1834370677988631
	pesos_i(61) := b"1111111111111111_1111111111111111_1110111100001001_1101010110000001"; -- -0.06625619509943043
	pesos_i(62) := b"1111111111111111_1111111111111111_1111010000011000_0101111111111010"; -- -0.04650306846369398
	pesos_i(63) := b"0000000000000000_0000000000000000_0000001000100011_0001101100111001"; -- 0.008348180297315738
	pesos_i(64) := b"0000000000000000_0000000000000000_0010011110111100_0111101111110001"; -- 0.15521978971990102
	pesos_i(65) := b"1111111111111111_1111111111111111_1110010111011001_0101100100000101"; -- -0.10215228674349465
	pesos_i(66) := b"1111111111111111_1111111111111111_1111010110000001_0111001010101010"; -- -0.04099353164793762
	pesos_i(67) := b"1111111111111111_1111111111111111_1100111101101000_0101011111011001"; -- -0.1898140998208054
	pesos_i(68) := b"1111111111111111_1111111111111111_1110011001100001_1000000111000000"; -- -0.10007466381502692
	pesos_i(69) := b"1111111111111111_1111111111111111_1101001101010110_1001110111000110"; -- -0.17445959013328563
	pesos_i(70) := b"1111111111111111_1111111111111111_1111101101011000_0111011111001100"; -- -0.01818133609192915
	pesos_i(71) := b"1111111111111111_1111111111111111_1101000000111011_0000011010100000"; -- -0.18659933660992317
	pesos_i(72) := b"1111111111111111_1111111111111111_1111110110000111_1110000111100100"; -- -0.009645349250009205
	pesos_i(73) := b"1111111111111111_1111111111111111_1111010011110001_0101011110110011"; -- -0.0431924045911351
	pesos_i(74) := b"0000000000000000_0000000000000000_0000000010000000_1010110000010000"; -- 0.0019633806841574675
	pesos_i(75) := b"0000000000000000_0000000000000000_0000111000101001_0001100111000110"; -- 0.055314646515159105
	pesos_i(76) := b"0000000000000000_0000000000000000_0000011001001100_1100001000111010"; -- 0.024608744774227614
	pesos_i(77) := b"0000000000000000_0000000000000000_0010100111110011_1100110001010111"; -- 0.1638763153978544
	pesos_i(78) := b"1111111111111111_1111111111111111_1101101101000110_0010110011110110"; -- -0.14346045489557732
	pesos_i(79) := b"0000000000000000_0000000000000000_0010110110010011_1001000101110101"; -- 0.17803296199465773
	pesos_i(80) := b"0000000000000000_0000000000000000_0010100100001000_1100100010111111"; -- 0.16029028571023912
	pesos_i(81) := b"1111111111111111_1111111111111111_1111010101010011_1100111001010110"; -- -0.04168997195958285
	pesos_i(82) := b"1111111111111111_1111111111111111_1111101010100110_0001000011111111"; -- -0.020903528085492007
	pesos_i(83) := b"0000000000000000_0000000000000000_0010000000111110_0100111011101100"; -- 0.12595074913027848
	pesos_i(84) := b"0000000000000000_0000000000000000_0010011110000101_1010101111000001"; -- 0.15438340631795078
	pesos_i(85) := b"1111111111111111_1111111111111111_1111000000000001_1110110011001101"; -- -0.062470626684343944
	pesos_i(86) := b"1111111111111111_1111111111111111_1111010110100010_0101010101011101"; -- -0.04049173820280458
	pesos_i(87) := b"1111111111111111_1111111111111111_1111010011011000_0011111101100001"; -- -0.0435753237931035
	pesos_i(88) := b"0000000000000000_0000000000000000_0001111011110111_0011111100001110"; -- 0.12096017927647501
	pesos_i(89) := b"0000000000000000_0000000000000000_0000010101010111_1010010011010101"; -- 0.02086858942388589
	pesos_i(90) := b"0000000000000000_0000000000000000_0001011111011110_0110110011101000"; -- 0.09323769251181796
	pesos_i(91) := b"0000000000000000_0000000000000000_0001111010111100_1011000001100011"; -- 0.12006666569614405
	pesos_i(92) := b"0000000000000000_0000000000000000_0000101100110000_0001001010010100"; -- 0.043702279286314594
	pesos_i(93) := b"1111111111111111_1111111111111111_1111111100010001_0110001000000001"; -- -0.003641009147561658
	pesos_i(94) := b"1111111111111111_1111111111111111_1111001111101011_1000101100010110"; -- -0.04718714435097432
	pesos_i(95) := b"0000000000000000_0000000000000000_0001101111011011_0110111100110011"; -- 0.10881705275710318
	pesos_i(96) := b"0000000000000000_0000000000000000_0011000011010000_0110011011010100"; -- 0.19067995710815927
	pesos_i(97) := b"1111111111111111_1111111111111111_1111000101111111_1101110100110011"; -- -0.05664269936169092
	pesos_i(98) := b"0000000000000000_0000000000000000_0010110111001111_1110011011111001"; -- 0.17895358638867692
	pesos_i(99) := b"1111111111111111_1111111111111111_1110100111010111_0011101001110011"; -- -0.086559626414586
	pesos_i(100) := b"0000000000000000_0000000000000000_0011010010000100_0101011010100001"; -- 0.20514432353739098
	pesos_i(101) := b"0000000000000000_0000000000000000_0010100110001111_0001000111111110"; -- 0.16233932926290007
	pesos_i(102) := b"0000000000000000_0000000000000000_0010110111011110_0100111010001010"; -- 0.17917338241758798
	pesos_i(103) := b"0000000000000000_0000000000000000_0000101011000011_0001101001101101"; -- 0.04203953893889788
	pesos_i(104) := b"0000000000000000_0000000000000000_0000010001011000_0010010101010111"; -- 0.016969998968789708
	pesos_i(105) := b"0000000000000000_0000000000000000_0010000110000110_1101001101010100"; -- 0.13096352392176056
	pesos_i(106) := b"0000000000000000_0000000000000000_0010011000110110_1111111000110110"; -- 0.14927662679394
	pesos_i(107) := b"0000000000000000_0000000000000000_0001010011110101_1110011110011100"; -- 0.08187720838803118
	pesos_i(108) := b"0000000000000000_0000000000000000_0010001101010100_0000111100100001"; -- 0.13800139012366322
	pesos_i(109) := b"0000000000000000_0000000000000000_0010011010011101_1000001011101010"; -- 0.15084093297609982
	pesos_i(110) := b"0000000000000000_0000000000000000_0000111000011101_1101111000110110"; -- 0.05514324968223026
	pesos_i(111) := b"1111111111111111_1111111111111111_1110010110100110_0110110001011011"; -- -0.10292933241590525
	pesos_i(112) := b"1111111111111111_1111111111111111_1111010000001111_1010110100101101"; -- -0.046635796170669715
	pesos_i(113) := b"0000000000000000_0000000000000000_0000111110111110_1000100111100100"; -- 0.061501138841832385
	pesos_i(114) := b"0000000000000000_0000000000000000_0010000000011011_0011110000111000"; -- 0.12541557662635452
	pesos_i(115) := b"0000000000000000_0000000000000000_0001110000101011_0011011111111010"; -- 0.11003446428676018
	pesos_i(116) := b"0000000000000000_0000000000000000_0010001001101101_1100110101011010"; -- 0.13448794788003512
	pesos_i(117) := b"1111111111111111_1111111111111111_1111001011100100_0010111001011110"; -- -0.051205732368351915
	pesos_i(118) := b"0000000000000000_0000000000000000_0000110011000000_1111101111100100"; -- 0.049819701363922685
	pesos_i(119) := b"0000000000000000_0000000000000000_0001111000000110_1010110001101010"; -- 0.11728932938353392
	pesos_i(120) := b"0000000000000000_0000000000000000_0001000010100110_1001010011000010"; -- 0.06504182572387802
	pesos_i(121) := b"1111111111111111_1111111111111111_1111101100101000_1100011100111101"; -- -0.018909022956747373
	pesos_i(122) := b"0000000000000000_0000000000000000_0010010001110011_1011011000110111"; -- 0.14239062155868276
	pesos_i(123) := b"0000000000000000_0000000000000000_0010101101010100_0010111001001000"; -- 0.1692532469044265
	pesos_i(124) := b"0000000000000000_0000000000000000_0001111000100001_0100010010010110"; -- 0.1176951281704944
	pesos_i(125) := b"1111111111111111_1111111111111111_1100111100010000_0000001011100100"; -- -0.19116193719390234
	pesos_i(126) := b"0000000000000000_0000000000000000_0000101100001001_1110100110001110"; -- 0.04311999999047865
	pesos_i(127) := b"1111111111111111_1111111111111111_1101100101111000_0110101100010101"; -- -0.15050631272970957
	pesos_i(128) := b"1111111111111111_1111111111111111_1111001011011001_0111100011001001"; -- -0.051369143518728906
	pesos_i(129) := b"0000000000000000_0000000000000000_0001001101110100_1110110000011010"; -- 0.07600284233039038
	pesos_i(130) := b"1111111111111111_1111111111111111_1101011111111111_0100000100011101"; -- -0.15626137782752408
	pesos_i(131) := b"0000000000000000_0000000000000000_0000110110011011_0011101011000101"; -- 0.05314986533040247
	pesos_i(132) := b"0000000000000000_0000000000000000_0001010110000110_1101100110110111"; -- 0.08408890465611753
	pesos_i(133) := b"0000000000000000_0000000000000000_0000101111001000_0000011001111101"; -- 0.0460208945434132
	pesos_i(134) := b"1111111111111111_1111111111111111_1101111101110001_1100101000011100"; -- -0.12716996007696202
	pesos_i(135) := b"1111111111111111_1111111111111111_1111001010111000_0001110101100011"; -- -0.051878131204544146
	pesos_i(136) := b"0000000000000000_0000000000000000_0010010101111111_1011111101100001"; -- 0.1464805232688651
	pesos_i(137) := b"0000000000000000_0000000000000000_0000110011000110_0000010111000010"; -- 0.04989658335812852
	pesos_i(138) := b"1111111111111111_1111111111111111_1111000000011110_0111111111110001"; -- -0.06203461052463575
	pesos_i(139) := b"0000000000000000_0000000000000000_0010110010010101_1001100101101100"; -- 0.1741577042371221
	pesos_i(140) := b"0000000000000000_0000000000000000_0000100011011110_0000001111011110"; -- 0.0346376816223031
	pesos_i(141) := b"0000000000000000_0000000000000000_0010001111000001_1010001001101111"; -- 0.13967337799155785
	pesos_i(142) := b"0000000000000000_0000000000000000_0001000111001011_1111000001110111"; -- 0.06951811692760329
	pesos_i(143) := b"1111111111111111_1111111111111111_1101000001110001_1110001101111010"; -- -0.1857621980694744
	pesos_i(144) := b"1111111111111111_1111111111111111_1110101010001111_0001001101110100"; -- -0.08375433365594655
	pesos_i(145) := b"0000000000000000_0000000000000000_0001011111110100_0010100101001011"; -- 0.0935693557027641
	pesos_i(146) := b"0000000000000000_0000000000000000_0000110110111000_0101111111100001"; -- 0.05359458206819538
	pesos_i(147) := b"1111111111111111_1111111111111111_1111011110011110_1101011000110000"; -- -0.03273259465151216
	pesos_i(148) := b"0000000000000000_0000000000000000_0011100001100001_1010000001010010"; -- 0.22023965843597104
	pesos_i(149) := b"0000000000000000_0000000000000000_0001101110000000_1101010100011111"; -- 0.10743457800455168
	pesos_i(150) := b"1111111111111111_1111111111111111_1111001101101010_0001000010011011"; -- -0.04916282870456059
	pesos_i(151) := b"1111111111111111_1111111111111111_1110101110101010_0010010000111010"; -- -0.07943509663724851
	pesos_i(152) := b"0000000000000000_0000000000000000_0010100000010001_1111101100111001"; -- 0.1565243734503522
	pesos_i(153) := b"1111111111111111_1111111111111111_1100111111111011_1000000011001100"; -- -0.1875686170951205
	pesos_i(154) := b"0000000000000000_0000000000000000_0001010001011110_1010111000101011"; -- 0.07956970743295955
	pesos_i(155) := b"0000000000000000_0000000000000000_0001101010100001_0001001011010010"; -- 0.1040202867362388
	pesos_i(156) := b"0000000000000000_0000000000000000_0101000000010111_0100100110110001"; -- 0.31285534446820723
	pesos_i(157) := b"0000000000000000_0000000000000000_0010101011010111_0010111110100010"; -- 0.16734597867977286
	pesos_i(158) := b"0000000000000000_0000000000000000_0000111110111100_0000100000101010"; -- 0.06146288886203145
	pesos_i(159) := b"1111111111111111_1111111111111111_1111110001111111_1110000000111100"; -- -0.013673768353132902
	pesos_i(160) := b"1111111111111111_1111111111111111_1101001110100100_0110000001111101"; -- -0.17327305750701483
	pesos_i(161) := b"1111111111111111_1111111111111111_1110000111100110_1001011111010101"; -- -0.11757517866377419
	pesos_i(162) := b"0000000000000000_0000000000000000_0001010111011100_1111111110010111"; -- 0.08540341792614023
	pesos_i(163) := b"0000000000000000_0000000000000000_0001110011111101_1001111000001010"; -- 0.11324489338094942
	pesos_i(164) := b"0000000000000000_0000000000000000_0010001010011110_1100110111000001"; -- 0.13523565255177816
	pesos_i(165) := b"1111111111111111_1111111111111111_1110100101100111_1111001100101100"; -- -0.08825760052214686
	pesos_i(166) := b"1111111111111111_1111111111111111_1101000100011011_1000110010010011"; -- -0.18317338377365122
	pesos_i(167) := b"1111111111111111_1111111111111111_1111010010111000_1010100001111011"; -- -0.04405734065704518
	pesos_i(168) := b"0000000000000000_0000000000000000_0000001010110010_0100100010110001"; -- 0.010532897102453588
	pesos_i(169) := b"0000000000000000_0000000000000000_0001011101100010_1111111101001100"; -- 0.09135432817858757
	pesos_i(170) := b"1111111111111111_1111111111111111_1110001000001101_0000001001110101"; -- -0.11698898918501931
	pesos_i(171) := b"0000000000000000_0000000000000000_0001000111010000_1110001101000010"; -- 0.06959362364718566
	pesos_i(172) := b"1111111111111111_1111111111111111_1111010100110001_0001001000111011"; -- -0.042219982661268744
	pesos_i(173) := b"0000000000000000_0000000000000000_0001101010101010_1111001101101110"; -- 0.10417100360169765
	pesos_i(174) := b"0000000000000000_0000000000000000_0000001110011011_1100011110010110"; -- 0.014095758559911575
	pesos_i(175) := b"0000000000000000_0000000000000000_0001101010111101_0000100101000011"; -- 0.10444696325702071
	pesos_i(176) := b"0000000000000000_0000000000000000_0001010111010011_0101011100100000"; -- 0.08525604761165721
	pesos_i(177) := b"1111111111111111_1111111111111111_1110001101100001_0011000010100001"; -- -0.11179824904070526
	pesos_i(178) := b"0000000000000000_0000000000000000_0001011010100010_1000001011100000"; -- 0.08841722448163254
	pesos_i(179) := b"0000000000000000_0000000000000000_0000100000111100_1001000100100011"; -- 0.03217417819922514
	pesos_i(180) := b"1111111111111111_1111111111111111_1111101111001001_1101101101101000"; -- -0.01645115570446645
	pesos_i(181) := b"1111111111111111_1111111111111111_1110001101010001_1111000011011010"; -- -0.11203093211783961
	pesos_i(182) := b"1111111111111111_1111111111111111_1101011011110111_1001011100110010"; -- -0.16028456708174238
	pesos_i(183) := b"0000000000000000_0000000000000000_0010000010111000_1101110001100011"; -- 0.1278207531803109
	pesos_i(184) := b"1111111111111111_1111111111111111_1111001111111110_1110000111101110"; -- -0.04689205120723
	pesos_i(185) := b"0000000000000000_0000000000000000_0010101100011011_1111100001100000"; -- 0.16839554163113066
	pesos_i(186) := b"0000000000000000_0000000000000000_0010000010110000_1100011001101111"; -- 0.12769737445363086
	pesos_i(187) := b"1111111111111111_1111111111111111_1110100101001000_0101100111110110"; -- -0.08873975507122983
	pesos_i(188) := b"1111111111111111_1111111111111111_1111000101111101_0100000000111010"; -- -0.05668257318516464
	pesos_i(189) := b"0000000000000000_0000000000000000_0000111000110011_0111010111100110"; -- 0.05547272544296984
	pesos_i(190) := b"0000000000000000_0000000000000000_0000100010001011_0110000010000111"; -- 0.03337672515566613
	pesos_i(191) := b"0000000000000000_0000000000000000_0000011101000011_0110000000011111"; -- 0.028371818105426584
	pesos_i(192) := b"0000000000000000_0000000000000000_0010100011001101_0100101000011011"; -- 0.15938246879183224
	pesos_i(193) := b"0000000000000000_0000000000000000_0001011101111011_1110010010100001"; -- 0.09173420835699407
	pesos_i(194) := b"0000000000000000_0000000000000000_0010110000111000_1000101000111111"; -- 0.17273773224060107
	pesos_i(195) := b"0000000000000000_0000000000000000_0000101101110011_0110001000000010"; -- 0.04472935252255246
	pesos_i(196) := b"0000000000000000_0000000000000000_0010011010011100_0001111110000110"; -- 0.1508197499237705
	pesos_i(197) := b"0000000000000000_0000000000000000_0000111000101011_0010011110110111"; -- 0.05534599512005403
	pesos_i(198) := b"0000000000000000_0000000000000000_0001100001011110_0100111010011100"; -- 0.09518901154059245
	pesos_i(199) := b"1111111111111111_1111111111111111_1110100011101110_1010011000000111"; -- -0.09010851229835498
	pesos_i(200) := b"0000000000000000_0000000000000000_0000111011011111_0111001000110101"; -- 0.05809701717213785
	pesos_i(201) := b"0000000000000000_0000000000000000_0001101100100010_1011001011000100"; -- 0.10599820411320848
	pesos_i(202) := b"0000000000000000_0000000000000000_0010010001111001_0111100110100000"; -- 0.14247856287213895
	pesos_i(203) := b"1111111111111111_1111111111111111_1111011010011011_1001111110101011"; -- -0.036687870831040956
	pesos_i(204) := b"1111111111111111_1111111111111111_1110111110111011_0010111110010100"; -- -0.06355002062867614
	pesos_i(205) := b"1111111111111111_1111111111111111_1101001001110101_1101111010011101"; -- -0.1778889529558613
	pesos_i(206) := b"1111111111111111_1111111111111111_1101111011001010_0011011110100000"; -- -0.12972690921450541
	pesos_i(207) := b"0000000000000000_0000000000000000_0010101100001101_1110010101001011"; -- 0.16818078121362567
	pesos_i(208) := b"1111111111111111_1111111111111111_1111001001011001_1000110110000111"; -- -0.05332103215731903
	pesos_i(209) := b"1111111111111111_1111111111111111_1101010110100101_1110011111000110"; -- -0.16543723503407315
	pesos_i(210) := b"1111111111111111_1111111111111111_1110010110000010_0001100110001011"; -- -0.10348358500281128
	pesos_i(211) := b"1111111111111111_1111111111111111_1101001000101001_0111100100110010"; -- -0.17905466577525828
	pesos_i(212) := b"0000000000000000_0000000000000000_0001110110000111_1011101101111100"; -- 0.11535236143191241
	pesos_i(213) := b"0000000000000000_0000000000000000_0010110001000101_0001000011011101"; -- 0.17292886160986973
	pesos_i(214) := b"1111111111111111_1111111111111111_1111010101101011_1111010100110100"; -- -0.04132144440621194
	pesos_i(215) := b"0000000000000000_0000000000000000_0010010101010100_1010011010110000"; -- 0.14582292374113345
	pesos_i(216) := b"0000000000000000_0000000000000000_0001000010010100_0001000110101001"; -- 0.06475935341189083
	pesos_i(217) := b"1111111111111111_1111111111111111_1101111000111111_1100100111001000"; -- -0.1318391692906531
	pesos_i(218) := b"1111111111111111_1111111111111111_1100100101100101_1011110011111111"; -- -0.2132913473497171
	pesos_i(219) := b"0000000000000000_0000000000000000_0001001101100101_0010110100111001"; -- 0.07576258319664586
	pesos_i(220) := b"0000000000000000_0000000000000000_0001110101001000_0111111101001111"; -- 0.11438747094254706
	pesos_i(221) := b"0000000000000000_0000000000000000_0001001000011110_1000101100011101"; -- 0.07077855535905375
	pesos_i(222) := b"1111111111111111_1111111111111111_1110111000110011_1011001101101101"; -- -0.06952360713893867
	pesos_i(223) := b"0000000000000000_0000000000000000_0000110100001011_0011101010100100"; -- 0.050952591845893784
	pesos_i(224) := b"1111111111111111_1111111111111111_1111000100010100_1011111001111001"; -- -0.05827722124880869
	pesos_i(225) := b"0000000000000000_0000000000000000_0010101110001011_1111101110100101"; -- 0.17010472084279699
	pesos_i(226) := b"1111111111111111_1111111111111111_1111010000110101_0111000010011111"; -- -0.04605957145240364
	pesos_i(227) := b"1111111111111111_1111111111111111_1101010010110010_1101110101111100"; -- -0.16914573408965078
	pesos_i(228) := b"1111111111111111_1111111111111111_1100101110111010_0111110000010010"; -- -0.20418572011336292
	pesos_i(229) := b"0000000000000000_0000000000000000_0001111111010000_1100000101111100"; -- 0.12427911078719492
	pesos_i(230) := b"1111111111111111_1111111111111111_1101011000011111_0001001011000111"; -- -0.16358835837308475
	pesos_i(231) := b"1111111111111111_1111111111111111_1110010000001111_0011010011001101"; -- -0.10914297089991663
	pesos_i(232) := b"0000000000000000_0000000000000000_0010011100010010_1110100000010101"; -- 0.15263224146032497
	pesos_i(233) := b"1111111111111111_1111111111111111_1101011110100001_0111010011011111"; -- -0.15769261888123073
	pesos_i(234) := b"0000000000000000_0000000000000000_0010010100111010_0110010001101111"; -- 0.145422245962118
	pesos_i(235) := b"0000000000000000_0000000000000000_0010011010111101_1011111111100110"; -- 0.1513328492714912
	pesos_i(236) := b"0000000000000000_0000000000000000_0000100110111110_0011001101111111"; -- 0.038058489231624706
	pesos_i(237) := b"0000000000000000_0000000000000000_0000111000010111_0101011110000110"; -- 0.05504366904178879
	pesos_i(238) := b"1111111111111111_1111111111111111_1101001000100111_0110011001001010"; -- -0.17908631023842048
	pesos_i(239) := b"0000000000000000_0000000000000000_0010010101001101_1101111001100010"; -- 0.145719431762318
	pesos_i(240) := b"1111111111111111_1111111111111111_1110101100010111_0011000011000111"; -- -0.08167739046053886
	pesos_i(241) := b"0000000000000000_0000000000000000_0010011101101111_0011011000000010"; -- 0.15404069473576146
	pesos_i(242) := b"1111111111111111_1111111111111111_1101100100101011_1111100001100100"; -- -0.15167281679749745
	pesos_i(243) := b"0000000000000000_0000000000000000_0001000001110100_0011001111000110"; -- 0.06427310551781444
	pesos_i(244) := b"1111111111111111_1111111111111111_1111001001100101_0111100001011101"; -- -0.053139188020565206
	pesos_i(245) := b"1111111111111111_1111111111111111_1111100000100111_0010110101011010"; -- -0.030652204105403164
	pesos_i(246) := b"0000000000000000_0000000000000000_0001111001100110_0101111000111000"; -- 0.11874951241502185
	pesos_i(247) := b"0000000000000000_0000000000000000_0010001010110000_0010111100000001"; -- 0.1355008485816227
	pesos_i(248) := b"1111111111111111_1111111111111111_1110000100111110_1111011011111001"; -- -0.12013298443187304
	pesos_i(249) := b"1111111111111111_1111111111111111_1110011111101011_1000110100100111"; -- -0.094062021196519
	pesos_i(250) := b"0000000000000000_0000000000000000_0001011001001011_0001100101111110"; -- 0.08708342874666915
	pesos_i(251) := b"0000000000000000_0000000000000000_0000101011110110_0100010010111101"; -- 0.04282025932874447
	pesos_i(252) := b"1111111111111111_1111111111111111_1111000110000001_1110010100111100"; -- -0.056611702773037405
	pesos_i(253) := b"1111111111111111_1111111111111111_1110010010001010_0010110100100000"; -- -0.10726659751816246
	pesos_i(254) := b"0000000000000000_0000000000000000_0010000100101100_0110111111011110"; -- 0.12958430440837443
	pesos_i(255) := b"0000000000000000_0000000000000000_0001000101110101_0111100010001001"; -- 0.06819871272234662
	pesos_i(256) := b"0000000000000000_0000000000000000_0011001011010001_1001100100101110"; -- 0.1985107170670049
	pesos_i(257) := b"1111111111111111_1111111111111111_1101011111010011_0111000111001110"; -- -0.15692986217671412
	pesos_i(258) := b"1111111111111111_1111111111111111_1101011010011111_1000001101101000"; -- -0.16162852002507308
	pesos_i(259) := b"1111111111111111_1111111111111111_1100101110111010_1110111111101000"; -- -0.20417881565933613
	pesos_i(260) := b"1111111111111111_1111111111111111_1110110100101110_0110000001000011"; -- -0.07351110810853022
	pesos_i(261) := b"1111111111111111_1111111111111111_1110010110001000_1110001011000111"; -- -0.10338003759615219
	pesos_i(262) := b"1111111111111111_1111111111111111_1101101101101010_1010011000110100"; -- -0.14290391189828167
	pesos_i(263) := b"0000000000000000_0000000000000000_0010110000000111_0100001010000110"; -- 0.17198577664216497
	pesos_i(264) := b"0000000000000000_0000000000000000_0000000000110101_0001000110010000"; -- 0.000809762580783872
	pesos_i(265) := b"1111111111111111_1111111111111111_1111101001110111_0101110111110111"; -- -0.021616103345549528
	pesos_i(266) := b"1111111111111111_1111111111111111_1101000101110110_1110111100001010"; -- -0.18177896501193072
	pesos_i(267) := b"1111111111111111_1111111111111111_1111100010111101_0110000101011100"; -- -0.028360285825877737
	pesos_i(268) := b"0000000000000000_0000000000000000_0001111011101111_1110110011111000"; -- 0.12084847492851532
	pesos_i(269) := b"1111111111111111_1111111111111111_1100100101111110_1000011011010001"; -- -0.21291310681647857
	pesos_i(270) := b"1111111111111111_1111111111111111_1110001011001100_0110000010011100"; -- -0.11406894872454694
	pesos_i(271) := b"1111111111111111_1111111111111111_1111011111010010_1011110101011100"; -- -0.03194061768333322
	pesos_i(272) := b"0000000000000000_0000000000000000_0000010001010111_0000101101100110"; -- 0.01695319411915222
	pesos_i(273) := b"0000000000000000_0000000000000000_0000111011000001_0100110011010110"; -- 0.057637026146141905
	pesos_i(274) := b"0000000000000000_0000000000000000_0001011111000000_0011110100011001"; -- 0.0927770792790976
	pesos_i(275) := b"1111111111111111_1111111111111111_1111000000101110_1100001010000001"; -- -0.061786502323798856
	pesos_i(276) := b"0000000000000000_0000000000000000_0010011001011010_1100100100011110"; -- 0.14982277852883033
	pesos_i(277) := b"0000000000000000_0000000000000000_0001010010001011_1000001011010100"; -- 0.08025376975585524
	pesos_i(278) := b"0000000000000000_0000000000000000_0000101100100001_0111001110111000"; -- 0.04347918750288701
	pesos_i(279) := b"0000000000000000_0000000000000000_0010101011100111_0001100100111011"; -- 0.16758878418792575
	pesos_i(280) := b"1111111111111111_1111111111111111_1111111111100010_1011001101000011"; -- -0.0004470788538627615
	pesos_i(281) := b"1111111111111111_1111111111111111_1101111111010110_0101101101111110"; -- -0.12563541575076875
	pesos_i(282) := b"0000000000000000_0000000000000000_0000111100110111_1010000001101101"; -- 0.0594425454699179
	pesos_i(283) := b"1111111111111111_1111111111111111_1111100101001001_1101111110011001"; -- -0.026216530962166504
	pesos_i(284) := b"1111111111111111_1111111111111111_1111101110001100_0000110111111010"; -- -0.017394186351501816
	pesos_i(285) := b"1111111111111111_1111111111111111_1111111000101010_1110011110001100"; -- -0.007157829680034682
	pesos_i(286) := b"0000000000000000_0000000000000000_0001110010011010_1110001000100110"; -- 0.11173833312189756
	pesos_i(287) := b"1111111111111111_1111111111111111_1101110100111001_1001011111110101"; -- -0.13583994178359812
	pesos_i(288) := b"0000000000000000_0000000000000000_0000100111011101_1001101001000000"; -- 0.03853763632942498
	pesos_i(289) := b"1111111111111111_1111111111111111_1111001111000001_1001110011010100"; -- -0.047826956091447645
	pesos_i(290) := b"0000000000000000_0000000000000000_0001011010010100_1110010100101111"; -- 0.08820946113747108
	pesos_i(291) := b"0000000000000000_0000000000000000_0000011000010011_0011010010000111"; -- 0.02373054790850648
	pesos_i(292) := b"0000000000000000_0000000000000000_0000100100011110_0001001010000010"; -- 0.035615116787761206
	pesos_i(293) := b"1111111111111111_1111111111111111_1101000010000111_1101100101000010"; -- -0.18542711400134484
	pesos_i(294) := b"0000000000000000_0000000000000000_0001100011100110_1000000010001000"; -- 0.09726718247737165
	pesos_i(295) := b"0000000000000000_0000000000000000_0000111001011100_1011111010011011"; -- 0.05610266962557008
	pesos_i(296) := b"1111111111111111_1111111111111111_1111001001011010_0010000010011101"; -- -0.05331226512167092
	pesos_i(297) := b"1111111111111111_1111111111111111_1110000111100011_1111011100100001"; -- -0.11761527477010278
	pesos_i(298) := b"1111111111111111_1111111111111111_1111001100010001_1001101000100101"; -- -0.05051266286115832
	pesos_i(299) := b"1111111111111111_1111111111111111_1111100001100010_1100111101010011"; -- -0.02974228120861474
	pesos_i(300) := b"1111111111111111_1111111111111111_1110101010100100_1101001101010001"; -- -0.0834224631963235
	pesos_i(301) := b"1111111111111111_1111111111111111_1110000111010000_0001110000101110"; -- -0.11791824228191468
	pesos_i(302) := b"0000000000000000_0000000000000000_0001000010000110_1010010011101100"; -- 0.06455450779815136
	pesos_i(303) := b"0000000000000000_0000000000000000_0010001100100001_0100101110100000"; -- 0.13722679754699324
	pesos_i(304) := b"0000000000000000_0000000000000000_0010001110101001_1001000001000110"; -- 0.13930608461693306
	pesos_i(305) := b"1111111111111111_1111111111111111_1110110110110111_1100111000111110"; -- -0.07141409857618987
	pesos_i(306) := b"1111111111111111_1111111111111111_1111100110111011_1100000101001100"; -- -0.024478835009813123
	pesos_i(307) := b"1111111111111111_1111111111111111_1111001111010000_0011001101110110"; -- -0.04760435451515926
	pesos_i(308) := b"1111111111111111_1111111111111111_1111011011001101_0101110000101100"; -- -0.035928954380227474
	pesos_i(309) := b"1111111111111111_1111111111111111_1111011111101011_1001101110110111"; -- -0.03156115319196052
	pesos_i(310) := b"0000000000000000_0000000000000000_0001111100101101_1110001110001010"; -- 0.12179395778953149
	pesos_i(311) := b"0000000000000000_0000000000000000_0001100011011101_1101111000000101"; -- 0.09713542579107437
	pesos_i(312) := b"1111111111111111_1111111111111111_1110100111110101_1111001101000011"; -- -0.08609084715241028
	pesos_i(313) := b"1111111111111111_1111111111111111_1110100111111001_1100011110110101"; -- -0.08603240811663405
	pesos_i(314) := b"1111111111111111_1111111111111111_1110011111100111_1100000110001101"; -- -0.09411993315905653
	pesos_i(315) := b"0000000000000000_0000000000000000_0000101000110110_1100100111001010"; -- 0.039898502136447626
	pesos_i(316) := b"1111111111111111_1111111111111111_1111110000001101_0101100100001010"; -- -0.015421328666609219
	pesos_i(317) := b"0000000000000000_0000000000000000_0000101000101001_1010000011011101"; -- 0.03969769845640898
	pesos_i(318) := b"0000000000000000_0000000000000000_0010001110101101_1101011101110110"; -- 0.13937136293991897
	pesos_i(319) := b"1111111111111111_1111111111111111_1111101101000101_1111101011010100"; -- -0.01846344293257573
	pesos_i(320) := b"0000000000000000_0000000000000000_0001000111110001_0000011001111101"; -- 0.07008400498816299
	pesos_i(321) := b"1111111111111111_1111111111111111_1101100000111100_0111101101111000"; -- -0.15532711330970664
	pesos_i(322) := b"1111111111111111_1111111111111111_1111110100101010_0000101110100101"; -- -0.01107718687583406
	pesos_i(323) := b"0000000000000000_0000000000000000_0000000100010000_1110111010111001"; -- 0.004164619492133201
	pesos_i(324) := b"0000000000000000_0000000000000000_0010100001100010_0011100010001100"; -- 0.15774873186278937
	pesos_i(325) := b"1111111111111111_1111111111111111_1110101111111111_1010111101000011"; -- -0.07812981238433479
	pesos_i(326) := b"0000000000000000_0000000000000000_0010000010000100_1110111101101100"; -- 0.12702843080644105
	pesos_i(327) := b"1111111111111111_1111111111111111_1111110100110111_1111001100011000"; -- -0.010865026974516795
	pesos_i(328) := b"0000000000000000_0000000000000000_0001011100000001_0111110001111010"; -- 0.08986642825973824
	pesos_i(329) := b"1111111111111111_1111111111111111_1110011001001001_0100110111011001"; -- -0.10044396840640937
	pesos_i(330) := b"0000000000000000_0000000000000000_0000101011101100_0001001111000101"; -- 0.04266475248205024
	pesos_i(331) := b"0000000000000000_0000000000000000_0010011001101101_0011010110001010"; -- 0.1501038991910391
	pesos_i(332) := b"0000000000000000_0000000000000000_0001010101101110_0101011011101011"; -- 0.08371489761356794
	pesos_i(333) := b"0000000000000000_0000000000000000_0001100010110000_1110100001110110"; -- 0.09644940252980203
	pesos_i(334) := b"0000000000000000_0000000000000000_0010000101000101_1000100110111001"; -- 0.12996731536986642
	pesos_i(335) := b"0000000000000000_0000000000000000_0010101101000001_0101001110101110"; -- 0.1689655590156828
	pesos_i(336) := b"0000000000000000_0000000000000000_0010001110000111_1100010111000011"; -- 0.13879047407596642
	pesos_i(337) := b"1111111111111111_1111111111111111_1101111011010001_0000111100110000"; -- -0.12962250788642582
	pesos_i(338) := b"1111111111111111_1111111111111111_1111100000100001_1001101100010001"; -- -0.030737217216770977
	pesos_i(339) := b"1111111111111111_1111111111111111_1111101111010110_1010000101110000"; -- -0.016256246629373465
	pesos_i(340) := b"1111111111111111_1111111111111111_1101100110001011_0110100001100101"; -- -0.15021655582675883
	pesos_i(341) := b"0000000000000000_0000000000000000_0000110000000011_0010011010001101"; -- 0.04692307423886525
	pesos_i(342) := b"0000000000000000_0000000000000000_0001110101011000_0001010101100101"; -- 0.11462529858956261
	pesos_i(343) := b"1111111111111111_1111111111111111_1111010010101111_0001101110110110"; -- -0.04420306012112959
	pesos_i(344) := b"1111111111111111_1111111111111111_1111110110101110_0011101111110110"; -- -0.009060146767401524
	pesos_i(345) := b"1111111111111111_1111111111111111_1110011001000101_1101101001000011"; -- -0.10049663422108672
	pesos_i(346) := b"0000000000000000_0000000000000000_0010001100100001_1010001110011001"; -- 0.13723204122870378
	pesos_i(347) := b"1111111111111111_1111111111111111_1111100110001011_0001101001001100"; -- -0.025221211001867458
	pesos_i(348) := b"0000000000000000_0000000000000000_0010010000001101_1001011011111000"; -- 0.14083236265103002
	pesos_i(349) := b"0000000000000000_0000000000000000_0001010001000010_1110100001100010"; -- 0.07914593124062295
	pesos_i(350) := b"1111111111111111_1111111111111111_1110100111100110_1101000111010111"; -- -0.08632172106829224
	pesos_i(351) := b"0000000000000000_0000000000000000_0001001001011100_0101010111100101"; -- 0.07172142819100513
	pesos_i(352) := b"0000000000000000_0000000000000000_0001101010011001_0000110101011011"; -- 0.10389789070585949
	pesos_i(353) := b"0000000000000000_0000000000000000_0001111010111001_0100100110011001"; -- 0.12001476284438649
	pesos_i(354) := b"0000000000000000_0000000000000000_0010010110011100_1011001001011100"; -- 0.14692225206668247
	pesos_i(355) := b"1111111111111111_1111111111111111_1111101011011101_1100100010111001"; -- -0.020053343572970603
	pesos_i(356) := b"1111111111111111_1111111111111111_1110111000011011_0011000001100100"; -- -0.0698976283494075
	pesos_i(357) := b"1111111111111111_1111111111111111_1101111001000101_0111111010000010"; -- -0.13175210299401602
	pesos_i(358) := b"0000000000000000_0000000000000000_0000001000111111_0001110001001010"; -- 0.008775489802126167
	pesos_i(359) := b"0000000000000000_0000000000000000_0010010101010011_1111011010011110"; -- 0.14581242892786442
	pesos_i(360) := b"1111111111111111_1111111111111111_1110011000010100_0111101100100100"; -- -0.10124998450740327
	pesos_i(361) := b"1111111111111111_1111111111111111_1111001010110100_1101110010111111"; -- -0.05192776048864982
	pesos_i(362) := b"0000000000000000_0000000000000000_0001110010101100_1110010111110101"; -- 0.11201321829104353
	pesos_i(363) := b"0000000000000000_0000000000000000_0010100001110111_1101101001101010"; -- 0.15807881436247456
	pesos_i(364) := b"1111111111111111_1111111111111111_1100101100100101_1101100001010101"; -- -0.20645378040373907
	pesos_i(365) := b"0000000000000000_0000000000000000_0011000000101001_1001010011110010"; -- 0.18813448814859476
	pesos_i(366) := b"1111111111111111_1111111111111111_1110110000000110_0111010110011111"; -- -0.07802643639559767
	pesos_i(367) := b"1111111111111111_1111111111111111_1101111111011011_0001011001000000"; -- -0.12556324909007294
	pesos_i(368) := b"0000000000000000_0000000000000000_0001101010101011_0011111011010110"; -- 0.10417549829885035
	pesos_i(369) := b"1111111111111111_1111111111111111_1111011100011000_0011010000100100"; -- -0.034786931233571135
	pesos_i(370) := b"1111111111111111_1111111111111111_1101101100100111_0100101110100001"; -- -0.14393164928373609
	pesos_i(371) := b"0000000000000000_0000000000000000_0010000100101000_0010000001010010"; -- 0.12951852804182773
	pesos_i(372) := b"0000000000000000_0000000000000000_0001000010100111_0111111101110111"; -- 0.06505581521928072
	pesos_i(373) := b"1111111111111111_1111111111111111_1111100101101011_0001001001101100"; -- -0.025709961573974326
	pesos_i(374) := b"0000000000000000_0000000000000000_0001101000101011_1110100000101000"; -- 0.10223246563193884
	pesos_i(375) := b"1111111111111111_1111111111111111_1101110000001100_1111001111001000"; -- -0.1404273639906977
	pesos_i(376) := b"1111111111111111_1111111111111111_1110100001101110_1011001010100011"; -- -0.09206088561706381
	pesos_i(377) := b"1111111111111111_1111111111111111_1110101110100001_1100001111100001"; -- -0.0795629097578375
	pesos_i(378) := b"0000000000000000_0000000000000000_0010000011001110_0010110011010111"; -- 0.12814598318754922
	pesos_i(379) := b"1111111111111111_1111111111111111_1101001101011001_1001110111010110"; -- -0.1744138099892435
	pesos_i(380) := b"1111111111111111_1111111111111111_1111000100000110_1001001001011110"; -- -0.05849347312771237
	pesos_i(381) := b"1111111111111111_1111111111111111_1111001100100100_0111001001001101"; -- -0.050225120634772816
	pesos_i(382) := b"1111111111111111_1111111111111111_1100111010010000_1110111111111100"; -- -0.19310093009589926
	pesos_i(383) := b"0000000000000000_0000000000000000_0000110001001101_1111110101100101"; -- 0.04806503016412514
	pesos_i(384) := b"1111111111111111_1111111111111111_1110000101100010_0011100111010011"; -- -0.11959494215972961
	pesos_i(385) := b"0000000000000000_0000000000000000_0001110001111001_1110000010010001"; -- 0.1112346986193767
	pesos_i(386) := b"0000000000000000_0000000000000000_0000110101001101_0110001001010010"; -- 0.05196203699461965
	pesos_i(387) := b"0000000000000000_0000000000000000_0011000110101111_1110110010111011"; -- 0.19409064823924174
	pesos_i(388) := b"0000000000000000_0000000000000000_0000010011111100_0110010000110000"; -- 0.019476186425562814
	pesos_i(389) := b"0000000000000000_0000000000000000_0001010100010010_0011001001100010"; -- 0.08230891130898306
	pesos_i(390) := b"0000000000000000_0000000000000000_0001111000101010_1000010010011111"; -- 0.11783627389737732
	pesos_i(391) := b"1111111111111111_1111111111111111_1111010101000101_1100100010101001"; -- -0.04190393334966121
	pesos_i(392) := b"0000000000000000_0000000000000000_0000100101100110_1000101100011101"; -- 0.03672093818542159
	pesos_i(393) := b"1111111111111111_1111111111111111_1111100010011001_1100110000111110"; -- -0.02890323159227716
	pesos_i(394) := b"1111111111111111_1111111111111111_1110101101000110_0011101110100001"; -- -0.08095958052574877
	pesos_i(395) := b"0000000000000000_0000000000000000_0001000010111110_1111010110100001"; -- 0.06541381057410549
	pesos_i(396) := b"1111111111111111_1111111111111111_1111001111110011_0110101011100101"; -- -0.04706699275946899
	pesos_i(397) := b"1111111111111111_1111111111111111_1111011001010110_0000100100011000"; -- -0.0377497021759719
	pesos_i(398) := b"1111111111111111_1111111111111111_1111010011011001_0001011111001011"; -- -0.043562424531009974
	pesos_i(399) := b"1111111111111111_1111111111111111_1110001001101000_1001001101101111"; -- -0.11559179818867356
	pesos_i(400) := b"0000000000000000_0000000000000000_0010010110001010_0000101011000100"; -- 0.14663760463824072
	pesos_i(401) := b"1111111111111111_1111111111111111_1111101111000100_1001100110110001"; -- -0.016531366727970596
	pesos_i(402) := b"1111111111111111_1111111111111111_1110110011110001_1111010100111010"; -- -0.07443301524306338
	pesos_i(403) := b"1111111111111111_1111111111111111_1110010100110011_1111001010010011"; -- -0.10467609309961766
	pesos_i(404) := b"1111111111111111_1111111111111111_1111011110011001_0100111001111000"; -- -0.03281697825386537
	pesos_i(405) := b"0000000000000000_0000000000000000_0000000011001011_0010011000110110"; -- 0.003099811645480302
	pesos_i(406) := b"1111111111111111_1111111111111111_1111110010001011_0101011010111111"; -- -0.013498857805972176
	pesos_i(407) := b"0000000000000000_0000000000000000_0000010101001110_1100011110011101"; -- 0.020733333536874548
	pesos_i(408) := b"1111111111111111_1111111111111111_1110000001100110_0011110010101001"; -- -0.12343998778071194
	pesos_i(409) := b"0000000000000000_0000000000000000_0000010111001001_0011101011001100"; -- 0.022601771099462827
	pesos_i(410) := b"0000000000000000_0000000000000000_0010101001011100_1000010111111010"; -- 0.16547429415290954
	pesos_i(411) := b"1111111111111111_1111111111111111_1101000000101000_1010000010111010"; -- -0.18688006832298917
	pesos_i(412) := b"0000000000000000_0000000000000000_0010011101010111_1010111100101110"; -- 0.15368170616520976
	pesos_i(413) := b"0000000000000000_0000000000000000_0010101110100100_1111100000011101"; -- 0.1704859801880722
	pesos_i(414) := b"1111111111111111_1111111111111111_1110001101000110_0110100001111001"; -- -0.11220690764877915
	pesos_i(415) := b"1111111111111111_1111111111111111_1110010101010010_0100100010101001"; -- -0.1042131984977148
	pesos_i(416) := b"1111111111111111_1111111111111111_1110100000010111_1101100111001010"; -- -0.09338606671802283
	pesos_i(417) := b"0000000000000000_0000000000000000_0010001001110111_1010111111011011"; -- 0.13463877775972363
	pesos_i(418) := b"1111111111111111_1111111111111111_1110011110100111_1110000110001000"; -- -0.09509458959135132
	pesos_i(419) := b"1111111111111111_1111111111111111_1100110010110110_1101001110011110"; -- -0.20033528699390926
	pesos_i(420) := b"0000000000000000_0000000000000000_0010101111101111_1000010101101011"; -- 0.17162355285273215
	pesos_i(421) := b"0000000000000000_0000000000000000_0010101001000110_0011111110101010"; -- 0.1651344099286917
	pesos_i(422) := b"1111111111111111_1111111111111111_1110011011011000_1100000001111111"; -- -0.09825512793301687
	pesos_i(423) := b"1111111111111111_1111111111111111_1111011000010010_1100100010111001"; -- -0.03877587788625928
	pesos_i(424) := b"0000000000000000_0000000000000000_0000011011100100_0110111010101111"; -- 0.02692310127145961
	pesos_i(425) := b"1111111111111111_1111111111111111_1110111000110000_0110110101101011"; -- -0.06957355631388641
	pesos_i(426) := b"1111111111111111_1111111111111111_1101011000010000_1110100011001000"; -- -0.16380448456188396
	pesos_i(427) := b"1111111111111111_1111111111111111_1100100010111100_1011011001011111"; -- -0.21587047745491278
	pesos_i(428) := b"0000000000000000_0000000000000000_0010001101000110_1111000100001111"; -- 0.1378012333413001
	pesos_i(429) := b"1111111111111111_1111111111111111_1111001111011000_1011010011110000"; -- -0.047474566755532396
	pesos_i(430) := b"0000000000000000_0000000000000000_0000100111110000_1101111111010111"; -- 0.03883170134217115
	pesos_i(431) := b"1111111111111111_1111111111111111_1111110001111001_0101101110110100"; -- -0.013773220637446827
	pesos_i(432) := b"0000000000000000_0000000000000000_0001100111000100_1000010001000000"; -- 0.1006548553360368
	pesos_i(433) := b"0000000000000000_0000000000000000_0001010000000100_1110111010100010"; -- 0.07820025883663928
	pesos_i(434) := b"0000000000000000_0000000000000000_0000111001001011_0100100100111101"; -- 0.05583627446670845
	pesos_i(435) := b"0000000000000000_0000000000000000_0001101010000000_1001110011110011"; -- 0.10352497996469587
	pesos_i(436) := b"0000000000000000_0000000000000000_0000100100100100_1010101110000100"; -- 0.035715789638983024
	pesos_i(437) := b"0000000000000000_0000000000000000_0010100010000000_0000100100101010"; -- 0.1582036712187354
	pesos_i(438) := b"1111111111111111_1111111111111111_1110010001000010_1000010101000011"; -- -0.10835997694227327
	pesos_i(439) := b"1111111111111111_1111111111111111_1110011001110100_0011000000111001"; -- -0.09978960620292388
	pesos_i(440) := b"1111111111111111_1111111111111111_1101010101101001_0100100100111001"; -- -0.16636221262648854
	pesos_i(441) := b"0000000000000000_0000000000000000_0001100100000101_0011010011011101"; -- 0.09773569494174761
	pesos_i(442) := b"1111111111111111_1111111111111111_1101001010101001_1101110010100010"; -- -0.17709561393893852
	pesos_i(443) := b"0000000000000000_0000000000000000_0000100000111111_1010100011100110"; -- 0.03222137093683114
	pesos_i(444) := b"0000000000000000_0000000000000000_0000010111000100_0110100011001111"; -- 0.022528219690978558
	pesos_i(445) := b"1111111111111111_1111111111111111_1100101110110000_1001001011011111"; -- -0.2043369488788118
	pesos_i(446) := b"0000000000000000_0000000000000000_0010011100000000_1110011001010010"; -- 0.15235747827004253
	pesos_i(447) := b"0000000000000000_0000000000000000_0000100011011100_1101110101011000"; -- 0.03462012664394338
	pesos_i(448) := b"0000000000000000_0000000000000000_0001011001110000_1010010111101110"; -- 0.08765637448898275
	pesos_i(449) := b"1111111111111111_1111111111111111_1111100100001000_0100110111100011"; -- -0.027217037180305312
	pesos_i(450) := b"0000000000000000_0000000000000000_0001110100011010_1001111001100011"; -- 0.11368741913874797
	pesos_i(451) := b"0000000000000000_0000000000000000_0001110111100101_0001100001011101"; -- 0.11677696480251759
	pesos_i(452) := b"0000000000000000_0000000000000000_0001000110100010_1111000011100000"; -- 0.06889253118084626
	pesos_i(453) := b"1111111111111111_1111111111111111_1111010110101010_1010010101010001"; -- -0.040364902135172596
	pesos_i(454) := b"1111111111111111_1111111111111111_1101111111100011_0111111101000011"; -- -0.1254349194350405
	pesos_i(455) := b"0000000000000000_0000000000000000_0000110100101100_1100001011001101"; -- 0.05146424769783568
	pesos_i(456) := b"1111111111111111_1111111111111111_1110010000011001_0011110000001111"; -- -0.10898995046146294
	pesos_i(457) := b"0000000000000000_0000000000000000_0000101111110100_1000100000010111"; -- 0.046700006029509904
	pesos_i(458) := b"0000000000000000_0000000000000000_0010100101000011_1010010011010100"; -- 0.1611884133202473
	pesos_i(459) := b"0000000000000000_0000000000000000_0001100110001001_1011011011110110"; -- 0.0997576095193897
	pesos_i(460) := b"1111111111111111_1111111111111111_1110111001011110_1010011010011010"; -- -0.06886824364953009
	pesos_i(461) := b"1111111111111111_1111111111111111_1110110000010100_0000100001101100"; -- -0.07781932231105493
	pesos_i(462) := b"1111111111111111_1111111111111111_1110101011001011_1111001010011011"; -- -0.08282550547059445
	pesos_i(463) := b"1111111111111111_1111111111111111_1111001010010001_1010100110001111"; -- -0.05246486901654336
	pesos_i(464) := b"0000000000000000_0000000000000000_0001011100001110_0000101100000001"; -- 0.09005802892333611
	pesos_i(465) := b"0000000000000000_0000000000000000_0001010011011000_0001101000011011"; -- 0.0814224544852956
	pesos_i(466) := b"1111111111111111_1111111111111111_1111010010010111_0010111111010010"; -- -0.04456807254408274
	pesos_i(467) := b"0000000000000000_0000000000000000_0010110110001100_1000100110000101"; -- 0.17792567726657776
	pesos_i(468) := b"0000000000000000_0000000000000000_0001011000000001_0000011110111001"; -- 0.08595321918499199
	pesos_i(469) := b"1111111111111111_1111111111111111_1111100101111010_0101010111001100"; -- -0.025477063808960806
	pesos_i(470) := b"0000000000000000_0000000000000000_0001000000101101_0011111111111100"; -- 0.06319045924582554
	pesos_i(471) := b"0000000000000000_0000000000000000_0000110001110110_0001000110111110"; -- 0.048676594517722396
	pesos_i(472) := b"1111111111111111_1111111111111111_1110100111001001_0001010101111101"; -- -0.08677545256225652
	pesos_i(473) := b"0000000000000000_0000000000000000_0000100011111010_1010010100000100"; -- 0.035074533063280906
	pesos_i(474) := b"1111111111111111_1111111111111111_1101011100101011_0000101101100110"; -- -0.1594994427638578
	pesos_i(475) := b"0000000000000000_0000000000000000_0010111010110000_0000011010100001"; -- 0.1823734419460625
	pesos_i(476) := b"0000000000000000_0000000000000000_0001010001100011_1100111111111011"; -- 0.07964801662977046
	pesos_i(477) := b"0000000000000000_0000000000000000_0010011010000011_1110101110001101"; -- 0.15045044126689186
	pesos_i(478) := b"1111111111111111_1111111111111111_1101100011100010_0000111000010110"; -- -0.1528006741955907
	pesos_i(479) := b"0000000000000000_0000000000000000_0001111010111110_1000010000100000"; -- 0.12009454515425332
	pesos_i(480) := b"0000000000000000_0000000000000000_0010101000000001_1110111101101100"; -- 0.1640920294388532
	pesos_i(481) := b"1111111111111111_1111111111111111_1101011011001101_0100101100000111"; -- -0.16092997618157476
	pesos_i(482) := b"0000000000000000_0000000000000000_0000010111011010_0001111111111110"; -- 0.022859572802887886
	pesos_i(483) := b"0000000000000000_0000000000000000_0001000011001101_1111100011111000"; -- 0.06564289135373126
	pesos_i(484) := b"1111111111111111_1111111111111111_1110001101101001_1101111000001011"; -- -0.11166584224707307
	pesos_i(485) := b"1111111111111111_1111111111111111_1110010110101110_0000110110010101"; -- -0.10281291106115052
	pesos_i(486) := b"1111111111111111_1111111111111111_1100111011011111_1101001110110101"; -- -0.1918971712627521
	pesos_i(487) := b"1111111111111111_1111111111111111_1101101100111001_1001000100101100"; -- -0.14365284605664538
	pesos_i(488) := b"0000000000000000_0000000000000000_0001001111111000_0001000011100011"; -- 0.07800393611550047
	pesos_i(489) := b"0000000000000000_0000000000000000_0001101011111101_1111000011111110"; -- 0.10543733783806578
	pesos_i(490) := b"1111111111111111_1111111111111111_1111110001011111_1010100110000100"; -- -0.014165311183096767
	pesos_i(491) := b"1111111111111111_1111111111111111_1110010101110011_0101011001110011"; -- -0.10370883650651633
	pesos_i(492) := b"1111111111111111_1111111111111111_1110101011010101_1111011110011001"; -- -0.08267262007073826
	pesos_i(493) := b"0000000000000000_0000000000000000_0001000001000001_0101100010100011"; -- 0.06349710435856126
	pesos_i(494) := b"1111111111111111_1111111111111111_1110000111100101_0110100011100110"; -- -0.11759323480289029
	pesos_i(495) := b"1111111111111111_1111111111111111_1101110100110110_1011001111001011"; -- -0.13588405884998317
	pesos_i(496) := b"1111111111111111_1111111111111111_1111000001000011_0011000011001011"; -- -0.061474752796456505
	pesos_i(497) := b"1111111111111111_1111111111111111_1101110011010100_1110100010110110"; -- -0.1373762661684855
	pesos_i(498) := b"0000000000000000_0000000000000000_0010001011010000_0000000101000010"; -- 0.13598640306925505
	pesos_i(499) := b"0000000000000000_0000000000000000_0001010111000101_1010111000010011"; -- 0.08504760716070756
	pesos_i(500) := b"1111111111111111_1111111111111111_1101110000111010_0010000110001010"; -- -0.13973799119360067
	pesos_i(501) := b"1111111111111111_1111111111111111_1111100010001101_0000110011111000"; -- -0.029097737814817122
	pesos_i(502) := b"1111111111111111_1111111111111111_1101101101001110_0101111000001001"; -- -0.14333545946594067
	pesos_i(503) := b"0000000000000000_0000000000000000_0001111111111001_1111110011000110"; -- 0.12490825500678569
	pesos_i(504) := b"0000000000000000_0000000000000000_0001101001001101_1111000101110100"; -- 0.10275181856609979
	pesos_i(505) := b"0000000000000000_0000000000000000_0000001110000111_1010011110000000"; -- 0.013788670307649454
	pesos_i(506) := b"1111111111111111_1111111111111111_1111100110010110_0111011110100001"; -- -0.02504780115115265
	pesos_i(507) := b"0000000000000000_0000000000000000_0000101111001011_0010100000100001"; -- 0.04606867613468099
	pesos_i(508) := b"0000000000000000_0000000000000000_0001111101100101_0100001111111101"; -- 0.12263894010614347
	pesos_i(509) := b"0000000000000000_0000000000000000_0000000001001111_0001101100000011"; -- 0.0012070544175971022
	pesos_i(510) := b"0000000000000000_0000000000000000_0010000011001001_1100111110100100"; -- 0.12807939287851103
	pesos_i(511) := b"0000000000000000_0000000000000000_0010101001001001_1100110011111011"; -- 0.16518860949669456
	pesos_i(512) := b"1111111111111111_1111111111111111_1101101101011011_0010111111110110"; -- -0.14313984153667125
	pesos_i(513) := b"0000000000000000_0000000000000000_0000010110011001_1000110001010111"; -- 0.021874209608510817
	pesos_i(514) := b"0000000000000000_0000000000000000_0001011011100110_0110000010000101"; -- 0.0894527746024575
	pesos_i(515) := b"1111111111111111_1111111111111111_1111000001100010_0101111001001011"; -- -0.060999018433166075
	pesos_i(516) := b"1111111111111111_1111111111111111_1101110110101000_0110110000111011"; -- -0.13414882244421802
	pesos_i(517) := b"1111111111111111_1111111111111111_1111101000001000_0110111110100101"; -- -0.023308775064952686
	pesos_i(518) := b"1111111111111111_1111111111111111_1101011011011110_1101001101100000"; -- -0.16066245000699697
	pesos_i(519) := b"1111111111111111_1111111111111111_1110000100111010_1010110001000000"; -- -0.12019847334558025
	pesos_i(520) := b"0000000000000000_0000000000000000_0000111101011100_0010110001100100"; -- 0.06000020450524255
	pesos_i(521) := b"1111111111111111_1111111111111111_1101010110000111_0100100011111010"; -- -0.16590446383286367
	pesos_i(522) := b"1111111111111111_1111111111111111_1111011000100100_0110111111010111"; -- -0.03850651735069441
	pesos_i(523) := b"0000000000000000_0000000000000000_0001100011001011_0011100000110000"; -- 0.09685088324917018
	pesos_i(524) := b"0000000000000000_0000000000000000_0001001110001001_1010111001110011"; -- 0.07631960214410398
	pesos_i(525) := b"1111111111111111_1111111111111111_1111110000010101_0100011010000100"; -- -0.015300362362227666
	pesos_i(526) := b"0000000000000000_0000000000000000_0010101110101000_0101110001011111"; -- 0.17053773221850874
	pesos_i(527) := b"1111111111111111_1111111111111111_1111011110011000_1011010111100010"; -- -0.03282607299366893
	pesos_i(528) := b"1111111111111111_1111111111111111_1111100101111011_1001101001111001"; -- -0.025457711606584433
	pesos_i(529) := b"1111111111111111_1111111111111111_1100110001100110_0110100100101111"; -- -0.20156233401999402
	pesos_i(530) := b"1111111111111111_1111111111111111_1111001000010100_0111001010010101"; -- -0.05437549461579931
	pesos_i(531) := b"0000000000000000_0000000000000000_0001110111001110_0011111000101101"; -- 0.11642826643581929
	pesos_i(532) := b"0000000000000000_0000000000000000_0000011010011010_0111100010110000"; -- 0.02579454706832258
	pesos_i(533) := b"1111111111111111_1111111111111111_1110000110000011_1111010101110010"; -- -0.11908021885981686
	pesos_i(534) := b"1111111111111111_1111111111111111_1111001110100011_0111010110101011"; -- -0.04828705391556589
	pesos_i(535) := b"0000000000000000_0000000000000000_0000110000001100_1010100000111011"; -- 0.04706813273459524
	pesos_i(536) := b"0000000000000000_0000000000000000_0010100000000111_0110111110110011"; -- 0.156363469401512
	pesos_i(537) := b"0000000000000000_0000000000000000_0000111110011010_0010100001110100"; -- 0.06094601472763867
	pesos_i(538) := b"0000000000000000_0000000000000000_0001110110001101_1000100000011010"; -- 0.11544085148363663
	pesos_i(539) := b"0000000000000000_0000000000000000_0001010001000000_0011101001101110"; -- 0.07910504511517578
	pesos_i(540) := b"1111111111111111_1111111111111111_1111110000000001_1100000110011111"; -- -0.015598200606382642
	pesos_i(541) := b"0000000000000000_0000000000000000_0000111001011001_1000110011100111"; -- 0.0560539307408402
	pesos_i(542) := b"1111111111111111_1111111111111111_1111000010100100_0100100000100001"; -- -0.059993259399649446
	pesos_i(543) := b"1111111111111111_1111111111111111_1110011110010100_1101001111011101"; -- -0.09538532115500842
	pesos_i(544) := b"0000000000000000_0000000000000000_0010001011001100_0001110011111011"; -- 0.13592702038076815
	pesos_i(545) := b"1111111111111111_1111111111111111_1111100100100100_1010111111010100"; -- -0.026783953533498987
	pesos_i(546) := b"0000000000000000_0000000000000000_0001110011000100_0001110110010101"; -- 0.11236748596009234
	pesos_i(547) := b"0000000000000000_0000000000000000_0010000000010010_1111111110100001"; -- 0.12528989493710166
	pesos_i(548) := b"0000000000000000_0000000000000000_0000100011011111_1001101101100111"; -- 0.03466197261541646
	pesos_i(549) := b"1111111111111111_1111111111111111_1101111001111000_0011111011010011"; -- -0.13097770067610495
	pesos_i(550) := b"1111111111111111_1111111111111111_1111000001010000_0000100111001001"; -- -0.06127871357471225
	pesos_i(551) := b"1111111111111111_1111111111111111_1110010101010100_1101010101010000"; -- -0.1041742973114718
	pesos_i(552) := b"0000000000000000_0000000000000000_0000101100101001_1111001000010000"; -- 0.0436087884339597
	pesos_i(553) := b"0000000000000000_0000000000000000_0001111111100010_0110100010010010"; -- 0.12454846913437287
	pesos_i(554) := b"0000000000000000_0000000000000000_0010101010101011_0100100101000111"; -- 0.16667612052268113
	pesos_i(555) := b"1111111111111111_1111111111111111_1111010111011111_1101101010001110"; -- -0.039553013097380185
	pesos_i(556) := b"1111111111111111_1111111111111111_1111011001010100_0010110111010011"; -- -0.03777803044273827
	pesos_i(557) := b"0000000000000000_0000000000000000_0000111110101100_1010010001111111"; -- 0.06122806654616528
	pesos_i(558) := b"1111111111111111_1111111111111111_1111010010111000_0110000101101010"; -- -0.04406157637128199
	pesos_i(559) := b"0000000000000000_0000000000000000_0001110001100110_1111100011001011"; -- 0.11094622563994802
	pesos_i(560) := b"1111111111111111_1111111111111111_1101111111111011_0101001011101100"; -- -0.12507135131837988
	pesos_i(561) := b"1111111111111111_1111111111111111_1101010001000101_1010111100101001"; -- -0.17081170320939146
	pesos_i(562) := b"0000000000000000_0000000000000000_0000000100001010_0100101010101101"; -- 0.004063289029498085
	pesos_i(563) := b"1111111111111111_1111111111111111_1100111010011111_1101011000110110"; -- -0.19287358460411697
	pesos_i(564) := b"1111111111111111_1111111111111111_1101110101011000_1001011000001011"; -- -0.13536703332772665
	pesos_i(565) := b"1111111111111111_1111111111111111_1100101111101001_0000111000101001"; -- -0.20347510813600467
	pesos_i(566) := b"0000000000000000_0000000000000000_0000011110111110_0010110101110110"; -- 0.03024562968810958
	pesos_i(567) := b"0000000000000000_0000000000000000_0000010011111111_1011100111110011"; -- 0.01952707454938866
	pesos_i(568) := b"1111111111111111_1111111111111111_1101111100000100_0101100001000011"; -- -0.12883995403801662
	pesos_i(569) := b"0000000000000000_0000000000000000_0000011011011101_0001100100100100"; -- 0.026811190845143468
	pesos_i(570) := b"1111111111111111_1111111111111111_1110101110101010_0000110111001011"; -- -0.07943643377746498
	pesos_i(571) := b"1111111111111111_1111111111111111_1110000100100001_0011101001011111"; -- -0.1205867306839288
	pesos_i(572) := b"0000000000000000_0000000000000000_0000101101010000_1100001101010100"; -- 0.044201095566661394
	pesos_i(573) := b"1111111111111111_1111111111111111_1101111111000101_1111100000001011"; -- -0.12588548399912683
	pesos_i(574) := b"0000000000000000_0000000000000000_0010000001001000_0110001000010101"; -- 0.12610447895475996
	pesos_i(575) := b"0000000000000000_0000000000000000_0000000000010101_1011001111111000"; -- 0.0003311615080060065
	pesos_i(576) := b"0000000000000000_0000000000000000_0000000100010111_0001100111011111"; -- 0.00425874424549578
	pesos_i(577) := b"1111111111111111_1111111111111111_1110101100100111_0010100110001100"; -- -0.08143368075476921
	pesos_i(578) := b"0000000000000000_0000000000000000_0001110010010010_1000001110010111"; -- 0.11161062666044033
	pesos_i(579) := b"0000000000000000_0000000000000000_0000001011000110_0010111110101000"; -- 0.010836580804197258
	pesos_i(580) := b"0000000000000000_0000000000000000_0010100010011010_1000110100010100"; -- 0.15860826239424572
	pesos_i(581) := b"1111111111111111_1111111111111111_1101110011010111_1001001111101000"; -- -0.1373355444198506
	pesos_i(582) := b"0000000000000000_0000000000000000_0000000001010111_1010100001111001"; -- 0.001337556475653311
	pesos_i(583) := b"1111111111111111_1111111111111111_1101100101011110_0101100100110000"; -- -0.15090410795326714
	pesos_i(584) := b"0000000000000000_0000000000000000_0010101101110110_1100111101101110"; -- 0.16978165079069316
	pesos_i(585) := b"0000000000000000_0000000000000000_0001010110001011_1011111011001111"; -- 0.08416359482684047
	pesos_i(586) := b"1111111111111111_1111111111111111_1101110111011100_0010011110101101"; -- -0.13335945156342607
	pesos_i(587) := b"1111111111111111_1111111111111111_1110111001001101_0111011010111100"; -- -0.06913049608582982
	pesos_i(588) := b"1111111111111111_1111111111111111_1110110110000111_0011100110101011"; -- -0.07215537621889183
	pesos_i(589) := b"1111111111111111_1111111111111111_1101011011111111_0110111111111100"; -- -0.16016483407861828
	pesos_i(590) := b"0000000000000000_0000000000000000_0000110010010111_1100011000000100"; -- 0.049190879864729094
	pesos_i(591) := b"0000000000000000_0000000000000000_0010101101100011_0000001001111001"; -- 0.169479517535149
	pesos_i(592) := b"1111111111111111_1111111111111111_1110000010011000_1011011010111111"; -- -0.12266977163724148
	pesos_i(593) := b"1111111111111111_1111111111111111_1110001010010100_1111000000010011"; -- -0.1149148896056219
	pesos_i(594) := b"1111111111111111_1111111111111111_1101011110101101_0000000011010000"; -- -0.15751643095980392
	pesos_i(595) := b"0000000000000000_0000000000000000_0001011010110010_0001001101110001"; -- 0.08865472322752371
	pesos_i(596) := b"1111111111111111_1111111111111111_1101010010011101_0100111111011010"; -- -0.16947461062779615
	pesos_i(597) := b"1111111111111111_1111111111111111_1101110001000101_1100110010101101"; -- -0.13955994402638588
	pesos_i(598) := b"1111111111111111_1111111111111111_1111010111000111_0111001011110000"; -- -0.039925400057021575
	pesos_i(599) := b"0000000000000000_0000000000000000_0010010010101001_1111010010001101"; -- 0.1432183116298898
	pesos_i(600) := b"0000000000000000_0000000000000000_0011010011101011_1011010010011000"; -- 0.20672157963352542
	pesos_i(601) := b"1111111111111111_1111111111111111_1110111011001000_0100111101010011"; -- -0.0672560141211189
	pesos_i(602) := b"0000000000000000_0000000000000000_0001101101111101_1111001011100010"; -- 0.10739057565527763
	pesos_i(603) := b"0000000000000000_0000000000000000_0001001111110111_0110100101011011"; -- 0.07799395067660242
	pesos_i(604) := b"0000000000000000_0000000000000000_0000000011101101_0100011000110111"; -- 0.0036205182507398704
	pesos_i(605) := b"0000000000000000_0000000000000000_0001001011111100_0011100010111100"; -- 0.07416109640458589
	pesos_i(606) := b"0000000000000000_0000000000000000_0000001011000010_1111001000101011"; -- 0.01078713946494204
	pesos_i(607) := b"0000000000000000_0000000000000000_0010001111000010_0101100001011101"; -- 0.13968422191462748
	pesos_i(608) := b"0000000000000000_0000000000000000_0001101100010000_1011000101001101"; -- 0.1057234586317536
	pesos_i(609) := b"1111111111111111_1111111111111111_1111010011010110_1010101111100110"; -- -0.04359937321264137
	pesos_i(610) := b"0000000000000000_0000000000000000_0001001011000101_0101100011010000"; -- 0.07332377518602708
	pesos_i(611) := b"1111111111111111_1111111111111111_1111100101000101_0111111010101110"; -- -0.026283342896315537
	pesos_i(612) := b"1111111111111111_1111111111111111_1101101011011010_0011000010111011"; -- -0.14510817953162614
	pesos_i(613) := b"1111111111111111_1111111111111111_1111010101110000_1010110110100100"; -- -0.041249415886423633
	pesos_i(614) := b"1111111111111111_1111111111111111_1111010000010011_0010011000010101"; -- -0.046582813076654905
	pesos_i(615) := b"1111111111111111_1111111111111111_1111100010111011_1010010100011001"; -- -0.028386765930213793
	pesos_i(616) := b"1111111111111111_1111111111111111_1101101101100100_0000110100100110"; -- -0.1430045874148533
	pesos_i(617) := b"0000000000000000_0000000000000000_0001011101100001_1110100110010000"; -- 0.09133777406420825
	pesos_i(618) := b"1111111111111111_1111111111111111_1101011101111010_1111110001111111"; -- -0.1582796278316019
	pesos_i(619) := b"1111111111111111_1111111111111111_1111110111100101_1110001001001110"; -- -0.008210998405754408
	pesos_i(620) := b"1111111111111111_1111111111111111_1110010000000111_0001000100010001"; -- -0.10926717124823015
	pesos_i(621) := b"0000000000000000_0000000000000000_0010000001000111_0111101000100000"; -- 0.1260906532073568
	pesos_i(622) := b"1111111111111111_1111111111111111_1110101010000110_1101101100100001"; -- -0.08387976117206086
	pesos_i(623) := b"1111111111111111_1111111111111111_1110110001101111_1000101010010110"; -- -0.07642301406603016
	pesos_i(624) := b"1111111111111111_1111111111111111_1110011110101001_0101101000000010"; -- -0.0950721496815206
	pesos_i(625) := b"1111111111111111_1111111111111111_1101100011100010_0101101100001111"; -- -0.15279608612251103
	pesos_i(626) := b"0000000000000000_0000000000000000_0000011000101110_1100110100110001"; -- 0.0241516347534065
	pesos_i(627) := b"1111111111111111_1111111111111111_1110001111000111_0111100010011010"; -- -0.11023756264615829
	pesos_i(628) := b"1111111111111111_1111111111111111_1101001110010001_1011011000101000"; -- -0.17355786816912952
	pesos_i(629) := b"1111111111111111_1111111111111111_1110000110001001_0101100111101010"; -- -0.1189979365719408
	pesos_i(630) := b"1111111111111111_1111111111111111_1111111000001111_0011111110001010"; -- -0.007579831005815213
	pesos_i(631) := b"1111111111111111_1111111111111111_1110111110010111_0001101001110101"; -- -0.06410059580557283
	pesos_i(632) := b"1111111111111111_1111111111111111_1101111100100101_0101100111100100"; -- -0.12833631686782224
	pesos_i(633) := b"1111111111111111_1111111111111111_1111010000001000_1010000001001010"; -- -0.04674337573453337
	pesos_i(634) := b"0000000000000000_0000000000000000_0000100010010011_0001100001001011"; -- 0.03349448996701489
	pesos_i(635) := b"0000000000000000_0000000000000000_0000000010100001_0000111011000111"; -- 0.002457545824311534
	pesos_i(636) := b"1111111111111111_1111111111111111_1101010011101001_1011010111010110"; -- -0.1683088639032655
	pesos_i(637) := b"1111111111111111_1111111111111111_1101011111011011_0111001111010101"; -- -0.1568076710285522
	pesos_i(638) := b"0000000000000000_0000000000000000_0000110010110101_1000011000001100"; -- 0.04964483074728823
	pesos_i(639) := b"1111111111111111_1111111111111111_1111100000010010_1110001010110101"; -- -0.030961829116139254
	pesos_i(640) := b"1111111111111111_1111111111111111_1101110011101100_1100101000000010"; -- -0.13701188527130892
	pesos_i(641) := b"1111111111111111_1111111111111111_1101110101000011_0110110111001001"; -- -0.13568986746553865
	pesos_i(642) := b"0000000000000000_0000000000000000_0000101000111011_0110000010011010"; -- 0.03996852639120013
	pesos_i(643) := b"0000000000000000_0000000000000000_0001100100010011_0011100101100110"; -- 0.09794958822525762
	pesos_i(644) := b"1111111111111111_1111111111111111_1111101001010111_1010111110111010"; -- -0.022099511342900294
	pesos_i(645) := b"1111111111111111_1111111111111111_1101101001111010_0101011100110000"; -- -0.14657073092805264
	pesos_i(646) := b"0000000000000000_0000000000000000_0001000010110011_0111001110111011"; -- 0.06523822140706784
	pesos_i(647) := b"1111111111111111_1111111111111111_1110101111111100_1101110111100011"; -- -0.07817280973087365
	pesos_i(648) := b"0000000000000000_0000000000000000_0000100001011100_0111001011101110"; -- 0.03266065884150258
	pesos_i(649) := b"0000000000000000_0000000000000000_0000110011101010_0110100000110001"; -- 0.05045176686996206
	pesos_i(650) := b"0000000000000000_0000000000000000_0100010011010001_0110010101010001"; -- 0.26882012587715104
	pesos_i(651) := b"0000000000000000_0000000000000000_0001010100011100_0100001001111000"; -- 0.08246245797636542
	pesos_i(652) := b"0000000000000000_0000000000000000_0000000100111110_0111001111100101"; -- 0.004859202841492065
	pesos_i(653) := b"0000000000000000_0000000000000000_0001000010110010_0100100001001011"; -- 0.0652203735395322
	pesos_i(654) := b"1111111111111111_1111111111111111_1101111000100111_1000010101110011"; -- -0.1322094530075436
	pesos_i(655) := b"0000000000000000_0000000000000000_0000011111010110_0001000100111010"; -- 0.03061015756595855
	pesos_i(656) := b"1111111111111111_1111111111111111_1110110010010100_1000111100011101"; -- -0.0758581689702538
	pesos_i(657) := b"1111111111111111_1111111111111111_1101110110011001_1010001110000000"; -- -0.1343744098009109
	pesos_i(658) := b"1111111111111111_1111111111111111_1110011011100010_0101011101000001"; -- -0.09810881296703615
	pesos_i(659) := b"1111111111111111_1111111111111111_1101001011111110_0111011000100001"; -- -0.17580472650202567
	pesos_i(660) := b"1111111111111111_1111111111111111_1110000011100010_0110010101110111"; -- -0.12154546593856752
	pesos_i(661) := b"0000000000000000_0000000000000000_0010100001000000_0101001111100111"; -- 0.1572315634009199
	pesos_i(662) := b"1111111111111111_1111111111111111_1111100110011001_0101010101111110"; -- -0.02500405964650106
	pesos_i(663) := b"1111111111111111_1111111111111111_1111100001110001_1000100111101001"; -- -0.029517536714410007
	pesos_i(664) := b"1111111111111111_1111111111111111_1101100110100110_0011000111010010"; -- -0.1498078214281784
	pesos_i(665) := b"0000000000000000_0000000000000000_0000010001110011_0000110010101100"; -- 0.017380516105838618
	pesos_i(666) := b"1111111111111111_1111111111111111_1110101110110011_1101010111111010"; -- -0.07928717271512596
	pesos_i(667) := b"1111111111111111_1111111111111111_1100000000001101_1110011000111000"; -- -0.24978791357246466
	pesos_i(668) := b"0000000000000000_0000000000000000_0000010101101101_1010101010100110"; -- 0.021204629536555723
	pesos_i(669) := b"1111111111111111_1111111111111111_1111001101101100_0000001111100011"; -- -0.04913306918976867
	pesos_i(670) := b"1111111111111111_1111111111111111_1110111101001111_1011000000011011"; -- -0.06519030903020884
	pesos_i(671) := b"1111111111111111_1111111111111111_1101100010100011_1010010100101001"; -- -0.15375297313662376
	pesos_i(672) := b"1111111111111111_1111111111111111_1111110010000010_1000111001000000"; -- -0.013632878670911255
	pesos_i(673) := b"1111111111111111_1111111111111111_1111110101010001_1010101001111111"; -- -0.010472625829957498
	pesos_i(674) := b"0000000000000000_0000000000000000_0001010010111001_1010100101011110"; -- 0.08095797104290613
	pesos_i(675) := b"0000000000000000_0000000000000000_0001010010101110_0000000011101001"; -- 0.08078008346560449
	pesos_i(676) := b"0000000000000000_0000000000000000_0000111111001111_1010001010101101"; -- 0.06176201558669629
	pesos_i(677) := b"0000000000000000_0000000000000000_0001011110101100_0001001001100101"; -- 0.09246935819776614
	pesos_i(678) := b"1111111111111111_1111111111111111_1101010011111010_0001101100110100"; -- -0.1680586813346377
	pesos_i(679) := b"0000000000000000_0000000000000000_0001111000000111_0100101101110111"; -- 0.1172988094888686
	pesos_i(680) := b"1111111111111111_1111111111111111_1110111100101000_0001110001100011"; -- -0.06579420655790733
	pesos_i(681) := b"1111111111111111_1111111111111111_1111001100001000_1101000101010010"; -- -0.05064670316502472
	pesos_i(682) := b"1111111111111111_1111111111111111_1101000111001111_1111001101011010"; -- -0.18042067586741733
	pesos_i(683) := b"0000000000000000_0000000000000000_0000010011110101_1110011011001100"; -- 0.01937715994769946
	pesos_i(684) := b"1111111111111111_1111111111111111_1110100110110000_1101011111111111"; -- -0.08714532868549787
	pesos_i(685) := b"1111111111111111_1111111111111111_1111100011101011_0111110010001100"; -- -0.02765676092214493
	pesos_i(686) := b"0000000000000000_0000000000000000_0010001011000010_1101101011001010"; -- 0.13578574602871477
	pesos_i(687) := b"0000000000000000_0000000000000000_0000010000111010_1101000101001000"; -- 0.016522483999146634
	pesos_i(688) := b"0000000000000000_0000000000000000_0010001110001101_1100110111101110"; -- 0.13888251359707238
	pesos_i(689) := b"0000000000000000_0000000000000000_0010000101100011_1000111110110110"; -- 0.13042543593232586
	pesos_i(690) := b"0000000000000000_0000000000000000_0001101111100000_1010001110100011"; -- 0.10889647237070268
	pesos_i(691) := b"1111111111111111_1111111111111111_1110101001101111_1011110010001001"; -- -0.0842325368188373
	pesos_i(692) := b"0000000000000000_0000000000000000_0010000011101000_1000011100110100"; -- 0.12854809785274693
	pesos_i(693) := b"0000000000000000_0000000000000000_0000001010011100_1111011111001001"; -- 0.010207640136954717
	pesos_i(694) := b"0000000000000000_0000000000000000_0000111011101111_0011000101001001"; -- 0.05833728832348187
	pesos_i(695) := b"0000000000000000_0000000000000000_0000000101000001_1100001110100011"; -- 0.004909732092643307
	pesos_i(696) := b"0000000000000000_0000000000000000_0000011011010000_1110001010001101"; -- 0.02662483168799437
	pesos_i(697) := b"0000000000000000_0000000000000000_0010110010001001_0011111110000011"; -- 0.17396923976542744
	pesos_i(698) := b"1111111111111111_1111111111111111_1111000100110001_0000011111001110"; -- -0.05784560424354493
	pesos_i(699) := b"1111111111111111_1111111111111111_1101110001001100_0101010110110100"; -- -0.13946022372843678
	pesos_i(700) := b"0000000000000000_0000000000000000_0000111100011010_1110011000001110"; -- 0.05900419087755903
	pesos_i(701) := b"1111111111111111_1111111111111111_1110100110111101_0010101001011001"; -- -0.08695731466820182
	pesos_i(702) := b"0000000000000000_0000000000000000_0010011110011100_1000110010100100"; -- 0.1547325039064936
	pesos_i(703) := b"0000000000000000_0000000000000000_0000011101111110_1011000000011000"; -- 0.029276853454713897
	pesos_i(704) := b"0000000000000000_0000000000000000_0001101011000010_0011000101011111"; -- 0.1045256478228111
	pesos_i(705) := b"1111111111111111_1111111111111111_1101011010001110_1101001000001011"; -- -0.16188323244808392
	pesos_i(706) := b"1111111111111111_1111111111111111_1111011100001000_0010011001000100"; -- -0.035031898954752255
	pesos_i(707) := b"1111111111111111_1111111111111111_1111111010101000_1111100000010010"; -- -0.005234237179312166
	pesos_i(708) := b"1111111111111111_1111111111111111_1110100111010100_0010110010111011"; -- -0.08660622064355467
	pesos_i(709) := b"1111111111111111_1111111111111111_1110001001011111_1111000001001110"; -- -0.11572359180760332
	pesos_i(710) := b"0000000000000000_0000000000000000_0001011011001110_0001110110111100"; -- 0.08908258280308642
	pesos_i(711) := b"1111111111111111_1111111111111111_1111001101110100_0101111000010111"; -- -0.049005622337001314
	pesos_i(712) := b"1111111111111111_1111111111111111_1110001001011111_1000110100001000"; -- -0.11572950894997022
	pesos_i(713) := b"0000000000000000_0000000000000000_0001011000111010_1010001000111101"; -- 0.08683217997659737
	pesos_i(714) := b"0000000000000000_0000000000000000_0000100100100100_1110111001010011"; -- 0.0357197716608052
	pesos_i(715) := b"1111111111111111_1111111111111111_1110011011100110_0001011001001110"; -- -0.0980516490597167
	pesos_i(716) := b"1111111111111111_1111111111111111_1111000011011010_0011011100100000"; -- -0.05917029837789005
	pesos_i(717) := b"1111111111111111_1111111111111111_1101111000101110_0101011100000011"; -- -0.13210540939773704
	pesos_i(718) := b"0000000000000000_0000000000000000_0001110001000101_1100111000000010"; -- 0.11044013540013815
	pesos_i(719) := b"1111111111111111_1111111111111111_1110011000011011_1000111110000001"; -- -0.1011419591255064
	pesos_i(720) := b"0000000000000000_0000000000000000_0000111110001011_1110001100110001"; -- 0.060728263427623816
	pesos_i(721) := b"1111111111111111_1111111111111111_1101100000001110_0010001100000100"; -- -0.15603428996149402
	pesos_i(722) := b"0000000000000000_0000000000000000_0010001010001101_0011010001110101"; -- 0.13496711593137745
	pesos_i(723) := b"0000000000000000_0000000000000000_0010111001011100_0011000110111100"; -- 0.18109427290313976
	pesos_i(724) := b"0000000000000000_0000000000000000_0010100110101101_1001001001111100"; -- 0.1628047515420909
	pesos_i(725) := b"1111111111111111_1111111111111111_1101101000111100_1000011010001111"; -- -0.14751395232298362
	pesos_i(726) := b"0000000000000000_0000000000000000_0000000101000011_0000111111110101"; -- 0.00492953987018949
	pesos_i(727) := b"0000000000000000_0000000000000000_0000011110010111_0100000010101100"; -- 0.02965168192875754
	pesos_i(728) := b"1111111111111111_1111111111111111_1111111110100100_0110001010011111"; -- -0.0013979303157617418
	pesos_i(729) := b"1111111111111111_1111111111111111_1101101111101110_1111001001000011"; -- -0.14088521831688677
	pesos_i(730) := b"1111111111111111_1111111111111111_1111000001110110_1100101110010100"; -- -0.060687328724770666
	pesos_i(731) := b"1111111111111111_1111111111111111_1110101111101101_0000010000101001"; -- -0.07841466899494867
	pesos_i(732) := b"0000000000000000_0000000000000000_0000011111001101_1101110001001100"; -- 0.03048493237493188
	pesos_i(733) := b"0000000000000000_0000000000000000_0000101001001010_1111111110000101"; -- 0.040206880438529505
	pesos_i(734) := b"0000000000000000_0000000000000000_0001000000010110_0110011101010010"; -- 0.06284185173773973
	pesos_i(735) := b"1111111111111111_1111111111111111_1110100110111011_0101011001101000"; -- -0.08698520620394563
	pesos_i(736) := b"0000000000000000_0000000000000000_0001111000110010_1100101001010000"; -- 0.11796249813947035
	pesos_i(737) := b"1111111111111111_1111111111111111_1111101101101110_0001100011111101"; -- -0.017851293713172123
	pesos_i(738) := b"0000000000000000_0000000000000000_0000000101101001_1111100001111110"; -- 0.005523234099626934
	pesos_i(739) := b"0000000000000000_0000000000000000_0001111101110010_1011000011101110"; -- 0.12284379768123767
	pesos_i(740) := b"0000000000000000_0000000000000000_0001010000110010_1011111011100110"; -- 0.07889931795622845
	pesos_i(741) := b"1111111111111111_1111111111111111_1100111110010100_0001111100000101"; -- -0.18914610024354336
	pesos_i(742) := b"1111111111111111_1111111111111111_1111010100110110_0110111000100001"; -- -0.042138211170341
	pesos_i(743) := b"1111111111111111_1111111111111111_1101010000001101_1100000111001101"; -- -0.17166508430308583
	pesos_i(744) := b"1111111111111111_1111111111111111_1111101100001011_0001011001000100"; -- -0.01936207627431319
	pesos_i(745) := b"0000000000000000_0000000000000000_0001011101100101_1101110100010000"; -- 0.09139806409974088
	pesos_i(746) := b"1111111111111111_1111111111111111_1101010010101011_0011010010011001"; -- -0.16926261200182582
	pesos_i(747) := b"1111111111111111_1111111111111111_1110001110110111_0010000101011000"; -- -0.11048690409243032
	pesos_i(748) := b"0000000000000000_0000000000000000_0010110101111111_1101101000110100"; -- 0.17773212223146503
	pesos_i(749) := b"1111111111111111_1111111111111111_1111111010011000_0100010000100011"; -- -0.005489102692550716
	pesos_i(750) := b"0000000000000000_0000000000000000_0000010110000010_1110000110000101"; -- 0.021528334503215292
	pesos_i(751) := b"1111111111111111_1111111111111111_1111111111000011_0000111100110011"; -- -0.0009298801754966729
	pesos_i(752) := b"0000000000000000_0000000000000000_0000000101111001_1010101000111001"; -- 0.0057627095844637755
	pesos_i(753) := b"0000000000000000_0000000000000000_0000000110100110_0111010000001011"; -- 0.00644612575372997
	pesos_i(754) := b"1111111111111111_1111111111111111_1101101000011011_0110100001100010"; -- -0.14801929092124574
	pesos_i(755) := b"1111111111111111_1111111111111111_1101110011001101_1101011100011111"; -- -0.13748412607082341
	pesos_i(756) := b"0000000000000000_0000000000000000_0010011011011100_1001110010000100"; -- 0.15180376275377772
	pesos_i(757) := b"1111111111111111_1111111111111111_1111111100000001_1100110101001000"; -- -0.0038787554005778836
	pesos_i(758) := b"0000000000000000_0000000000000000_0001010100011100_0101110111010001"; -- 0.08246408803243334
	pesos_i(759) := b"0000000000000000_0000000000000000_0001110110111011_0000101001111100"; -- 0.11613526842341722
	pesos_i(760) := b"0000000000000000_0000000000000000_0000010111000011_0010110101101110"; -- 0.022509421623687215
	pesos_i(761) := b"0000000000000000_0000000000000000_0001110110001001_0010011100111011"; -- 0.11537404243052779
	pesos_i(762) := b"0000000000000000_0000000000000000_0000101110011111_1101000010110110"; -- 0.04540733757254806
	pesos_i(763) := b"1111111111111111_1111111111111111_1111111011110101_1000101000101001"; -- -0.004065861804042151
	pesos_i(764) := b"0000000000000000_0000000000000000_0000001000111101_1011100001111111"; -- 0.008754283059868417
	pesos_i(765) := b"1111111111111111_1111111111111111_1100111011011011_0111010000001011"; -- -0.19196390844731517
	pesos_i(766) := b"0000000000000000_0000000000000000_0001010001110110_1001001101110100"; -- 0.07993432589264587
	pesos_i(767) := b"0000000000000000_0000000000000000_0010100111010010_0110111010001011"; -- 0.16336718453594523
	pesos_i(768) := b"0000000000000000_0000000000000000_0001100100100101_1110010000000010"; -- 0.09823441556650517
	pesos_i(769) := b"1111111111111111_1111111111111111_1110111001010010_0000111001001011"; -- -0.06906042730902104
	pesos_i(770) := b"0000000000000000_0000000000000000_0010001001011010_1101111010110111"; -- 0.13419906586982988
	pesos_i(771) := b"0000000000000000_0000000000000000_0010001110110010_1010011110010001"; -- 0.1394448021317237
	pesos_i(772) := b"1111111111111111_1111111111111111_1101110001010111_0100000011011101"; -- -0.1392936190901022
	pesos_i(773) := b"1111111111111111_1111111111111111_1110110010110001_0000000110100101"; -- -0.07542409634177248
	pesos_i(774) := b"1111111111111111_1111111111111111_1101010101001001_0011100111001000"; -- -0.166851414468342
	pesos_i(775) := b"1111111111111111_1111111111111111_1111101010000100_1100000000010011"; -- -0.021411891383002576
	pesos_i(776) := b"0000000000000000_0000000000000000_0000001001101101_0011110100011010"; -- 0.00947934995357557
	pesos_i(777) := b"0000000000000000_0000000000000000_0010001010001011_0001110001100101"; -- 0.13493516404775543
	pesos_i(778) := b"0000000000000000_0000000000000000_0001000100000011_1111010101101110"; -- 0.06646665517405043
	pesos_i(779) := b"0000000000000000_0000000000000000_0001000100100110_0000011100100100"; -- 0.06698650966661532
	pesos_i(780) := b"0000000000000000_0000000000000000_0000100010101100_0010001011011001"; -- 0.033876588898760655
	pesos_i(781) := b"0000000000000000_0000000000000000_0011001111101101_0011010111010000"; -- 0.20283829052420274
	pesos_i(782) := b"1111111111111111_1111111111111111_1101111000010000_0011011110000001"; -- -0.13256505104380192
	pesos_i(783) := b"1111111111111111_1111111111111111_1101010011100100_1001011010010100"; -- -0.16838702083532506
	pesos_i(784) := b"1111111111111111_1111111111111111_1110101010010101_1010000011110110"; -- -0.08365434647402692
	pesos_i(785) := b"1111111111111111_1111111111111111_1111010111101000_0001111000001100"; -- -0.03942692000926121
	pesos_i(786) := b"0000000000000000_0000000000000000_0001000010001101_1000101101010110"; -- 0.06465979442461102
	pesos_i(787) := b"0000000000000000_0000000000000000_0000010111110011_0100110111101010"; -- 0.023243779706706384
	pesos_i(788) := b"0000000000000000_0000000000000000_0001100011011010_0110001010101110"; -- 0.0970822978949391
	pesos_i(789) := b"1111111111111111_1111111111111111_1110000101011010_0110110110001101"; -- -0.11971392922440253
	pesos_i(790) := b"1111111111111111_1111111111111111_1110000111101111_1001011010100011"; -- -0.11743792079928286
	pesos_i(791) := b"1111111111111111_1111111111111111_1111010100110111_0100001110101011"; -- -0.04212548326430317
	pesos_i(792) := b"0000000000000000_0000000000000000_0001111011011111_0100000000011101"; -- 0.12059403141237438
	pesos_i(793) := b"0000000000000000_0000000000000000_0010001110101111_0010111101000010"; -- 0.13939185494690473
	pesos_i(794) := b"0000000000000000_0000000000000000_0000110100100000_0100110001101110"; -- 0.051274086904901095
	pesos_i(795) := b"0000000000000000_0000000000000000_0010010000111010_1001110100011101"; -- 0.14151937445937646
	pesos_i(796) := b"1111111111111111_1111111111111111_1101101110100111_1110110111011011"; -- -0.14196885492470895
	pesos_i(797) := b"1111111111111111_1111111111111111_1111100100101100_0100111101111011"; -- -0.026667625849363413
	pesos_i(798) := b"0000000000000000_0000000000000000_0010000011110100_1010001100111110"; -- 0.12873287461560026
	pesos_i(799) := b"0000000000000000_0000000000000000_0000010001011011_0100110001001111"; -- 0.017018098073797512
	pesos_i(800) := b"1111111111111111_1111111111111111_1100111110001011_1110100101010110"; -- -0.18927137035892322
	pesos_i(801) := b"0000000000000000_0000000000000000_0001111100011101_1100101010001011"; -- 0.12154832748641453
	pesos_i(802) := b"1111111111111111_1111111111111111_1111111001100100_0001111011000100"; -- -0.006284787319608631
	pesos_i(803) := b"1111111111111111_1111111111111111_1110101101100001_0111010110111110"; -- -0.08054412940175143
	pesos_i(804) := b"1111111111111111_1111111111111111_1101110110111000_0110110000110111"; -- -0.13390468271714717
	pesos_i(805) := b"0000000000000000_0000000000000000_0001011101001000_0110111110101110"; -- 0.09094903946899553
	pesos_i(806) := b"1111111111111111_1111111111111111_1110010010000110_1000000000001011"; -- -0.10732269030564132
	pesos_i(807) := b"0000000000000000_0000000000000000_0001111110111110_1000101111101110"; -- 0.12400126039513991
	pesos_i(808) := b"1111111111111111_1111111111111111_1101000000011100_0000111010001011"; -- -0.18707188706627603
	pesos_i(809) := b"1111111111111111_1111111111111111_1100111111111101_0100001011111111"; -- -0.18754178313257588
	pesos_i(810) := b"1111111111111111_1111111111111111_1101001010011110_1001011000010101"; -- -0.1772676657483637
	pesos_i(811) := b"1111111111111111_1111111111111111_1101100001110010_1110001010011000"; -- -0.15449699197362152
	pesos_i(812) := b"0000000000000000_0000000000000000_0010101001101010_0110110011000011"; -- 0.16568641430004674
	pesos_i(813) := b"0000000000000000_0000000000000000_0011010001011101_0000100101010100"; -- 0.20454462341011226
	pesos_i(814) := b"0000000000000000_0000000000000000_0000011010100111_0000011000011111"; -- 0.02598608271715609
	pesos_i(815) := b"0000000000000000_0000000000000000_0010101001011110_1111011110011000"; -- 0.16551158396167512
	pesos_i(816) := b"0000000000000000_0000000000000000_0000000110110101_0001101010011011"; -- 0.006669676526432628
	pesos_i(817) := b"0000000000000000_0000000000000000_0000111011100000_0111001110111000"; -- 0.05811236606758195
	pesos_i(818) := b"0000000000000000_0000000000000000_0001000011111110_1001110010011101"; -- 0.06638506721858785
	pesos_i(819) := b"1111111111111111_1111111111111111_1110101001111110_1011100010101001"; -- -0.08400388608272837
	pesos_i(820) := b"0000000000000000_0000000000000000_0100001000101000_1011111000111111"; -- 0.25843419109564464
	pesos_i(821) := b"0000000000000000_0000000000000000_0000100010101111_1011110111100011"; -- 0.033931606253834234
	pesos_i(822) := b"1111111111111111_1111111111111111_1101111110000010_1111101000001001"; -- -0.12690770426819536
	pesos_i(823) := b"0000000000000000_0000000000000000_0000111001001001_1000000110111111"; -- 0.05580912507276298
	pesos_i(824) := b"1111111111111111_1111111111111111_1101100000111000_0001100101000111"; -- -0.15539400118423297
	pesos_i(825) := b"0000000000000000_0000000000000000_0000001001111100_0010000100001111"; -- 0.009706560290730545
	pesos_i(826) := b"1111111111111111_1111111111111111_1111110111101111_1100011110000101"; -- -0.00806000722288273
	pesos_i(827) := b"0000000000000000_0000000000000000_0010101110110110_0010111110000111"; -- 0.17074868246902317
	pesos_i(828) := b"0000000000000000_0000000000000000_0000011001011001_0000011101101101"; -- 0.02479597475876415
	pesos_i(829) := b"0000000000000000_0000000000000000_0001000010111110_0010000100111100"; -- 0.06540115088355852
	pesos_i(830) := b"1111111111111111_1111111111111111_1110101101010000_0111010011001110"; -- -0.08080358470041922
	pesos_i(831) := b"0000000000000000_0000000000000000_0000100110011001_1000011110010011"; -- 0.03749892564239235
	pesos_i(832) := b"1111111111111111_1111111111111111_1110010001110010_0001000100000111"; -- -0.10763448303261403
	pesos_i(833) := b"1111111111111111_1111111111111111_1111000100101110_0000100100111000"; -- -0.057891296334115216
	pesos_i(834) := b"0000000000000000_0000000000000000_0010010000001010_0110101000111010"; -- 0.14078391947640245
	pesos_i(835) := b"0000000000000000_0000000000000000_0000010001111100_0000100110101100"; -- 0.01751766644121555
	pesos_i(836) := b"0000000000000000_0000000000000000_0011110101000100_1111001001101001"; -- 0.23933329637852344
	pesos_i(837) := b"1111111111111111_1111111111111111_1110000011000100_1001101110010010"; -- -0.12200000453677075
	pesos_i(838) := b"1111111111111111_1111111111111111_1110111001110100_1111011110101011"; -- -0.06852771828628659
	pesos_i(839) := b"0000000000000000_0000000000000000_0001001111001000_1011110000001100"; -- 0.07728171632536814
	pesos_i(840) := b"1111111111111111_1111111111111111_1110000000111000_1101101110111001"; -- -0.12413241134721632
	pesos_i(841) := b"1111111111111111_1111111111111111_1110010100010111_1100010000011010"; -- -0.10510610917932439
	pesos_i(842) := b"0000000000000000_0000000000000000_0000000101000000_0000100110101110"; -- 0.004883389356520218
	pesos_i(843) := b"1111111111111111_1111111111111111_1110101110010111_0010000000110001"; -- -0.07972525413815412
	pesos_i(844) := b"0000000000000000_0000000000000000_0100100000110110_0011111101101111"; -- 0.28207775558321296
	pesos_i(845) := b"0000000000000000_0000000000000000_0010100100010011_1110001100110100"; -- 0.1604597093329172
	pesos_i(846) := b"1111111111111111_1111111111111111_1111110000000000_1110011101011100"; -- -0.0156112098263432
	pesos_i(847) := b"0000000000000000_0000000000000000_0000011000010011_0000001101101000"; -- 0.023727620031442964
	pesos_i(848) := b"0000000000000000_0000000000000000_0100000010000001_0101111100100100"; -- 0.25197405465606637
	pesos_i(849) := b"0000000000000000_0000000000000000_0000101000011001_0110101100000000"; -- 0.039450347328524954
	pesos_i(850) := b"1111111111111111_1111111111111111_1111000101101010_1000001011001001"; -- -0.056968523055268346
	pesos_i(851) := b"1111111111111111_1111111111111111_1111010010110110_1110101100111101"; -- -0.04408387920458581
	pesos_i(852) := b"1111111111111111_1111111111111111_1110110001110001_0010111001111000"; -- -0.07639798709120689
	pesos_i(853) := b"0000000000000000_0000000000000000_0001101010111011_1011111010110100"; -- 0.10442726045259992
	pesos_i(854) := b"1111111111111111_1111111111111111_1101110001010001_1111011100111111"; -- -0.1393743009566103
	pesos_i(855) := b"1111111111111111_1111111111111111_1100111110110010_0110000101110011"; -- -0.18868437714539202
	pesos_i(856) := b"0000000000000000_0000000000000000_0101110101000110_1111111010111101"; -- 0.3643645488740019
	pesos_i(857) := b"0000000000000000_0000000000000000_0011101100111111_1101011010110101"; -- 0.23144285119233984
	pesos_i(858) := b"1111111111111111_1111111111111111_1111001111111001_0011100100101010"; -- -0.046978404329393486
	pesos_i(859) := b"1111111111111111_1111111111111111_1101110000100000_0001101000000110"; -- -0.14013516760575961
	pesos_i(860) := b"0000000000000000_0000000000000000_0001010101001000_0000100011101001"; -- 0.08313041383053386
	pesos_i(861) := b"1111111111111111_1111111111111111_1110001101111000_1010110100000100"; -- -0.11143988287502586
	pesos_i(862) := b"0000000000000000_0000000000000000_0011010010100111_0100010011110001"; -- 0.2056773270491923
	pesos_i(863) := b"0000000000000000_0000000000000000_0000011000000110_0011010101110100"; -- 0.023532238802838883
	pesos_i(864) := b"1111111111111111_1111111111111111_1011100010101110_0101100110110000"; -- -0.2785896249486602
	pesos_i(865) := b"1111111111111111_1111111111111111_1110111110100101_0101100001100011"; -- -0.06388328145482573
	pesos_i(866) := b"1111111111111111_1111111111111111_1110000110111000_0111101111011111"; -- -0.1182787494407501
	pesos_i(867) := b"1111111111111111_1111111111111111_1110100111000010_1101000101100100"; -- -0.08687106423078757
	pesos_i(868) := b"0000000000000000_0000000000000000_0011011000110101_0110110000101101"; -- 0.2117526636760747
	pesos_i(869) := b"1111111111111111_1111111111111111_1101100111010010_1110000010010001"; -- -0.14912601911879922
	pesos_i(870) := b"0000000000000000_0000000000000000_0000010100011010_1111111010001010"; -- 0.019943150187681197
	pesos_i(871) := b"0000000000000000_0000000000000000_0001001101010101_0110101010111101"; -- 0.07552210905647345
	pesos_i(872) := b"1111111111111111_1111111111111111_1101011001000111_0101010110111101"; -- -0.16297401546747414
	pesos_i(873) := b"0000000000000000_0000000000000000_0011101111110101_1110010111100011"; -- 0.23422085565089873
	pesos_i(874) := b"1111111111111111_1111111111111111_1111010110010110_0011010100001111"; -- -0.040676769167969695
	pesos_i(875) := b"1111111111111111_1111111111111111_1110000101011100_0111110101101111"; -- -0.11968246498951282
	pesos_i(876) := b"0000000000000000_0000000000000000_0011000100100010_0100010111101111"; -- 0.19192921724077555
	pesos_i(877) := b"0000000000000000_0000000000000000_0001001100101111_1010001011111000"; -- 0.07494562689250217
	pesos_i(878) := b"1111111111111111_1111111111111111_1110011000111001_0110100110000010"; -- -0.10068646035620406
	pesos_i(879) := b"1111111111111111_1111111111111111_1111000111111000_1111010001000100"; -- -0.05479501098083859
	pesos_i(880) := b"0000000000000000_0000000000000000_0010111001110011_1100010000101100"; -- 0.1814539535600408
	pesos_i(881) := b"1111111111111111_1111111111111111_1110111111110010_0111010101101001"; -- -0.06270662492008158
	pesos_i(882) := b"1111111111111111_1111111111111111_1100111110001000_1010110110101100"; -- -0.18932070313728855
	pesos_i(883) := b"1111111111111111_1111111111111111_1110111000110111_0011010011110101"; -- -0.069470110140529
	pesos_i(884) := b"0000000000000000_0000000000000000_0010101101110000_0100110110101011"; -- 0.16968236369844747
	pesos_i(885) := b"1111111111111111_1111111111111111_1111101110111010_0110110001111101"; -- -0.01668664883540154
	pesos_i(886) := b"1111111111111111_1111111111111111_1110000001110001_1010111101110000"; -- -0.12326529991427608
	pesos_i(887) := b"0000000000000000_0000000000000000_0011100001110011_1001011001100100"; -- 0.22051372482491677
	pesos_i(888) := b"1111111111111111_1111111111111111_1101011110010000_1101100111100001"; -- -0.15794599783453428
	pesos_i(889) := b"1111111111111111_1111111111111111_1101110000110001_0100011100111110"; -- -0.13987307301351037
	pesos_i(890) := b"1111111111111111_1111111111111111_1111110110100101_1100110110101001"; -- -0.009188791532648358
	pesos_i(891) := b"0000000000000000_0000000000000000_0110000110011100_0000000011000110"; -- 0.38128666720978777
	pesos_i(892) := b"0000000000000000_0000000000000000_0011000110110000_1110100110111000"; -- 0.19410572755711347
	pesos_i(893) := b"1111111111111111_1111111111111111_1101111010001101_0000001101011101"; -- -0.1306608103716434
	pesos_i(894) := b"1111111111111111_1111111111111111_1111100001000101_1010001000110011"; -- -0.03018747565837193
	pesos_i(895) := b"0000000000000000_0000000000000000_0000111101110101_0101100000101101"; -- 0.060384283988692555
	pesos_i(896) := b"0000000000000000_0000000000000000_0000110111011000_1101010101110110"; -- 0.054089871651812976
	pesos_i(897) := b"1111111111111111_1111111111111111_1110010100000011_1100000111111000"; -- -0.10541141225094537
	pesos_i(898) := b"1111111111111111_1111111111111111_1110110000001000_1010001111000011"; -- -0.07799316883414838
	pesos_i(899) := b"0000000000000000_0000000000000000_0000110111011101_1001001011010010"; -- 0.05416219352700393
	pesos_i(900) := b"0000000000000000_0000000000000000_0000111000110110_1101100100110100"; -- 0.055524421024628685
	pesos_i(901) := b"0000000000000000_0000000000000000_0000000100001001_1110001001010101"; -- 0.0040570695730386425
	pesos_i(902) := b"1111111111111111_1111111111111111_1111000010111110_0100000000000110"; -- -0.05959701408109592
	pesos_i(903) := b"1111111111111111_1111111111111111_1101111101101100_0101011010100110"; -- -0.12725313610180194
	pesos_i(904) := b"1111111111111111_1111111111111111_1110111001011000_0100000110101101"; -- -0.06896581192205938
	pesos_i(905) := b"0000000000000000_0000000000000000_0010010101111000_1110101000010011"; -- 0.14637625657207967
	pesos_i(906) := b"1111111111111111_1111111111111111_1111110001011010_0101111110100100"; -- -0.014246008314085304
	pesos_i(907) := b"0000000000000000_0000000000000000_0001101001001110_1101110100101110"; -- 0.10276586881393303
	pesos_i(908) := b"0000000000000000_0000000000000000_0011001110000011_1001001111110101"; -- 0.2012264702111569
	pesos_i(909) := b"1111111111111111_1111111111111111_1110011000101100_0000010010000010"; -- -0.1008908446145905
	pesos_i(910) := b"0000000000000000_0000000000000000_0010000110001111_0010000101011111"; -- 0.1310902458408097
	pesos_i(911) := b"0000000000000000_0000000000000000_0001011011110111_0111001100010101"; -- 0.08971328031509312
	pesos_i(912) := b"0000000000000000_0000000000000000_0000100011111110_1000001101001110"; -- 0.03513355874570188
	pesos_i(913) := b"1111111111111111_1111111111111111_1111101001010010_0010101111101001"; -- -0.022183662049596726
	pesos_i(914) := b"0000000000000000_0000000000000000_0001111110011100_0010110101011000"; -- 0.1234768238489146
	pesos_i(915) := b"0000000000000000_0000000000000000_0010011011100111_1101010011101000"; -- 0.15197497041958177
	pesos_i(916) := b"0000000000000000_0000000000000000_0010001110111101_0110010000101111"; -- 0.13960863262522916
	pesos_i(917) := b"0000000000000000_0000000000000000_0010000001000011_1011100101010100"; -- 0.12603338533876637
	pesos_i(918) := b"0000000000000000_0000000000000000_0001110111110110_0000111100010001"; -- 0.11703581021680752
	pesos_i(919) := b"1111111111111111_1111111111111111_1101011101011111_1001100001000011"; -- -0.1586975895799547
	pesos_i(920) := b"1111111111111111_1111111111111111_1101111110111011_0101111010101100"; -- -0.12604721357755536
	pesos_i(921) := b"1111111111111111_1111111111111111_1110100101111100_1010111101001001"; -- -0.08794121226095064
	pesos_i(922) := b"0000000000000000_0000000000000000_0000010111000100_1000100000101111"; -- 0.022530089863186914
	pesos_i(923) := b"0000000000000000_0000000000000000_0000100000001110_0011101100111010"; -- 0.0314671531346513
	pesos_i(924) := b"0000000000000000_0000000000000000_0000011111011100_1001001100001100"; -- 0.0307094482454243
	pesos_i(925) := b"1111111111111111_1111111111111111_1110001111000111_0110101001001001"; -- -0.11023841598666904
	pesos_i(926) := b"1111111111111111_1111111111111111_1110101101101001_0001001011111111"; -- -0.08042794495880617
	pesos_i(927) := b"1111111111111111_1111111111111111_1110011000001101_1011011000010001"; -- -0.10135328384985823
	pesos_i(928) := b"0000000000000000_0000000000000000_0000110111010000_1010000110011011"; -- 0.05396471059684677
	pesos_i(929) := b"0000000000000000_0000000000000000_0000000000101001_1110001000010011"; -- 0.0006390854226211302
	pesos_i(930) := b"1111111111111111_1111111111111111_1110010100100111_1001000010000000"; -- -0.10486504426426482
	pesos_i(931) := b"0000000000000000_0000000000000000_0010111010001011_1010101010010000"; -- 0.18181863799580503
	pesos_i(932) := b"1111111111111111_1111111111111111_1111001111001001_1000100001100111"; -- -0.04770610322764605
	pesos_i(933) := b"0000000000000000_0000000000000000_0001110100011111_1101100111000100"; -- 0.11376725241517881
	pesos_i(934) := b"1111111111111111_1111111111111111_1110101101111100_1111000100110000"; -- -0.08012478416880216
	pesos_i(935) := b"0000000000000000_0000000000000000_0001110010000001_0001100100000100"; -- 0.11134487490652356
	pesos_i(936) := b"0000000000000000_0000000000000000_0010110010100010_1000110000101010"; -- 0.17435527822575175
	pesos_i(937) := b"1111111111111111_1111111111111111_1111111010010001_1100111010110010"; -- -0.005587655500888438
	pesos_i(938) := b"1111111111111111_1111111111111111_1111101101001001_0100000110010100"; -- -0.018413449697194512
	pesos_i(939) := b"0000000000000000_0000000000000000_0010101001100111_0010011011001010"; -- 0.1656364672457341
	pesos_i(940) := b"1111111111111111_1111111111111111_1110011101010001_1001011101010101"; -- -0.09641126798753775
	pesos_i(941) := b"1111111111111111_1111111111111111_1101111101010111_0101100001000001"; -- -0.1275734749446981
	pesos_i(942) := b"0000000000000000_0000000000000000_0001111111010100_0100101100010010"; -- 0.12433308782508107
	pesos_i(943) := b"1111111111111111_1111111111111111_1101011101001010_1001111101111011"; -- -0.15901759374096963
	pesos_i(944) := b"1111111111111111_1111111111111111_1111110110000100_0000010000110101"; -- -0.00970433901823644
	pesos_i(945) := b"0000000000000000_0000000000000000_0001001011111011_1111011101010010"; -- 0.0741571974692554
	pesos_i(946) := b"0000000000000000_0000000000000000_0000001000101111_0010001001000110"; -- 0.00853170587862896
	pesos_i(947) := b"1111111111111111_1111111111111111_1110110101010100_0010011011101001"; -- -0.07293469255633667
	pesos_i(948) := b"1111111111111111_1111111111111111_1110110001101011_1001011011000111"; -- -0.0764833224597649
	pesos_i(949) := b"0000000000000000_0000000000000000_0000001100010101_0110011100100111"; -- 0.012045332861857539
	pesos_i(950) := b"1111111111111111_1111111111111111_1111011000011000_0001100001010110"; -- -0.038694838572338006
	pesos_i(951) := b"1111111111111111_1111111111111111_1110001111010100_0100111110010111"; -- -0.11004164277643351
	pesos_i(952) := b"1111111111111111_1111111111111111_1100000000110000_1010101010100010"; -- -0.24925740767115295
	pesos_i(953) := b"1111111111111111_1111111111111111_1110010100111111_0100010111110110"; -- -0.10450327620160581
	pesos_i(954) := b"0000000000000000_0000000000000000_0010100001010111_1110101000011111"; -- 0.1575914694305104
	pesos_i(955) := b"0000000000000000_0000000000000000_0000001110101110_0100001100111101"; -- 0.014377787049420587
	pesos_i(956) := b"0000000000000000_0000000000000000_0001001010010010_0011110001110010"; -- 0.0725438860988442
	pesos_i(957) := b"1111111111111111_1111111111111111_1110101001011110_1100000010001000"; -- -0.08449169814811228
	pesos_i(958) := b"1111111111111111_1111111111111111_1111101100010100_0100011010101111"; -- -0.019221861123735
	pesos_i(959) := b"0000000000000000_0000000000000000_0001110000101000_1100100011110011"; -- 0.10999732913586732
	pesos_i(960) := b"0000000000000000_0000000000000000_0001101001100001_0001100011000100"; -- 0.10304407860542443
	pesos_i(961) := b"0000000000000000_0000000000000000_0000101100001001_0111101110100101"; -- 0.04311344891641528
	pesos_i(962) := b"1111111111111111_1111111111111111_1110101101101111_0111110010011110"; -- -0.08033009671842735
	pesos_i(963) := b"1111111111111111_1111111111111111_1100111000001000_0111010011001101"; -- -0.19518346785232
	pesos_i(964) := b"0000000000000000_0000000000000000_0001011111011011_1101000000110001"; -- 0.09319783401945608
	pesos_i(965) := b"1111111111111111_1111111111111111_1110011100011000_1001011001011010"; -- -0.09728107740475896
	pesos_i(966) := b"1111111111111111_1111111111111111_1101011010101101_0000000100011100"; -- -0.16142266347504763
	pesos_i(967) := b"1111111111111111_1111111111111111_1101101011011111_0000011010001110"; -- -0.14503439927060932
	pesos_i(968) := b"1111111111111111_1111111111111111_1111111001101100_0011101110101101"; -- -0.006160993730725348
	pesos_i(969) := b"0000000000000000_0000000000000000_0010100000111111_0111001110110001"; -- 0.15721819940159412
	pesos_i(970) := b"1111111111111111_1111111111111111_1101110001101110_0101000011010111"; -- -0.1389417147236991
	pesos_i(971) := b"0000000000000000_0000000000000000_0010000100011110_1011110001000111"; -- 0.12937523588697059
	pesos_i(972) := b"0000000000000000_0000000000000000_0010000010110010_0011110110000101"; -- 0.12771973122556562
	pesos_i(973) := b"1111111111111111_1111111111111111_1111111000101010_0110001001000111"; -- -0.007165773024311174
	pesos_i(974) := b"1111111111111111_1111111111111111_1111011011001100_1001011101111011"; -- -0.03594067811560509
	pesos_i(975) := b"1111111111111111_1111111111111111_1111101110100001_0110000110010110"; -- -0.017068768430172392
	pesos_i(976) := b"1111111111111111_1111111111111111_1101101000110001_0001100101011001"; -- -0.1476883085354258
	pesos_i(977) := b"0000000000000000_0000000000000000_0010101101110101_1011100001110000"; -- 0.1697650216676266
	pesos_i(978) := b"1111111111111111_1111111111111111_1110011101110101_0001000001000111"; -- -0.09587000147142505
	pesos_i(979) := b"0000000000000000_0000000000000000_0001100111011001_0001011110011001"; -- 0.10096881374705516
	pesos_i(980) := b"0000000000000000_0000000000000000_0001001101011001_1000101001100101"; -- 0.07558503128806278
	pesos_i(981) := b"1111111111111111_1111111111111111_1110101110001000_1010011101000011"; -- -0.07994608515138893
	pesos_i(982) := b"1111111111111111_1111111111111111_1101010110101110_0111010110110101"; -- -0.16530670484036686
	pesos_i(983) := b"1111111111111111_1111111111111111_1101000010100010_1101110101000110"; -- -0.18501488726566923
	pesos_i(984) := b"1111111111111111_1111111111111111_1101100001011000_1111100100111011"; -- -0.15489237134065376
	pesos_i(985) := b"1111111111111111_1111111111111111_1101010010010000_0000100011101011"; -- -0.16967720293365585
	pesos_i(986) := b"1111111111111111_1111111111111111_1111011000010101_1100001011000100"; -- -0.038730456570982355
	pesos_i(987) := b"0000000000000000_0000000000000000_0010000001110111_1111010010000111"; -- 0.12683037089219798
	pesos_i(988) := b"1111111111111111_1111111111111111_1111110101001100_0010000001101001"; -- -0.01055715031603362
	pesos_i(989) := b"1111111111111111_1111111111111111_1101110110000101_0010000000100100"; -- -0.13468741526420291
	pesos_i(990) := b"0000000000000000_0000000000000000_0001110010001111_1100111010101111"; -- 0.11156932613059393
	pesos_i(991) := b"1111111111111111_1111111111111111_1111110110010111_1110100010100001"; -- -0.009400807109048611
	pesos_i(992) := b"1111111111111111_1111111111111111_1101010100110010_1110000000001110"; -- -0.16719245583457565
	pesos_i(993) := b"0000000000000000_0000000000000000_0000000001010011_1111111011011011"; -- 0.0012816701602736255
	pesos_i(994) := b"1111111111111111_1111111111111111_1111010000101111_0100110100111100"; -- -0.04615323340965985
	pesos_i(995) := b"0000000000000000_0000000000000000_0000111000000101_1101010100110000"; -- 0.05477650091776303
	pesos_i(996) := b"0000000000000000_0000000000000000_0001111010101100_1000001001110111"; -- 0.11981978791571446
	pesos_i(997) := b"1111111111111111_1111111111111111_1110100101010001_1111101110010110"; -- -0.08859279233694871
	pesos_i(998) := b"1111111111111111_1111111111111111_1101010001100001_0000011001110110"; -- -0.1703945122831376
	pesos_i(999) := b"0000000000000000_0000000000000000_0010100101000001_1100101100100011"; -- 0.16116017928735157
	pesos_i(1000) := b"0000000000000000_0000000000000000_0000101000111000_1010010110110011"; -- 0.039926868531219184
	pesos_i(1001) := b"1111111111111111_1111111111111111_1110111101101001_1100001001101001"; -- -0.06479248936134
	pesos_i(1002) := b"1111111111111111_1111111111111111_1101000000110100_1110100110000001"; -- -0.18669262494845193
	pesos_i(1003) := b"0000000000000000_0000000000000000_0001010110010100_1001001001011100"; -- 0.08429827448447128
	pesos_i(1004) := b"0000000000000000_0000000000000000_0010110011010010_0111101001111011"; -- 0.17508664610038535
	pesos_i(1005) := b"1111111111111111_1111111111111111_1111101101110011_1001110100010010"; -- -0.01776712725110558
	pesos_i(1006) := b"0000000000000000_0000000000000000_0000000000001010_0010011000100100"; -- 0.00015486123904500428
	pesos_i(1007) := b"1111111111111111_1111111111111111_1111100000111111_0101101011001001"; -- -0.030283285104282943
	pesos_i(1008) := b"0000000000000000_0000000000000000_0001010010110000_0110000000111000"; -- 0.08081628196345358
	pesos_i(1009) := b"0000000000000000_0000000000000000_0010000100010101_1101110100001010"; -- 0.12923985952293937
	pesos_i(1010) := b"1111111111111111_1111111111111111_1111101111000001_0001001111000100"; -- -0.01658512556679329
	pesos_i(1011) := b"1111111111111111_1111111111111111_1110011101111110_1011110000100000"; -- -0.09572242952705667
	pesos_i(1012) := b"0000000000000000_0000000000000000_0001000000011001_1111001101001111"; -- 0.062895972072153
	pesos_i(1013) := b"0000000000000000_0000000000000000_0010101100001000_0010110011011110"; -- 0.16809349469710957
	pesos_i(1014) := b"0000000000000000_0000000000000000_0010100000000110_1100111011100100"; -- 0.15635388441620351
	pesos_i(1015) := b"0000000000000000_0000000000000000_0001011010010110_0011111000010000"; -- 0.08823001768377384
	pesos_i(1016) := b"1111111111111111_1111111111111111_1111111100111011_1110101101111100"; -- -0.0029919453993258894
	pesos_i(1017) := b"1111111111111111_1111111111111111_1111111010010101_0010110010000011"; -- -0.005536287300305675
	pesos_i(1018) := b"0000000000000000_0000000000000000_0001001001100000_0010001010101011"; -- 0.071779410060635
	pesos_i(1019) := b"0000000000000000_0000000000000000_0010110010011010_1110010100001110"; -- 0.1742385062755094
	pesos_i(1020) := b"1111111111111111_1111111111111111_1110111101011101_1011001011011011"; -- -0.06497652204838167
	pesos_i(1021) := b"1111111111111111_1111111111111111_1111001110011110_1001111110100011"; -- -0.048360846311469044
	pesos_i(1022) := b"1111111111111111_1111111111111111_1110111001011101_1111110111101110"; -- -0.06887829724363373
	pesos_i(1023) := b"1111111111111111_1111111111111111_1101010101001010_0111000101010010"; -- -0.1668328450822599
	pesos_i(1024) := b"1111111111111111_1111111111111111_1111101110000000_0100101000011000"; -- -0.017573708740257505
	pesos_i(1025) := b"0000000000000000_0000000000000000_0010001001000101_1011000100100110"; -- 0.1338759152426841
	pesos_i(1026) := b"0000000000000000_0000000000000000_0001000010101110_0110001010000100"; -- 0.06516090117008427
	pesos_i(1027) := b"1111111111111111_1111111111111111_1111001010101111_1110001111100001"; -- -0.052003629349450686
	pesos_i(1028) := b"0000000000000000_0000000000000000_0000101110001100_0000101010011000"; -- 0.04510561180709961
	pesos_i(1029) := b"1111111111111111_1111111111111111_1110011110001110_0000010111011101"; -- -0.09548915253629053
	pesos_i(1030) := b"0000000000000000_0000000000000000_0001011001001101_1001001110001001"; -- 0.08712122059947883
	pesos_i(1031) := b"1111111111111111_1111111111111111_1110111101000010_1111011001010011"; -- -0.06538448777563068
	pesos_i(1032) := b"0000000000000000_0000000000000000_0000011011101100_0011011100110100"; -- 0.027041864696011688
	pesos_i(1033) := b"0000000000000000_0000000000000000_0010000101100001_1110100001100101"; -- 0.13040020437003746
	pesos_i(1034) := b"0000000000000000_0000000000000000_0010001011000001_1001000001100000"; -- 0.13576605165878214
	pesos_i(1035) := b"1111111111111111_1111111111111111_1110101001000000_0110100101100001"; -- -0.08495465645800547
	pesos_i(1036) := b"0000000000000000_0000000000000000_0000001010101001_0101100010000110"; -- 0.010396511649315652
	pesos_i(1037) := b"0000000000000000_0000000000000000_0000111110010001_0110110111000110"; -- 0.060812817305775264
	pesos_i(1038) := b"1111111111111111_1111111111111111_1110110011100001_0111100111111101"; -- -0.07468450142739995
	pesos_i(1039) := b"1111111111111111_1111111111111111_1110000101101110_0110101000100101"; -- -0.11940895655697174
	pesos_i(1040) := b"1111111111111111_1111111111111111_1111111010001110_0010100010111100"; -- -0.0056433239537065595
	pesos_i(1041) := b"1111111111111111_1111111111111111_1111111011000101_1100010000111101"; -- -0.004794821733780583
	pesos_i(1042) := b"1111111111111111_1111111111111111_1101110000101010_1110011000100100"; -- -0.13997041333596377
	pesos_i(1043) := b"0000000000000000_0000000000000000_0010001101000101_0011110110101110"; -- 0.13777528274048056
	pesos_i(1044) := b"1111111111111111_1111111111111111_1111000010111010_1100111001001110"; -- -0.05964956848353861
	pesos_i(1045) := b"0000000000000000_0000000000000000_0010010010100000_1100111001101001"; -- 0.14307870933695463
	pesos_i(1046) := b"1111111111111111_1111111111111111_1111001101101100_0100110010011000"; -- -0.049128735514708755
	pesos_i(1047) := b"0000000000000000_0000000000000000_0010001111111100_0001100101000100"; -- 0.140565470709839
	pesos_i(1048) := b"0000000000000000_0000000000000000_0000011011100001_0101000010000101"; -- 0.02687552685047454
	pesos_i(1049) := b"0000000000000000_0000000000000000_0000110010110000_1011000011110111"; -- 0.04957109484955247
	pesos_i(1050) := b"0000000000000000_0000000000000000_0001111010010111_1110110001100111"; -- 0.11950566779663745
	pesos_i(1051) := b"0000000000000000_0000000000000000_0001010100011000_0100110001101110"; -- 0.08240201639058578
	pesos_i(1052) := b"1111111111111111_1111111111111111_1110001010110110_0111111010010100"; -- -0.11440285574381705
	pesos_i(1053) := b"1111111111111111_1111111111111111_1101011001011100_0100000101011001"; -- -0.16265479629011118
	pesos_i(1054) := b"0000000000000000_0000000000000000_0000011100100001_0011011000100000"; -- 0.02785051606593185
	pesos_i(1055) := b"1111111111111111_1111111111111111_1101000001101100_1010011000000011"; -- -0.1858421556228057
	pesos_i(1056) := b"1111111111111111_1111111111111111_1110111110001010_0011010011101110"; -- -0.06429738222575183
	pesos_i(1057) := b"1111111111111111_1111111111111111_1111010110101110_1100101011100100"; -- -0.0403016275160954
	pesos_i(1058) := b"1111111111111111_1111111111111111_1111011111111001_0010001011011001"; -- -0.03135473447127987
	pesos_i(1059) := b"1111111111111111_1111111111111111_1111000011101110_0100110000010101"; -- -0.058863873428451396
	pesos_i(1060) := b"1111111111111111_1111111111111111_1110001100100100_1001101000100011"; -- -0.11272274628985339
	pesos_i(1061) := b"0000000000000000_0000000000000000_0001110110010000_1101110011101000"; -- 0.11549168263418719
	pesos_i(1062) := b"1111111111111111_1111111111111111_1110011001110100_0011100110101010"; -- -0.09978904351824681
	pesos_i(1063) := b"0000000000000000_0000000000000000_0001100000000011_1110001000110110"; -- 0.09380925951253691
	pesos_i(1064) := b"0000000000000000_0000000000000000_0001101101100010_1000001110111011"; -- 0.10697196301328336
	pesos_i(1065) := b"1111111111111111_1111111111111111_1111110011100111_1001000001110000"; -- -0.012091610549248451
	pesos_i(1066) := b"0000000000000000_0000000000000000_0010000011001010_1001000110110111"; -- 0.12809096068028725
	pesos_i(1067) := b"0000000000000000_0000000000000000_0001101101100001_0011000000011000"; -- 0.10695171908894925
	pesos_i(1068) := b"1111111111111111_1111111111111111_1101111011000100_1001011010011000"; -- -0.12981280117150248
	pesos_i(1069) := b"1111111111111111_1111111111111111_1111010100110010_1100100011100111"; -- -0.04219383585513706
	pesos_i(1070) := b"1111111111111111_1111111111111111_1110001000111010_1011100011000100"; -- -0.11629147732076844
	pesos_i(1071) := b"1111111111111111_1111111111111111_1110111111100110_1111011101001100"; -- -0.06288198838412387
	pesos_i(1072) := b"1111111111111111_1111111111111111_1111001111010001_1101010100010000"; -- -0.047579463650167686
	pesos_i(1073) := b"0000000000000000_0000000000000000_0001001000111111_0011100010010000"; -- 0.07127717506584898
	pesos_i(1074) := b"0000000000000000_0000000000000000_0010001011001010_1010110001011100"; -- 0.13590504869532
	pesos_i(1075) := b"1111111111111111_1111111111111111_1111100011010000_0110100101011000"; -- -0.028069892860289988
	pesos_i(1076) := b"0000000000000000_0000000000000000_0001000111000010_0100010010011100"; -- 0.06937054443111904
	pesos_i(1077) := b"1111111111111111_1111111111111111_1111100000011101_1000010010111000"; -- -0.030799584515722768
	pesos_i(1078) := b"1111111111111111_1111111111111111_1110000101011111_1111101100100101"; -- -0.119629195758838
	pesos_i(1079) := b"0000000000000000_0000000000000000_0000001011111000_1101111111010100"; -- 0.01161002091996893
	pesos_i(1080) := b"1111111111111111_1111111111111111_1111100000110001_1110001111100100"; -- -0.03048873591861743
	pesos_i(1081) := b"0000000000000000_0000000000000000_0000001010000110_0110001110011111"; -- 0.009863115602280158
	pesos_i(1082) := b"1111111111111111_1111111111111111_1111001100001111_0011110001110001"; -- -0.05054876550737709
	pesos_i(1083) := b"0000000000000000_0000000000000000_0000010100010010_0010000100111010"; -- 0.019807888705636406
	pesos_i(1084) := b"1111111111111111_1111111111111111_1101101010000010_1100010000010101"; -- -0.14644217008643762
	pesos_i(1085) := b"1111111111111111_1111111111111111_1111101001100100_1101000001000001"; -- -0.02189920828440572
	pesos_i(1086) := b"0000000000000000_0000000000000000_0001111011110011_1011100001011101"; -- 0.12090637468159508
	pesos_i(1087) := b"0000000000000000_0000000000000000_0010110011000010_1000111001110011"; -- 0.17484369580554637
	pesos_i(1088) := b"0000000000000000_0000000000000000_0000110001100010_0111110010101110"; -- 0.04837779275149017
	pesos_i(1089) := b"1111111111111111_1111111111111111_1110000100000000_1010010101011101"; -- -0.12108389353452495
	pesos_i(1090) := b"1111111111111111_1111111111111111_1101111110100100_1110000011010011"; -- -0.12639040792747563
	pesos_i(1091) := b"0000000000000000_0000000000000000_0010111101110011_1101110110110001"; -- 0.1853617246757321
	pesos_i(1092) := b"1111111111111111_1111111111111111_1110101001100110_1100010001111010"; -- -0.08436939255914926
	pesos_i(1093) := b"0000000000000000_0000000000000000_0000010001100000_0011100010010101"; -- 0.0170932163473352
	pesos_i(1094) := b"1111111111111111_1111111111111111_1101101111100001_1001001111110010"; -- -0.141089204138043
	pesos_i(1095) := b"1111111111111111_1111111111111111_1110001010110001_1100001000001001"; -- -0.11447512884186221
	pesos_i(1096) := b"1111111111111111_1111111111111111_1110101100111110_0111000101010011"; -- -0.08107845038473685
	pesos_i(1097) := b"1111111111111111_1111111111111111_1111101100011001_1101111100011100"; -- -0.019136481907331887
	pesos_i(1098) := b"1111111111111111_1111111111111111_1101100011010101_0000110111000101"; -- -0.1529990573079779
	pesos_i(1099) := b"0000000000000000_0000000000000000_0010011001010000_0101010001101111"; -- 0.14966323570970988
	pesos_i(1100) := b"1111111111111111_1111111111111111_1111110000011000_1111010011001110"; -- -0.01524419752195783
	pesos_i(1101) := b"1111111111111111_1111111111111111_1100110100111100_1011101000100000"; -- -0.19829212871146767
	pesos_i(1102) := b"1111111111111111_1111111111111111_1100111010000010_0011001111111000"; -- -0.1933257598939817
	pesos_i(1103) := b"0000000000000000_0000000000000000_0001111111000100_1001000110111111"; -- 0.12409315969969618
	pesos_i(1104) := b"1111111111111111_1111111111111111_1110101001010011_1110100001000110"; -- -0.08465717590459833
	pesos_i(1105) := b"1111111111111111_1111111111111111_1110000000010011_0000000011010101"; -- -0.1247100334237039
	pesos_i(1106) := b"1111111111111111_1111111111111111_1110111111010000_0110010011111000"; -- -0.06322640375740125
	pesos_i(1107) := b"0000000000000000_0000000000000000_0000100011111000_1100000110011110"; -- 0.03504572008456968
	pesos_i(1108) := b"1111111111111111_1111111111111111_1110001001000000_0010110000011101"; -- -0.11620830806430539
	pesos_i(1109) := b"1111111111111111_1111111111111111_1101110011000101_1101001010000111"; -- -0.13760647011673938
	pesos_i(1110) := b"0000000000000000_0000000000000000_0010011010010111_1110101011110110"; -- 0.15075558199565042
	pesos_i(1111) := b"1111111111111111_1111111111111111_1111000010110001_0000001001100100"; -- -0.05979905190161727
	pesos_i(1112) := b"1111111111111111_1111111111111111_1110001011000100_0000000111100011"; -- -0.11419666478980912
	pesos_i(1113) := b"1111111111111111_1111111111111111_1110000011010101_1101000111111010"; -- -0.12173736237213581
	pesos_i(1114) := b"0000000000000000_0000000000000000_0001001011001011_1110111000000011"; -- 0.07342422087512018
	pesos_i(1115) := b"1111111111111111_1111111111111111_1101111011011110_0000011101110011"; -- -0.129424604774253
	pesos_i(1116) := b"0000000000000000_0000000000000000_0010010000010000_1100010001010000"; -- 0.1408808417636294
	pesos_i(1117) := b"1111111111111111_1111111111111111_1111011001101101_1010010110111100"; -- -0.0373894133717196
	pesos_i(1118) := b"0000000000000000_0000000000000000_0000111011010010_0111110000100100"; -- 0.057899245072498266
	pesos_i(1119) := b"1111111111111111_1111111111111111_1111001000110110_0001000101100001"; -- -0.05386248962058111
	pesos_i(1120) := b"0000000000000000_0000000000000000_0011000001110111_0010011100101111"; -- 0.1893181313499338
	pesos_i(1121) := b"0000000000000000_0000000000000000_0000000101010101_1010010101110000"; -- 0.005213107808418855
	pesos_i(1122) := b"1111111111111111_1111111111111111_1101111010011011_1101001011111110"; -- -0.1304348116826108
	pesos_i(1123) := b"0000000000000000_0000000000000000_0000100001000010_0111010000000001"; -- 0.03226399455697021
	pesos_i(1124) := b"0000000000000000_0000000000000000_0000100011011011_0010001010000010"; -- 0.034593731648561325
	pesos_i(1125) := b"0000000000000000_0000000000000000_0000110000001011_0101011111101011"; -- 0.04704808689112678
	pesos_i(1126) := b"0000000000000000_0000000000000000_0010111001101001_1100000010100011"; -- 0.18130115477845038
	pesos_i(1127) := b"1111111111111111_1111111111111111_1110010101000101_0101111110011100"; -- -0.10441019488646516
	pesos_i(1128) := b"1111111111111111_1111111111111111_1110111110111100_0011111100110000"; -- -0.06353383136432285
	pesos_i(1129) := b"1111111111111111_1111111111111111_1101110000001101_0011010111111101"; -- -0.14042341779984613
	pesos_i(1130) := b"0000000000000000_0000000000000000_0001110011000101_1010001111000110"; -- 0.11239074309811067
	pesos_i(1131) := b"0000000000000000_0000000000000000_0000010110111110_0000111011100101"; -- 0.022431307655004836
	pesos_i(1132) := b"0000000000000000_0000000000000000_0000001001010000_0111100110100011"; -- 0.009040453222223091
	pesos_i(1133) := b"0000000000000000_0000000000000000_0010011000110011_1011111011000001"; -- 0.14922706809636596
	pesos_i(1134) := b"0000000000000000_0000000000000000_0001111110000110_0110100000100001"; -- 0.12314463427757932
	pesos_i(1135) := b"0000000000000000_0000000000000000_0000101110010010_1001110101001100"; -- 0.04520590872418496
	pesos_i(1136) := b"0000000000000000_0000000000000000_0001001011011101_1011001010011011"; -- 0.07369533811552252
	pesos_i(1137) := b"1111111111111111_1111111111111111_1110110100111100_0000011110101111"; -- -0.07330276476526001
	pesos_i(1138) := b"1111111111111111_1111111111111111_1111010100010100_0101001000111001"; -- -0.04265867338081075
	pesos_i(1139) := b"1111111111111111_1111111111111111_1101111011110110_0011100001110000"; -- -0.1290554739553762
	pesos_i(1140) := b"0000000000000000_0000000000000000_0001001101110101_0011110100011010"; -- 0.07600767033691765
	pesos_i(1141) := b"1111111111111111_1111111111111111_1111001110000111_1011011000111110"; -- -0.048710451047129344
	pesos_i(1142) := b"0000000000000000_0000000000000000_0000011011111100_1100100110001000"; -- 0.027294726993445872
	pesos_i(1143) := b"0000000000000000_0000000000000000_0010011010111110_1001000000001001"; -- 0.1513452550652324
	pesos_i(1144) := b"1111111111111111_1111111111111111_1111100001011111_1001011111001111"; -- -0.029791366574999752
	pesos_i(1145) := b"0000000000000000_0000000000000000_0000110110000011_0011110001111100"; -- 0.05278375659058613
	pesos_i(1146) := b"1111111111111111_1111111111111111_1101101011000110_0011100001111100"; -- -0.14541289302059407
	pesos_i(1147) := b"0000000000000000_0000000000000000_0001001111011000_0010110000110111"; -- 0.07751728391970146
	pesos_i(1148) := b"0000000000000000_0000000000000000_0000101000100011_1001110000000110"; -- 0.03960585723659202
	pesos_i(1149) := b"1111111111111111_1111111111111111_1111110010111111_0111100101110010"; -- -0.012703332496479397
	pesos_i(1150) := b"0000000000000000_0000000000000000_0010011100010110_0100010110110001"; -- 0.1526835973637648
	pesos_i(1151) := b"0000000000000000_0000000000000000_0000111100010001_1000111101111100"; -- 0.058861701827660984
	pesos_i(1152) := b"0000000000000000_0000000000000000_0010111000100100_0000111110001111"; -- 0.1802377437471374
	pesos_i(1153) := b"1111111111111111_1111111111111111_1110000100100011_1000101100001110"; -- -0.12055140396404615
	pesos_i(1154) := b"1111111111111111_1111111111111111_1111010000110011_0101011001011101"; -- -0.04609165406880106
	pesos_i(1155) := b"1111111111111111_1111111111111111_1101000000000111_1101101110111000"; -- -0.18738009231034958
	pesos_i(1156) := b"0000000000000000_0000000000000000_0000011111001010_1100100111011011"; -- 0.03043805699089029
	pesos_i(1157) := b"0000000000000000_0000000000000000_0010000111000111_0111111011001011"; -- 0.13195030640078212
	pesos_i(1158) := b"1111111111111111_1111111111111111_1101001001010111_0000010110101111"; -- -0.17835964657473666
	pesos_i(1159) := b"1111111111111111_1111111111111111_1110100111001101_0001110101001100"; -- -0.0867139519549987
	pesos_i(1160) := b"1111111111111111_1111111111111111_1101011101110011_1101000001110110"; -- -0.1583890639404641
	pesos_i(1161) := b"0000000000000000_0000000000000000_0000000111001010_0011110101001101"; -- 0.006992179119181924
	pesos_i(1162) := b"1111111111111111_1111111111111111_1111110110101010_0011001110101101"; -- -0.00912167568138534
	pesos_i(1163) := b"0000000000000000_0000000000000000_0000101010011111_0111110010001110"; -- 0.04149607140668297
	pesos_i(1164) := b"0000000000000000_0000000000000000_0001010100100101_1101010001111000"; -- 0.08260848932112484
	pesos_i(1165) := b"0000000000000000_0000000000000000_0010000110001111_0000001010001110"; -- 0.13108840902854918
	pesos_i(1166) := b"1111111111111111_1111111111111111_1101010111101001_1001101101110100"; -- -0.16440418643859694
	pesos_i(1167) := b"0000000000000000_0000000000000000_0001000110100101_0101101010000110"; -- 0.06892934571526452
	pesos_i(1168) := b"1111111111111111_1111111111111111_1101110101010111_0111010001111101"; -- -0.13538429218754544
	pesos_i(1169) := b"0000000000000000_0000000000000000_0000001110110000_0110011010000110"; -- 0.014410407675130153
	pesos_i(1170) := b"1111111111111111_1111111111111111_1101110001111000_0101001111000000"; -- -0.13878895337233607
	pesos_i(1171) := b"0000000000000000_0000000000000000_0000111000001010_0001011000110100"; -- 0.0548414114099905
	pesos_i(1172) := b"0000000000000000_0000000000000000_0001101100100111_0101000001000110"; -- 0.10606862736523145
	pesos_i(1173) := b"1111111111111111_1111111111111111_1111001111110110_1000011000001111"; -- -0.04701959730762972
	pesos_i(1174) := b"1111111111111111_1111111111111111_1110100010001010_1111111011010011"; -- -0.09162909842273197
	pesos_i(1175) := b"1111111111111111_1111111111111111_1111110110000101_0000101101100011"; -- -0.009688652394409757
	pesos_i(1176) := b"0000000000000000_0000000000000000_0001000110010000_0000010001101000"; -- 0.06860377814292654
	pesos_i(1177) := b"1111111111111111_1111111111111111_1110000101101110_1000111010111010"; -- -0.11940677614674802
	pesos_i(1178) := b"1111111111111111_1111111111111111_1100110000101001_1000101100101101"; -- -0.20249109416349323
	pesos_i(1179) := b"1111111111111111_1111111111111111_1111100011000111_0010010000010101"; -- -0.028211350404382385
	pesos_i(1180) := b"0000000000000000_0000000000000000_0000100010011000_0010111011110111"; -- 0.03357213525969846
	pesos_i(1181) := b"1111111111111111_1111111111111111_1111100011011100_1110110100000110"; -- -0.027878938688408992
	pesos_i(1182) := b"0000000000000000_0000000000000000_0001011010111111_1110011011111101"; -- 0.08886569673748691
	pesos_i(1183) := b"1111111111111111_1111111111111111_1101100111111101_0110111000101100"; -- -0.14847670951859046
	pesos_i(1184) := b"1111111111111111_1111111111111111_1111100111100100_0001011100110000"; -- -0.02386336405467459
	pesos_i(1185) := b"1111111111111111_1111111111111111_1110001101101100_0110011111000010"; -- -0.11162711629332418
	pesos_i(1186) := b"1111111111111111_1111111111111111_1110110101000110_1100111011000010"; -- -0.0731383109577483
	pesos_i(1187) := b"0000000000000000_0000000000000000_0001101111110110_1011001101111010"; -- 0.10923310984434509
	pesos_i(1188) := b"1111111111111111_1111111111111111_1110110100111111_1001001111010001"; -- -0.07324863577828976
	pesos_i(1189) := b"1111111111111111_1111111111111111_1111001111011101_0110110110000010"; -- -0.04740253050178981
	pesos_i(1190) := b"1111111111111111_1111111111111111_1110001111101000_0000111001010010"; -- -0.10974035741357734
	pesos_i(1191) := b"1111111111111111_1111111111111111_1110001000011100_1011111101110111"; -- -0.11674884175859185
	pesos_i(1192) := b"1111111111111111_1111111111111111_1111000010101111_0000010101111001"; -- -0.059829385815950854
	pesos_i(1193) := b"0000000000000000_0000000000000000_0001100001001001_0010111110100011"; -- 0.09486673097461687
	pesos_i(1194) := b"0000000000000000_0000000000000000_0000101100010100_0100111110011101"; -- 0.04327867100682367
	pesos_i(1195) := b"1111111111111111_1111111111111111_1111101101000100_0011000011001000"; -- -0.018490744650012814
	pesos_i(1196) := b"1111111111111111_1111111111111111_1101100011101101_1100010111111101"; -- -0.15262186590439342
	pesos_i(1197) := b"1111111111111111_1111111111111111_1101101110001001_1101111001100000"; -- -0.14242754124062493
	pesos_i(1198) := b"0000000000000000_0000000000000000_0010101001001111_1110000001001011"; -- 0.16528131322568215
	pesos_i(1199) := b"0000000000000000_0000000000000000_0001010111110011_0000000111011110"; -- 0.08573924713567338
	pesos_i(1200) := b"0000000000000000_0000000000000000_0010001010010000_0011010110111001"; -- 0.13501296777544466
	pesos_i(1201) := b"0000000000000000_0000000000000000_0010110100000010_1011111110010001"; -- 0.17582318576167613
	pesos_i(1202) := b"1111111111111111_1111111111111111_1111111100000001_0011100111001110"; -- -0.0038875458065319663
	pesos_i(1203) := b"0000000000000000_0000000000000000_0001010001110001_0011001110101011"; -- 0.0798523228383899
	pesos_i(1204) := b"1111111111111111_1111111111111111_1101010111110100_0100110111111001"; -- -0.1642409578992805
	pesos_i(1205) := b"0000000000000000_0000000000000000_0001000111010001_1110101010101000"; -- 0.06960932358630824
	pesos_i(1206) := b"0000000000000000_0000000000000000_0001101100100011_0010111101111001"; -- 0.10600563726635892
	pesos_i(1207) := b"0000000000000000_0000000000000000_0010000110111101_1100010101110000"; -- 0.13180192941399937
	pesos_i(1208) := b"1111111111111111_1111111111111111_1111011111001011_0001001101100111"; -- -0.032057559381668786
	pesos_i(1209) := b"0000000000000000_0000000000000000_0001000100011111_1001100100111101"; -- 0.06688840628056505
	pesos_i(1210) := b"0000000000000000_0000000000000000_0010011000101001_0001011100010101"; -- 0.14906448603466943
	pesos_i(1211) := b"1111111111111111_1111111111111111_1111101000000011_0100011100100100"; -- -0.023387483237617107
	pesos_i(1212) := b"0000000000000000_0000000000000000_0000011000101011_1111111001111110"; -- 0.02410879694980521
	pesos_i(1213) := b"1111111111111111_1111111111111111_1101111110100100_0110010000110110"; -- -0.12639783556641457
	pesos_i(1214) := b"0000000000000000_0000000000000000_0010101100010110_0101010001110100"; -- 0.16830947725850012
	pesos_i(1215) := b"0000000000000000_0000000000000000_0000110101111100_1101100001000110"; -- 0.05268623085954895
	pesos_i(1216) := b"0000000000000000_0000000000000000_0000111001110010_1101011011101010"; -- 0.05643981193117767
	pesos_i(1217) := b"1111111111111111_1111111111111111_1111001010000101_1000011000100010"; -- -0.052650086212308406
	pesos_i(1218) := b"0000000000000000_0000000000000000_0000011010000111_1001010100010100"; -- 0.025506322195704225
	pesos_i(1219) := b"0000000000000000_0000000000000000_0000011001110010_0101110000010010"; -- 0.025182489870778015
	pesos_i(1220) := b"1111111111111111_1111111111111111_1110011100010101_0111010010010111"; -- -0.09732886604941468
	pesos_i(1221) := b"1111111111111111_1111111111111111_1100110100100010_0000011100111000"; -- -0.19869952089641746
	pesos_i(1222) := b"1111111111111111_1111111111111111_1110010000101110_1000000011010010"; -- -0.10866541734405287
	pesos_i(1223) := b"1111111111111111_1111111111111111_1111101111100111_0110100110111111"; -- -0.016000166869215172
	pesos_i(1224) := b"1111111111111111_1111111111111111_1110110010100110_0110001100010001"; -- -0.07558613615558138
	pesos_i(1225) := b"1111111111111111_1111111111111111_1101000000100010_0110011110111010"; -- -0.18697501856702417
	pesos_i(1226) := b"0000000000000000_0000000000000000_0001010000001110_0101011010010001"; -- 0.07834378279241117
	pesos_i(1227) := b"0000000000000000_0000000000000000_0001010100011111_1000000111010011"; -- 0.08251201054621507
	pesos_i(1228) := b"0000000000000000_0000000000000000_0001111110011000_0011000111100100"; -- 0.12341605976420456
	pesos_i(1229) := b"0000000000000000_0000000000000000_0010110010111101_1110000010101100"; -- 0.1747723027357845
	pesos_i(1230) := b"0000000000000000_0000000000000000_0001010100010110_0101000011011111"; -- 0.08237176354452617
	pesos_i(1231) := b"0000000000000000_0000000000000000_0010010110101101_0010010001101010"; -- 0.14717319106304197
	pesos_i(1232) := b"1111111111111111_1111111111111111_1110011010101110_1000110001011110"; -- -0.0988991041842174
	pesos_i(1233) := b"1111111111111111_1111111111111111_1110001100110010_1000110111001100"; -- -0.11250985886613518
	pesos_i(1234) := b"1111111111111111_1111111111111111_1101101010110101_1110110010000110"; -- -0.14566156118135806
	pesos_i(1235) := b"1111111111111111_1111111111111111_1110010000100100_0010110111101010"; -- -0.10882294689783777
	pesos_i(1236) := b"0000000000000000_0000000000000000_0000011101111110_1111101111110110"; -- 0.029281375391743268
	pesos_i(1237) := b"1111111111111111_1111111111111111_1110001101010011_0101010111110010"; -- -0.11200964787343479
	pesos_i(1238) := b"1111111111111111_1111111111111111_1111111010110101_1111000011101111"; -- -0.005036298534664473
	pesos_i(1239) := b"0000000000000000_0000000000000000_0000001010011011_0010001000010001"; -- 0.010179642809731564
	pesos_i(1240) := b"1111111111111111_1111111111111111_1100110100110000_0010111011100010"; -- -0.19848353380503364
	pesos_i(1241) := b"0000000000000000_0000000000000000_0010100000100100_0100011110010111"; -- 0.1568035835980174
	pesos_i(1242) := b"0000000000000000_0000000000000000_0000111000111111_0000110011110001"; -- 0.055649575011584185
	pesos_i(1243) := b"1111111111111111_1111111111111111_1111000101101101_0111011000111100"; -- -0.05692349466469589
	pesos_i(1244) := b"1111111111111111_1111111111111111_1101001111001110_0011011101001110"; -- -0.17263464304923865
	pesos_i(1245) := b"1111111111111111_1111111111111111_1101000111100001_0001011000010100"; -- -0.1801592066176957
	pesos_i(1246) := b"0000000000000000_0000000000000000_0010001110011100_1000101001001011"; -- 0.13910736388096595
	pesos_i(1247) := b"1111111111111111_1111111111111111_1110110101010111_0000111100110110"; -- -0.07289032879121193
	pesos_i(1248) := b"1111111111111111_1111111111111111_1111111111010110_1101111001010000"; -- -0.0006276182500162189
	pesos_i(1249) := b"1111111111111111_1111111111111111_1101100010000100_0000110100011111"; -- -0.15423505777524968
	pesos_i(1250) := b"1111111111111111_1111111111111111_1101101100010100_1011110010100110"; -- -0.1442148299143223
	pesos_i(1251) := b"1111111111111111_1111111111111111_1101011011010011_1000010000101100"; -- -0.16083501738569006
	pesos_i(1252) := b"0000000000000000_0000000000000000_0000100110001111_0111100001001100"; -- 0.03734542697943152
	pesos_i(1253) := b"0000000000000000_0000000000000000_0000101100110111_0111101111110011"; -- 0.043815371233213864
	pesos_i(1254) := b"0000000000000000_0000000000000000_0011000110001000_1101111101010000"; -- 0.19349475576803635
	pesos_i(1255) := b"0000000000000000_0000000000000000_0001100111101111_1101011111100101"; -- 0.10131596882230111
	pesos_i(1256) := b"1111111111111111_1111111111111111_1110110001101001_1110110110111101"; -- -0.07650865685020453
	pesos_i(1257) := b"0000000000000000_0000000000000000_0010100011010110_1000000011011010"; -- 0.1595230610628767
	pesos_i(1258) := b"0000000000000000_0000000000000000_0001000110010110_1011001110001110"; -- 0.06870577063838722
	pesos_i(1259) := b"1111111111111111_1111111111111111_1110110001110111_0011101101011000"; -- -0.07630566688771119
	pesos_i(1260) := b"1111111111111111_1111111111111111_1101100000010000_0010100010001010"; -- -0.1560034430500194
	pesos_i(1261) := b"0000000000000000_0000000000000000_0000001000001111_1100010110110010"; -- 0.008053165284656863
	pesos_i(1262) := b"1111111111111111_1111111111111111_1101100010100001_1111000101011110"; -- -0.15377894827956498
	pesos_i(1263) := b"1111111111111111_1111111111111111_1111011010101000_0001101111010000"; -- -0.03649736560904917
	pesos_i(1264) := b"1111111111111111_1111111111111111_1110111001111000_0000110011001111"; -- -0.06848068182239633
	pesos_i(1265) := b"0000000000000000_0000000000000000_0011000001011111_1011011011100101"; -- 0.18896048622509767
	pesos_i(1266) := b"1111111111111111_1111111111111111_1111011000111000_0010110011011001"; -- -0.03820533459982764
	pesos_i(1267) := b"0000000000000000_0000000000000000_0000011110110110_0000111101111101"; -- 0.03012177272099955
	pesos_i(1268) := b"0000000000000000_0000000000000000_0011010010011100_1001101101010001"; -- 0.20551462861315686
	pesos_i(1269) := b"1111111111111111_1111111111111111_1110101101110101_0110000000000100"; -- -0.08024024861595234
	pesos_i(1270) := b"1111111111111111_1111111111111111_1101011111110111_0111111001000001"; -- -0.15637980381780048
	pesos_i(1271) := b"0000000000000000_0000000000000000_0000100111010000_0011000000110011"; -- 0.0383329511158921
	pesos_i(1272) := b"1111111111111111_1111111111111111_1110001111010010_1100011110011100"; -- -0.11006500662074413
	pesos_i(1273) := b"0000000000000000_0000000000000000_0010100110010101_1110000011100010"; -- 0.16244321365773176
	pesos_i(1274) := b"1111111111111111_1111111111111111_1100110111110101_1011110101010011"; -- -0.19546906211900997
	pesos_i(1275) := b"1111111111111111_1111111111111111_1101010111110110_0110101010011010"; -- -0.16420873390500704
	pesos_i(1276) := b"1111111111111111_1111111111111111_1101101110100111_1001010100001100"; -- -0.14197414829315277
	pesos_i(1277) := b"1111111111111111_1111111111111111_1110000011011100_0111110001000000"; -- -0.1216356604683233
	pesos_i(1278) := b"0000000000000000_0000000000000000_0000001010101111_1000100101000100"; -- 0.010490969690927351
	pesos_i(1279) := b"1111111111111111_1111111111111111_1110001010001101_0111101110010100"; -- -0.11502864495238885
	pesos_i(1280) := b"0000000000000000_0000000000000000_0001111010111110_0011001101101010"; -- 0.12008973454223887
	pesos_i(1281) := b"0000000000000000_0000000000000000_0010110010101010_1011110000011110"; -- 0.1744802068380064
	pesos_i(1282) := b"1111111111111111_1111111111111111_1110001010110101_0010111101110101"; -- -0.11442283046021458
	pesos_i(1283) := b"1111111111111111_1111111111111111_1110010111111100_1111011010001110"; -- -0.10160883945465296
	pesos_i(1284) := b"0000000000000000_0000000000000000_0000110010110000_0001111111111100"; -- 0.04956245328865995
	pesos_i(1285) := b"0000000000000000_0000000000000000_0000100101101101_1000110000011110"; -- 0.036827809542556204
	pesos_i(1286) := b"0000000000000000_0000000000000000_0001010101011000_1101011110000011"; -- 0.08338686894477251
	pesos_i(1287) := b"1111111111111111_1111111111111111_1111100111000010_0111000100101010"; -- -0.024376799857139295
	pesos_i(1288) := b"1111111111111111_1111111111111111_1111110011010111_1011110101010100"; -- -0.012333075470960391
	pesos_i(1289) := b"0000000000000000_0000000000000000_0010011011000111_0010010110100101"; -- 0.15147624271444177
	pesos_i(1290) := b"0000000000000000_0000000000000000_0000110001000110_1100001111000101"; -- 0.047954783982272854
	pesos_i(1291) := b"0000000000000000_0000000000000000_0000110111110001_0010010100101110"; -- 0.0544608343281893
	pesos_i(1292) := b"0000000000000000_0000000000000000_0001010101010010_1010110010000110"; -- 0.08329275387324149
	pesos_i(1293) := b"1111111111111111_1111111111111111_1110011110011001_1011110000111111"; -- -0.09531043493325032
	pesos_i(1294) := b"1111111111111111_1111111111111111_1101101111101000_0011111101100000"; -- -0.1409874333968828
	pesos_i(1295) := b"0000000000000000_0000000000000000_0000110010001010_0100110001111111"; -- 0.04898527241762204
	pesos_i(1296) := b"1111111111111111_1111111111111111_1110000101011111_0101111110101111"; -- -0.1196384619224708
	pesos_i(1297) := b"1111111111111111_1111111111111111_1101110100000101_0101100010001000"; -- -0.13663717913108844
	pesos_i(1298) := b"0000000000000000_0000000000000000_0010011100111010_1011101010011110"; -- 0.15323988310227166
	pesos_i(1299) := b"0000000000000000_0000000000000000_0010010011010111_0010011101110001"; -- 0.1439079905286907
	pesos_i(1300) := b"1111111111111111_1111111111111111_1111100011011101_1111001000110001"; -- -0.02786337176976869
	pesos_i(1301) := b"1111111111111111_1111111111111111_1101111110101011_0010111110100110"; -- -0.1262941571039115
	pesos_i(1302) := b"1111111111111111_1111111111111111_1110110011010011_0110101001000001"; -- -0.07489906227754428
	pesos_i(1303) := b"0000000000000000_0000000000000000_0001010101101010_1100110101000001"; -- 0.08366091577372226
	pesos_i(1304) := b"1111111111111111_1111111111111111_1111110000000110_0010000010000010"; -- -0.015531509650195051
	pesos_i(1305) := b"0000000000000000_0000000000000000_0000101110000101_1110110000110011"; -- 0.04501224745513444
	pesos_i(1306) := b"0000000000000000_0000000000000000_0010011100001110_1111111101111001"; -- 0.152572600431228
	pesos_i(1307) := b"1111111111111111_1111111111111111_1110000111001010_0001000111111011"; -- -0.11801040286575697
	pesos_i(1308) := b"1111111111111111_1111111111111111_1111100100111001_0000010111010101"; -- -0.026473651485428403
	pesos_i(1309) := b"0000000000000000_0000000000000000_0010000100010011_1110110110000001"; -- 0.12921032328456258
	pesos_i(1310) := b"1111111111111111_1111111111111111_1111010110101011_0000101001001100"; -- -0.040358883214295045
	pesos_i(1311) := b"1111111111111111_1111111111111111_1111001001111010_0111000100000001"; -- -0.05281919211032521
	pesos_i(1312) := b"1111111111111111_1111111111111111_1101101000001100_0101010001010010"; -- -0.14824936875513067
	pesos_i(1313) := b"0000000000000000_0000000000000000_0000101001111101_0111101011101111"; -- 0.040977176132524246
	pesos_i(1314) := b"1111111111111111_1111111111111111_1101111101001001_1111011110001000"; -- -0.12777760442647124
	pesos_i(1315) := b"1111111111111111_1111111111111111_1110001111010000_0110100101101010"; -- -0.11010113875900862
	pesos_i(1316) := b"0000000000000000_0000000000000000_0001000111100100_0001111011111010"; -- 0.06988710015896799
	pesos_i(1317) := b"1111111111111111_1111111111111111_1111001101111001_1111110110000111"; -- -0.04891982508643806
	pesos_i(1318) := b"1111111111111111_1111111111111111_1110110101101000_1110001101100101"; -- -0.07261828209616887
	pesos_i(1319) := b"1111111111111111_1111111111111111_1110111001110101_1010010000010010"; -- -0.0685174422236139
	pesos_i(1320) := b"1111111111111111_1111111111111111_1110001000000100_0110110010010101"; -- -0.11711999293779456
	pesos_i(1321) := b"0000000000000000_0000000000000000_0000010000011111_0011011110101110"; -- 0.01610134120714938
	pesos_i(1322) := b"1111111111111111_1111111111111111_1110001111100011_1110101010101110"; -- -0.10980351698630125
	pesos_i(1323) := b"0000000000000000_0000000000000000_0000010011100011_0000010000001000"; -- 0.01908898546941775
	pesos_i(1324) := b"1111111111111111_1111111111111111_1101101001000010_0001111000101000"; -- -0.14742862258039066
	pesos_i(1325) := b"1111111111111111_1111111111111111_1110110001000011_1101011000110001"; -- -0.07708989427110659
	pesos_i(1326) := b"1111111111111111_1111111111111111_1110000111010000_0000100101011110"; -- -0.11791936357417493
	pesos_i(1327) := b"0000000000000000_0000000000000000_0000110110101001_0000111101100000"; -- 0.053360901704711514
	pesos_i(1328) := b"1111111111111111_1111111111111111_1101100010110110_1011101011101110"; -- -0.15346175854150762
	pesos_i(1329) := b"1111111111111111_1111111111111111_1110011010000100_1010001001111001"; -- -0.0995386557693542
	pesos_i(1330) := b"1111111111111111_1111111111111111_1111101011001100_1111101010110010"; -- -0.020309764373350733
	pesos_i(1331) := b"0000000000000000_0000000000000000_0000011011110101_0011111000011010"; -- 0.02717960495141187
	pesos_i(1332) := b"0000000000000000_0000000000000000_0000110000100111_1111111011111011"; -- 0.0474852909057795
	pesos_i(1333) := b"1111111111111111_1111111111111111_1110110101101100_1010110111100101"; -- -0.07256043582213496
	pesos_i(1334) := b"0000000000000000_0000000000000000_0001111011110011_1111001101010001"; -- 0.12090988842139298
	pesos_i(1335) := b"0000000000000000_0000000000000000_0010111111011010_0101010010101011"; -- 0.1869252126476874
	pesos_i(1336) := b"0000000000000000_0000000000000000_0010011100100101_0010100000101000"; -- 0.152910718609285
	pesos_i(1337) := b"1111111111111111_1111111111111111_1110001011100011_1111001001001101"; -- -0.11370931257243787
	pesos_i(1338) := b"1111111111111111_1111111111111111_1101011110101000_1100000110001001"; -- -0.15758123786575357
	pesos_i(1339) := b"1111111111111111_1111111111111111_1101110111011110_0100101000100110"; -- -0.1333268792584303
	pesos_i(1340) := b"1111111111111111_1111111111111111_1111100100111101_0111000010010100"; -- -0.026406253661848067
	pesos_i(1341) := b"0000000000000000_0000000000000000_0010011100000001_0010011110011111"; -- 0.15236137039701672
	pesos_i(1342) := b"1111111111111111_1111111111111111_1110001000110110_0000110011111010"; -- -0.11636275201034067
	pesos_i(1343) := b"1111111111111111_1111111111111111_1100010000101111_0100011011000100"; -- -0.23365361890251066
	pesos_i(1344) := b"1111111111111111_1111111111111111_1110011110000000_0101110001101111"; -- -0.09569761542098001
	pesos_i(1345) := b"1111111111111111_1111111111111111_1110110111001001_1110100101100010"; -- -0.07113782273301947
	pesos_i(1346) := b"0000000000000000_0000000000000000_0000000010110011_1110101000011000"; -- 0.0027452762692480627
	pesos_i(1347) := b"0000000000000000_0000000000000000_0010101101001000_1000000010111101"; -- 0.16907505610614362
	pesos_i(1348) := b"1111111111111111_1111111111111111_1111111010101100_1010110111001110"; -- -0.00517762874547296
	pesos_i(1349) := b"1111111111111111_1111111111111111_1111011011010111_1101101011000101"; -- -0.03576882062124582
	pesos_i(1350) := b"0000000000000000_0000000000000000_0000000001100010_1111101010100111"; -- 0.0015103014523437216
	pesos_i(1351) := b"1111111111111111_1111111111111111_1100101110101000_1111111110101101"; -- -0.2044525338857174
	pesos_i(1352) := b"0000000000000000_0000000000000000_0001001110111000_0110100010010100"; -- 0.07703260051334573
	pesos_i(1353) := b"1111111111111111_1111111111111111_1110100011111100_1001010111111011"; -- -0.08989584573304432
	pesos_i(1354) := b"1111111111111111_1111111111111111_1101010001010101_1010111100101001"; -- -0.1705675625740309
	pesos_i(1355) := b"0000000000000000_0000000000000000_0001011101000101_0000100010110110"; -- 0.09089712557537645
	pesos_i(1356) := b"0000000000000000_0000000000000000_0001111100001101_0010011111101110"; -- 0.12129449414246504
	pesos_i(1357) := b"0000000000000000_0000000000000000_0010101100110000_0001001011100110"; -- 0.16870229829966532
	pesos_i(1358) := b"1111111111111111_1111111111111111_1111111010000010_0100101111111111"; -- -0.005824327666657648
	pesos_i(1359) := b"1111111111111111_1111111111111111_1110000110001111_1001001110001110"; -- -0.11890294824920009
	pesos_i(1360) := b"0000000000000000_0000000000000000_0000001001000111_0011001010111011"; -- 0.008898897705737993
	pesos_i(1361) := b"0000000000000000_0000000000000000_0001001101100111_0000011100001101"; -- 0.07579082552922238
	pesos_i(1362) := b"1111111111111111_1111111111111111_1111101000111101_0000101000111100"; -- -0.022506103880360624
	pesos_i(1363) := b"1111111111111111_1111111111111111_1101110010100101_1101010101110000"; -- -0.13809457790611845
	pesos_i(1364) := b"1111111111111111_1111111111111111_1101001110011101_0010100001110101"; -- -0.1733832087997597
	pesos_i(1365) := b"0000000000000000_0000000000000000_0001101111110100_0101011101010011"; -- 0.10919709948753684
	pesos_i(1366) := b"0000000000000000_0000000000000000_0001111100011000_0101110001001001"; -- 0.12146546151764538
	pesos_i(1367) := b"0000000000000000_0000000000000000_0001100000110001_1001000100101100"; -- 0.09450633361562084
	pesos_i(1368) := b"0000000000000000_0000000000000000_0000110101010010_0101101001110110"; -- 0.05203786269357868
	pesos_i(1369) := b"0000000000000000_0000000000000000_0010111011001010_0100000001100100"; -- 0.18277361343554724
	pesos_i(1370) := b"1111111111111111_1111111111111111_1110100111110010_1110110110011011"; -- -0.08613696056146292
	pesos_i(1371) := b"1111111111111111_1111111111111111_1111001111010001_1100101101100001"; -- -0.047580040677519725
	pesos_i(1372) := b"0000000000000000_0000000000000000_0001011110101111_1000111101001100"; -- 0.09252257918651488
	pesos_i(1373) := b"1111111111111111_1111111111111111_1111000111011101_0011010001010000"; -- -0.05521843946187924
	pesos_i(1374) := b"0000000000000000_0000000000000000_0001110101111011_1001110101001000"; -- 0.1151674556429392
	pesos_i(1375) := b"1111111111111111_1111111111111111_1111111001000100_1001110110001111"; -- -0.006765511106576627
	pesos_i(1376) := b"0000000000000000_0000000000000000_0010101111100111_0001011000100011"; -- 0.17149484975878898
	pesos_i(1377) := b"0000000000000000_0000000000000000_0010010101000110_1000111001000000"; -- 0.14560784394807608
	pesos_i(1378) := b"1111111111111111_1111111111111111_1111000101011011_0100000001110111"; -- -0.057201357826386245
	pesos_i(1379) := b"0000000000000000_0000000000000000_0010110111011011_0010101101011011"; -- 0.17912550895880525
	pesos_i(1380) := b"1111111111111111_1111111111111111_1111101111111110_0001001001111110"; -- -0.015654415270736577
	pesos_i(1381) := b"1111111111111111_1111111111111111_1101011000111001_1001110101110001"; -- -0.16318336472980102
	pesos_i(1382) := b"1111111111111111_1111111111111111_1101000110110001_1110100000001101"; -- -0.18087911295326572
	pesos_i(1383) := b"1111111111111111_1111111111111111_1110110010001101_0000111100111011"; -- -0.07597260295665646
	pesos_i(1384) := b"1111111111111111_1111111111111111_1111000000101110_1101001111010110"; -- -0.06178546928550974
	pesos_i(1385) := b"1111111111111111_1111111111111111_1110001100101111_1100101000010010"; -- -0.11255204258882794
	pesos_i(1386) := b"0000000000000000_0000000000000000_0001011000000101_0111100101000011"; -- 0.08602102160181162
	pesos_i(1387) := b"1111111111111111_1111111111111111_1111111101000011_0101110011110110"; -- -0.0028783702535408674
	pesos_i(1388) := b"0000000000000000_0000000000000000_0010100000001010_0010101001001101"; -- 0.1564051092478142
	pesos_i(1389) := b"1111111111111111_1111111111111111_1111011111001111_0001110010010000"; -- -0.03199597812729773
	pesos_i(1390) := b"1111111111111111_1111111111111111_1111010100100100_1010001110000110"; -- -0.04240968687807239
	pesos_i(1391) := b"1111111111111111_1111111111111111_1111001110100011_1111110001000001"; -- -0.048279031803688206
	pesos_i(1392) := b"0000000000000000_0000000000000000_0000111111101001_0010011000111011"; -- 0.06215132661572957
	pesos_i(1393) := b"0000000000000000_0000000000000000_0000001110001101_0010010010001101"; -- 0.013872417844683823
	pesos_i(1394) := b"1111111111111111_1111111111111111_1111000110000110_1100000100110101"; -- -0.05653755625094767
	pesos_i(1395) := b"0000000000000000_0000000000000000_0010100001101111_0100100001011001"; -- 0.1579480378463519
	pesos_i(1396) := b"0000000000000000_0000000000000000_0000000011000110_0001001100100101"; -- 0.0030223814226998935
	pesos_i(1397) := b"1111111111111111_1111111111111111_1110010010000001_1001111011110001"; -- -0.10739714253266175
	pesos_i(1398) := b"1111111111111111_1111111111111111_1101100010001001_0110010010100000"; -- -0.15415354812823373
	pesos_i(1399) := b"0000000000000000_0000000000000000_0010101000001010_1011100000101110"; -- 0.16422606587772964
	pesos_i(1400) := b"1111111111111111_1111111111111111_1101011110111011_1011110011000110"; -- -0.15729160464069708
	pesos_i(1401) := b"0000000000000000_0000000000000000_0000111100110000_1110100110000100"; -- 0.05934009055405724
	pesos_i(1402) := b"0000000000000000_0000000000000000_0000101001110011_1101010011010110"; -- 0.040829946856741274
	pesos_i(1403) := b"0000000000000000_0000000000000000_0010100000111101_1110111101110001"; -- 0.15719505787562232
	pesos_i(1404) := b"1111111111111111_1111111111111111_1100111111111011_1100000100001111"; -- -0.18756478671478416
	pesos_i(1405) := b"0000000000000000_0000000000000000_0001001100000101_1111010111001000"; -- 0.07430969354490069
	pesos_i(1406) := b"0000000000000000_0000000000000000_0001101110001111_0010001001101000"; -- 0.10765280758945157
	pesos_i(1407) := b"0000000000000000_0000000000000000_0010010100111101_1001001001011100"; -- 0.14547075988720767
	pesos_i(1408) := b"0000000000000000_0000000000000000_0000000110110001_0111101101111100"; -- 0.006614415943477672
	pesos_i(1409) := b"0000000000000000_0000000000000000_0001010111000111_0111110001101000"; -- 0.0850751641734524
	pesos_i(1410) := b"1111111111111111_1111111111111111_1110001000010001_0111000000011110"; -- -0.11692141783651623
	pesos_i(1411) := b"1111111111111111_1111111111111111_1101110001111100_1001000111101001"; -- -0.13872421320828782
	pesos_i(1412) := b"0000000000000000_0000000000000000_0000010101110101_1001101110101011"; -- 0.021325806782521488
	pesos_i(1413) := b"0000000000000000_0000000000000000_0001111110101100_0011000001101000"; -- 0.1237211470070671
	pesos_i(1414) := b"1111111111111111_1111111111111111_1111010001110111_1110001111010101"; -- -0.045045624366486646
	pesos_i(1415) := b"0000000000000000_0000000000000000_0100001010101111_1000001001101001"; -- 0.2604905610632978
	pesos_i(1416) := b"0000000000000000_0000000000000000_0010010111001110_0001011011100011"; -- 0.14767592471079194
	pesos_i(1417) := b"0000000000000000_0000000000000000_0000110000100110_0001101011001111"; -- 0.047456431989950844
	pesos_i(1418) := b"0000000000000000_0000000000000000_0000000001111001_0000001101101101"; -- 0.0018465177685772416
	pesos_i(1419) := b"1111111111111111_1111111111111111_1111001001010110_1101000110111001"; -- -0.05336274360556075
	pesos_i(1420) := b"1111111111111111_1111111111111111_1110011100010010_0100011110000010"; -- -0.09737732968915877
	pesos_i(1421) := b"1111111111111111_1111111111111111_1101000101010000_0101100101011101"; -- -0.18236772037139054
	pesos_i(1422) := b"0000000000000000_0000000000000000_0010011110101111_0011111001001100"; -- 0.15501775132163803
	pesos_i(1423) := b"0000000000000000_0000000000000000_0010100001001101_0111111100001011"; -- 0.1574324991898634
	pesos_i(1424) := b"1111111111111111_1111111111111111_1111000111000001_1011011000101111"; -- -0.05563794479210766
	pesos_i(1425) := b"1111111111111111_1111111111111111_1110010101101101_1001000111000001"; -- -0.10379685433107828
	pesos_i(1426) := b"0000000000000000_0000000000000000_0010000000010000_1110011110101111"; -- 0.12525795007210924
	pesos_i(1427) := b"0000000000000000_0000000000000000_0001110111011100_1110110010011100"; -- 0.11665228650120642
	pesos_i(1428) := b"0000000000000000_0000000000000000_0001101111011010_0010111111101010"; -- 0.10879802184136615
	pesos_i(1429) := b"0000000000000000_0000000000000000_0010010110001000_0010100001101101"; -- 0.14660885487256614
	pesos_i(1430) := b"0000000000000000_0000000000000000_0001100000011000_1000100001100110"; -- 0.09412434092524187
	pesos_i(1431) := b"1111111111111111_1111111111111111_1111111000000001_0011010111100111"; -- -0.007794028326965611
	pesos_i(1432) := b"0000000000000000_0000000000000000_0000010101010000_1100001110010111"; -- 0.020763611262043142
	pesos_i(1433) := b"0000000000000000_0000000000000000_0000000011000111_1011001000000001"; -- 0.003047108787682378
	pesos_i(1434) := b"0000000000000000_0000000000000000_0000011100111001_0100000001001111"; -- 0.028217334111785765
	pesos_i(1435) := b"0000000000000000_0000000000000000_0001101111011100_1110001010010111"; -- 0.10883918936068
	pesos_i(1436) := b"1111111111111111_1111111111111111_1101001100011000_0111111001011011"; -- -0.17540750760255241
	pesos_i(1437) := b"1111111111111111_1111111111111111_1101100001101011_0000110111101111"; -- -0.1546164791527786
	pesos_i(1438) := b"0000000000000000_0000000000000000_0000101011010000_1000000111000010"; -- 0.04224406232868698
	pesos_i(1439) := b"0000000000000000_0000000000000000_0010100100000110_0110010110000010"; -- 0.16025385299094316
	pesos_i(1440) := b"1111111111111111_1111111111111111_1110000111110100_1100001011110011"; -- -0.11735898567687343
	pesos_i(1441) := b"1111111111111111_1111111111111111_1111000000100100_0011011101001011"; -- -0.06194738783634935
	pesos_i(1442) := b"1111111111111111_1111111111111111_1110100011101110_1100000101001111"; -- -0.0901068860357905
	pesos_i(1443) := b"0000000000000000_0000000000000000_0000000101001100_1101011101101001"; -- 0.005078757497354183
	pesos_i(1444) := b"1111111111111111_1111111111111111_1111011110011000_1110100011010011"; -- -0.03282303666817639
	pesos_i(1445) := b"1111111111111111_1111111111111111_1110001011011011_0000111010111110"; -- -0.11384494653081274
	pesos_i(1446) := b"0000000000000000_0000000000000000_0010000100001111_1101011110110100"; -- 0.12914798874627875
	pesos_i(1447) := b"0000000000000000_0000000000000000_0001000000000001_1000000011111011"; -- 0.06252294652462384
	pesos_i(1448) := b"1111111111111111_1111111111111111_1100101110111111_0110101001000110"; -- -0.20411048700990317
	pesos_i(1449) := b"1111111111111111_1111111111111111_1110011010101110_1111011101000100"; -- -0.09889273261725616
	pesos_i(1450) := b"0000000000000000_0000000000000000_0000001011001101_0111010010101101"; -- 0.010947506265038107
	pesos_i(1451) := b"0000000000000000_0000000000000000_0000110100111000_1101011101010110"; -- 0.05164857710975675
	pesos_i(1452) := b"0000000000000000_0000000000000000_0000010110111110_1011100010110111"; -- 0.022441429853858642
	pesos_i(1453) := b"0000000000000000_0000000000000000_0001110110110000_0001100101000010"; -- 0.11596830231586851
	pesos_i(1454) := b"0000000000000000_0000000000000000_0001011110010010_0010011110000001"; -- 0.09207388784145218
	pesos_i(1455) := b"0000000000000000_0000000000000000_0001010101011101_0000110000010111"; -- 0.083451038073085
	pesos_i(1456) := b"0000000000000000_0000000000000000_0010110010110011_0010000001110010"; -- 0.17460825709922384
	pesos_i(1457) := b"1111111111111111_1111111111111111_1111001111100101_0110010011110110"; -- -0.04728096960645117
	pesos_i(1458) := b"1111111111111111_1111111111111111_1111010010010111_1110001010010101"; -- -0.04455741740411457
	pesos_i(1459) := b"0000000000000000_0000000000000000_0010101011110010_1001100011111101"; -- 0.1677642457793847
	pesos_i(1460) := b"1111111111111111_1111111111111111_1101000000010100_1011100110111111"; -- -0.1871837528995118
	pesos_i(1461) := b"0000000000000000_0000000000000000_0000111100001101_0011010111111101"; -- 0.058795332210844854
	pesos_i(1462) := b"1111111111111111_1111111111111111_1110011010000011_1111100110100111"; -- -0.09954871822295515
	pesos_i(1463) := b"1111111111111111_1111111111111111_1100101100001100_1000010110010000"; -- -0.20684018357087136
	pesos_i(1464) := b"1111111111111111_1111111111111111_1100111001010001_1010000111011010"; -- -0.19406689107609296
	pesos_i(1465) := b"0000000000000000_0000000000000000_0001110101000000_0101100111110100"; -- 0.11426317420583264
	pesos_i(1466) := b"1111111111111111_1111111111111111_1101101011100111_0101001001011011"; -- -0.14490781096086916
	pesos_i(1467) := b"0000000000000000_0000000000000000_0000010101110110_0101101010110010"; -- 0.02133719307761977
	pesos_i(1468) := b"0000000000000000_0000000000000000_0011010010100110_1110101010110011"; -- 0.20567194809587153
	pesos_i(1469) := b"0000000000000000_0000000000000000_0001101111101101_0100110110110101"; -- 0.10908971482142218
	pesos_i(1470) := b"0000000000000000_0000000000000000_0010001011101101_0011010010111111"; -- 0.136431977016639
	pesos_i(1471) := b"0000000000000000_0000000000000000_0001011111001110_0110011111101101"; -- 0.09299325499183822
	pesos_i(1472) := b"1111111111111111_1111111111111111_1111110101100011_1000010001111100"; -- -0.01020023325159787
	pesos_i(1473) := b"1111111111111111_1111111111111111_1111011100010101_0011001111100111"; -- -0.03483272181216936
	pesos_i(1474) := b"1111111111111111_1111111111111111_1100111100110111_0100000101011010"; -- -0.19056312132311887
	pesos_i(1475) := b"1111111111111111_1111111111111111_1101010011000011_0110010111001110"; -- -0.16889346803565886
	pesos_i(1476) := b"1111111111111111_1111111111111111_1111011111100110_1001010110100100"; -- -0.031637809270277366
	pesos_i(1477) := b"1111111111111111_1111111111111111_1111010101101011_0111001010011110"; -- -0.041329227767070875
	pesos_i(1478) := b"0000000000000000_0000000000000000_0000101010010101_0001000100100000"; -- 0.041337080377430405
	pesos_i(1479) := b"1111111111111111_1111111111111111_1111010100011111_1011000100011100"; -- -0.04248517089782061
	pesos_i(1480) := b"1111111111111111_1111111111111111_1101001101011100_0100011010111101"; -- -0.17437322517023002
	pesos_i(1481) := b"0000000000000000_0000000000000000_0000010101110111_1101110011010111"; -- 0.021360209006723987
	pesos_i(1482) := b"1111111111111111_1111111111111111_1110011000011011_0010011101101111"; -- -0.10114816216693251
	pesos_i(1483) := b"0000000000000000_0000000000000000_0001101011000010_1000101011000000"; -- 0.10453097516669062
	pesos_i(1484) := b"1111111111111111_1111111111111111_1101010010000100_1010110011010100"; -- -0.1698505384696356
	pesos_i(1485) := b"1111111111111111_1111111111111111_1100101101001001_0100100110010001"; -- -0.20591297343815412
	pesos_i(1486) := b"0000000000000000_0000000000000000_0001111110011111_0010101100100000"; -- 0.12352246784885182
	pesos_i(1487) := b"0000000000000000_0000000000000000_0000001110111011_0000110001100110"; -- 0.014572882458072707
	pesos_i(1488) := b"1111111111111111_1111111111111111_1110111110000001_0110011110100000"; -- -0.06443168969009773
	pesos_i(1489) := b"0000000000000000_0000000000000000_0000011110010101_0100010010110100"; -- 0.02962140459731802
	pesos_i(1490) := b"1111111111111111_1111111111111111_1110110110110000_1011000101000001"; -- -0.07152263788320776
	pesos_i(1491) := b"1111111111111111_1111111111111111_1111001000001110_0010001001110110"; -- -0.054471823002373285
	pesos_i(1492) := b"1111111111111111_1111111111111111_1101111000111100_0010011011111101"; -- -0.1318946487667075
	pesos_i(1493) := b"0000000000000000_0000000000000000_0010011000110111_0111010001111101"; -- 0.1492836766338771
	pesos_i(1494) := b"1111111111111111_1111111111111111_1110001100100100_1010000010001011"; -- -0.11272236439049269
	pesos_i(1495) := b"0000000000000000_0000000000000000_0000110110110101_0001111011101000"; -- 0.05354493294835045
	pesos_i(1496) := b"1111111111111111_1111111111111111_1110011101001010_0110100011101011"; -- -0.09652084598094196
	pesos_i(1497) := b"1111111111111111_1111111111111111_1111110010100100_1001001011100110"; -- -0.013113802851441259
	pesos_i(1498) := b"0000000000000000_0000000000000000_0001110100000000_1111010011100111"; -- 0.11329584741951237
	pesos_i(1499) := b"0000000000000000_0000000000000000_0010100001110100_1010000010001001"; -- 0.15802958824652846
	pesos_i(1500) := b"0000000000000000_0000000000000000_0001111111101001_0110001111111000"; -- 0.1246550064698748
	pesos_i(1501) := b"1111111111111111_1111111111111111_1111000011011111_0000011000010001"; -- -0.05909692847180584
	pesos_i(1502) := b"1111111111111111_1111111111111111_1101000001101110_0100101010000110"; -- -0.18581709135543076
	pesos_i(1503) := b"0000000000000000_0000000000000000_0000011001010011_1001000110110100"; -- 0.024712664150001677
	pesos_i(1504) := b"1111111111111111_1111111111111111_1110100001110000_1000110110011110"; -- -0.09203257460122698
	pesos_i(1505) := b"1111111111111111_1111111111111111_1110111100110001_0000001000011111"; -- -0.06565844301273148
	pesos_i(1506) := b"0000000000000000_0000000000000000_0001110100110100_1001100000111110"; -- 0.1140837813323563
	pesos_i(1507) := b"0000000000000000_0000000000000000_0000001011001111_0001001100011111"; -- 0.010972209020451757
	pesos_i(1508) := b"1111111111111111_1111111111111111_1100001111100110_0100010110100000"; -- -0.234767578515109
	pesos_i(1509) := b"1111111111111111_1111111111111111_1111010011001010_1010110001100110"; -- -0.04378244896933586
	pesos_i(1510) := b"0000000000000000_0000000000000000_0010001110011011_0001000000101110"; -- 0.13908482660622826
	pesos_i(1511) := b"0000000000000000_0000000000000000_0001101110110010_1010010110101111"; -- 0.10819469007532384
	pesos_i(1512) := b"1111111111111111_1111111111111111_1110110011111100_1110111010111111"; -- -0.07426555483450616
	pesos_i(1513) := b"0000000000000000_0000000000000000_0010001100110110_1001110111001110"; -- 0.1375521304946164
	pesos_i(1514) := b"0000000000000000_0000000000000000_0000101010110001_0101001011010001"; -- 0.041768241955718315
	pesos_i(1515) := b"1111111111111111_1111111111111111_1110111011100101_0000100011010010"; -- -0.06681771166822793
	pesos_i(1516) := b"1111111111111111_1111111111111111_1110100010001000_0011011010001011"; -- -0.09167155367870014
	pesos_i(1517) := b"0000000000000000_0000000000000000_0001111101001000_0100011011011111"; -- 0.12219660701880271
	pesos_i(1518) := b"1111111111111111_1111111111111111_1110101001111010_1010001110010111"; -- -0.0840661769376985
	pesos_i(1519) := b"0000000000000000_0000000000000000_0010110010010000_1111110110101000"; -- 0.1740873846228851
	pesos_i(1520) := b"1111111111111111_1111111111111111_1101111011000100_0001101100111101"; -- -0.12982015375216716
	pesos_i(1521) := b"0000000000000000_0000000000000000_0000011011100000_0110011010010101"; -- 0.026861583203306783
	pesos_i(1522) := b"1111111111111111_1111111111111111_1111101111001011_0100000110110000"; -- -0.016429800465665084
	pesos_i(1523) := b"0000000000000000_0000000000000000_0011001100001001_1011000110101011"; -- 0.19936666888760482
	pesos_i(1524) := b"0000000000000000_0000000000000000_0000100100011011_1010011001101110"; -- 0.03557815735007322
	pesos_i(1525) := b"1111111111111111_1111111111111111_1110110100100101_1001100010100000"; -- -0.07364507756225339
	pesos_i(1526) := b"1111111111111111_1111111111111111_1110001101110001_1001100001111111"; -- -0.11154791733012966
	pesos_i(1527) := b"1111111111111111_1111111111111111_1101000111010110_1110101101010100"; -- -0.18031434243431488
	pesos_i(1528) := b"1111111111111111_1111111111111111_1111000011100101_0011111000010111"; -- -0.0590020365358169
	pesos_i(1529) := b"0000000000000000_0000000000000000_0001010101101110_0110000110100110"; -- 0.08371553701230777
	pesos_i(1530) := b"0000000000000000_0000000000000000_0010100100010011_0110110100000001"; -- 0.16045266405368114
	pesos_i(1531) := b"0000000000000000_0000000000000000_0001000000111011_1111101101010110"; -- 0.06341524943250747
	pesos_i(1532) := b"0000000000000000_0000000000000000_0001100101011011_0011001111001100"; -- 0.09904788721431149
	pesos_i(1533) := b"0000000000000000_0000000000000000_0000010100100000_0010011011010111"; -- 0.020021846271731526
	pesos_i(1534) := b"1111111111111111_1111111111111111_1101110010101000_1110110001101000"; -- -0.13804743251504023
	pesos_i(1535) := b"0000000000000000_0000000000000000_0010010000110010_1011011111101101"; -- 0.14139890221861548
	pesos_i(1536) := b"1111111111111111_1111111111111111_1101101111010010_0100010101111101"; -- -0.14132276242654593
	pesos_i(1537) := b"1111111111111111_1111111111111111_1111111010100011_0111100111010111"; -- -0.005318055049811032
	pesos_i(1538) := b"1111111111111111_1111111111111111_1111011111000100_0100100110011010"; -- -0.03216114024775979
	pesos_i(1539) := b"0000000000000000_0000000000000000_0000010000011001_1110010010000000"; -- 0.016020089309691832
	pesos_i(1540) := b"0000000000000000_0000000000000000_0010110101100000_1111000000001000"; -- 0.17726040071908933
	pesos_i(1541) := b"0000000000000000_0000000000000000_0000111101101010_1000111000010101"; -- 0.06021965048347054
	pesos_i(1542) := b"0000000000000000_0000000000000000_0010101000111101_0111101000011110"; -- 0.16500056495472587
	pesos_i(1543) := b"1111111111111111_1111111111111111_1111110100000000_0110100111100110"; -- -0.011712438058501867
	pesos_i(1544) := b"0000000000000000_0000000000000000_0001000110010010_0111110101101100"; -- 0.06864150895989869
	pesos_i(1545) := b"1111111111111111_1111111111111111_1101110001000110_1010011110011111"; -- -0.1395468936549818
	pesos_i(1546) := b"1111111111111111_1111111111111111_1111110111010011_0001100010110110"; -- -0.008497672629476566
	pesos_i(1547) := b"0000000000000000_0000000000000000_0001000000000000_1001011110111000"; -- 0.06250904302781506
	pesos_i(1548) := b"1111111111111111_1111111111111111_1101101100111011_0110110100011100"; -- -0.14362447813212567
	pesos_i(1549) := b"1111111111111111_1111111111111111_1101001000100111_1100111100001001"; -- -0.17908006699244777
	pesos_i(1550) := b"0000000000000000_0000000000000000_0010100001000101_0010101001111101"; -- 0.15730538905545027
	pesos_i(1551) := b"1111111111111111_1111111111111111_1101110110100101_0101110011011011"; -- -0.13419551526243756
	pesos_i(1552) := b"1111111111111111_1111111111111111_1100001010011101_1011011111110101"; -- -0.2397809054628716
	pesos_i(1553) := b"0000000000000000_0000000000000000_0000011100110101_1010011110110000"; -- 0.028162460757060304
	pesos_i(1554) := b"1111111111111111_1111111111111111_1111000111010000_0010111111111100"; -- -0.05541706182901948
	pesos_i(1555) := b"0000000000000000_0000000000000000_0000100000001011_1000010110110010"; -- 0.03142581552111062
	pesos_i(1556) := b"1111111111111111_1111111111111111_1110001001110100_1110101011010000"; -- -0.11540348455770517
	pesos_i(1557) := b"0000000000000000_0000000000000000_0001011110111101_1011101010011111"; -- 0.09273878473084474
	pesos_i(1558) := b"0000000000000000_0000000000000000_0000010101001101_1000101011000100"; -- 0.020714447856477206
	pesos_i(1559) := b"0000000000000000_0000000000000000_0011000101011001_1010010000100011"; -- 0.1927740654542677
	pesos_i(1560) := b"0000000000000000_0000000000000000_0001011110110011_0111010100001011"; -- 0.09258204955769384
	pesos_i(1561) := b"1111111111111111_1111111111111111_1111011101001100_0110011111011101"; -- -0.033990391303590745
	pesos_i(1562) := b"0000000000000000_0000000000000000_0000011011001100_0100110100010110"; -- 0.026554887714743514
	pesos_i(1563) := b"1111111111111111_1111111111111111_1110001010101001_0011111100010110"; -- -0.11460500448754038
	pesos_i(1564) := b"1111111111111111_1111111111111111_1110101100001111_1011110100001010"; -- -0.08179110057022378
	pesos_i(1565) := b"0000000000000000_0000000000000000_0000011100011001_1001011011100101"; -- 0.02773421365875754
	pesos_i(1566) := b"0000000000000000_0000000000000000_0000001101001100_0010011000010111"; -- 0.01288068832072023
	pesos_i(1567) := b"0000000000000000_0000000000000000_0001011111001100_0110101100000001"; -- 0.09296292085679157
	pesos_i(1568) := b"1111111111111111_1111111111111111_1101011110110101_0010101110010000"; -- -0.1573918127567736
	pesos_i(1569) := b"1111111111111111_1111111111111111_1110101110111011_0010110010101011"; -- -0.07917519405872966
	pesos_i(1570) := b"0000000000000000_0000000000000000_0010111000100010_1111001001110011"; -- 0.18022074998899662
	pesos_i(1571) := b"0000000000000000_0000000000000000_0000010100011110_0010001111110100"; -- 0.01999115666035415
	pesos_i(1572) := b"0000000000000000_0000000000000000_0000000101000100_1111100001100100"; -- 0.004958652794674304
	pesos_i(1573) := b"1111111111111111_1111111111111111_1111110111010010_0110101010101110"; -- -0.008508045653760163
	pesos_i(1574) := b"1111111111111111_1111111111111111_1111001110001100_0101111101101001"; -- -0.04863933261972264
	pesos_i(1575) := b"0000000000000000_0000000000000000_0001011010010000_0000010100011100"; -- 0.08813507024958571
	pesos_i(1576) := b"0000000000000000_0000000000000000_0001111000010110_0000110001110111"; -- 0.11752393624893709
	pesos_i(1577) := b"0000000000000000_0000000000000000_0001111111000000_1100111011101100"; -- 0.12403577094895527
	pesos_i(1578) := b"0000000000000000_0000000000000000_0011000010000101_0011101100000010"; -- 0.18953293619940337
	pesos_i(1579) := b"0000000000000000_0000000000000000_0001000011010110_0010111111001011"; -- 0.06576822949723327
	pesos_i(1580) := b"1111111111111111_1111111111111111_1101101010001110_0001001110001000"; -- -0.14626958783538202
	pesos_i(1581) := b"1111111111111111_1111111111111111_1101001111001000_0011011000011000"; -- -0.17272626789761228
	pesos_i(1582) := b"1111111111111111_1111111111111111_1101101111111110_1000011100100111"; -- -0.1406474619793785
	pesos_i(1583) := b"0000000000000000_0000000000000000_0001110111010110_0001011100110111"; -- 0.11654801457265777
	pesos_i(1584) := b"0000000000000000_0000000000000000_0011000011110010_0011110100101111"; -- 0.19119627367248015
	pesos_i(1585) := b"1111111111111111_1111111111111111_1110010000000001_1001110010101011"; -- -0.10935040301104702
	pesos_i(1586) := b"0000000000000000_0000000000000000_0000010011110001_1000001011001101"; -- 0.01931016443527992
	pesos_i(1587) := b"0000000000000000_0000000000000000_0001100001101000_1111100101100000"; -- 0.09535177795704868
	pesos_i(1588) := b"0000000000000000_0000000000000000_0001001011110101_1100100000010010"; -- 0.07406282842084429
	pesos_i(1589) := b"1111111111111111_1111111111111111_1110111111010000_0000011001111101"; -- -0.06323203516777166
	pesos_i(1590) := b"1111111111111111_1111111111111111_1110001000011001_1100101111111101"; -- -0.11679387168617557
	pesos_i(1591) := b"0000000000000000_0000000000000000_0000001111000110_0110111100010101"; -- 0.01474661128080226
	pesos_i(1592) := b"1111111111111111_1111111111111111_1110000110001111_0111110101111100"; -- -0.11890426373826393
	pesos_i(1593) := b"0000000000000000_0000000000000000_0001010101101101_0011000001111100"; -- 0.08369734786351335
	pesos_i(1594) := b"1111111111111111_1111111111111111_1110011111100100_0010101110011101"; -- -0.09417464653810574
	pesos_i(1595) := b"0000000000000000_0000000000000000_0010011001100001_1001000001010111"; -- 0.14992620593409128
	pesos_i(1596) := b"0000000000000000_0000000000000000_0001001000100110_1100100000110001"; -- 0.07090426631594066
	pesos_i(1597) := b"1111111111111111_1111111111111111_1110000000100001_1111100100101101"; -- -0.12448160802407265
	pesos_i(1598) := b"0000000000000000_0000000000000000_0011000001110011_1011100110101010"; -- 0.1892658272990472
	pesos_i(1599) := b"0000000000000000_0000000000000000_0001111011011100_0010010101111111"; -- 0.120546668528385
	pesos_i(1600) := b"0000000000000000_0000000000000000_0001111100100100_0000000111011010"; -- 0.12164317683892767
	pesos_i(1601) := b"0000000000000000_0000000000000000_0010111000001001_0000100000011111"; -- 0.17982531305703697
	pesos_i(1602) := b"0000000000000000_0000000000000000_0011000010010100_0010101010001011"; -- 0.18976083661981535
	pesos_i(1603) := b"0000000000000000_0000000000000000_0010000111111010_1011101110000010"; -- 0.13273212355245184
	pesos_i(1604) := b"1111111111111111_1111111111111111_1101110001110100_0010111110111101"; -- -0.13885213514720435
	pesos_i(1605) := b"1111111111111111_1111111111111111_1101000111011100_0111000001100100"; -- -0.18023011730530122
	pesos_i(1606) := b"0000000000000000_0000000000000000_0001010001110101_1101110101000100"; -- 0.0799234668792827
	pesos_i(1607) := b"0000000000000000_0000000000000000_0001101010000100_1101111111011001"; -- 0.10359000261460716
	pesos_i(1608) := b"1111111111111111_1111111111111111_1111111011100001_1011010001111001"; -- -0.0043685153906891094
	pesos_i(1609) := b"1111111111111111_1111111111111111_1101010011100111_1111100001110010"; -- -0.16833541127972682
	pesos_i(1610) := b"1111111111111111_1111111111111111_1111100110101111_1110101000001110"; -- -0.024659511213615815
	pesos_i(1611) := b"1111111111111111_1111111111111111_1101110001100110_1011011000011010"; -- -0.13905774947160165
	pesos_i(1612) := b"0000000000000000_0000000000000000_0001110011001010_1001100000001001"; -- 0.11246633750851953
	pesos_i(1613) := b"1111111111111111_1111111111111111_1111111010000111_0111111110010111"; -- -0.005744958545663786
	pesos_i(1614) := b"1111111111111111_1111111111111111_1110100111101110_0111101001011111"; -- -0.0862048643790483
	pesos_i(1615) := b"0000000000000000_0000000000000000_0010011001010101_0110000011100011"; -- 0.14974027192596195
	pesos_i(1616) := b"1111111111111111_1111111111111111_1111101101100110_0100111001111110"; -- -0.017970175007170464
	pesos_i(1617) := b"1111111111111111_1111111111111111_1110000000101010_0110110100000010"; -- -0.12435263355842095
	pesos_i(1618) := b"1111111111111111_1111111111111111_1101110111011110_1111010100000100"; -- -0.13331669478144006
	pesos_i(1619) := b"1111111111111111_1111111111111111_1101000000100010_0100101010010100"; -- -0.1869767559530988
	pesos_i(1620) := b"0000000000000000_0000000000000000_0001111001001111_1001000000111110"; -- 0.11840154178243295
	pesos_i(1621) := b"1111111111111111_1111111111111111_1111010000001001_1110100100001010"; -- -0.04672378074909961
	pesos_i(1622) := b"1111111111111111_1111111111111111_1101001000010001_1011011011011000"; -- -0.17941720216809157
	pesos_i(1623) := b"1111111111111111_1111111111111111_1101110011010001_0011100000011001"; -- -0.13743256931560988
	pesos_i(1624) := b"1111111111111111_1111111111111111_1101001001101111_1010110101011011"; -- -0.177983441723784
	pesos_i(1625) := b"1111111111111111_1111111111111111_1110110001000100_0001111111001111"; -- -0.07708550644287698
	pesos_i(1626) := b"1111111111111111_1111111111111111_1111110011011100_1110110111000011"; -- -0.012253894603438259
	pesos_i(1627) := b"1111111111111111_1111111111111111_1110111100100011_0011010001010001"; -- -0.06586907411875739
	pesos_i(1628) := b"1111111111111111_1111111111111111_1111011000000111_0110101110111011"; -- -0.038949267292397144
	pesos_i(1629) := b"1111111111111111_1111111111111111_1101010101000110_1001011000110110"; -- -0.16689168152376851
	pesos_i(1630) := b"1111111111111111_1111111111111111_1111011010010100_0001100010000111"; -- -0.03680273734915118
	pesos_i(1631) := b"0000000000000000_0000000000000000_0001110001111111_0011001111000011"; -- 0.11131595150781404
	pesos_i(1632) := b"1111111111111111_1111111111111111_1101100110000011_0101101001100010"; -- -0.15033946141702098
	pesos_i(1633) := b"0000000000000000_0000000000000000_0001001101000010_0010100000111111"; -- 0.07522822897716347
	pesos_i(1634) := b"0000000000000000_0000000000000000_0000110101000011_1110010010100100"; -- 0.05181721692389682
	pesos_i(1635) := b"1111111111111111_1111111111111111_1111111001001001_1001001110110010"; -- -0.00668980514678566
	pesos_i(1636) := b"1111111111111111_1111111111111111_1101001110000101_0110010110101010"; -- -0.17374577134687416
	pesos_i(1637) := b"0000000000000000_0000000000000000_0001000010111001_0110101011100001"; -- 0.06532924645941462
	pesos_i(1638) := b"0000000000000000_0000000000000000_0010111111110000_0111101101000010"; -- 0.18726320610750435
	pesos_i(1639) := b"0000000000000000_0000000000000000_0000111101111101_0010111100000101"; -- 0.060503901280105965
	pesos_i(1640) := b"0000000000000000_0000000000000000_0000100010101011_1100000001000101"; -- 0.03387071304172312
	pesos_i(1641) := b"0000000000000000_0000000000000000_0000010111111010_1110011100100110"; -- 0.023359724725031422
	pesos_i(1642) := b"0000000000000000_0000000000000000_0001001100100101_0010010100111111"; -- 0.07478554525212816
	pesos_i(1643) := b"0000000000000000_0000000000000000_0001001001000010_1111111001111110"; -- 0.07133474890166536
	pesos_i(1644) := b"1111111111111111_1111111111111111_1111011010010011_1110011100000110"; -- -0.03680568786862645
	pesos_i(1645) := b"1111111111111111_1111111111111111_1101000001101101_0000111110110101"; -- -0.1858358557542454
	pesos_i(1646) := b"0000000000000000_0000000000000000_0000010110001100_1100100011111101"; -- 0.021679460413530832
	pesos_i(1647) := b"1111111111111111_1111111111111111_1111011000011011_0011110011101010"; -- -0.038646881839236036
	pesos_i(1648) := b"0000000000000000_0000000000000000_0000110100111101_1001000110001110"; -- 0.05172071179466159
	pesos_i(1649) := b"1111111111111111_1111111111111111_1100111111111101_1010110100001101"; -- -0.18753546166867582
	pesos_i(1650) := b"1111111111111111_1111111111111111_1111101010010101_0000000000101011"; -- -0.02116393037500114
	pesos_i(1651) := b"1111111111111111_1111111111111111_1110010100110000_0000001111111010"; -- -0.10473609117715907
	pesos_i(1652) := b"1111111111111111_1111111111111111_1111001100001110_1111101011110111"; -- -0.05055266839312944
	pesos_i(1653) := b"0000000000000000_0000000000000000_0010010011001001_1001001101001010"; -- 0.1437007958052443
	pesos_i(1654) := b"1111111111111111_1111111111111111_1101110000101010_1111101010010111"; -- -0.13996919455487983
	pesos_i(1655) := b"1111111111111111_1111111111111111_1111101101101001_1010100010011111"; -- -0.017919026591430992
	pesos_i(1656) := b"0000000000000000_0000000000000000_0001110000101010_1100101011111111"; -- 0.11002796862461678
	pesos_i(1657) := b"1111111111111111_1111111111111111_1110001001001100_1100111001011111"; -- -0.11601553125540306
	pesos_i(1658) := b"0000000000000000_0000000000000000_0001101110111001_0101110100110101"; -- 0.10829718149037654
	pesos_i(1659) := b"0000000000000000_0000000000000000_0000100001001001_0111001111010000"; -- 0.03237079457706729
	pesos_i(1660) := b"1111111111111111_1111111111111111_1101000000100100_0011001110110110"; -- -0.18694760149498987
	pesos_i(1661) := b"1111111111111111_1111111111111111_1101001101110011_0110101111011000"; -- -0.17402006116945107
	pesos_i(1662) := b"1111111111111111_1111111111111111_1101111100110110_0110101110000111"; -- -0.12807586628896694
	pesos_i(1663) := b"0000000000000000_0000000000000000_0000010111000001_1001111101101110"; -- 0.022485698978478103
	pesos_i(1664) := b"1111111111111111_1111111111111111_1111000000101001_1010000110111011"; -- -0.061864749696020405
	pesos_i(1665) := b"1111111111111111_1111111111111111_1101111111000110_0111101110100011"; -- -0.1258776405171193
	pesos_i(1666) := b"1111111111111111_1111111111111111_1101011101100101_0010101001111001"; -- -0.15861258066798473
	pesos_i(1667) := b"0000000000000000_0000000000000000_0001110010011101_1011110101101101"; -- 0.11178192042429269
	pesos_i(1668) := b"0000000000000000_0000000000000000_0001000010101000_1011101100000010"; -- 0.06507462316176083
	pesos_i(1669) := b"1111111111111111_1111111111111111_1111010111110110_1111100010010010"; -- -0.03920027192458381
	pesos_i(1670) := b"0000000000000000_0000000000000000_0001100001111001_1101011000001001"; -- 0.09560907097485388
	pesos_i(1671) := b"1111111111111111_1111111111111111_1110010110011101_0011001000110011"; -- -0.10307012802764237
	pesos_i(1672) := b"0000000000000000_0000000000000000_0000110000000101_0010110110101101"; -- 0.04695401640816377
	pesos_i(1673) := b"0000000000000000_0000000000000000_0001110010000111_0100100101110000"; -- 0.11143931368392423
	pesos_i(1674) := b"0000000000000000_0000000000000000_0001100001011010_1010010111010011"; -- 0.09513317487913758
	pesos_i(1675) := b"0000000000000000_0000000000000000_0010111110001000_0001111011011111"; -- 0.18567078529601355
	pesos_i(1676) := b"1111111111111111_1111111111111111_1101110111111000_0101101010110110"; -- -0.13292916355366152
	pesos_i(1677) := b"1111111111111111_1111111111111111_1101101010001011_1010010110101110"; -- -0.14630665297438408
	pesos_i(1678) := b"1111111111111111_1111111111111111_1110101100011111_0110100101001011"; -- -0.08155195165578767
	pesos_i(1679) := b"1111111111111111_1111111111111111_1111110110110100_0110111100011000"; -- -0.00896554636614108
	pesos_i(1680) := b"0000000000000000_0000000000000000_0000110100101100_0101111101111010"; -- 0.051458327536464926
	pesos_i(1681) := b"0000000000000000_0000000000000000_0010001011000000_0100000111100001"; -- 0.13574611422786415
	pesos_i(1682) := b"1111111111111111_1111111111111111_1110010011111010_0010001110010000"; -- -0.10555818311727744
	pesos_i(1683) := b"0000000000000000_0000000000000000_0001011001101011_0011110100010011"; -- 0.0875738308507143
	pesos_i(1684) := b"0000000000000000_0000000000000000_0010101101010110_1001011010110101"; -- 0.16928998860158817
	pesos_i(1685) := b"0000000000000000_0000000000000000_0000101001111110_0011010000010110"; -- 0.04098821191915747
	pesos_i(1686) := b"0000000000000000_0000000000000000_0010001100101111_1011010011100111"; -- 0.13744669581384966
	pesos_i(1687) := b"0000000000000000_0000000000000000_0000101101100011_1100111001010000"; -- 0.04449166733777249
	pesos_i(1688) := b"1111111111111111_1111111111111111_1110010000111100_1011100100011110"; -- -0.10844843882920442
	pesos_i(1689) := b"1111111111111111_1111111111111111_1101111001100110_1111000111101001"; -- -0.13124168452379148
	pesos_i(1690) := b"1111111111111111_1111111111111111_1110111101001101_0111101001001100"; -- -0.06522403387288442
	pesos_i(1691) := b"1111111111111111_1111111111111111_1101100100000111_0010000110001011"; -- -0.15223493917491868
	pesos_i(1692) := b"0000000000000000_0000000000000000_0001001100000110_0111101111010010"; -- 0.07431768305351788
	pesos_i(1693) := b"1111111111111111_1111111111111111_1111111111001110_1101000101010001"; -- -0.0007504632119270382
	pesos_i(1694) := b"0000000000000000_0000000000000000_0000011011011100_1110101100101000"; -- 0.026808450103856796
	pesos_i(1695) := b"1111111111111111_1111111111111111_1111000110101000_0110100000010101"; -- -0.05602406955594266
	pesos_i(1696) := b"1111111111111111_1111111111111111_1101010010110101_1101001001110111"; -- -0.16910061455035558
	pesos_i(1697) := b"0000000000000000_0000000000000000_0000110101010001_0010000110111101"; -- 0.05201922287823382
	pesos_i(1698) := b"1111111111111111_1111111111111111_1111101111010011_0100100001000101"; -- -0.01630733779787155
	pesos_i(1699) := b"1111111111111111_1111111111111111_1101110111000111_0011101001010101"; -- -0.1336787740039001
	pesos_i(1700) := b"0000000000000000_0000000000000000_0010110100000010_0000011100101001"; -- 0.17581219445470006
	pesos_i(1701) := b"0000000000000000_0000000000000000_0010110000001010_1001000101100011"; -- 0.17203625352444338
	pesos_i(1702) := b"0000000000000000_0000000000000000_0001110001010101_0000010111010110"; -- 0.11067234492124123
	pesos_i(1703) := b"1111111111111111_1111111111111111_1101011110110011_1110101110001110"; -- -0.15741088654216415
	pesos_i(1704) := b"0000000000000000_0000000000000000_0001101111000100_1010001001101000"; -- 0.10846915277803713
	pesos_i(1705) := b"0000000000000000_0000000000000000_0001000000001001_0110011001011010"; -- 0.06264342979995095
	pesos_i(1706) := b"1111111111111111_1111111111111111_1111010111101101_0010001101001011"; -- -0.03935031338695799
	pesos_i(1707) := b"0000000000000000_0000000000000000_0010000001011011_0000111011101101"; -- 0.1263894393899177
	pesos_i(1708) := b"0000000000000000_0000000000000000_0010110100100010_0111101101011101"; -- 0.17630740191565702
	pesos_i(1709) := b"1111111111111111_1111111111111111_1110110110011011_0000101111101101"; -- -0.07185292684828691
	pesos_i(1710) := b"0000000000000000_0000000000000000_0000110011101001_0101000000011001"; -- 0.050435072072146446
	pesos_i(1711) := b"1111111111111111_1111111111111111_1111100100010111_0001110110010001"; -- -0.026991035634294502
	pesos_i(1712) := b"0000000000000000_0000000000000000_0010010011100001_0111011011110011"; -- 0.14406531747155246
	pesos_i(1713) := b"1111111111111111_1111111111111111_1110110010001101_0011010000000000"; -- -0.07597041122446369
	pesos_i(1714) := b"0000000000000000_0000000000000000_0000110010001100_0011111001100101"; -- 0.04901494945968543
	pesos_i(1715) := b"1111111111111111_1111111111111111_1110011001110100_1010010000101101"; -- -0.09978269472879388
	pesos_i(1716) := b"1111111111111111_1111111111111111_1111001000011111_1011111000100011"; -- -0.05420314445482885
	pesos_i(1717) := b"0000000000000000_0000000000000000_0001100000001010_1011001001001011"; -- 0.09391321489184859
	pesos_i(1718) := b"0000000000000000_0000000000000000_0000100011011011_1011110101100000"; -- 0.034602962524140586
	pesos_i(1719) := b"0000000000000000_0000000000000000_0000101101001011_1111111010000111"; -- 0.044128330199397645
	pesos_i(1720) := b"0000000000000000_0000000000000000_0000010101001010_1001110101010000"; -- 0.020669776952888172
	pesos_i(1721) := b"1111111111111111_1111111111111111_1110000010111100_0000111100101101"; -- -0.12213044302740175
	pesos_i(1722) := b"1111111111111111_1111111111111111_1111000010001101_0001100000011111"; -- -0.060347072927743994
	pesos_i(1723) := b"1111111111111111_1111111111111111_1111011110100011_1101111111101010"; -- -0.03265572111352758
	pesos_i(1724) := b"1111111111111111_1111111111111111_1101010010010111_1111011110011111"; -- -0.16955616349569017
	pesos_i(1725) := b"1111111111111111_1111111111111111_1111110100010110_1001011111110001"; -- -0.011374000135083436
	pesos_i(1726) := b"1111111111111111_1111111111111111_1101111101000111_1100001101001011"; -- -0.12781123553586016
	pesos_i(1727) := b"0000000000000000_0000000000000000_0001101111001100_1111001010001001"; -- 0.10859599929139703
	pesos_i(1728) := b"0000000000000000_0000000000000000_0001001011000000_0100000001110011"; -- 0.0732460288669527
	pesos_i(1729) := b"0000000000000000_0000000000000000_0001011111111100_0001001111110110"; -- 0.09369015451361194
	pesos_i(1730) := b"0000000000000000_0000000000000000_0001101001100100_1011011111110000"; -- 0.10309934238449374
	pesos_i(1731) := b"0000000000000000_0000000000000000_0010100001101101_0100100011011110"; -- 0.15791755133410576
	pesos_i(1732) := b"1111111111111111_1111111111111111_1110111100000000_1101100010010011"; -- -0.06639334113156264
	pesos_i(1733) := b"0000000000000000_0000000000000000_0000010110000010_0100110011001001"; -- 0.021519469309006816
	pesos_i(1734) := b"0000000000000000_0000000000000000_0001000111001000_1010101100001011"; -- 0.06946820279092895
	pesos_i(1735) := b"1111111111111111_1111111111111111_1111010110001000_1011111100101110"; -- -0.04088215952898135
	pesos_i(1736) := b"0000000000000000_0000000000000000_0000001101100001_1011100110110011"; -- 0.01320992102857552
	pesos_i(1737) := b"0000000000000000_0000000000000000_0010000100010101_0000100011000111"; -- 0.1292272076266321
	pesos_i(1738) := b"0000000000000000_0000000000000000_0001010101000110_0010010010110001"; -- 0.08310155229659878
	pesos_i(1739) := b"0000000000000000_0000000000000000_0000000101001110_1110101010111010"; -- 0.0051104264306137594
	pesos_i(1740) := b"1111111111111111_1111111111111111_1110111001111110_1111110110111011"; -- -0.06837476913096142
	pesos_i(1741) := b"1111111111111111_1111111111111111_1111111101111011_1111111110111011"; -- -0.002014176133507817
	pesos_i(1742) := b"0000000000000000_0000000000000000_0001100000110111_0001011010110100"; -- 0.09459058652957514
	pesos_i(1743) := b"1111111111111111_1111111111111111_1100010101100101_0000000001111101"; -- -0.22892758328375484
	pesos_i(1744) := b"0000000000000000_0000000000000000_0000101100110100_1100101001011010"; -- 0.043774268177223234
	pesos_i(1745) := b"1111111111111111_1111111111111111_1101011101011001_0101011110100111"; -- -0.15879299325832708
	pesos_i(1746) := b"1111111111111111_1111111111111111_1111111110001110_1100011010011100"; -- -0.001727663838341752
	pesos_i(1747) := b"1111111111111111_1111111111111111_1111111000010000_1111110000101000"; -- -0.007553329684258536
	pesos_i(1748) := b"0000000000000000_0000000000000000_0010101100011101_0001001000111100"; -- 0.16841234176837822
	pesos_i(1749) := b"1111111111111111_1111111111111111_1111101011011101_0000001101010100"; -- -0.020065109216970734
	pesos_i(1750) := b"0000000000000000_0000000000000000_0000110001111101_1101001011010011"; -- 0.04879491472039107
	pesos_i(1751) := b"1111111111111111_1111111111111111_1111011011001111_0000101101010111"; -- -0.03590325466049313
	pesos_i(1752) := b"0000000000000000_0000000000000000_0001010011001100_0100111101101100"; -- 0.08124252685842005
	pesos_i(1753) := b"1111111111111111_1111111111111111_1101110011101111_0010111000010100"; -- -0.1369754030514223
	pesos_i(1754) := b"0000000000000000_0000000000000000_0001010101000100_1111111101111010"; -- 0.08308407530807858
	pesos_i(1755) := b"0000000000000000_0000000000000000_0001001110001111_1111110001110010"; -- 0.07641580376919921
	pesos_i(1756) := b"1111111111111111_1111111111111111_1111010011000001_1010001010101111"; -- -0.043920357041360256
	pesos_i(1757) := b"0000000000000000_0000000000000000_0001010101101011_0111000111001010"; -- 0.08367072275367629
	pesos_i(1758) := b"0000000000000000_0000000000000000_0001000010001001_0011001110010100"; -- 0.06459352845981914
	pesos_i(1759) := b"1111111111111111_1111111111111111_1101100101011111_1000011110000011"; -- -0.15088608801232622
	pesos_i(1760) := b"0000000000000000_0000000000000000_0010000100100001_0111000000001010"; -- 0.12941646815207267
	pesos_i(1761) := b"1111111111111111_1111111111111111_1110101010111110_0110000000110111"; -- -0.0830325952995767
	pesos_i(1762) := b"0000000000000000_0000000000000000_0001110110100011_0010101010111010"; -- 0.11577097921443996
	pesos_i(1763) := b"1111111111111111_1111111111111111_1111001100100010_0011100010001110"; -- -0.05025908019805372
	pesos_i(1764) := b"0000000000000000_0000000000000000_0001011011010010_0000011001101011"; -- 0.08914222834979221
	pesos_i(1765) := b"1111111111111111_1111111111111111_1110011110001110_0010111010101100"; -- -0.09548672009246716
	pesos_i(1766) := b"0000000000000000_0000000000000000_0000011000011101_1010011111010110"; -- 0.023890008688898616
	pesos_i(1767) := b"1111111111111111_1111111111111111_1110110110100001_1110010101001101"; -- -0.07174841766140153
	pesos_i(1768) := b"1111111111111111_1111111111111111_1111110000101101_1110111110110011"; -- -0.014924067309912489
	pesos_i(1769) := b"1111111111111111_1111111111111111_1101110010110001_1110011010101000"; -- -0.13791044608080594
	pesos_i(1770) := b"1111111111111111_1111111111111111_1111000111000011_1100001111110110"; -- -0.05560660593181174
	pesos_i(1771) := b"1111111111111111_1111111111111111_1101101010010111_1100011011100000"; -- -0.1461215688878196
	pesos_i(1772) := b"0000000000000000_0000000000000000_0010100010010111_1100000100001101"; -- 0.15856558386104497
	pesos_i(1773) := b"0000000000000000_0000000000000000_0000100011001011_1010111111111001"; -- 0.034358023047673276
	pesos_i(1774) := b"1111111111111111_1111111111111111_1111101110001100_1110100111010001"; -- -0.01738108309262693
	pesos_i(1775) := b"0000000000000000_0000000000000000_0001100010010011_0110101101111010"; -- 0.095999448033584
	pesos_i(1776) := b"1111111111111111_1111111111111111_1111101011100000_1110011000100101"; -- -0.020005813488428795
	pesos_i(1777) := b"1111111111111111_1111111111111111_1100011000100011_0001100010001101"; -- -0.22602697896851362
	pesos_i(1778) := b"0000000000000000_0000000000000000_0000110010011011_1100011111100101"; -- 0.04925202685907654
	pesos_i(1779) := b"1111111111111111_1111111111111111_1101011100011011_0000000010111000"; -- -0.1597442197533712
	pesos_i(1780) := b"1111111111111111_1111111111111111_1101010100001010_1101000100000111"; -- -0.16780370305936682
	pesos_i(1781) := b"0000000000000000_0000000000000000_0010001101110110_1011101001100000"; -- 0.13853039584176136
	pesos_i(1782) := b"0000000000000000_0000000000000000_0010001100000101_0110010101110010"; -- 0.13680109060109216
	pesos_i(1783) := b"1111111111111111_1111111111111111_1101010001010100_1001101000010101"; -- -0.17058407765919675
	pesos_i(1784) := b"0000000000000000_0000000000000000_0010010001101001_1100011110001010"; -- 0.1422390662880553
	pesos_i(1785) := b"1111111111111111_1111111111111111_1111101000101101_1110010010000111"; -- -0.02273723309431939
	pesos_i(1786) := b"1111111111111111_1111111111111111_1111011001001000_0000110110010101"; -- -0.037963057710153125
	pesos_i(1787) := b"0000000000000000_0000000000000000_0001101001111100_0110011101000011"; -- 0.10346074471861649
	pesos_i(1788) := b"1111111111111111_1111111111111111_1111111110010011_1110011001110010"; -- -0.0016494725022848876
	pesos_i(1789) := b"0000000000000000_0000000000000000_0001000010000011_0001000100100001"; -- 0.06449992238599091
	pesos_i(1790) := b"1111111111111111_1111111111111111_1111000111001010_0110001010000010"; -- -0.05550560297640891
	pesos_i(1791) := b"0000000000000000_0000000000000000_0000011010001111_0011010001110110"; -- 0.025622633861319632
	pesos_i(1792) := b"0000000000000000_0000000000000000_0010011100001100_0000100010000000"; -- 0.15252736206809275
	pesos_i(1793) := b"0000000000000000_0000000000000000_0000110011001111_0111011110110000"; -- 0.050040703216261605
	pesos_i(1794) := b"0000000000000000_0000000000000000_0010001110100101_1101010111100111"; -- 0.13924919974808014
	pesos_i(1795) := b"1111111111111111_1111111111111111_1100111110010110_0101110101001000"; -- -0.18911187171473137
	pesos_i(1796) := b"1111111111111111_1111111111111111_1101011101101011_1111101000101001"; -- -0.1585086489681316
	pesos_i(1797) := b"0000000000000000_0000000000000000_0001100001101011_1111101100010101"; -- 0.09539765617919616
	pesos_i(1798) := b"0000000000000000_0000000000000000_0001000010001010_0010001111001011"; -- 0.06460784631864817
	pesos_i(1799) := b"0000000000000000_0000000000000000_0001010010010000_1111111111100111"; -- 0.08033751856713278
	pesos_i(1800) := b"1111111111111111_1111111111111111_1101010110110100_0011101001100000"; -- -0.16521868860231534
	pesos_i(1801) := b"1111111111111111_1111111111111111_1110011110001000_0001011010000010"; -- -0.09557971304912864
	pesos_i(1802) := b"0000000000000000_0000000000000000_0000101011110100_1110110011101100"; -- 0.042799766252935266
	pesos_i(1803) := b"1111111111111111_1111111111111111_1110100010111110_0001000111001000"; -- -0.09084977031727594
	pesos_i(1804) := b"0000000000000000_0000000000000000_0000011111001111_0010011010110100"; -- 0.030504626319919372
	pesos_i(1805) := b"0000000000000000_0000000000000000_0001001000111111_0111110000011010"; -- 0.07128120078515807
	pesos_i(1806) := b"1111111111111111_1111111111111111_1101111111000101_1000001000101101"; -- -0.12589250955281084
	pesos_i(1807) := b"1111111111111111_1111111111111111_1111110000100101_0111110101010101"; -- -0.015052954545810064
	pesos_i(1808) := b"0000000000000000_0000000000000000_0000101110011000_0010000111000000"; -- 0.04529009769745657
	pesos_i(1809) := b"1111111111111111_1111111111111111_1101111100100100_1010000001010011"; -- -0.1283473776102594
	pesos_i(1810) := b"0000000000000000_0000000000000000_0010000001111110_1010010100000010"; -- 0.12693244274875276
	pesos_i(1811) := b"1111111111111111_1111111111111111_1111011010111011_0111111000100001"; -- -0.0362015886908984
	pesos_i(1812) := b"1111111111111111_1111111111111111_1111100100110111_1111110010011001"; -- -0.026489460591991396
	pesos_i(1813) := b"0000000000000000_0000000000000000_0010010000100110_1101101010110000"; -- 0.14121786878205192
	pesos_i(1814) := b"0000000000000000_0000000000000000_0000001111100000_0011101100001111"; -- 0.015140239009103943
	pesos_i(1815) := b"1111111111111111_1111111111111111_1101000001111101_1000111010001001"; -- -0.18558415561452093
	pesos_i(1816) := b"1111111111111111_1111111111111111_1111010001101111_0011011111000101"; -- -0.04517795038556497
	pesos_i(1817) := b"1111111111111111_1111111111111111_1110001100110000_1010111011011010"; -- -0.11253840618594892
	pesos_i(1818) := b"1111111111111111_1111111111111111_1110110000101111_1100010110010001"; -- -0.07739606100831198
	pesos_i(1819) := b"1111111111111111_1111111111111111_1111011100010110_1001000001101111"; -- -0.034811947737197375
	pesos_i(1820) := b"0000000000000000_0000000000000000_0001110011101101_0001100001100110"; -- 0.11299278725236328
	pesos_i(1821) := b"0000000000000000_0000000000000000_0000001010100001_1010111101010000"; -- 0.010279614474114695
	pesos_i(1822) := b"1111111111111111_1111111111111111_1110001110111100_1101101111000101"; -- -0.11039949840056307
	pesos_i(1823) := b"0000000000000000_0000000000000000_0000110101001101_0010001010000001"; -- 0.05195823342248779
	pesos_i(1824) := b"1111111111111111_1111111111111111_1101011100001111_0101111010110101"; -- -0.15992172310552108
	pesos_i(1825) := b"0000000000000000_0000000000000000_0010000101000110_0011011111011101"; -- 0.12997769488337388
	pesos_i(1826) := b"0000000000000000_0000000000000000_0010001111010101_1111001011011100"; -- 0.13998334761172104
	pesos_i(1827) := b"0000000000000000_0000000000000000_0000001110011001_1000111110100000"; -- 0.01406190547432376
	pesos_i(1828) := b"1111111111111111_1111111111111111_1101001100000010_1100111110101010"; -- -0.17573835465844317
	pesos_i(1829) := b"0000000000000000_0000000000000000_0000000000001110_0001110001011100"; -- 0.00021531343365385975
	pesos_i(1830) := b"1111111111111111_1111111111111111_1101110000000110_1010001001101111"; -- -0.14052376550278117
	pesos_i(1831) := b"0000000000000000_0000000000000000_0001000101000010_0010011011001101"; -- 0.06741564277468587
	pesos_i(1832) := b"1111111111111111_1111111111111111_1111101100011100_1111001010101010"; -- -0.019089539907026155
	pesos_i(1833) := b"1111111111111111_1111111111111111_1101110000111000_0101000010110101"; -- -0.1397656972066511
	pesos_i(1834) := b"1111111111111111_1111111111111111_1110111001110011_1010110100101000"; -- -0.06854741831377988
	pesos_i(1835) := b"1111111111111111_1111111111111111_1101000010011000_0010110010111110"; -- -0.18517799729006656
	pesos_i(1836) := b"0000000000000000_0000000000000000_0010111101011110_1100001110001101"; -- 0.1850397319873465
	pesos_i(1837) := b"1111111111111111_1111111111111111_1101010100011011_1011111000100010"; -- -0.16754543000675923
	pesos_i(1838) := b"1111111111111111_1111111111111111_1100010000101110_1101001011110010"; -- -0.23366052236794813
	pesos_i(1839) := b"0000000000000000_0000000000000000_0001010111111100_1010001001100110"; -- 0.08588614452902751
	pesos_i(1840) := b"1111111111111111_1111111111111111_1111100110011010_0001001100100110"; -- -0.024992755116935654
	pesos_i(1841) := b"0000000000000000_0000000000000000_0010110111001100_1010110111000001"; -- 0.17890439943894912
	pesos_i(1842) := b"1111111111111111_1111111111111111_1101010011000110_1111101110011001"; -- -0.16883876346722246
	pesos_i(1843) := b"0000000000000000_0000000000000000_0001101001000010_1110101110011011"; -- 0.10258362320579943
	pesos_i(1844) := b"0000000000000000_0000000000000000_0000010001100111_0101010111101000"; -- 0.017201775786482458
	pesos_i(1845) := b"1111111111111111_1111111111111111_1110101000000011_1000110011000100"; -- -0.08588333340373809
	pesos_i(1846) := b"1111111111111111_1111111111111111_1110011000110010_0000100010101000"; -- -0.10079904465201409
	pesos_i(1847) := b"1111111111111111_1111111111111111_1101101011000110_1110101110010100"; -- -0.14540221831006045
	pesos_i(1848) := b"1111111111111111_1111111111111111_1110001011000010_0110011011110100"; -- -0.11422115835604368
	pesos_i(1849) := b"0000000000000000_0000000000000000_0010011101011111_0010110110001001"; -- 0.15379604912301115
	pesos_i(1850) := b"1111111111111111_1111111111111111_1111001111000111_0111000111001110"; -- -0.04773796764888318
	pesos_i(1851) := b"0000000000000000_0000000000000000_0000111000111010_1111010010001110"; -- 0.05558708643758509
	pesos_i(1852) := b"1111111111111111_1111111111111111_1111101011000101_1100101011111101"; -- -0.020419419600498867
	pesos_i(1853) := b"0000000000000000_0000000000000000_0010000010001110_1011001101010100"; -- 0.1271774367774028
	pesos_i(1854) := b"0000000000000000_0000000000000000_0001001110010101_0001110001000100"; -- 0.07649399435554759
	pesos_i(1855) := b"1111111111111111_1111111111111111_1101101110001101_0100011111000110"; -- -0.14237548271384098
	pesos_i(1856) := b"0000000000000000_0000000000000000_0001101110110110_0001100001111011"; -- 0.10824730882680385
	pesos_i(1857) := b"0000000000000000_0000000000000000_0001011111001000_0101100010000101"; -- 0.09290078401526258
	pesos_i(1858) := b"1111111111111111_1111111111111111_1101000010010100_1000000000101011"; -- -0.18523405982273847
	pesos_i(1859) := b"0000000000000000_0000000000000000_0010000100100000_1110011111010111"; -- 0.1294083500298358
	pesos_i(1860) := b"0000000000000000_0000000000000000_0000101010001010_1001101111011001"; -- 0.041177502141659716
	pesos_i(1861) := b"1111111111111111_1111111111111111_1101000101000001_1001110011110110"; -- -0.1825925731292346
	pesos_i(1862) := b"0000000000000000_0000000000000000_0010000011110110_1101100101001000"; -- 0.12876661309112525
	pesos_i(1863) := b"1111111111111111_1111111111111111_1111001011001000_0000111110011101"; -- -0.05163481164358838
	pesos_i(1864) := b"0000000000000000_0000000000000000_0001111101100101_0101000010100111"; -- 0.12263969501712244
	pesos_i(1865) := b"1111111111111111_1111111111111111_1111000011110000_1111100001100000"; -- -0.05882308630210319
	pesos_i(1866) := b"0000000000000000_0000000000000000_0000111110000010_0001101011000100"; -- 0.06057898785044435
	pesos_i(1867) := b"1111111111111111_1111111111111111_1111111111010011_0000001100001101"; -- -0.0006864636812313142
	pesos_i(1868) := b"1111111111111111_1111111111111111_1101000110011011_1001101100000111"; -- -0.18121939726144146
	pesos_i(1869) := b"1111111111111111_1111111111111111_1101100010011111_0010000110010010"; -- -0.15382185157461434
	pesos_i(1870) := b"1111111111111111_1111111111111111_1101101011001011_0000110001000100"; -- -0.14533923474927482
	pesos_i(1871) := b"1111111111111111_1111111111111111_1111111101010100_1110010101011100"; -- -0.0026108409375736417
	pesos_i(1872) := b"0000000000000000_0000000000000000_0010000001011110_1100010111110111"; -- 0.12644612586453968
	pesos_i(1873) := b"1111111111111111_1111111111111111_1101100000010110_1100001100110110"; -- -0.15590267127833657
	pesos_i(1874) := b"1111111111111111_1111111111111111_1110010111000110_1000000100111101"; -- -0.10243980658499474
	pesos_i(1875) := b"1111111111111111_1111111111111111_1111010101000001_0110100010011000"; -- -0.04197069439168951
	pesos_i(1876) := b"1111111111111111_1111111111111111_1111001111111010_1101011100000011"; -- -0.046953736924266576
	pesos_i(1877) := b"1111111111111111_1111111111111111_1110101111110111_0110010101111011"; -- -0.07825628044399034
	pesos_i(1878) := b"0000000000000000_0000000000000000_0000010110111000_1000010010000100"; -- 0.022346765660797466
	pesos_i(1879) := b"0000000000000000_0000000000000000_0010001100010101_0010000111110011"; -- 0.13704120821464913
	pesos_i(1880) := b"1111111111111111_1111111111111111_1111110100110111_0101110100110110"; -- -0.010873960827469576
	pesos_i(1881) := b"1111111111111111_1111111111111111_1101110100011111_1101000000010101"; -- -0.13623332480023548
	pesos_i(1882) := b"0000000000000000_0000000000000000_0001101101000001_0110100011100000"; -- 0.1064668223714898
	pesos_i(1883) := b"1111111111111111_1111111111111111_1101011001001100_1011001010011111"; -- -0.16289218540059414
	pesos_i(1884) := b"1111111111111111_1111111111111111_1101010111110011_1000110100101001"; -- -0.16425245038966602
	pesos_i(1885) := b"0000000000000000_0000000000000000_0010001100111101_1011111011100010"; -- 0.1376609136043655
	pesos_i(1886) := b"1111111111111111_1111111111111111_1101101110111011_0100100000100001"; -- -0.1416735571419622
	pesos_i(1887) := b"1111111111111111_1111111111111111_1111111001110101_1010010010000001"; -- -0.0060174165219140825
	pesos_i(1888) := b"0000000000000000_0000000000000000_0000100001011110_0011100101100111"; -- 0.03268774759417972
	pesos_i(1889) := b"1111111111111111_1111111111111111_1110100100010010_0110100100110001"; -- -0.08956282195812756
	pesos_i(1890) := b"0000000000000000_0000000000000000_0001000010010011_1101010001010010"; -- 0.06475569729860443
	pesos_i(1891) := b"1111111111111111_1111111111111111_1100111101100101_0100010011011100"; -- -0.18986100803360734
	pesos_i(1892) := b"0000000000000000_0000000000000000_0010001100101010_1001001010001110"; -- 0.1373683545832614
	pesos_i(1893) := b"0000000000000000_0000000000000000_0001001100001001_0100011111001100"; -- 0.07436035854279201
	pesos_i(1894) := b"1111111111111111_1111111111111111_1111101110111010_1001010010100000"; -- -0.016684256489408716
	pesos_i(1895) := b"1111111111111111_1111111111111111_1100101111110001_1101111111100100"; -- -0.20334053681960954
	pesos_i(1896) := b"0000000000000000_0000000000000000_0000010011111101_0011011110010111"; -- 0.019488787033027005
	pesos_i(1897) := b"1111111111111111_1111111111111111_1101100111100010_0101010101101000"; -- -0.14889017298113247
	pesos_i(1898) := b"0000000000000000_0000000000000000_0001010010110110_1110001110011000"; -- 0.08091566522028001
	pesos_i(1899) := b"1111111111111111_1111111111111111_1111101000101110_1000100001000011"; -- -0.022727473814319336
	pesos_i(1900) := b"0000000000000000_0000000000000000_0000001001001001_1100010100111010"; -- 0.00893814724155951
	pesos_i(1901) := b"0000000000000000_0000000000000000_0010011001001110_1110010011011110"; -- 0.1496413271236311
	pesos_i(1902) := b"1111111111111111_1111111111111111_1111110011111011_0001000111000110"; -- -0.011793984508529606
	pesos_i(1903) := b"0000000000000000_0000000000000000_0010010010110101_1000000110100000"; -- 0.14339456711649318
	pesos_i(1904) := b"1111111111111111_1111111111111111_1110110000010010_1001000101011101"; -- -0.0778416775554202
	pesos_i(1905) := b"1111111111111111_1111111111111111_1110001110011000_1101110110110000"; -- -0.11094870050986083
	pesos_i(1906) := b"0000000000000000_0000000000000000_0001011001110111_0000000100001001"; -- 0.08775335768723243
	pesos_i(1907) := b"0000000000000000_0000000000000000_0010100000101010_0111010001001000"; -- 0.15689780000866718
	pesos_i(1908) := b"0000000000000000_0000000000000000_0000000001010010_1111010001001110"; -- 0.0012657824851931845
	pesos_i(1909) := b"0000000000000000_0000000000000000_0001010101000000_1010100101011111"; -- 0.08301790787780643
	pesos_i(1910) := b"0000000000000000_0000000000000000_0001101111000011_1100010100001001"; -- 0.10845595806893375
	pesos_i(1911) := b"0000000000000000_0000000000000000_0001111111001100_0110011010010010"; -- 0.12421265672582177
	pesos_i(1912) := b"1111111111111111_1111111111111111_1101011101010001_1000000101100011"; -- -0.15891257609323522
	pesos_i(1913) := b"0000000000000000_0000000000000000_0010100001000100_0100100000001111"; -- 0.15729189268754284
	pesos_i(1914) := b"0000000000000000_0000000000000000_0000000000000010_0101101001011110"; -- 3.590378888037879e-05
	pesos_i(1915) := b"1111111111111111_1111111111111111_1100111010001110_0100100100110010"; -- -0.1931413892513329
	pesos_i(1916) := b"0000000000000000_0000000000000000_0010010110110101_1010100111011111"; -- 0.147303215971968
	pesos_i(1917) := b"0000000000000000_0000000000000000_0001111010000111_0101011011111111"; -- 0.11925262197817212
	pesos_i(1918) := b"1111111111111111_1111111111111111_1111001000001110_1001011110001001"; -- -0.05446484469994223
	pesos_i(1919) := b"0000000000000000_0000000000000000_0001011001000011_0011011110101000"; -- 0.086963156180638
	pesos_i(1920) := b"1111111111111111_1111111111111111_1111011110001011_1111110000100110"; -- -0.03302024904183724
	pesos_i(1921) := b"1111111111111111_1111111111111111_1101101001110111_0011110001010011"; -- -0.14661810847633877
	pesos_i(1922) := b"1111111111111111_1111111111111111_1101001110110100_1000010110111011"; -- -0.17302669708141785
	pesos_i(1923) := b"1111111111111111_1111111111111111_1110010110101100_0100010111011000"; -- -0.10284007522065712
	pesos_i(1924) := b"1111111111111111_1111111111111111_1110101000110100_0111001110101111"; -- -0.08513714773649791
	pesos_i(1925) := b"0000000000000000_0000000000000000_0010010110001001_0101001110000001"; -- 0.14662668122736075
	pesos_i(1926) := b"0000000000000000_0000000000000000_0001100001000101_0101000001010101"; -- 0.09480764456546907
	pesos_i(1927) := b"1111111111111111_1111111111111111_1101000010011101_0110110011101110"; -- -0.18509787750271187
	pesos_i(1928) := b"1111111111111111_1111111111111111_1101110110110111_0100111001010110"; -- -0.13392172235193514
	pesos_i(1929) := b"1111111111111111_1111111111111111_1101000110010101_1010010010001110"; -- -0.18131038214480738
	pesos_i(1930) := b"1111111111111111_1111111111111111_1110101011111100_1101111011001010"; -- -0.0820790058278395
	pesos_i(1931) := b"0000000000000000_0000000000000000_0001110001111101_0100100001000111"; -- 0.11128665674922415
	pesos_i(1932) := b"1111111111111111_1111111111111111_1101101011011111_0001101110000101"; -- -0.1450331497560526
	pesos_i(1933) := b"0000000000000000_0000000000000000_0001000001010001_0100100110100100"; -- 0.06374035119589191
	pesos_i(1934) := b"1111111111111111_1111111111111111_1101010010011110_0101010010111100"; -- -0.16945906073049133
	pesos_i(1935) := b"1111111111111111_1111111111111111_1110101011000011_1101111010111010"; -- -0.08294876065082898
	pesos_i(1936) := b"0000000000000000_0000000000000000_0010001110111001_0100011111101000"; -- 0.13954591192663937
	pesos_i(1937) := b"1111111111111111_1111111111111111_1111111001100101_0101100010010110"; -- -0.006266082057414171
	pesos_i(1938) := b"0000000000000000_0000000000000000_0010000110010001_0001010111011101"; -- 0.13112007765398256
	pesos_i(1939) := b"0000000000000000_0000000000000000_0001100000011001_0110000110110000"; -- 0.09413729240036457
	pesos_i(1940) := b"1111111111111111_1111111111111111_1101101100001111_0100001010010010"; -- -0.14429840016141965
	pesos_i(1941) := b"0000000000000000_0000000000000000_0001100111010001_0001001001100000"; -- 0.10084643203358702
	pesos_i(1942) := b"1111111111111111_1111111111111111_1111011111111001_0000000010101110"; -- -0.03135677094304756
	pesos_i(1943) := b"1111111111111111_1111111111111111_1101001011100000_0010101110001101"; -- -0.1762669354197246
	pesos_i(1944) := b"1111111111111111_1111111111111111_1111011101100010_0011101011101111"; -- -0.033657375914944714
	pesos_i(1945) := b"0000000000000000_0000000000000000_0000011101110011_0011010000001101"; -- 0.029101613322463103
	pesos_i(1946) := b"1111111111111111_1111111111111111_1110010011100010_1101011011111001"; -- -0.10591370034430833
	pesos_i(1947) := b"1111111111111111_1111111111111111_1110100001110110_1000100010001001"; -- -0.09194132473444035
	pesos_i(1948) := b"0000000000000000_0000000000000000_0001011001011000_0101101011110001"; -- 0.0872856940114134
	pesos_i(1949) := b"0000000000000000_0000000000000000_0010100111100000_0101111110110000"; -- 0.16357992214358774
	pesos_i(1950) := b"1111111111111111_1111111111111111_1111111001010011_0011010001001110"; -- -0.00654290291811401
	pesos_i(1951) := b"1111111111111111_1111111111111111_1101110000000011_1101011010100101"; -- -0.14056642992029889
	pesos_i(1952) := b"0000000000000000_0000000000000000_0000000110001101_1111101100111010"; -- 0.006072713503345255
	pesos_i(1953) := b"0000000000000000_0000000000000000_0001101000000110_1101010010111011"; -- 0.10166673244800158
	pesos_i(1954) := b"1111111111111111_1111111111111111_1101101111011110_0000100000111110"; -- -0.14114330760157698
	pesos_i(1955) := b"1111111111111111_1111111111111111_1111011111011010_1001000001011011"; -- -0.0318212297793955
	pesos_i(1956) := b"0000000000000000_0000000000000000_0001110110110010_0000100011011110"; -- 0.11599784308493537
	pesos_i(1957) := b"0000000000000000_0000000000000000_0001001101010110_1110100001101110"; -- 0.07554485986035973
	pesos_i(1958) := b"1111111111111111_1111111111111111_1110001110111110_1001101100010100"; -- -0.11037283667005097
	pesos_i(1959) := b"1111111111111111_1111111111111111_1101011100111111_0101110011000010"; -- -0.15918941740984838
	pesos_i(1960) := b"0000000000000000_0000000000000000_0010101111011110_0010110111101011"; -- 0.17135893810367886
	pesos_i(1961) := b"1111111111111111_1111111111111111_1111100010100100_0100001001010110"; -- -0.028743604660564442
	pesos_i(1962) := b"0000000000000000_0000000000000000_0000011000101010_1100101000110011"; -- 0.024090421229212722
	pesos_i(1963) := b"1111111111111111_1111111111111111_1111011000011110_1110101001111111"; -- -0.03859075920689747
	pesos_i(1964) := b"1111111111111111_1111111111111111_1101010111010000_0101101101010111"; -- -0.16478947758396598
	pesos_i(1965) := b"1111111111111111_1111111111111111_1110110110001101_1000001010000010"; -- -0.07205948178907692
	pesos_i(1966) := b"1111111111111111_1111111111111111_1110001010001101_0000001001001111"; -- -0.11503587305504132
	pesos_i(1967) := b"0000000000000000_0000000000000000_0000000110111110_1011110001100111"; -- 0.0068166496283932005
	pesos_i(1968) := b"1111111111111111_1111111111111111_1110110011010111_1111001100110111"; -- -0.07482986358826839
	pesos_i(1969) := b"0000000000000000_0000000000000000_0000011000000111_1010111010011011"; -- 0.023554718817385172
	pesos_i(1970) := b"1111111111111111_1111111111111111_1110010101110100_0110010011010101"; -- -0.1036927203932584
	pesos_i(1971) := b"0000000000000000_0000000000000000_0000001111110101_1000000011100100"; -- 0.015464835894016187
	pesos_i(1972) := b"0000000000000000_0000000000000000_0000010000110101_1111011110001101"; -- 0.01644847089256277
	pesos_i(1973) := b"0000000000000000_0000000000000000_0000100101001011_1110101101100111"; -- 0.03631469020400218
	pesos_i(1974) := b"0000000000000000_0000000000000000_0001011010001100_1001010010110000"; -- 0.0880825928279133
	pesos_i(1975) := b"1111111111111111_1111111111111111_1111100001100111_0100011001111111"; -- -0.029674142899831772
	pesos_i(1976) := b"1111111111111111_1111111111111111_1101101000110101_0010000110110111"; -- -0.14762677456467807
	pesos_i(1977) := b"0000000000000000_0000000000000000_0001011001011001_1001101000110110"; -- 0.08730472388012037
	pesos_i(1978) := b"0000000000000000_0000000000000000_0010110010001000_0100011001001110"; -- 0.17395438571719724
	pesos_i(1979) := b"1111111111111111_1111111111111111_1111010100011000_1101001100111110"; -- -0.04258994814898526
	pesos_i(1980) := b"0000000000000000_0000000000000000_0001000011111001_1011101111101010"; -- 0.06631063914388215
	pesos_i(1981) := b"0000000000000000_0000000000000000_0000010010001101_1111010000111001"; -- 0.017791046025947856
	pesos_i(1982) := b"1111111111111111_1111111111111111_1100101011010110_0100010010111100"; -- -0.2076680223284642
	pesos_i(1983) := b"0000000000000000_0000000000000000_0001110000110001_0100100001100001"; -- 0.11012699485151076
	pesos_i(1984) := b"1111111111111111_1111111111111111_1101000111000111_1100110001001110"; -- -0.18054507352610438
	pesos_i(1985) := b"0000000000000000_0000000000000000_0000101011110001_1011010100011010"; -- 0.04275066265070474
	pesos_i(1986) := b"0000000000000000_0000000000000000_0001000010000010_1101110011001000"; -- 0.06449680217244202
	pesos_i(1987) := b"0000000000000000_0000000000000000_0000100110100100_1111010110011001"; -- 0.03767333006916857
	pesos_i(1988) := b"0000000000000000_0000000000000000_0010010010001011_1010000001010010"; -- 0.14275552745798017
	pesos_i(1989) := b"1111111111111111_1111111111111111_1101110000100110_1100100111000100"; -- -0.14003313986640728
	pesos_i(1990) := b"1111111111111111_1111111111111111_1110111110001010_1001010111101001"; -- -0.06429160168090836
	pesos_i(1991) := b"1111111111111111_1111111111111111_1110011010111110_0101000000101111"; -- -0.0986585506696355
	pesos_i(1992) := b"0000000000000000_0000000000000000_0010010100101111_0101011000111110"; -- 0.1452535534574473
	pesos_i(1993) := b"1111111111111111_1111111111111111_1101100100001001_1010011011010000"; -- -0.15219647813610046
	pesos_i(1994) := b"1111111111111111_1111111111111111_1110000110011110_1001001101111011"; -- -0.11867407075653132
	pesos_i(1995) := b"1111111111111111_1111111111111111_1110110100000101_0100000111011101"; -- -0.0741385303501794
	pesos_i(1996) := b"1111111111111111_1111111111111111_1101100001001001_1110000001010001"; -- -0.15512273815149624
	pesos_i(1997) := b"1111111111111111_1111111111111111_1111101101100101_0000001101100100"; -- -0.017989910210061577
	pesos_i(1998) := b"0000000000000000_0000000000000000_0001101101100110_1001111101000110"; -- 0.10703463983732298
	pesos_i(1999) := b"0000000000000000_0000000000000000_0010101001110101_0101100011111011"; -- 0.1658530819108115
	pesos_i(2000) := b"0000000000000000_0000000000000000_0001001001011111_1100101110111011"; -- 0.07177422819100525
	pesos_i(2001) := b"0000000000000000_0000000000000000_0001000010001110_0101010001001011"; -- 0.06467177229338263
	pesos_i(2002) := b"0000000000000000_0000000000000000_0001000001000111_1111110000011010"; -- 0.0635984005397873
	pesos_i(2003) := b"1111111111111111_1111111111111111_1110110000010010_0100010010010001"; -- -0.07784625485985519
	pesos_i(2004) := b"1111111111111111_1111111111111111_1110000101000000_1011110101010111"; -- -0.12010590195478965
	pesos_i(2005) := b"1111111111111111_1111111111111111_1110100101111100_0111000100001110"; -- -0.08794492146938959
	pesos_i(2006) := b"1111111111111111_1111111111111111_1111000111001010_1000101001010101"; -- -0.055503229453281025
	pesos_i(2007) := b"1111111111111111_1111111111111111_1110010101101100_0010110111001011"; -- -0.10381807134975378
	pesos_i(2008) := b"1111111111111111_1111111111111111_1101111001100010_0010000001101110"; -- -0.13131520574359848
	pesos_i(2009) := b"0000000000000000_0000000000000000_0000010110010001_1011011011111001"; -- 0.02175468044500288
	pesos_i(2010) := b"0000000000000000_0000000000000000_0001011001111001_1100110100000111"; -- 0.08779603409808547
	pesos_i(2011) := b"1111111111111111_1111111111111111_1111101000101101_0101110011010111"; -- -0.022745320770278105
	pesos_i(2012) := b"1111111111111111_1111111111111111_1101100111001110_1000011011001111"; -- -0.14919240423804198
	pesos_i(2013) := b"1111111111111111_1111111111111111_1111111000001111_1101100010001101"; -- -0.007570710816069163
	pesos_i(2014) := b"1111111111111111_1111111111111111_1110111011111111_0010111010011000"; -- -0.06641873169827024
	pesos_i(2015) := b"0000000000000000_0000000000000000_0010011001110000_0001011001011000"; -- 0.15014781617615947
	pesos_i(2016) := b"1111111111111111_1111111111111111_1110000010011000_0011110101100000"; -- -0.12267700584019917
	pesos_i(2017) := b"0000000000000000_0000000000000000_0001000110000010_1111101001010001"; -- 0.0684048126307168
	pesos_i(2018) := b"0000000000000000_0000000000000000_0001010100001111_1101011000000110"; -- 0.08227288861619843
	pesos_i(2019) := b"1111111111111111_1111111111111111_1101111000101111_0001101101000100"; -- -0.13209371180572207
	pesos_i(2020) := b"0000000000000000_0000000000000000_0011001111101000_0001110011000101"; -- 0.2027605038388044
	pesos_i(2021) := b"0000000000000000_0000000000000000_0000111111000000_1110010010010000"; -- 0.061537060832752746
	pesos_i(2022) := b"0000000000000000_0000000000000000_0010011010010110_1000111001100100"; -- 0.15073480557657776
	pesos_i(2023) := b"1111111111111111_1111111111111111_1111010001101110_1000011100100100"; -- -0.04518847817910607
	pesos_i(2024) := b"1111111111111111_1111111111111111_1110111011011101_0111111100011001"; -- -0.06693273211680521
	pesos_i(2025) := b"1111111111111111_1111111111111111_1100101101100011_0000000111111010"; -- -0.20552051199339966
	pesos_i(2026) := b"0000000000000000_0000000000000000_0000110011011001_1100101110000111"; -- 0.05019828849129658
	pesos_i(2027) := b"1111111111111111_1111111111111111_1110111001100001_0101000001101100"; -- -0.06882760384023084
	pesos_i(2028) := b"1111111111111111_1111111111111111_1111111110110011_1110101000101000"; -- -0.001160969991262472
	pesos_i(2029) := b"1111111111111111_1111111111111111_1100111001001010_1101111111001001"; -- -0.1941700108908181
	pesos_i(2030) := b"0000000000000000_0000000000000000_0000101110101001_0001001001001001"; -- 0.04554857518963537
	pesos_i(2031) := b"1111111111111111_1111111111111111_1101000000010010_0011100000001010"; -- -0.18722200150564944
	pesos_i(2032) := b"1111111111111111_1111111111111111_1110111101001110_0000100101111011"; -- -0.06521549926919339
	pesos_i(2033) := b"0000000000000000_0000000000000000_0001110101001011_1111000011001101"; -- 0.11444001202468948
	pesos_i(2034) := b"0000000000000000_0000000000000000_0000010011001100_1111100001110010"; -- 0.018752601505073435
	pesos_i(2035) := b"1111111111111111_1111111111111111_1101111110000000_1000001010010010"; -- -0.12694534235190744
	pesos_i(2036) := b"0000000000000000_0000000000000000_0010011101100101_1111111001010010"; -- 0.15390004648331684
	pesos_i(2037) := b"0000000000000000_0000000000000000_0000111110010000_0101110111001011"; -- 0.060796606150015274
	pesos_i(2038) := b"0000000000000000_0000000000000000_0011001111101000_0110110010101101"; -- 0.20276526653915494
	pesos_i(2039) := b"0000000000000000_0000000000000000_0001100100011111_1100010000111001"; -- 0.09814096817109219
	pesos_i(2040) := b"0000000000000000_0000000000000000_0010010110011001_0111111001001100"; -- 0.14687337260261357
	pesos_i(2041) := b"1111111111111111_1111111111111111_1111000000110110_1011001100111101"; -- -0.06166534190823984
	pesos_i(2042) := b"1111111111111111_1111111111111111_1110101010010101_0000100000110111"; -- -0.08366345084849407
	pesos_i(2043) := b"0000000000000000_0000000000000000_0010100110010001_0101000010001101"; -- 0.1623735755582357
	pesos_i(2044) := b"1111111111111111_1111111111111111_1110001001101000_1000001100001111"; -- -0.11559277430032082
	pesos_i(2045) := b"0000000000000000_0000000000000000_0000000010110010_0001000001100011"; -- 0.0027170410696079673
	pesos_i(2046) := b"0000000000000000_0000000000000000_0001010001101001_1010101010101000"; -- 0.07973734478401709
	pesos_i(2047) := b"0000000000000000_0000000000000000_0000111000101000_1111010000101010"; -- 0.0553124047756968
	pesos_i(2048) := b"0000000000000000_0000000000000000_0001111011100001_1010011000001000"; -- 0.12063062387639673
	pesos_i(2049) := b"0000000000000000_0000000000000000_0001110001111000_0011101111110111"; -- 0.1112096288074207
	pesos_i(2050) := b"1111111111111111_1111111111111111_1101001110110010_0110101110001111"; -- -0.17305877447704754
	pesos_i(2051) := b"0000000000000000_0000000000000000_0010011000001001_0011101011111010"; -- 0.1485783442746316
	pesos_i(2052) := b"0000000000000000_0000000000000000_0001010011000101_1110111101001100"; -- 0.0811452447148435
	pesos_i(2053) := b"0000000000000000_0000000000000000_0000101101000100_1001010000110000"; -- 0.04401518035915278
	pesos_i(2054) := b"0000000000000000_0000000000000000_0011000110001001_1110110110101100"; -- 0.19351087036017228
	pesos_i(2055) := b"1111111111111111_1111111111111111_1111100001011110_1100010010101110"; -- -0.02980395070749284
	pesos_i(2056) := b"0000000000000000_0000000000000000_0011010000110001_1111110101101101"; -- 0.20388778604201374
	pesos_i(2057) := b"0000000000000000_0000000000000000_0000010001011101_0010000110001001"; -- 0.017046066133533377
	pesos_i(2058) := b"1111111111111111_1111111111111111_1101000100111111_0101001110010010"; -- -0.18262746512990916
	pesos_i(2059) := b"0000000000000000_0000000000000000_0001010010001100_0110010011010111"; -- 0.08026724105585005
	pesos_i(2060) := b"0000000000000000_0000000000000000_0000110010101111_0011110001111111"; -- 0.04954889397746673
	pesos_i(2061) := b"0000000000000000_0000000000000000_0000000111101111_0101101001101000"; -- 0.007558489114594062
	pesos_i(2062) := b"1111111111111111_1111111111111111_1111001000000111_1100000001000010"; -- -0.05456922895200046
	pesos_i(2063) := b"0000000000000000_0000000000000000_0001100000011111_1101000010110011"; -- 0.09423546193762766
	pesos_i(2064) := b"1111111111111111_1111111111111111_1100111101011110_0101010100011111"; -- -0.18996685025811674
	pesos_i(2065) := b"1111111111111111_1111111111111111_1110000111010001_0010101110110111"; -- -0.1179020574472229
	pesos_i(2066) := b"0000000000000000_0000000000000000_0001011001110010_1000110101111110"; -- 0.08768543566079769
	pesos_i(2067) := b"0000000000000000_0000000000000000_0001100101110001_1011110110101011"; -- 0.09939179815138743
	pesos_i(2068) := b"0000000000000000_0000000000000000_0001101010101110_0011111001101011"; -- 0.10422124967330852
	pesos_i(2069) := b"1111111111111111_1111111111111111_1110111000011010_1000001100100011"; -- -0.06990795517510931
	pesos_i(2070) := b"1111111111111111_1111111111111111_1111100010111011_1010111000100000"; -- -0.028386227810139848
	pesos_i(2071) := b"1111111111111111_1111111111111111_1111100000111010_1011110010100110"; -- -0.030353745980570432
	pesos_i(2072) := b"1111111111111111_1111111111111111_1110011001110011_0011011111010110"; -- -0.09980441109236428
	pesos_i(2073) := b"0000000000000000_0000000000000000_0001100000000110_0110000101001101"; -- 0.0938473522304579
	pesos_i(2074) := b"1111111111111111_1111111111111111_1110110010110100_0111011111111010"; -- -0.07537126672166293
	pesos_i(2075) := b"0000000000000000_0000000000000000_0001100000001001_0000110001100001"; -- 0.09388806700424096
	pesos_i(2076) := b"0000000000000000_0000000000000000_0000110000001101_1011011111101110"; -- 0.04708432727957177
	pesos_i(2077) := b"0000000000000000_0000000000000000_0000010000111000_1111000010011110"; -- 0.016493834057875956
	pesos_i(2078) := b"0000000000000000_0000000000000000_0000110111010110_1010001100001101"; -- 0.054056349338792054
	pesos_i(2079) := b"0000000000000000_0000000000000000_0000010011101101_0100011010001100"; -- 0.019245538045172653
	pesos_i(2080) := b"1111111111111111_1111111111111111_1101101001100101_1111100110100011"; -- -0.14688148272592502
	pesos_i(2081) := b"1111111111111111_1111111111111111_1110111101111110_0001010110110001"; -- -0.06448234972773599
	pesos_i(2082) := b"1111111111111111_1111111111111111_1111100110011010_0110001000001111"; -- -0.02498805180110867
	pesos_i(2083) := b"1111111111111111_1111111111111111_1110101000010011_1001001011010011"; -- -0.08563883167563421
	pesos_i(2084) := b"0000000000000000_0000000000000000_0001011001111010_1101011001001110"; -- 0.0878118459079236
	pesos_i(2085) := b"0000000000000000_0000000000000000_0010010011100100_0111011010110101"; -- 0.14411107941251552
	pesos_i(2086) := b"1111111111111111_1111111111111111_1101011010010101_0111101100011001"; -- -0.16178160326629532
	pesos_i(2087) := b"1111111111111111_1111111111111111_1110010010010010_1010101110111101"; -- -0.10713698034034586
	pesos_i(2088) := b"1111111111111111_1111111111111111_1111100011011000_0110010011011011"; -- -0.027948090095624645
	pesos_i(2089) := b"0000000000000000_0000000000000000_0000100110011001_1011110001111000"; -- 0.037502078250031566
	pesos_i(2090) := b"0000000000000000_0000000000000000_0001000011001000_0111010111111111"; -- 0.06555879083572405
	pesos_i(2091) := b"0000000000000000_0000000000000000_0000100111001001_0011010110111010"; -- 0.038226468859287814
	pesos_i(2092) := b"1111111111111111_1111111111111111_1111011000001010_1101010011101101"; -- -0.03889722067414216
	pesos_i(2093) := b"0000000000000000_0000000000000000_0011011100010101_1000010010011010"; -- 0.2151720881914884
	pesos_i(2094) := b"1111111111111111_1111111111111111_1101111011001001_0100110110011111"; -- -0.12974085676410613
	pesos_i(2095) := b"1111111111111111_1111111111111111_1110001111011110_0010010111000000"; -- -0.10989154871444895
	pesos_i(2096) := b"0000000000000000_0000000000000000_0010001111100101_0000101001101110"; -- 0.14021363441300538
	pesos_i(2097) := b"1111111111111111_1111111111111111_1101110011101011_1110001101110010"; -- -0.13702562782854927
	pesos_i(2098) := b"0000000000000000_0000000000000000_0001111100100010_0010001001010010"; -- 0.12161459441635539
	pesos_i(2099) := b"0000000000000000_0000000000000000_0010100101000100_1100010011100011"; -- 0.16120558295019438
	pesos_i(2100) := b"0000000000000000_0000000000000000_0001101001101110_0100100111101011"; -- 0.1032453727663412
	pesos_i(2101) := b"0000000000000000_0000000000000000_0001000110010110_0001011010010110"; -- 0.06869641448333486
	pesos_i(2102) := b"0000000000000000_0000000000000000_0001100100110000_1101101010001111"; -- 0.09840169899813743
	pesos_i(2103) := b"0000000000000000_0000000000000000_0000101101100110_0010000000011111"; -- 0.044527061102962846
	pesos_i(2104) := b"1111111111111111_1111111111111111_1101111110000011_0110100100110101"; -- -0.12690107776139975
	pesos_i(2105) := b"0000000000000000_0000000000000000_0001111011100011_1011110000011110"; -- 0.1206624576878156
	pesos_i(2106) := b"0000000000000000_0000000000000000_0010101110101111_0110101111001000"; -- 0.17064546239533743
	pesos_i(2107) := b"0000000000000000_0000000000000000_0010110110011101_0011010001000110"; -- 0.17817999571350207
	pesos_i(2108) := b"0000000000000000_0000000000000000_0001011111101011_0110011111010011"; -- 0.09343575390461344
	pesos_i(2109) := b"1111111111111111_1111111111111111_1110100000111000_0000111001100100"; -- -0.09289465002886846
	pesos_i(2110) := b"1111111111111111_1111111111111111_1111111011101110_1111000001001111"; -- -0.004166584798075866
	pesos_i(2111) := b"1111111111111111_1111111111111111_1101010000011000_1000101000111001"; -- -0.17150055041092702
	pesos_i(2112) := b"1111111111111111_1111111111111111_1101101000010111_1110111001011000"; -- -0.14807234145724857
	pesos_i(2113) := b"0000000000000000_0000000000000000_0000110001000011_1001111001100100"; -- 0.04790677962880189
	pesos_i(2114) := b"1111111111111111_1111111111111111_1111010000110101_1100010000101111"; -- -0.04605459061578621
	pesos_i(2115) := b"0000000000000000_0000000000000000_0000011111111111_1110010110100011"; -- 0.03124842858902223
	pesos_i(2116) := b"0000000000000000_0000000000000000_0010111101110110_1111100011011011"; -- 0.185409120052775
	pesos_i(2117) := b"0000000000000000_0000000000000000_0000101000011100_1011001010000010"; -- 0.03950038606654598
	pesos_i(2118) := b"0000000000000000_0000000000000000_0000110001011001_0000111000010101"; -- 0.04823387158972951
	pesos_i(2119) := b"0000000000000000_0000000000000000_0000110010110000_1111011000001011"; -- 0.04957521220041022
	pesos_i(2120) := b"1111111111111111_1111111111111111_1111100110000111_1100111110011000"; -- -0.02527143985239445
	pesos_i(2121) := b"1111111111111111_1111111111111111_1110010011011101_0110000111100111"; -- -0.10599697223430672
	pesos_i(2122) := b"0000000000000000_0000000000000000_0000000000000001_0100001111101101"; -- 1.9307474859925344e-05
	pesos_i(2123) := b"1111111111111111_1111111111111111_1100110011001101_0001100000001111"; -- -0.19999551420045097
	pesos_i(2124) := b"1111111111111111_1111111111111111_1110011100100101_0010011010100011"; -- -0.09708937194207302
	pesos_i(2125) := b"1111111111111111_1111111111111111_1100101000101101_1000110110001101"; -- -0.2102424174762178
	pesos_i(2126) := b"0000000000000000_0000000000000000_0010111111110111_0100111111101010"; -- 0.18736743410215917
	pesos_i(2127) := b"1111111111111111_1111111111111111_1111010110100100_1111111110111001"; -- -0.04045106628402731
	pesos_i(2128) := b"1111111111111111_1111111111111111_1101011101011000_1101000100111110"; -- -0.15880100486164103
	pesos_i(2129) := b"0000000000000000_0000000000000000_0000011110111000_0011000011111110"; -- 0.030154287380658007
	pesos_i(2130) := b"1111111111111111_1111111111111111_1110000001110000_0101111110100101"; -- -0.1232853147787749
	pesos_i(2131) := b"0000000000000000_0000000000000000_0000001101010100_1110010001010111"; -- 0.01301409849777557
	pesos_i(2132) := b"0000000000000000_0000000000000000_0001010000011111_1011001101110101"; -- 0.07860871904835816
	pesos_i(2133) := b"1111111111111111_1111111111111111_1110100100101111_0100110111011001"; -- -0.08912194673501392
	pesos_i(2134) := b"1111111111111111_1111111111111111_1100110000110010_1001011001100000"; -- -0.20235309738543988
	pesos_i(2135) := b"0000000000000000_0000000000000000_0001000111100110_1100010001011100"; -- 0.06992747537327787
	pesos_i(2136) := b"0000000000000000_0000000000000000_0010001011010111_0100110010100010"; -- 0.1360977073894193
	pesos_i(2137) := b"1111111111111111_1111111111111111_1111010100110000_1110011011100010"; -- -0.042222566469060266
	pesos_i(2138) := b"1111111111111111_1111111111111111_1101100010111100_0010101001010100"; -- -0.15337882477285492
	pesos_i(2139) := b"0000000000000000_0000000000000000_0010001111110001_0110011000011000"; -- 0.14040220338819384
	pesos_i(2140) := b"1111111111111111_1111111111111111_1101100011101001_1011100100000000"; -- -0.1526836753914998
	pesos_i(2141) := b"1111111111111111_1111111111111111_1110101010101100_0001010101001011"; -- -0.08331171918202944
	pesos_i(2142) := b"1111111111111111_1111111111111111_1101001101101000_1101000111111000"; -- -0.1741818207942314
	pesos_i(2143) := b"1111111111111111_1111111111111111_1101100011100010_0101100011011110"; -- -0.15279621688187117
	pesos_i(2144) := b"1111111111111111_1111111111111111_1110100110000011_0100010111101111"; -- -0.08784068023031157
	pesos_i(2145) := b"1111111111111111_1111111111111111_1101001001111101_1001010100101011"; -- -0.17777126037827945
	pesos_i(2146) := b"0000000000000000_0000000000000000_0010100100001101_0000110101110001"; -- 0.16035541533185463
	pesos_i(2147) := b"0000000000000000_0000000000000000_0010001101110000_1011010001001101"; -- 0.13843848102980816
	pesos_i(2148) := b"0000000000000000_0000000000000000_0001011110111001_0101011010010001"; -- 0.09267178579031737
	pesos_i(2149) := b"0000000000000000_0000000000000000_0010100011011001_0101101011001100"; -- 0.15956656922373322
	pesos_i(2150) := b"0000000000000000_0000000000000000_0001000100010100_1001000011100110"; -- 0.06672006232489043
	pesos_i(2151) := b"1111111111111111_1111111111111111_1111000111010010_1100111011000111"; -- -0.05537707940358525
	pesos_i(2152) := b"0000000000000000_0000000000000000_0000010011011111_1001010100010111"; -- 0.019036596482742304
	pesos_i(2153) := b"1111111111111111_1111111111111111_1111110100111100_0001001111111111"; -- -0.01080203072227769
	pesos_i(2154) := b"0000000000000000_0000000000000000_0001000100110000_1010100000000100"; -- 0.06714868627967671
	pesos_i(2155) := b"1111111111111111_1111111111111111_1111010001111100_0111101000000010"; -- -0.04497563782527209
	pesos_i(2156) := b"0000000000000000_0000000000000000_0001000010111100_1000110000010101"; -- 0.06537700199377977
	pesos_i(2157) := b"1111111111111111_1111111111111111_1110001010110011_0110000011001010"; -- -0.11445040759652936
	pesos_i(2158) := b"0000000000000000_0000000000000000_0000101000011110_0001101111101011"; -- 0.0395219276681876
	pesos_i(2159) := b"1111111111111111_1111111111111111_1110010000011000_0011011001111011"; -- -0.10900554177051566
	pesos_i(2160) := b"1111111111111111_1111111111111111_1110110010011010_1101011101110101"; -- -0.07576230418182678
	pesos_i(2161) := b"1111111111111111_1111111111111111_1101111010011001_0110001001010000"; -- -0.13047204533130427
	pesos_i(2162) := b"0000000000000000_0000000000000000_0000011011001010_0010111100010100"; -- 0.026522581542055734
	pesos_i(2163) := b"0000000000000000_0000000000000000_0000010001100010_1100101011111101"; -- 0.017132460447526754
	pesos_i(2164) := b"1111111111111111_1111111111111111_1101010101001100_0110010010110110"; -- -0.16680307917790482
	pesos_i(2165) := b"0000000000000000_0000000000000000_0000010111100001_1001011101100010"; -- 0.022973500765027032
	pesos_i(2166) := b"1111111111111111_1111111111111111_1110111010101101_1011010011110010"; -- -0.06766194430961073
	pesos_i(2167) := b"1111111111111111_1111111111111111_1111101001110101_1000111010101110"; -- -0.021643717210707944
	pesos_i(2168) := b"0000000000000000_0000000000000000_0001001100000100_1000101010111111"; -- 0.0742880551688372
	pesos_i(2169) := b"1111111111111111_1111111111111111_1110011010001111_0000001001011001"; -- -0.09938035313889519
	pesos_i(2170) := b"1111111111111111_1111111111111111_1110010110010100_1111010101111011"; -- -0.10319581752011613
	pesos_i(2171) := b"1111111111111111_1111111111111111_1101100001100011_0111110000011111"; -- -0.15473198159389503
	pesos_i(2172) := b"1111111111111111_1111111111111111_1111100000000010_1011110101110100"; -- -0.031208190066768886
	pesos_i(2173) := b"0000000000000000_0000000000000000_0001010100010001_1111110100011110"; -- 0.08230573641571493
	pesos_i(2174) := b"1111111111111111_1111111111111111_1101010001001010_1101100110000010"; -- -0.17073288515978835
	pesos_i(2175) := b"0000000000000000_0000000000000000_0001111011111100_1010000101000010"; -- 0.12104232654481532
	pesos_i(2176) := b"1111111111111111_1111111111111111_1110011010111111_1101101100011110"; -- -0.09863501096598096
	pesos_i(2177) := b"1111111111111111_1111111111111111_1111001110001011_1011001101011011"; -- -0.048649587794153626
	pesos_i(2178) := b"0000000000000000_0000000000000000_0001001001010000_0001101001011000"; -- 0.07153477332066988
	pesos_i(2179) := b"0000000000000000_0000000000000000_0000000100110110_1000101100000000"; -- 0.004738509613852652
	pesos_i(2180) := b"0000000000000000_0000000000000000_0000001000001111_0110000011110001"; -- 0.008047160051531974
	pesos_i(2181) := b"0000000000000000_0000000000000000_0000100001010011_1101011111001001"; -- 0.032529341274301245
	pesos_i(2182) := b"1111111111111111_1111111111111111_1110100010011100_0101000101111110"; -- -0.09136477155714719
	pesos_i(2183) := b"1111111111111111_1111111111111111_1111011001011100_1011010011111001"; -- -0.03764790460294963
	pesos_i(2184) := b"0000000000000000_0000000000000000_0010110111011010_1010100000101110"; -- 0.17911769024615531
	pesos_i(2185) := b"1111111111111111_1111111111111111_1101010100001001_0000101101000001"; -- -0.16783075016645269
	pesos_i(2186) := b"0000000000000000_0000000000000000_0000100100111000_0111111011101001"; -- 0.036018306685602124
	pesos_i(2187) := b"0000000000000000_0000000000000000_0001000001010111_1000001101001110"; -- 0.06383534096251511
	pesos_i(2188) := b"1111111111111111_1111111111111111_1110111101010110_0100110001111010"; -- -0.06508943572302975
	pesos_i(2189) := b"1111111111111111_1111111111111111_1110100000101100_0101101001111000"; -- -0.09307322090943425
	pesos_i(2190) := b"1111111111111111_1111111111111111_1110011110000010_1011110101001001"; -- -0.09566132508041014
	pesos_i(2191) := b"0000000000000000_0000000000000000_0000110010110110_0111011100101110"; -- 0.04965920334546131
	pesos_i(2192) := b"0000000000000000_0000000000000000_0000100010011101_0101001111011111"; -- 0.03365062888751528
	pesos_i(2193) := b"0000000000000000_0000000000000000_0001100000011010_0011111000001010"; -- 0.09415042640507522
	pesos_i(2194) := b"1111111111111111_1111111111111111_1110000000101001_1000110011100101"; -- -0.12436599156487121
	pesos_i(2195) := b"0000000000000000_0000000000000000_0010101111111100_1001100100100111"; -- 0.17182309354166148
	pesos_i(2196) := b"0000000000000000_0000000000000000_0010101100111111_0110001010011110"; -- 0.16893593170143184
	pesos_i(2197) := b"1111111111111111_1111111111111111_1101101110011011_0011100011101111"; -- -0.142162744170324
	pesos_i(2198) := b"0000000000000000_0000000000000000_0000000001011011_0011101111011111"; -- 0.001392118316431925
	pesos_i(2199) := b"0000000000000000_0000000000000000_0000100001000011_0001011001100111"; -- 0.03227367417486151
	pesos_i(2200) := b"1111111111111111_1111111111111111_1101000011011110_1000100011001110"; -- -0.1841043947101924
	pesos_i(2201) := b"1111111111111111_1111111111111111_1110001110101101_1111100000110101"; -- -0.1106266852024806
	pesos_i(2202) := b"0000000000000000_0000000000000000_0010011000111001_0101000001000110"; -- 0.1493120357028314
	pesos_i(2203) := b"0000000000000000_0000000000000000_0000110010001111_0000111101101100"; -- 0.04905792600395245
	pesos_i(2204) := b"0000000000000000_0000000000000000_0001110101101111_0010010000111111"; -- 0.11497713613384151
	pesos_i(2205) := b"0000000000000000_0000000000000000_0000100010010010_0110000101111100"; -- 0.033483593722265066
	pesos_i(2206) := b"0000000000000000_0000000000000000_0001011011110001_0111000111001011"; -- 0.08962165078419974
	pesos_i(2207) := b"0000000000000000_0000000000000000_0011001000100000_0001111011010111"; -- 0.19580261936949625
	pesos_i(2208) := b"0000000000000000_0000000000000000_0010100000101010_1011101001100010"; -- 0.15690197839084527
	pesos_i(2209) := b"1111111111111111_1111111111111111_1101010111001000_0111000001111011"; -- -0.16491028792508305
	pesos_i(2210) := b"0000000000000000_0000000000000000_0000011001001100_0001000011101000"; -- 0.0245981756267581
	pesos_i(2211) := b"1111111111111111_1111111111111111_1111110011100100_0100011000001010"; -- -0.012141821539364744
	pesos_i(2212) := b"1111111111111111_1111111111111111_1111010101101110_1110000000111010"; -- -0.04127691832265634
	pesos_i(2213) := b"1111111111111111_1111111111111111_1110101011001010_1100101100011100"; -- -0.0828431183783923
	pesos_i(2214) := b"1111111111111111_1111111111111111_1100111010111110_1011001001110110"; -- -0.19240269292589304
	pesos_i(2215) := b"1111111111111111_1111111111111111_1111010001001100_0111001000111001"; -- -0.045708523827427884
	pesos_i(2216) := b"0000000000000000_0000000000000000_0011000110110000_1101101101000010"; -- 0.19410486559477846
	pesos_i(2217) := b"1111111111111111_1111111111111111_1110111101010010_0111001011011011"; -- -0.06514818343869763
	pesos_i(2218) := b"0000000000000000_0000000000000000_0010000001000010_0101000011100101"; -- 0.1260119016750551
	pesos_i(2219) := b"0000000000000000_0000000000000000_0010100100110000_0110011110101011"; -- 0.1608948509066411
	pesos_i(2220) := b"1111111111111111_1111111111111111_1110111110110011_0110101101111000"; -- -0.06366852109351218
	pesos_i(2221) := b"0000000000000000_0000000000000000_0010011111110110_1001111001000100"; -- 0.1561068453990811
	pesos_i(2222) := b"1111111111111111_1111111111111111_1101101100001010_0010101100000101"; -- -0.14437609796320322
	pesos_i(2223) := b"0000000000000000_0000000000000000_0000100000011010_0000100001010010"; -- 0.031647224557577826
	pesos_i(2224) := b"1111111111111111_1111111111111111_1111100011011001_0000111001100111"; -- -0.027937984412059427
	pesos_i(2225) := b"1111111111111111_1111111111111111_1101110011111011_1100000001110110"; -- -0.1367835722909083
	pesos_i(2226) := b"0000000000000000_0000000000000000_0000110111000110_1010000011011011"; -- 0.05381207805545728
	pesos_i(2227) := b"1111111111111111_1111111111111111_1111000111000011_1001010011110010"; -- -0.05560940823968439
	pesos_i(2228) := b"1111111111111111_1111111111111111_1100111010100111_1100101001010110"; -- -0.19275222201614264
	pesos_i(2229) := b"1111111111111111_1111111111111111_1111101100001101_1100111110011100"; -- -0.019320511349187254
	pesos_i(2230) := b"1111111111111111_1111111111111111_1100111101110110_0100001100001101"; -- -0.18960171623673244
	pesos_i(2231) := b"0000000000000000_0000000000000000_0001100100001000_1100011001011010"; -- 0.09779014289421781
	pesos_i(2232) := b"0000000000000000_0000000000000000_0000100100000110_1010001100101010"; -- 0.035257528043378256
	pesos_i(2233) := b"1111111111111111_1111111111111111_1101101001110001_1100101110111011"; -- -0.14670111359412089
	pesos_i(2234) := b"0000000000000000_0000000000000000_0000101110001101_1001010011110111"; -- 0.045129118297905196
	pesos_i(2235) := b"0000000000000000_0000000000000000_0010011000001010_0010100010100100"; -- 0.1485925102763175
	pesos_i(2236) := b"0000000000000000_0000000000000000_0001001011100010_0100010100101101"; -- 0.07376510949929695
	pesos_i(2237) := b"1111111111111111_1111111111111111_1110101100011110_0001100001101101"; -- -0.08157203035908359
	pesos_i(2238) := b"1111111111111111_1111111111111111_1111100000010011_0000001001000010"; -- -0.03095994851710438
	pesos_i(2239) := b"0000000000000000_0000000000000000_0000001100011000_0010010111011010"; -- 0.012087217065024948
	pesos_i(2240) := b"1111111111111111_1111111111111111_1101101011100010_1010001010110100"; -- -0.1449793158550018
	pesos_i(2241) := b"1111111111111111_1111111111111111_1111100100000100_0101010000111001"; -- -0.02727769468746882
	pesos_i(2242) := b"0000000000000000_0000000000000000_0001101110110100_1100111101011101"; -- 0.10822769194468285
	pesos_i(2243) := b"0000000000000000_0000000000000000_0000101010100100_0001111100110110"; -- 0.041566801740766365
	pesos_i(2244) := b"1111111111111111_1111111111111111_1110101101000111_0011110110110101"; -- -0.0809441979676278
	pesos_i(2245) := b"0000000000000000_0000000000000000_0010100011100001_0101001110001101"; -- 0.15968820753655116
	pesos_i(2246) := b"0000000000000000_0000000000000000_0001100110001110_1000001000011010"; -- 0.09983075268020679
	pesos_i(2247) := b"0000000000000000_0000000000000000_0000010111001001_1001100011100011"; -- 0.022607379255511924
	pesos_i(2248) := b"1111111111111111_1111111111111111_1110010101101010_1100001111001001"; -- -0.10383964854763256
	pesos_i(2249) := b"1111111111111111_1111111111111111_1111101110011001_1011000011011010"; -- -0.01718611399979856
	pesos_i(2250) := b"1111111111111111_1111111111111111_1110010110110011_0010101010000111"; -- -0.10273489196545918
	pesos_i(2251) := b"0000000000000000_0000000000000000_0000010111000000_1001111101001111"; -- 0.022470433141760462
	pesos_i(2252) := b"0000000000000000_0000000000000000_0010000110000001_0110010110110001"; -- 0.1308806950763628
	pesos_i(2253) := b"1111111111111111_1111111111111111_1110100001010000_0111101011000010"; -- -0.0925219799726214
	pesos_i(2254) := b"1111111111111111_1111111111111111_1111011011001011_0100010001101101"; -- -0.03596088739578942
	pesos_i(2255) := b"1111111111111111_1111111111111111_1111101010100101_0010101100000101"; -- -0.02091723569533303
	pesos_i(2256) := b"1111111111111111_1111111111111111_1111001010001000_1011100001001111"; -- -0.05260131910203014
	pesos_i(2257) := b"0000000000000000_0000000000000000_0000001010111110_0000001101011000"; -- 0.010711869335971671
	pesos_i(2258) := b"1111111111111111_1111111111111111_1100111101000100_1000000010000101"; -- -0.19036099203472415
	pesos_i(2259) := b"0000000000000000_0000000000000000_0000111000101110_0000110000101011"; -- 0.055390129621293305
	pesos_i(2260) := b"1111111111111111_1111111111111111_1110001101001100_0001011001111011"; -- -0.1121202420456952
	pesos_i(2261) := b"0000000000000000_0000000000000000_0000010111001111_1000100110010111"; -- 0.022698020383840733
	pesos_i(2262) := b"1111111111111111_1111111111111111_1101011010000110_1110100001100000"; -- -0.1620039716957516
	pesos_i(2263) := b"0000000000000000_0000000000000000_0001100000110001_0101011001110011"; -- 0.09450283335589103
	pesos_i(2264) := b"1111111111111111_1111111111111111_1101111111000011_1110111011111000"; -- -0.12591654241188988
	pesos_i(2265) := b"1111111111111111_1111111111111111_1111011000000000_0110011100010101"; -- -0.039056355838664784
	pesos_i(2266) := b"1111111111111111_1111111111111111_1110000111100001_1101101010011111"; -- -0.11764749154630644
	pesos_i(2267) := b"1111111111111111_1111111111111111_1110110011011111_0000111100100011"; -- -0.07472138786147767
	pesos_i(2268) := b"0000000000000000_0000000000000000_0001110101000111_0101001101010010"; -- 0.11436959037247028
	pesos_i(2269) := b"0000000000000000_0000000000000000_0000111000010110_1001110111001110"; -- 0.05503259929007736
	pesos_i(2270) := b"1111111111111111_1111111111111111_1110010000110011_1010100111001100"; -- -0.10858668113307621
	pesos_i(2271) := b"1111111111111111_1111111111111111_1110010111101110_1110000011011011"; -- -0.10182375578017823
	pesos_i(2272) := b"1111111111111111_1111111111111111_1101100111010010_1100001101101001"; -- -0.14912775692879915
	pesos_i(2273) := b"1111111111111111_1111111111111111_1110111110111110_1010110100001011"; -- -0.06349676600786817
	pesos_i(2274) := b"0000000000000000_0000000000000000_0010010010011111_1010111010010001"; -- 0.14306155253590985
	pesos_i(2275) := b"0000000000000000_0000000000000000_0000000000110111_1000100111001001"; -- 0.0008474459250116864
	pesos_i(2276) := b"1111111111111111_1111111111111111_1110110010000010_1001110010001001"; -- -0.0761320271630738
	pesos_i(2277) := b"0000000000000000_0000000000000000_0000111011010101_1000001111111101"; -- 0.05794548927580855
	pesos_i(2278) := b"1111111111111111_1111111111111111_1110001001011010_1101011010001010"; -- -0.11580142150951625
	pesos_i(2279) := b"1111111111111111_1111111111111111_1110111001111101_0100101101001111"; -- -0.06840066258569291
	pesos_i(2280) := b"1111111111111111_1111111111111111_1101101010010000_1001100010010110"; -- -0.1462311396564232
	pesos_i(2281) := b"0000000000000000_0000000000000000_0000001000111000_0001111011110010"; -- 0.00866883675583521
	pesos_i(2282) := b"1111111111111111_1111111111111111_1110110000010010_1011110010100011"; -- -0.07783909808333093
	pesos_i(2283) := b"1111111111111111_1111111111111111_1111100011101111_1011100011011000"; -- -0.027592131800113544
	pesos_i(2284) := b"1111111111111111_1111111111111111_1110110000110111_1111001101111001"; -- -0.07727125449526578
	pesos_i(2285) := b"1111111111111111_1111111111111111_1110100011001011_1100110111100010"; -- -0.0906401942799611
	pesos_i(2286) := b"0000000000000000_0000000000000000_0001110010101110_1100111011000001"; -- 0.11204235268187875
	pesos_i(2287) := b"1111111111111111_1111111111111111_1111110100100010_0000101010100010"; -- -0.011199317318563077
	pesos_i(2288) := b"1111111111111111_1111111111111111_1110101101010010_1001100010010100"; -- -0.08077093492640822
	pesos_i(2289) := b"1111111111111111_1111111111111111_1110011001000100_0011001010111111"; -- -0.10052187771678267
	pesos_i(2290) := b"1111111111111111_1111111111111111_1111000111111001_0111011000010001"; -- -0.054787274232026256
	pesos_i(2291) := b"1111111111111111_1111111111111111_1111100100001010_0000100100111101"; -- -0.027190611394036432
	pesos_i(2292) := b"0000000000000000_0000000000000000_0010001011101000_0110001010110011"; -- 0.13635842209672858
	pesos_i(2293) := b"0000000000000000_0000000000000000_0000100110000010_1011011110010111"; -- 0.037150835299521866
	pesos_i(2294) := b"0000000000000000_0000000000000000_0001100011110010_0110110000000101"; -- 0.09744906550717736
	pesos_i(2295) := b"0000000000000000_0000000000000000_0010001010110001_0101110011101111"; -- 0.13551884483090285
	pesos_i(2296) := b"1111111111111111_1111111111111111_1110011010010110_1000100111011100"; -- -0.09926546460130593
	pesos_i(2297) := b"1111111111111111_1111111111111111_1110011110111010_1100010100000000"; -- -0.09480637301758299
	pesos_i(2298) := b"1111111111111111_1111111111111111_1111000110001001_1011101110000111"; -- -0.056492118513830014
	pesos_i(2299) := b"0000000000000000_0000000000000000_0000100100010100_0011010010111000"; -- 0.035464568024383525
	pesos_i(2300) := b"0000000000000000_0000000000000000_0001011100100100_1011010010110111"; -- 0.09040383778274341
	pesos_i(2301) := b"0000000000000000_0000000000000000_0000000110110110_1000000010111000"; -- 0.006691021925755769
	pesos_i(2302) := b"1111111111111111_1111111111111111_1111010110110011_0101101011111000"; -- -0.04023200455427022
	pesos_i(2303) := b"0000000000000000_0000000000000000_0001011001101110_1011110110001010"; -- 0.08762726413937982
	pesos_i(2304) := b"1111111111111111_1111111111111111_1110001101100010_0100100001010110"; -- -0.1117815770062623
	pesos_i(2305) := b"0000000000000000_0000000000000000_0011001111100101_0111111100101011"; -- 0.20272059245280924
	pesos_i(2306) := b"0000000000000000_0000000000000000_0001010110101110_0101101101010111"; -- 0.08469172357021681
	pesos_i(2307) := b"1111111111111111_1111111111111111_1101001010100101_1110001110011001"; -- -0.17715623385367477
	pesos_i(2308) := b"0000000000000000_0000000000000000_0001010011110011_1010000101101101"; -- 0.08184250736759943
	pesos_i(2309) := b"0000000000000000_0000000000000000_0010010101000010_0100010101000010"; -- 0.14554245815644068
	pesos_i(2310) := b"1111111111111111_1111111111111111_1101011001010001_1011011100000010"; -- -0.16281563006000052
	pesos_i(2311) := b"0000000000000000_0000000000000000_0010100001000111_1000010000100101"; -- 0.15734125052776832
	pesos_i(2312) := b"0000000000000000_0000000000000000_0000000010100000_1110011111011101"; -- 0.0024552263857918477
	pesos_i(2313) := b"1111111111111111_1111111111111111_1101010110110101_0001010111110010"; -- -0.1652056011916991
	pesos_i(2314) := b"1111111111111111_1111111111111111_1110001011110011_1111101010101000"; -- -0.11346467404034585
	pesos_i(2315) := b"0000000000000000_0000000000000000_0000011110010011_0001011010110000"; -- 0.02958814427581124
	pesos_i(2316) := b"0000000000000000_0000000000000000_0010101000111101_1011000100011000"; -- 0.16500384170000526
	pesos_i(2317) := b"1111111111111111_1111111111111111_1110101010100000_1011111110110110"; -- -0.08348466691824716
	pesos_i(2318) := b"0000000000000000_0000000000000000_0001010000011101_1100110001001011"; -- 0.07857968174893544
	pesos_i(2319) := b"0000000000000000_0000000000000000_0010001001110110_1011111010011100"; -- 0.13462439820206926
	pesos_i(2320) := b"0000000000000000_0000000000000000_0000110010011111_1111110011001100"; -- 0.0493162152775563
	pesos_i(2321) := b"1111111111111111_1111111111111111_1110001101011100_0011001111000100"; -- -0.11187435592451499
	pesos_i(2322) := b"0000000000000000_0000000000000000_0000111000111101_0110111110111111"; -- 0.05562494681262242
	pesos_i(2323) := b"0000000000000000_0000000000000000_0000011101000000_0000111110001100"; -- 0.028321239218626393
	pesos_i(2324) := b"0000000000000000_0000000000000000_0010010010110111_0000010110000101"; -- 0.14341768747950784
	pesos_i(2325) := b"0000000000000000_0000000000000000_0001011000011001_1100100000100000"; -- 0.0863308980454184
	pesos_i(2326) := b"0000000000000000_0000000000000000_0000001011010001_0010011000100111"; -- 0.011003860969858855
	pesos_i(2327) := b"1111111111111111_1111111111111111_1110111111000000_1010111111001001"; -- -0.06346608487943128
	pesos_i(2328) := b"1111111111111111_1111111111111111_1101111110110000_1110101001010001"; -- -0.126206736857939
	pesos_i(2329) := b"0000000000000000_0000000000000000_0010011001111010_1001011111101111"; -- 0.1503081281979406
	pesos_i(2330) := b"0000000000000000_0000000000000000_0000110001111100_0001000010110001"; -- 0.04876808473777529
	pesos_i(2331) := b"1111111111111111_1111111111111111_1111000110101100_0001010101101110"; -- -0.05596796099331922
	pesos_i(2332) := b"0000000000000000_0000000000000000_0001101110110111_0100000110000110"; -- 0.10826501391775513
	pesos_i(2333) := b"1111111111111111_1111111111111111_1101010111110111_1100010111100001"; -- -0.16418803456596956
	pesos_i(2334) := b"0000000000000000_0000000000000000_0101000011011110_0001001110001010"; -- 0.31588861588571815
	pesos_i(2335) := b"1111111111111111_1111111111111111_1100000100001111_1000101100111010"; -- -0.2458565696832411
	pesos_i(2336) := b"0000000000000000_0000000000000000_0000000101000101_1000111101100011"; -- 0.004967652902082336
	pesos_i(2337) := b"0000000000000000_0000000000000000_0010000011111111_0001001011101101"; -- 0.12889211936422834
	pesos_i(2338) := b"1111111111111111_1111111111111111_1111101011010000_1111100100011001"; -- -0.020248824425593115
	pesos_i(2339) := b"1111111111111111_1111111111111111_1111000001010101_0000010000000111"; -- -0.061202762805382525
	pesos_i(2340) := b"1111111111111111_1111111111111111_1111010100010101_1110110001111001"; -- -0.04263422057511246
	pesos_i(2341) := b"0000000000000000_0000000000000000_0001010011100111_1101010010100000"; -- 0.0816624537648416
	pesos_i(2342) := b"0000000000000000_0000000000000000_0001000000100000_0111011011111110"; -- 0.06299537363271379
	pesos_i(2343) := b"0000000000000000_0000000000000000_0001100111010111_0011001011001011"; -- 0.10093991714237045
	pesos_i(2344) := b"1111111111111111_1111111111111111_1111101110100100_1100000010110010"; -- -0.01701732305201629
	pesos_i(2345) := b"0000000000000000_0000000000000000_0000001011110100_1101010010001011"; -- 0.011548313114064039
	pesos_i(2346) := b"1111111111111111_1111111111111111_1111101100110011_0100000111100101"; -- -0.018749124100265895
	pesos_i(2347) := b"1111111111111111_1111111111111111_1101011000101001_1111010010100111"; -- -0.1634223072337138
	pesos_i(2348) := b"1111111111111111_1111111111111111_1101111110101101_1010110000100011"; -- -0.12625621932953168
	pesos_i(2349) := b"0000000000000000_0000000000000000_0000010010010110_1111000001100101"; -- 0.017928147049912416
	pesos_i(2350) := b"0000000000000000_0000000000000000_0001001011001111_0100011101111101"; -- 0.07347533044656211
	pesos_i(2351) := b"1111111111111111_1111111111111111_1111110111000110_1001111110100101"; -- -0.008687994165218302
	pesos_i(2352) := b"0000000000000000_0000000000000000_0001100000000101_1000000011110101"; -- 0.09383398036456156
	pesos_i(2353) := b"0000000000000000_0000000000000000_0001001111101001_0100110000010110"; -- 0.07777858294439732
	pesos_i(2354) := b"0000000000000000_0000000000000000_0000101010111101_0000100000010010"; -- 0.04194689211783609
	pesos_i(2355) := b"0000000000000000_0000000000000000_0010000101101111_1001111100011000"; -- 0.13060945836966414
	pesos_i(2356) := b"0000000000000000_0000000000000000_0100010100100111_0011110100001000"; -- 0.2701299806222936
	pesos_i(2357) := b"1111111111111111_1111111111111111_1111110110001100_1000000110100100"; -- -0.009574792419658964
	pesos_i(2358) := b"1111111111111111_1111111111111111_1111001110110011_1000110010011110"; -- -0.04804154537039485
	pesos_i(2359) := b"0000000000000000_0000000000000000_0000001001001111_1110111111101101"; -- 0.009032245107222288
	pesos_i(2360) := b"0000000000000000_0000000000000000_0011000001111111_1101011000000100"; -- 0.18945062242817323
	pesos_i(2361) := b"1111111111111111_1111111111111111_1101101101000100_1100100010011011"; -- -0.14348169537241698
	pesos_i(2362) := b"0000000000000000_0000000000000000_0000101000110010_1111111110000001"; -- 0.03984066861863825
	pesos_i(2363) := b"1111111111111111_1111111111111111_1101011000001100_0011111101100101"; -- -0.16387561583062737
	pesos_i(2364) := b"0000000000000000_0000000000000000_0001010110100100_0101100100010111"; -- 0.08453900160770578
	pesos_i(2365) := b"1111111111111111_1111111111111111_1011010011010110_0110011011001101"; -- -0.29360349184159884
	pesos_i(2366) := b"1111111111111111_1111111111111111_1101011001000001_1010011011101101"; -- -0.1630607291024861
	pesos_i(2367) := b"1111111111111111_1111111111111111_1001111001010010_0001101110110111"; -- -0.38155962731802223
	pesos_i(2368) := b"0000000000000000_0000000000000000_0000000010010001_0011110111010101"; -- 0.002216209971452923
	pesos_i(2369) := b"0000000000000000_0000000000000000_0001111111110111_1010001110011010"; -- 0.12487242225832151
	pesos_i(2370) := b"0000000000000000_0000000000000000_0010000011010000_1111100111101010"; -- 0.1281887241736302
	pesos_i(2371) := b"0000000000000000_0000000000000000_0011001100110000_1010111101101000"; -- 0.1999616269860485
	pesos_i(2372) := b"0000000000000000_0000000000000000_0001000010100100_1011100011111011"; -- 0.06501346718879152
	pesos_i(2373) := b"1111111111111111_1111111111111111_1110000010011010_1101010110011100"; -- -0.12263741429359125
	pesos_i(2374) := b"1111111111111111_1111111111111111_1110100110000100_1110101001100101"; -- -0.0878156187696362
	pesos_i(2375) := b"1111111111111111_1111111111111111_1110001100111011_1111000001100101"; -- -0.1123666526985326
	pesos_i(2376) := b"1111111111111111_1111111111111111_1101001001110000_1011111101110101"; -- -0.17796710382695627
	pesos_i(2377) := b"0000000000000000_0000000000000000_0010010011010110_1010001100110010"; -- 0.1439001081199493
	pesos_i(2378) := b"0000000000000000_0000000000000000_0001100011010101_1010100010110110"; -- 0.0970101779740864
	pesos_i(2379) := b"0000000000000000_0000000000000000_0001101000011011_0010001111100111"; -- 0.10197662735953544
	pesos_i(2380) := b"0000000000000000_0000000000000000_0010000000010111_0010011100101011"; -- 0.1253532866588474
	pesos_i(2381) := b"1111111111111111_1111111111111111_1101111000011010_0100000011010000"; -- -0.13241190838067213
	pesos_i(2382) := b"0000000000000000_0000000000000000_0001001011010100_0000001010100100"; -- 0.07354752056534725
	pesos_i(2383) := b"0000000000000000_0000000000000000_0010101100010001_0100110010101001"; -- 0.16823271876531196
	pesos_i(2384) := b"1111111111111111_1111111111111111_1110000011001110_1111010010000100"; -- -0.12184211516228316
	pesos_i(2385) := b"1111111111111111_1111111111111111_1111110101010110_1001110111001101"; -- -0.010397088389708022
	pesos_i(2386) := b"1111111111111111_1111111111111111_1110110001101000_0011010001101110"; -- -0.07653496091376069
	pesos_i(2387) := b"0000000000000000_0000000000000000_0010110110000100_1000010101011000"; -- 0.17780335812210582
	pesos_i(2388) := b"1111111111111111_1111111111111111_1100000000101000_0110111110101101"; -- -0.2493829921158892
	pesos_i(2389) := b"0000000000000000_0000000000000000_0001010001010011_1100111000101110"; -- 0.07940376881949522
	pesos_i(2390) := b"1111111111111111_1111111111111111_1100000110010001_0010010100011011"; -- -0.24387901382188773
	pesos_i(2391) := b"0000000000000000_0000000000000000_0011111010100011_1111001110110100"; -- 0.24468920853299883
	pesos_i(2392) := b"1111111111111111_1111111111111111_1111111010100001_0000110101111110"; -- -0.005355030823295591
	pesos_i(2393) := b"1111111111111111_1111111111111111_1111010100111100_0111101001111010"; -- -0.04204592256246807
	pesos_i(2394) := b"1111111111111111_1111111111111111_1111010100000101_1101011101010001"; -- -0.042879622238174736
	pesos_i(2395) := b"1111111111111111_1111111111111111_1100110101110010_0010011011010101"; -- -0.1974769335020119
	pesos_i(2396) := b"0000000000000000_0000000000000000_0010101011111101_1000011100101101"; -- 0.16793103070260856
	pesos_i(2397) := b"0000000000000000_0000000000000000_0000101011011000_0110101110010000"; -- 0.04236480954632188
	pesos_i(2398) := b"0000000000000000_0000000000000000_0001100010010100_0010000011010111"; -- 0.0960102582600562
	pesos_i(2399) := b"0000000000000000_0000000000000000_0011111011001100_0101010100100011"; -- 0.24530536746262216
	pesos_i(2400) := b"0000000000000000_0000000000000000_0000011110110101_1100010000111010"; -- 0.030117286940800445
	pesos_i(2401) := b"1111111111111111_1111111111111111_1111010000000111_1000000000110011"; -- -0.0467605473066077
	pesos_i(2402) := b"1111111111111111_1111111111111111_1101001001010110_1110111000001101"; -- -0.1783610552875022
	pesos_i(2403) := b"0000000000000000_0000000000000000_0001101001001110_0100001111000110"; -- 0.10275672512440596
	pesos_i(2404) := b"1111111111111111_1111111111111111_1101110101010001_1100010111101101"; -- -0.13547099069648383
	pesos_i(2405) := b"0000000000000000_0000000000000000_0001100000100010_1100000010101000"; -- 0.09428028203367496
	pesos_i(2406) := b"1111111111111111_1111111111111111_1111110110101011_1010010000110111"; -- -0.009099709078768559
	pesos_i(2407) := b"0000000000000000_0000000000000000_0000100001110101_1100100100010001"; -- 0.03304726291320777
	pesos_i(2408) := b"0000000000000000_0000000000000000_0010100101000011_0011011000111110"; -- 0.16118182203425757
	pesos_i(2409) := b"1111111111111111_1111111111111111_1101101011010100_1000101110100111"; -- -0.1451943128045234
	pesos_i(2410) := b"0000000000000000_0000000000000000_0000011110101101_1010001011010100"; -- 0.02999322580700178
	pesos_i(2411) := b"0000000000000000_0000000000000000_0010110111001111_1000011011100111"; -- 0.17894786011877412
	pesos_i(2412) := b"0000000000000000_0000000000000000_0000101101110111_0011010001010111"; -- 0.04478766548477922
	pesos_i(2413) := b"1111111111111111_1111111111111111_1110011010111011_1110000010011001"; -- -0.09869571937104238
	pesos_i(2414) := b"1111111111111111_1111111111111111_1100111101000001_1001100111010010"; -- -0.19040526026466653
	pesos_i(2415) := b"1111111111111111_1111111111111111_1101011011011010_0101000000011001"; -- -0.16073130971706068
	pesos_i(2416) := b"1111111111111111_1111111111111111_1110101100100100_1011001010110000"; -- -0.08147128304891063
	pesos_i(2417) := b"0000000000000000_0000000000000000_0001011110001000_1000110100110011"; -- 0.09192736149934107
	pesos_i(2418) := b"1111111111111111_1111111111111111_1100111100010110_1000001100000111"; -- -0.19106274669786527
	pesos_i(2419) := b"1111111111111111_1111111111111111_1111100101111011_0010011010000001"; -- -0.0254646238278467
	pesos_i(2420) := b"1111111111111111_1111111111111111_1111011001110010_1010011010011001"; -- -0.03731306809533657
	pesos_i(2421) := b"1111111111111111_1111111111111111_1110000101011100_1011100001100011"; -- -0.11967895102388715
	pesos_i(2422) := b"1111111111111111_1111111111111111_1111111011100011_1001111110111111"; -- -0.004339233178391688
	pesos_i(2423) := b"1111111111111111_1111111111111111_1111011001111111_0110101000001001"; -- -0.037118313706239636
	pesos_i(2424) := b"1111111111111111_1111111111111111_1110001001010110_1101010111000000"; -- -0.11586250366491961
	pesos_i(2425) := b"1111111111111111_1111111111111111_1101111000001011_0001110110111000"; -- -0.13264288185772774
	pesos_i(2426) := b"0000000000000000_0000000000000000_0011011001111001_0000010101110011"; -- 0.21278413837340865
	pesos_i(2427) := b"1111111111111111_1111111111111111_1111010000111100_1100101101001011"; -- -0.04594735538895282
	pesos_i(2428) := b"1111111111111111_1111111111111111_1111111011101010_1010000111000011"; -- -0.004232301540669524
	pesos_i(2429) := b"1111111111111111_1111111111111111_1101011100010001_0010111000011011"; -- -0.1598941025933051
	pesos_i(2430) := b"0000000000000000_0000000000000000_0000000100000011_0111111011000111"; -- 0.003959582910432976
	pesos_i(2431) := b"1111111111111111_1111111111111111_1111100111101010_1101011100100101"; -- -0.023760369768564032
	pesos_i(2432) := b"0000000000000000_0000000000000000_0000001110000010_0011010010010110"; -- 0.01370552690911514
	pesos_i(2433) := b"0000000000000000_0000000000000000_0101001011010010_1010000011001001"; -- 0.3235264291677548
	pesos_i(2434) := b"0000000000000000_0000000000000000_0001101111100010_1101100101100100"; -- 0.10893019386649169
	pesos_i(2435) := b"0000000000000000_0000000000000000_0000000000011101_1000000100100111"; -- 0.00045020301889128755
	pesos_i(2436) := b"0000000000000000_0000000000000000_0000000100011110_0011011001010001"; -- 0.004367251115431082
	pesos_i(2437) := b"1111111111111111_1111111111111111_1101110111000000_0100011111011111"; -- -0.13378477872484767
	pesos_i(2438) := b"0000000000000000_0000000000000000_0000010111100001_1111101000110000"; -- 0.02297938986934836
	pesos_i(2439) := b"1111111111111111_1111111111111111_1100111011110010_0111111110110000"; -- -0.1916122622773175
	pesos_i(2440) := b"0000000000000000_0000000000000000_0010011101000111_0010100100001101"; -- 0.15342957095188187
	pesos_i(2441) := b"0000000000000000_0000000000000000_0000010010001011_0000100011000100"; -- 0.01774649419664261
	pesos_i(2442) := b"1111111111111111_1111111111111111_1101110000000010_0110110011100111"; -- -0.14058799133442504
	pesos_i(2443) := b"1111111111111111_1111111111111111_1101001011010111_1011101000010001"; -- -0.17639576996176018
	pesos_i(2444) := b"0000000000000000_0000000000000000_0001010111110010_0011111111110010"; -- 0.08572768846341185
	pesos_i(2445) := b"1111111111111111_1111111111111111_1101001101101000_1101101101000000"; -- -0.17418126770359219
	pesos_i(2446) := b"0000000000000000_0000000000000000_0000111101100101_0111110010101010"; -- 0.06014231818218731
	pesos_i(2447) := b"1111111111111111_1111111111111111_1110110001000100_1001110001110101"; -- -0.07707807676445463
	pesos_i(2448) := b"1111111111111111_1111111111111111_1111011101111101_0010010101101000"; -- -0.03324667174087615
	pesos_i(2449) := b"0000000000000000_0000000000000000_0001100010010110_0100110010110101"; -- 0.09604339048076559
	pesos_i(2450) := b"0000000000000000_0000000000000000_0000100110110100_1100001101010101"; -- 0.037914474660632094
	pesos_i(2451) := b"0000000000000000_0000000000000000_0001100011000111_1011001101100000"; -- 0.0967971907048821
	pesos_i(2452) := b"0000000000000000_0000000000000000_0000010100110011_0010000000011001"; -- 0.02031136132471781
	pesos_i(2453) := b"1111111111111111_1111111111111111_1110110010111011_0111001101010010"; -- -0.07526473277560923
	pesos_i(2454) := b"0000000000000000_0000000000000000_0001001110100000_0001101011001110"; -- 0.07666175389014784
	pesos_i(2455) := b"0000000000000000_0000000000000000_0010011011101000_0010101000100111"; -- 0.15198005151172334
	pesos_i(2456) := b"1111111111111111_1111111111111111_1101010000101010_1101010011101101"; -- -0.17122143955607347
	pesos_i(2457) := b"0000000000000000_0000000000000000_0000110100001101_1100100001010000"; -- 0.05099155379033442
	pesos_i(2458) := b"0000000000000000_0000000000000000_0010111000101110_1000010010000101"; -- 0.1803973029960056
	pesos_i(2459) := b"0000000000000000_0000000000000000_0000011000101010_1000011111101000"; -- 0.02408646973800032
	pesos_i(2460) := b"1111111111111111_1111111111111111_1101011010010110_0010001101011010"; -- -0.16177157461714992
	pesos_i(2461) := b"1111111111111111_1111111111111111_1101001010111001_1100000011101111"; -- -0.17685312420694002
	pesos_i(2462) := b"0000000000000000_0000000000000000_0000010110000010_1111000011001111"; -- 0.021529245971021876
	pesos_i(2463) := b"1111111111111111_1111111111111111_1100000101111001_1010111110111110"; -- -0.24423696143523455
	pesos_i(2464) := b"1111111111111111_1111111111111111_1110000111100001_1100100000110110"; -- -0.11764858899720494
	pesos_i(2465) := b"0000000000000000_0000000000000000_0001100101101111_1000000001101110"; -- 0.09935763058146982
	pesos_i(2466) := b"1111111111111111_1111111111111111_1110100111101001_0110001010000011"; -- -0.08628258043495851
	pesos_i(2467) := b"0000000000000000_0000000000000000_0100000100000101_1001010000100111"; -- 0.25399137459830734
	pesos_i(2468) := b"0000000000000000_0000000000000000_0011111011111101_1111101101001110"; -- 0.24606295249414212
	pesos_i(2469) := b"0000000000000000_0000000000000000_0001010110100101_1100001000010000"; -- 0.08456051714930662
	pesos_i(2470) := b"1111111111111111_1111111111111111_1110111100101001_1110011100100101"; -- -0.06576686239484644
	pesos_i(2471) := b"1111111111111111_1111111111111111_1110000011101101_1011110000000001"; -- -0.12137246106084285
	pesos_i(2472) := b"1111111111111111_1111111111111111_1100010111000101_0101011110010110"; -- -0.22745754798443693
	pesos_i(2473) := b"0000000000000000_0000000000000000_0010000110001001_1010000000001000"; -- 0.13100624281557624
	pesos_i(2474) := b"0000000000000000_0000000000000000_0000000101101011_0100000100001011"; -- 0.005542817209564704
	pesos_i(2475) := b"1111111111111111_1111111111111111_1101111001010111_1111100001111011"; -- -0.13147017478540957
	pesos_i(2476) := b"0000000000000000_0000000000000000_0001011000100000_0100000001001100"; -- 0.0864296136568638
	pesos_i(2477) := b"0000000000000000_0000000000000000_0010110001101001_0010100000011101"; -- 0.17347956380968363
	pesos_i(2478) := b"0000000000000000_0000000000000000_0001100101101111_1010110010110011"; -- 0.09936026929376485
	pesos_i(2479) := b"0000000000000000_0000000000000000_0011111000101110_1110011110110001"; -- 0.2429032141535785
	pesos_i(2480) := b"0000000000000000_0000000000000000_0001000110010000_1101010011111110"; -- 0.06861621095308475
	pesos_i(2481) := b"1111111111111111_1111111111111111_1110101010111000_1010110110101101"; -- -0.08311953097454415
	pesos_i(2482) := b"1111111111111111_1111111111111111_1110000001010011_0011011011000100"; -- -0.12373025629138941
	pesos_i(2483) := b"0000000000000000_0000000000000000_0000101111101001_0110011011011011"; -- 0.04653017844471431
	pesos_i(2484) := b"0000000000000000_0000000000000000_0010000100011101_0100010100100011"; -- 0.12935287565896894
	pesos_i(2485) := b"0000000000000000_0000000000000000_0000010101010111_1010010001100011"; -- 0.0208685627906971
	pesos_i(2486) := b"1111111111111111_1111111111111111_1111010000010010_1101111011011000"; -- -0.046587059265129016
	pesos_i(2487) := b"0000000000000000_0000000000000000_0001000001101000_0001111011100000"; -- 0.06408875446096507
	pesos_i(2488) := b"1111111111111111_1111111111111111_1100000110100000_1111101010001110"; -- -0.24363740947836768
	pesos_i(2489) := b"1111111111111111_1111111111111111_1100011101000001_0011010100100000"; -- -0.2216612621411959
	pesos_i(2490) := b"0000000000000000_0000000000000000_0001001001111111_0010000001010111"; -- 0.07225229375769768
	pesos_i(2491) := b"0000000000000000_0000000000000000_0010001000101110_1011101001111110"; -- 0.13352552014709523
	pesos_i(2492) := b"1111111111111111_1111111111111111_1110001110100100_1101000010101111"; -- -0.11076637013508633
	pesos_i(2493) := b"1111111111111111_1111111111111111_1111011001111101_0101111111100000"; -- -0.03714943681934391
	pesos_i(2494) := b"0000000000000000_0000000000000000_0001101010000100_0000001011100001"; -- 0.10357683181501315
	pesos_i(2495) := b"0000000000000000_0000000000000000_0010010001010110_0000101111010000"; -- 0.14193795989852875
	pesos_i(2496) := b"0000000000000000_0000000000000000_0000010011001001_1100001101110101"; -- 0.018703666796001134
	pesos_i(2497) := b"1111111111111111_1111111111111111_1110010001011010_0100111100100011"; -- -0.10799699210758029
	pesos_i(2498) := b"1111111111111111_1111111111111111_1111011111111100_1101111010100101"; -- -0.031297764429208015
	pesos_i(2499) := b"1111111111111111_1111111111111111_1101110110100100_1010001101011101"; -- -0.134206571386329
	pesos_i(2500) := b"0000000000000000_0000000000000000_0000110111111111_1111000110011011"; -- 0.054686642056660274
	pesos_i(2501) := b"1111111111111111_1111111111111111_1111100111010101_0100011000110000"; -- -0.024089444398299104
	pesos_i(2502) := b"1111111111111111_1111111111111111_1110100110101000_0111100111101110"; -- -0.08727300584921183
	pesos_i(2503) := b"0000000000000000_0000000000000000_0000010111110100_1101000101001111"; -- 0.023266870286132894
	pesos_i(2504) := b"0000000000000000_0000000000000000_0000100111001110_0001100000000110"; -- 0.03830099255960282
	pesos_i(2505) := b"0000000000000000_0000000000000000_0000010111000001_0100110110011111"; -- 0.02248082284855416
	pesos_i(2506) := b"1111111111111111_1111111111111111_1110011101001010_1100101011001000"; -- -0.09651501285878732
	pesos_i(2507) := b"0000000000000000_0000000000000000_0001011111000001_0110111101001001"; -- 0.0927953293602552
	pesos_i(2508) := b"0000000000000000_0000000000000000_0000011111001111_0011100110100001"; -- 0.030505754381134627
	pesos_i(2509) := b"0000000000000000_0000000000000000_0000111000001000_0000011110011011"; -- 0.054810023617633825
	pesos_i(2510) := b"0000000000000000_0000000000000000_0000110101110001_0001101010011001"; -- 0.05250707849086593
	pesos_i(2511) := b"1111111111111111_1111111111111111_1111111101110011_1001110100100011"; -- -0.0021421231603503954
	pesos_i(2512) := b"0000000000000000_0000000000000000_0000111110010110_0011100000101011"; -- 0.060885916199593174
	pesos_i(2513) := b"0000000000000000_0000000000000000_0001100100000010_1010001111111111"; -- 0.09769654243586336
	pesos_i(2514) := b"1111111111111111_1111111111111111_1101011110011000_1001010111100100"; -- -0.15782797997360853
	pesos_i(2515) := b"0000000000000000_0000000000000000_0010000001110110_1100001101011110"; -- 0.12681218198057614
	pesos_i(2516) := b"0000000000000000_0000000000000000_0001101110110010_0111100101110010"; -- 0.10819205307302987
	pesos_i(2517) := b"1111111111111111_1111111111111111_1111010110111001_0110111111101010"; -- -0.040139203477581945
	pesos_i(2518) := b"1111111111111111_1111111111111111_1111000011001101_1110110000101110"; -- -0.05935787081006495
	pesos_i(2519) := b"0000000000000000_0000000000000000_0001010001010111_1011111110111011"; -- 0.07946394268930311
	pesos_i(2520) := b"1111111111111111_1111111111111111_1110100110110100_0111110000000100"; -- -0.08708977611874558
	pesos_i(2521) := b"0000000000000000_0000000000000000_0001100100110001_1100100000100110"; -- 0.09841586036051414
	pesos_i(2522) := b"1111111111111111_1111111111111111_1101101001100110_1101101011010100"; -- -0.1468680603922519
	pesos_i(2523) := b"0000000000000000_0000000000000000_0000110010000111_0111001010110100"; -- 0.048941773293501065
	pesos_i(2524) := b"0000000000000000_0000000000000000_0000111100010101_0010101011001100"; -- 0.058916735503750366
	pesos_i(2525) := b"0000000000000000_0000000000000000_0010001101011110_0000110101001001"; -- 0.13815386813495129
	pesos_i(2526) := b"1111111111111111_1111111111111111_1110010111000110_0000110011000100"; -- -0.10244674876156144
	pesos_i(2527) := b"0000000000000000_0000000000000000_0001001001011101_1110010111010101"; -- 0.0717452663960671
	pesos_i(2528) := b"1111111111111111_1111111111111111_1110100001101110_0110101000110101"; -- -0.09206520282338251
	pesos_i(2529) := b"1111111111111111_1111111111111111_1100111100101001_0011001010110000"; -- -0.19077761853153485
	pesos_i(2530) := b"1111111111111111_1111111111111111_1110101101010010_1101001101011100"; -- -0.08076743139003759
	pesos_i(2531) := b"1111111111111111_1111111111111111_1110101001100010_0110011100100101"; -- -0.08443599085518004
	pesos_i(2532) := b"1111111111111111_1111111111111111_1100011100000010_0111100001000010"; -- -0.22261856445433847
	pesos_i(2533) := b"0000000000000000_0000000000000000_0010001000110010_0000000000111010"; -- 0.13357545286685654
	pesos_i(2534) := b"1111111111111111_1111111111111111_1111111110010110_0010010010111001"; -- -0.0016152428074596068
	pesos_i(2535) := b"1111111111111111_1111111111111111_1110001010111110_0000101000111101"; -- -0.11428771975069457
	pesos_i(2536) := b"1111111111111111_1111111111111111_1111101100100010_1011111011100000"; -- -0.019001074198922722
	pesos_i(2537) := b"1111111111111111_1111111111111111_1110001110101000_0011111010011101"; -- -0.11071404134142354
	pesos_i(2538) := b"1111111111111111_1111111111111111_1110100001100011_0100110001010111"; -- -0.0922348296459829
	pesos_i(2539) := b"1111111111111111_1111111111111111_1110110010011000_1111000110101000"; -- -0.07579126019040824
	pesos_i(2540) := b"1111111111111111_1111111111111111_1111010001011000_0110010000101000"; -- -0.04552625670290301
	pesos_i(2541) := b"1111111111111111_1111111111111111_1110100100011110_1101111111011001"; -- -0.08937264390980944
	pesos_i(2542) := b"0000000000000000_0000000000000000_0010111100110010_1101101110000001"; -- 0.18436977300757212
	pesos_i(2543) := b"0000000000000000_0000000000000000_0001000001101011_0110000001111010"; -- 0.06413844090615783
	pesos_i(2544) := b"1111111111111111_1111111111111111_1110110010001000_1010001111100101"; -- -0.07604003590303562
	pesos_i(2545) := b"1111111111111111_1111111111111111_1110110101100000_1000111011100110"; -- -0.0727453887410506
	pesos_i(2546) := b"1111111111111111_1111111111111111_1110011100111111_0010001010000010"; -- -0.09669288956037093
	pesos_i(2547) := b"0000000000000000_0000000000000000_0001011100000000_0111111111110111"; -- 0.08985137733942898
	pesos_i(2548) := b"0000000000000000_0000000000000000_0000111001110011_0111110101111110"; -- 0.05644974075185936
	pesos_i(2549) := b"1111111111111111_1111111111111111_1110111111100011_0100110011101101"; -- -0.06293791980625438
	pesos_i(2550) := b"1111111111111111_1111111111111111_1101011101101001_1101001001011001"; -- -0.1585415395566731
	pesos_i(2551) := b"0000000000000000_0000000000000000_0001001110100011_0100101001000100"; -- 0.07671035921748183
	pesos_i(2552) := b"1111111111111111_1111111111111111_1111011010110011_1011111001100101"; -- -0.03631982829626764
	pesos_i(2553) := b"0000000000000000_0000000000000000_0000100110110001_1011100101001011"; -- 0.03786809987264399
	pesos_i(2554) := b"1111111111111111_1111111111111111_1101110000101010_0100110100000100"; -- -0.13997954029692145
	pesos_i(2555) := b"1111111111111111_1111111111111111_1111101101011111_1000110001010001"; -- -0.018073301630746226
	pesos_i(2556) := b"1111111111111111_1111111111111111_1111000110110000_0011011100111111"; -- -0.05590491014999744
	pesos_i(2557) := b"0000000000000000_0000000000000000_0001000011011110_1110110101000110"; -- 0.06590159368082399
	pesos_i(2558) := b"0000000000000000_0000000000000000_0000111011110011_0100100001110010"; -- 0.05839970386624267
	pesos_i(2559) := b"0000000000000000_0000000000000000_0001011111011101_0010010000110110"; -- 0.09321810083669489
	pesos_i(2560) := b"0000000000000000_0000000000000000_0011000110010110_1001110000111010"; -- 0.1937043801896795
	pesos_i(2561) := b"0000000000000000_0000000000000000_0000111010001110_1001001010100110"; -- 0.05686298898128781
	pesos_i(2562) := b"0000000000000000_0000000000000000_0000100010000010_0110100001101001"; -- 0.033239865973997314
	pesos_i(2563) := b"0000000000000000_0000000000000000_0010010010000110_1001101011011110"; -- 0.1426789085440744
	pesos_i(2564) := b"1111111111111111_1111111111111111_1101011010111001_0001110010101101"; -- -0.16123791485087716
	pesos_i(2565) := b"0000000000000000_0000000000000000_0001101111101000_0100000111010111"; -- 0.10901271338902485
	pesos_i(2566) := b"1111111111111111_1111111111111111_1110001001011000_0100100001111110"; -- -0.11584040562819145
	pesos_i(2567) := b"0000000000000000_0000000000000000_0001110110010001_0101101100000101"; -- 0.11549919953874101
	pesos_i(2568) := b"1111111111111111_1111111111111111_1101100000100001_0001000111100111"; -- -0.15574539289493258
	pesos_i(2569) := b"0000000000000000_0000000000000000_0001110111001110_0000101101100001"; -- 0.11642523868277055
	pesos_i(2570) := b"1111111111111111_1111111111111111_1111111000100100_0011011111101010"; -- -0.007259850758446401
	pesos_i(2571) := b"1111111111111111_1111111111111111_1111000110010111_1110110111101111"; -- -0.05627549084584592
	pesos_i(2572) := b"1111111111111111_1111111111111111_1111011110101101_1101100101000001"; -- -0.032503530047815796
	pesos_i(2573) := b"0000000000000000_0000000000000000_0000100010001001_0010011100000011"; -- 0.03334277942429403
	pesos_i(2574) := b"1111111111111111_1111111111111111_1111100001000100_0111001000101110"; -- -0.030205596807771053
	pesos_i(2575) := b"1111111111111111_1111111111111111_1111110100001000_0100000101100010"; -- -0.011592782493248851
	pesos_i(2576) := b"1111111111111111_1111111111111111_1111010000001010_1000101001000111"; -- -0.046714170133665384
	pesos_i(2577) := b"1111111111111111_1111111111111111_1110100000010110_0000110101101111"; -- -0.09341350598848469
	pesos_i(2578) := b"1111111111111111_1111111111111111_1101101100100110_0100110000101100"; -- -0.14394687580457532
	pesos_i(2579) := b"1111111111111111_1111111111111111_1110001100110111_0001111110101110"; -- -0.11244012824122981
	pesos_i(2580) := b"1111111111111111_1111111111111111_1101110010100111_0010111001010111"; -- -0.13807402011834324
	pesos_i(2581) := b"1111111111111111_1111111111111111_1110010110010110_1001110111011100"; -- -0.10317052248940205
	pesos_i(2582) := b"0000000000000000_0000000000000000_0000110011101011_1011001100011011"; -- 0.05047149099510681
	pesos_i(2583) := b"1111111111111111_1111111111111111_1110011010100111_0011010110001110"; -- -0.09901109010819702
	pesos_i(2584) := b"0000000000000000_0000000000000000_0001001100110101_0001011010101100"; -- 0.0750288170752913
	pesos_i(2585) := b"1111111111111111_1111111111111111_1101010101101011_1111111011111001"; -- -0.16632086197533977
	pesos_i(2586) := b"1111111111111111_1111111111111111_1111000000001101_0110101110001001"; -- -0.06229522622411377
	pesos_i(2587) := b"0000000000000000_0000000000000000_0000001000000111_1001110010100100"; -- 0.007928648052298481
	pesos_i(2588) := b"0000000000000000_0000000000000000_0001011110100011_0101010111101111"; -- 0.09233605462445775
	pesos_i(2589) := b"1111111111111111_1111111111111111_1110101010100010_1000000111011010"; -- -0.08345783631987176
	pesos_i(2590) := b"1111111111111111_1111111111111111_1110100000010101_1111000011111100"; -- -0.09341520156905482
	pesos_i(2591) := b"1111111111111111_1111111111111111_1100100100100100_0000101101111100"; -- -0.21429374903302092
	pesos_i(2592) := b"1111111111111111_1111111111111111_1110011001111100_1000110101111000"; -- -0.09966197799277225
	pesos_i(2593) := b"1111111111111111_1111111111111111_1111100010001111_0111001000000000"; -- -0.02906119832855766
	pesos_i(2594) := b"0000000000000000_0000000000000000_0000000111001011_0001000110110001"; -- 0.007004838699003257
	pesos_i(2595) := b"0000000000000000_0000000000000000_0001111100111111_0100001110100000"; -- 0.12205908438281221
	pesos_i(2596) := b"0000000000000000_0000000000000000_0001111111111001_0010101111101100"; -- 0.12489580637728936
	pesos_i(2597) := b"0000000000000000_0000000000000000_0000001001011011_1111001010010101"; -- 0.009215508834814284
	pesos_i(2598) := b"0000000000000000_0000000000000000_0000001110110110_1010011111001010"; -- 0.014505850574054633
	pesos_i(2599) := b"1111111111111111_1111111111111111_1110100000011011_1001000010110111"; -- -0.0933293869809781
	pesos_i(2600) := b"1111111111111111_1111111111111111_1110110110100111_1101001101111110"; -- -0.07165792631962527
	pesos_i(2601) := b"1111111111111111_1111111111111111_1110111100101111_1000110100000000"; -- -0.06568068258800085
	pesos_i(2602) := b"1111111111111111_1111111111111111_1101000101110010_1000001001110100"; -- -0.18184647238286228
	pesos_i(2603) := b"0000000000000000_0000000000000000_0010000100110000_1000110110001101"; -- 0.12964710906665594
	pesos_i(2604) := b"1111111111111111_1111111111111111_1101000011110010_1100011011010001"; -- -0.18379552271873242
	pesos_i(2605) := b"1111111111111111_1111111111111111_1101100100011001_1111100011001101"; -- -0.1519474506276784
	pesos_i(2606) := b"1111111111111111_1111111111111111_1101100110110000_1101110011010001"; -- -0.14964504149653204
	pesos_i(2607) := b"0000000000000000_0000000000000000_0000000010101011_0000111110011101"; -- 0.0026101835521394434
	pesos_i(2608) := b"1111111111111111_1111111111111111_1100111001111001_0010001000001100"; -- -0.19346415721149993
	pesos_i(2609) := b"1111111111111111_1111111111111111_1110111000110010_1010111101001010"; -- -0.06953911260979163
	pesos_i(2610) := b"0000000000000000_0000000000000000_0001100110001111_0110100010010101"; -- 0.09984449042527474
	pesos_i(2611) := b"1111111111111111_1111111111111111_1111000010000111_1000000100110011"; -- -0.06043236259768417
	pesos_i(2612) := b"0000000000000000_0000000000000000_0000100011101000_1110000010010000"; -- 0.034803424018815504
	pesos_i(2613) := b"0000000000000000_0000000000000000_0010100010110111_1101110100110000"; -- 0.1590555420895016
	pesos_i(2614) := b"1111111111111111_1111111111111111_1111100111101101_1101000111011100"; -- -0.023714908454156435
	pesos_i(2615) := b"1111111111111111_1111111111111111_1110011101110111_0011101111011111"; -- -0.09583688546329037
	pesos_i(2616) := b"1111111111111111_1111111111111111_1100111010110110_0011110100010100"; -- -0.19253175979106568
	pesos_i(2617) := b"0000000000000000_0000000000000000_0000001001101000_1000000110111000"; -- 0.009407145959432019
	pesos_i(2618) := b"0000000000000000_0000000000000000_0010011010101100_0000010110010111"; -- 0.15106234485877593
	pesos_i(2619) := b"0000000000000000_0000000000000000_0000000010000101_0011111000000011"; -- 0.002033115175696327
	pesos_i(2620) := b"1111111111111111_1111111111111111_1110101100101000_1000000101111011"; -- -0.08141318072942277
	pesos_i(2621) := b"0000000000000000_0000000000000000_0001000010100101_0100101101110111"; -- 0.06502219822992666
	pesos_i(2622) := b"1111111111111111_1111111111111111_1101001001111100_1101100100100011"; -- -0.1777824677185466
	pesos_i(2623) := b"0000000000000000_0000000000000000_0010101101100000_1001000010010101"; -- 0.16944221152650157
	pesos_i(2624) := b"1111111111111111_1111111111111111_1110011100100000_1000000111101111"; -- -0.09716022421331354
	pesos_i(2625) := b"0000000000000000_0000000000000000_0000010111110101_0000110000001011"; -- 0.023270371185092287
	pesos_i(2626) := b"1111111111111111_1111111111111111_1111101110011101_1110101010011001"; -- -0.01712163697220567
	pesos_i(2627) := b"0000000000000000_0000000000000000_0010100100000110_0111111010110111"; -- 0.16025535552167078
	pesos_i(2628) := b"1111111111111111_1111111111111111_1110100111010101_1110110001000110"; -- -0.08657954487407775
	pesos_i(2629) := b"1111111111111111_1111111111111111_1111010101100010_0001100111101001"; -- -0.04147184422757176
	pesos_i(2630) := b"1111111111111111_1111111111111111_1111101010110100_1111100001111000"; -- -0.020676108088582067
	pesos_i(2631) := b"1111111111111111_1111111111111111_1110001001110011_0100001101011110"; -- -0.11542872377454837
	pesos_i(2632) := b"1111111111111111_1111111111111111_1111101010111001_1010001100100010"; -- -0.020604900596432937
	pesos_i(2633) := b"1111111111111111_1111111111111111_1111001111100100_1110011111100000"; -- -0.04728842536552307
	pesos_i(2634) := b"0000000000000000_0000000000000000_0000000010000000_1110100010101111"; -- 0.0019669939215408903
	pesos_i(2635) := b"0000000000000000_0000000000000000_0000111010010100_1001000000110011"; -- 0.05695439568325591
	pesos_i(2636) := b"1111111111111111_1111111111111111_1110101010100001_0010000101000011"; -- -0.08347885230245665
	pesos_i(2637) := b"0000000000000000_0000000000000000_0001001001101011_0110111011101010"; -- 0.07195180152437741
	pesos_i(2638) := b"0000000000000000_0000000000000000_0001100101011011_1010110011010010"; -- 0.09905510062331838
	pesos_i(2639) := b"0000000000000000_0000000000000000_0010000001100000_1100000010110100"; -- 0.1264763296352626
	pesos_i(2640) := b"0000000000000000_0000000000000000_0000100011001000_0000110011001100"; -- 0.03430252046825801
	pesos_i(2641) := b"1111111111111111_1111111111111111_1110100110010000_0001100010100101"; -- -0.08764501554419857
	pesos_i(2642) := b"0000000000000000_0000000000000000_0000100000111110_1001000001010001"; -- 0.03220464681967908
	pesos_i(2643) := b"0000000000000000_0000000000000000_0001101111001110_0111001011011011"; -- 0.10861890643299775
	pesos_i(2644) := b"0000000000000000_0000000000000000_0001010001110011_1001001010001110"; -- 0.07988849606251737
	pesos_i(2645) := b"0000000000000000_0000000000000000_0010010100011111_0110001010110101"; -- 0.14501015575854734
	pesos_i(2646) := b"1111111111111111_1111111111111111_1111110110001100_0110110111111100"; -- -0.009575963923206338
	pesos_i(2647) := b"1111111111111111_1111111111111111_1110101001101010_0111101010000000"; -- -0.08431276679957483
	pesos_i(2648) := b"0000000000000000_0000000000000000_0001010100111101_0011001010101110"; -- 0.08296505689534486
	pesos_i(2649) := b"0000000000000000_0000000000000000_0001011111000011_1110100001011110"; -- 0.09283306405330313
	pesos_i(2650) := b"0000000000000000_0000000000000000_0001000100001110_0011101101000001"; -- 0.06662340479093158
	pesos_i(2651) := b"0000000000000000_0000000000000000_0000100001101100_1000111000101110"; -- 0.032906423744993245
	pesos_i(2652) := b"1111111111111111_1111111111111111_1110111011011111_1010010010100011"; -- -0.06689997696203198
	pesos_i(2653) := b"0000000000000000_0000000000000000_0010001111101000_1000000000100101"; -- 0.1402664269722052
	pesos_i(2654) := b"0000000000000000_0000000000000000_0010001010110100_0010110101011001"; -- 0.13556178506327385
	pesos_i(2655) := b"0000000000000000_0000000000000000_0001001111011100_0110111000000001"; -- 0.07758224024660192
	pesos_i(2656) := b"0000000000000000_0000000000000000_0001110000110000_1100000101010101"; -- 0.11011894535184459
	pesos_i(2657) := b"1111111111111111_1111111111111111_1110000110010111_0010101101111110"; -- -0.11878708055601812
	pesos_i(2658) := b"0000000000000000_0000000000000000_0001100000001001_1000100100001110"; -- 0.09389549814072279
	pesos_i(2659) := b"1111111111111111_1111111111111111_1101100100100111_0100100110000000"; -- -0.15174427619792671
	pesos_i(2660) := b"1111111111111111_1111111111111111_1101011000010111_1111100101101101"; -- -0.16369668097157164
	pesos_i(2661) := b"0000000000000000_0000000000000000_0010101100111111_1010101101000000"; -- 0.16894026095542783
	pesos_i(2662) := b"1111111111111111_1111111111111111_1101111001000110_1110001001111011"; -- -0.13173088556186963
	pesos_i(2663) := b"1111111111111111_1111111111111111_1111000100000110_1100001110011010"; -- -0.05849053856982869
	pesos_i(2664) := b"1111111111111111_1111111111111111_1111001100011111_1010001101010000"; -- -0.05029849341915448
	pesos_i(2665) := b"1111111111111111_1111111111111111_1110000110110101_1100001100101110"; -- -0.1183202754953644
	pesos_i(2666) := b"1111111111111111_1111111111111111_1101111000101000_1000010100001001"; -- -0.13219421899800107
	pesos_i(2667) := b"1111111111111111_1111111111111111_1110111000000101_0110110111111111"; -- -0.07022964985529266
	pesos_i(2668) := b"1111111111111111_1111111111111111_1111111001000001_0001011010011010"; -- -0.006819331649871235
	pesos_i(2669) := b"1111111111111111_1111111111111111_1111111001101010_1011001000100101"; -- -0.0061844501500998095
	pesos_i(2670) := b"1111111111111111_1111111111111111_1101001110000111_0000001110100000"; -- -0.17372109752251974
	pesos_i(2671) := b"1111111111111111_1111111111111111_1100111000000111_0011001101101100"; -- -0.1952026235303022
	pesos_i(2672) := b"0000000000000000_0000000000000000_0001000001111101_1011000011100101"; -- 0.06441789237684845
	pesos_i(2673) := b"0000000000000000_0000000000000000_0001111100110000_0001000110100100"; -- 0.12182722332927648
	pesos_i(2674) := b"1111111111111111_1111111111111111_1101011111111100_0101001100111010"; -- -0.1563060745024125
	pesos_i(2675) := b"1111111111111111_1111111111111111_1111110000111011_1111111010101111"; -- -0.014709551100658427
	pesos_i(2676) := b"0000000000000000_0000000000000000_0010111000000101_1101000100001000"; -- 0.179776253209416
	pesos_i(2677) := b"0000000000000000_0000000000000000_0010100011110011_0100101100011001"; -- 0.15996236196968056
	pesos_i(2678) := b"1111111111111111_1111111111111111_1101000101110001_1000101110101011"; -- -0.181861182040675
	pesos_i(2679) := b"0000000000000000_0000000000000000_0001000001101010_1100101010110111"; -- 0.06412951449891675
	pesos_i(2680) := b"0000000000000000_0000000000000000_0001111011000001_0000001011100011"; -- 0.12013261828385789
	pesos_i(2681) := b"1111111111111111_1111111111111111_1101111110101101_0110011000001110"; -- -0.1262603965236791
	pesos_i(2682) := b"0000000000000000_0000000000000000_0000101010001111_1001010100000101"; -- 0.0412533890828945
	pesos_i(2683) := b"0000000000000000_0000000000000000_0001001000011100_0000111110001001"; -- 0.07074067213783337
	pesos_i(2684) := b"0000000000000000_0000000000000000_0010101000010001_1111100101100110"; -- 0.16433676483173976
	pesos_i(2685) := b"0000000000000000_0000000000000000_0000011001010100_1101100111000001"; -- 0.024732217316379198
	pesos_i(2686) := b"1111111111111111_1111111111111111_1100111000010000_1001100011111110"; -- -0.1950592404442112
	pesos_i(2687) := b"0000000000000000_0000000000000000_0000110110110010_1010010001100000"; -- 0.053507111958172954
	pesos_i(2688) := b"0000000000000000_0000000000000000_0010001011100000_1011010101111011"; -- 0.13624128582584671
	pesos_i(2689) := b"0000000000000000_0000000000000000_0000111000011101_0100100111101000"; -- 0.05513440993809252
	pesos_i(2690) := b"0000000000000000_0000000000000000_0011000011110010_0111101100001101"; -- 0.19119996129090389
	pesos_i(2691) := b"0000000000000000_0000000000000000_0001010100111101_0011001000010011"; -- 0.08296502078312311
	pesos_i(2692) := b"1111111111111111_1111111111111111_1110101010110001_0001000111111111"; -- -0.08323562172019687
	pesos_i(2693) := b"0000000000000000_0000000000000000_0010110101011010_1111110111110111"; -- 0.177169678449193
	pesos_i(2694) := b"1111111111111111_1111111111111111_1101101101101101_1000100111110101"; -- -0.1428598190275875
	pesos_i(2695) := b"1111111111111111_1111111111111111_1111111110001110_0001000100010110"; -- -0.0017384835537636364
	pesos_i(2696) := b"0000000000000000_0000000000000000_0000010110001010_0111111000011011"; -- 0.02164447946785314
	pesos_i(2697) := b"1111111111111111_1111111111111111_1110010001110000_0110101111110011"; -- -0.10765958145612005
	pesos_i(2698) := b"0000000000000000_0000000000000000_0010101001010001_0100000111010111"; -- 0.16530238638025646
	pesos_i(2699) := b"0000000000000000_0000000000000000_0010010011001101_1100000101100100"; -- 0.14376457875319112
	pesos_i(2700) := b"1111111111111111_1111111111111111_1111111000000100_1010101011000111"; -- -0.007741285694932277
	pesos_i(2701) := b"0000000000000000_0000000000000000_0001001101101000_0001000110011000"; -- 0.0758067126741974
	pesos_i(2702) := b"0000000000000000_0000000000000000_0000100010110001_0101010100111011"; -- 0.03395588571898836
	pesos_i(2703) := b"0000000000000000_0000000000000000_0000100010110001_1001111001110101"; -- 0.03396025053010314
	pesos_i(2704) := b"1111111111111111_1111111111111111_1100111011001101_0101100100111000"; -- -0.19217913035512396
	pesos_i(2705) := b"0000000000000000_0000000000000000_0010111001101110_0011001010000101"; -- 0.18136897798885127
	pesos_i(2706) := b"1111111111111111_1111111111111111_1111000111001010_0101101101111000"; -- -0.055506022753739594
	pesos_i(2707) := b"1111111111111111_1111111111111111_1101010111101000_0110011110010100"; -- -0.16442253731530457
	pesos_i(2708) := b"1111111111111111_1111111111111111_1101000000111011_1010000101000000"; -- -0.1865901201884925
	pesos_i(2709) := b"1111111111111111_1111111111111111_1101011110101101_1101100100010111"; -- -0.15750354004304837
	pesos_i(2710) := b"1111111111111111_1111111111111111_1101011100101010_1111111000110111"; -- -0.1595002283711599
	pesos_i(2711) := b"0000000000000000_0000000000000000_0010001010101100_0100111010101110"; -- 0.13544170137382017
	pesos_i(2712) := b"0000000000000000_0000000000000000_0001010010001001_0110011011101100"; -- 0.08022158881514671
	pesos_i(2713) := b"1111111111111111_1111111111111111_1101010110110000_1000010101010001"; -- -0.1652752569021301
	pesos_i(2714) := b"1111111111111111_1111111111111111_1110110110011010_1101111101110000"; -- -0.07185557850243912
	pesos_i(2715) := b"0000000000000000_0000000000000000_0000101101011010_0111111100111101"; -- 0.04434962504789357
	pesos_i(2716) := b"1111111111111111_1111111111111111_1111110101100101_1110010101110010"; -- -0.010163936396137125
	pesos_i(2717) := b"1111111111111111_1111111111111111_1111001011100010_1000010101001011"; -- -0.05123106868100109
	pesos_i(2718) := b"1111111111111111_1111111111111111_1111110111011001_0000011000001011"; -- -0.008407232501609765
	pesos_i(2719) := b"0000000000000000_0000000000000000_0001010011001011_0000000000101100"; -- 0.0812225443250839
	pesos_i(2720) := b"0000000000000000_0000000000000000_0000100110010110_0110000100101101"; -- 0.0374508605822914
	pesos_i(2721) := b"1111111111111111_1111111111111111_1101111110101100_0000101101011001"; -- -0.12628106186158755
	pesos_i(2722) := b"0000000000000000_0000000000000000_0000011100110110_0001110100110000"; -- 0.02816946430838904
	pesos_i(2723) := b"1111111111111111_1111111111111111_1111010110110100_1100011111111011"; -- -0.04021024827074646
	pesos_i(2724) := b"0000000000000000_0000000000000000_0001000101110001_0011011110111010"; -- 0.06813381472249286
	pesos_i(2725) := b"1111111111111111_1111111111111111_1111000011111110_0100101011101101"; -- -0.05861980172333743
	pesos_i(2726) := b"0000000000000000_0000000000000000_0000011010001010_0110111000101001"; -- 0.025549778983931747
	pesos_i(2727) := b"0000000000000000_0000000000000000_0010101000110011_0110010010101111"; -- 0.16484669945368802
	pesos_i(2728) := b"1111111111111111_1111111111111111_1111100000011110_0111011001110011"; -- -0.030785176184134413
	pesos_i(2729) := b"0000000000000000_0000000000000000_0001011010100001_0110100000101111"; -- 0.08840037487001821
	pesos_i(2730) := b"0000000000000000_0000000000000000_0001100110000110_0000010111110110"; -- 0.09970128296089062
	pesos_i(2731) := b"0000000000000000_0000000000000000_0001110101101000_1110001000111010"; -- 0.11488164828521269
	pesos_i(2732) := b"0000000000000000_0000000000000000_0001111111111101_1001001100011110"; -- 0.12496299250678394
	pesos_i(2733) := b"0000000000000000_0000000000000000_0010000011011100_1011110000000110"; -- 0.12836814064389976
	pesos_i(2734) := b"1111111111111111_1111111111111111_1101010001011101_0011100111101000"; -- -0.1704524812277325
	pesos_i(2735) := b"0000000000000000_0000000000000000_0000101000110011_1111111001000110"; -- 0.03985585418088363
	pesos_i(2736) := b"0000000000000000_0000000000000000_0010011011100001_0111111101001101"; -- 0.15187831519951178
	pesos_i(2737) := b"1111111111111111_1111111111111111_1110000111011110_1101010110100000"; -- -0.11769356571773015
	pesos_i(2738) := b"0000000000000000_0000000000000000_0001110011100010_0011101011010101"; -- 0.11282699302923074
	pesos_i(2739) := b"0000000000000000_0000000000000000_0000010100010110_0100110110010001"; -- 0.019871566671223678
	pesos_i(2740) := b"1111111111111111_1111111111111111_1110100000011000_1010110101101010"; -- -0.0933734528669517
	pesos_i(2741) := b"0000000000000000_0000000000000000_0001010001111100_1010001111001110"; -- 0.08002685346287502
	pesos_i(2742) := b"0000000000000000_0000000000000000_0010100111101001_0100100101011001"; -- 0.16371591964654825
	pesos_i(2743) := b"1111111111111111_1111111111111111_1101001001011110_1000010101000000"; -- -0.17824523156750563
	pesos_i(2744) := b"0000000000000000_0000000000000000_0000001101000011_0101010000110010"; -- 0.012746107389884648
	pesos_i(2745) := b"1111111111111111_1111111111111111_1100101010010001_1000100110010000"; -- -0.20871677631951258
	pesos_i(2746) := b"1111111111111111_1111111111111111_1110110101000111_1110011100001011"; -- -0.07312160472532377
	pesos_i(2747) := b"0000000000000000_0000000000000000_0001001101011000_0101000000111100"; -- 0.07556630572067598
	pesos_i(2748) := b"1111111111111111_1111111111111111_1101101101010110_1000011011111010"; -- -0.14321094888577107
	pesos_i(2749) := b"1111111111111111_1111111111111111_1111001100010100_1011001010010111"; -- -0.0504654294120877
	pesos_i(2750) := b"0000000000000000_0000000000000000_0000110001111011_0110110000011001"; -- 0.04875827414652032
	pesos_i(2751) := b"1111111111111111_1111111111111111_1111110101000100_1011011100100100"; -- -0.010670236244934307
	pesos_i(2752) := b"1111111111111111_1111111111111111_1111110001100010_1011101111111111"; -- -0.014118433212804059
	pesos_i(2753) := b"1111111111111111_1111111111111111_1101010101111110_0011111001110011"; -- -0.16604242038547037
	pesos_i(2754) := b"0000000000000000_0000000000000000_0000010000111100_0111100101011100"; -- 0.016547760996702698
	pesos_i(2755) := b"1111111111111111_1111111111111111_1110111111000001_1101110010000001"; -- -0.06344816062425399
	pesos_i(2756) := b"0000000000000000_0000000000000000_0010101010011011_1000110100100111"; -- 0.16643602554318712
	pesos_i(2757) := b"1111111111111111_1111111111111111_1101101101110001_1100011101011111"; -- -0.14279512332147812
	pesos_i(2758) := b"1111111111111111_1111111111111111_1100111011001010_1110110111011001"; -- -0.1922160477510198
	pesos_i(2759) := b"1111111111111111_1111111111111111_1101111001010011_0111110101101010"; -- -0.13153854525937178
	pesos_i(2760) := b"1111111111111111_1111111111111111_1100111011000001_1101111010000011"; -- -0.19235429102307944
	pesos_i(2761) := b"0000000000000000_0000000000000000_0010001111011101_1011011000011111"; -- 0.1401017975953913
	pesos_i(2762) := b"0000000000000000_0000000000000000_0010101011000000_0110011100100111"; -- 0.1669983359597894
	pesos_i(2763) := b"1111111111111111_1111111111111111_1110000101101011_1000010111110000"; -- -0.11945307619227666
	pesos_i(2764) := b"0000000000000000_0000000000000000_0001110000110011_0110100110010001"; -- 0.11015949054403792
	pesos_i(2765) := b"0000000000000000_0000000000000000_0001001011101011_1101001100111101"; -- 0.07391090619957447
	pesos_i(2766) := b"0000000000000000_0000000000000000_0010000100001011_1101100001101001"; -- 0.12908699578171529
	pesos_i(2767) := b"0000000000000000_0000000000000000_0000001111111011_0011000101111110"; -- 0.01555165595620218
	pesos_i(2768) := b"0000000000000000_0000000000000000_0010010011101000_0001001000100100"; -- 0.1441661202718329
	pesos_i(2769) := b"1111111111111111_1111111111111111_1101001001010001_1101010101101001"; -- -0.1784388178650825
	pesos_i(2770) := b"0000000000000000_0000000000000000_0000100010001101_1000111011000011"; -- 0.0334099984313637
	pesos_i(2771) := b"0000000000000000_0000000000000000_0001110010111111_1011001011000100"; -- 0.11230008390452763
	pesos_i(2772) := b"0000000000000000_0000000000000000_0000011111001110_0001110101111101"; -- 0.030488818094978838
	pesos_i(2773) := b"1111111111111111_1111111111111111_1101011100110111_1100010100011000"; -- -0.15930526880766682
	pesos_i(2774) := b"0000000000000000_0000000000000000_0001000001111010_0011010101000101"; -- 0.06436474748286299
	pesos_i(2775) := b"0000000000000000_0000000000000000_0000001110101110_0111001000011000"; -- 0.014380579723976676
	pesos_i(2776) := b"0000000000000000_0000000000000000_0001110001110010_1010000101010101"; -- 0.11112411801633168
	pesos_i(2777) := b"1111111111111111_1111111111111111_1101101000001111_1101000100101001"; -- -0.1481961512349387
	pesos_i(2778) := b"1111111111111111_1111111111111111_1110011000000001_1100101000010110"; -- -0.10153519597290074
	pesos_i(2779) := b"0000000000000000_0000000000000000_0001101110001110_1000010001111110"; -- 0.10764339521924231
	pesos_i(2780) := b"0000000000000000_0000000000000000_0000100111111111_0110111110010010"; -- 0.039053891319067835
	pesos_i(2781) := b"0000000000000000_0000000000000000_0000101101010101_0001111000001010"; -- 0.044267537488325265
	pesos_i(2782) := b"1111111111111111_1111111111111111_1110110010001110_0010111111100100"; -- -0.07595539739526988
	pesos_i(2783) := b"1111111111111111_1111111111111111_1101100111010010_1100111110010101"; -- -0.14912703149716974
	pesos_i(2784) := b"0000000000000000_0000000000000000_0001110000101000_0110000101110110"; -- 0.10999116076274863
	pesos_i(2785) := b"0000000000000000_0000000000000000_0001111101010001_0010011111111111"; -- 0.12233209587010486
	pesos_i(2786) := b"0000000000000000_0000000000000000_0000001011111010_0010101111001010"; -- 0.01162980740990802
	pesos_i(2787) := b"0000000000000000_0000000000000000_0001001001101100_1010110010011100"; -- 0.07197073760462341
	pesos_i(2788) := b"0000000000000000_0000000000000000_0001011010011110_1111100001110100"; -- 0.08836319756187726
	pesos_i(2789) := b"1111111111111111_1111111111111111_1111011010100100_1100010001010110"; -- -0.03654835597511876
	pesos_i(2790) := b"1111111111111111_1111111111111111_1110000001111001_1010001011110001"; -- -0.12314397436839811
	pesos_i(2791) := b"0000000000000000_0000000000000000_0010001101111101_1110100111001011"; -- 0.13864003385150456
	pesos_i(2792) := b"0000000000000000_0000000000000000_0010001000011001_0001100100100010"; -- 0.13319546774521762
	pesos_i(2793) := b"1111111111111111_1111111111111111_1101110011111010_1011001001001110"; -- -0.1367996748701125
	pesos_i(2794) := b"0000000000000000_0000000000000000_0001011000111101_1100101111101111"; -- 0.0868804416384159
	pesos_i(2795) := b"0000000000000000_0000000000000000_0000101000001100_1010110000010010"; -- 0.039255861568854584
	pesos_i(2796) := b"1111111111111111_1111111111111111_1110011100111110_1110010011111100"; -- -0.0966965564408238
	pesos_i(2797) := b"1111111111111111_1111111111111111_1111110000000101_0010000100000110"; -- -0.015546737736999133
	pesos_i(2798) := b"1111111111111111_1111111111111111_1101100000101110_0110101100111000"; -- -0.15554170497776273
	pesos_i(2799) := b"1111111111111111_1111111111111111_1110110100111110_0111110011000010"; -- -0.07326526898885771
	pesos_i(2800) := b"0000000000000000_0000000000000000_0000010000000111_1110000100011000"; -- 0.01574522819377548
	pesos_i(2801) := b"1111111111111111_1111111111111111_1100111000111001_0110010101011011"; -- -0.19443670769794216
	pesos_i(2802) := b"0000000000000000_0000000000000000_0001001110000001_0100000100101011"; -- 0.07619101799866691
	pesos_i(2803) := b"0000000000000000_0000000000000000_0001000011111111_0011111111000011"; -- 0.0663947917939728
	pesos_i(2804) := b"1111111111111111_1111111111111111_1111101000101101_0001100110001101"; -- -0.02274933152634854
	pesos_i(2805) := b"1111111111111111_1111111111111111_1101101101100100_1111111110100110"; -- -0.14299013323783047
	pesos_i(2806) := b"1111111111111111_1111111111111111_1111101100001000_0111111101000110"; -- -0.019401593658753033
	pesos_i(2807) := b"0000000000000000_0000000000000000_0000000101010110_0010100110001001"; -- 0.005220981531506597
	pesos_i(2808) := b"1111111111111111_1111111111111111_1110001010010101_0101011111110000"; -- -0.11490869902168793
	pesos_i(2809) := b"0000000000000000_0000000000000000_0000100010100100_0001111011010110"; -- 0.03375427938094175
	pesos_i(2810) := b"1111111111111111_1111111111111111_1111000100000100_0001100111000101"; -- -0.05853117874489838
	pesos_i(2811) := b"0000000000000000_0000000000000000_0000001000011111_0101010010111100"; -- 0.008290573125275258
	pesos_i(2812) := b"1111111111111111_1111111111111111_1111001110001000_1001111101101011"; -- -0.04869655271185541
	pesos_i(2813) := b"1111111111111111_1111111111111111_1110010011101001_0011000111101011"; -- -0.10581672688378668
	pesos_i(2814) := b"1111111111111111_1111111111111111_1110011110001000_1100010100110100"; -- -0.09556930055860807
	pesos_i(2815) := b"0000000000000000_0000000000000000_0001010011001010_0101101011001110"; -- 0.08121268777080631
	pesos_i(2816) := b"0000000000000000_0000000000000000_0000010000010101_1000011011110101"; -- 0.01595347858554572
	pesos_i(2817) := b"0000000000000000_0000000000000000_0000100001011000_1111101001001100"; -- 0.03260769223121994
	pesos_i(2818) := b"1111111111111111_1111111111111111_1110111100011101_1110111001000010"; -- -0.06594954382395318
	pesos_i(2819) := b"1111111111111111_1111111111111111_1100110100101100_1000001000111110"; -- -0.19853960019985614
	pesos_i(2820) := b"0000000000000000_0000000000000000_0010101001010111_1111011110001110"; -- 0.1654047699759354
	pesos_i(2821) := b"1111111111111111_1111111111111111_1111000111010101_1111010100010100"; -- -0.055329020186333594
	pesos_i(2822) := b"0000000000000000_0000000000000000_0010000010000011_1011100111001111"; -- 0.12700997630746957
	pesos_i(2823) := b"1111111111111111_1111111111111111_1110001110011101_0100100001010110"; -- -0.11088130864223951
	pesos_i(2824) := b"1111111111111111_1111111111111111_1101101000010111_1000000000010000"; -- -0.14807891467452441
	pesos_i(2825) := b"0000000000000000_0000000000000000_0010101010000001_0000101001010000"; -- 0.16603149837008704
	pesos_i(2826) := b"1111111111111111_1111111111111111_1101101011010100_1111000001110000"; -- -0.14518830543620717
	pesos_i(2827) := b"0000000000000000_0000000000000000_0010000001010010_0101110010111100"; -- 0.12625674803392686
	pesos_i(2828) := b"0000000000000000_0000000000000000_0001101011100011_0101110010000010"; -- 0.1050317590448688
	pesos_i(2829) := b"1111111111111111_1111111111111111_1110101111000101_0111110001111110"; -- -0.07901784832339181
	pesos_i(2830) := b"1111111111111111_1111111111111111_1110111100111011_0100111000010010"; -- -0.06550132797919313
	pesos_i(2831) := b"0000000000000000_0000000000000000_0001111010010111_0101000011001110"; -- 0.1194963935634985
	pesos_i(2832) := b"0000000000000000_0000000000000000_0001001011101010_1101110100111000"; -- 0.07389624226257459
	pesos_i(2833) := b"0000000000000000_0000000000000000_0010101000100010_1001110111101001"; -- 0.16459071103564685
	pesos_i(2834) := b"1111111111111111_1111111111111111_1101000001001001_0001000100101100"; -- -0.18638508493857925
	pesos_i(2835) := b"0000000000000000_0000000000000000_0010001110100001_1101101111011001"; -- 0.13918851907710267
	pesos_i(2836) := b"1111111111111111_1111111111111111_1101011101111001_0000110001001111"; -- -0.15830920285621172
	pesos_i(2837) := b"0000000000000000_0000000000000000_0000111000001010_1101100011100101"; -- 0.05485301583637145
	pesos_i(2838) := b"0000000000000000_0000000000000000_0000111000001000_0101000001000111"; -- 0.05481435511675705
	pesos_i(2839) := b"0000000000000000_0000000000000000_0010011110010111_1110100111111110"; -- 0.15466177412312532
	pesos_i(2840) := b"1111111111111111_1111111111111111_1101011111101100_1001110111011110"; -- -0.15654576626073602
	pesos_i(2841) := b"1111111111111111_1111111111111111_1101111101001001_1111000011010101"; -- -0.12777800374723028
	pesos_i(2842) := b"1111111111111111_1111111111111111_1111011111001101_1110011100000011"; -- -0.03201442883543196
	pesos_i(2843) := b"0000000000000000_0000000000000000_0000001000111010_0011010010111100"; -- 0.008700652994015309
	pesos_i(2844) := b"0000000000000000_0000000000000000_0011000011101111_0100100000000000"; -- 0.19115114201579353
	pesos_i(2845) := b"0000000000000000_0000000000000000_0010001110001100_0110000100000001"; -- 0.1388607623922345
	pesos_i(2846) := b"1111111111111111_1111111111111111_1110110000110110_1101100111001101"; -- -0.07728804352991998
	pesos_i(2847) := b"1111111111111111_1111111111111111_1101111111100000_1010001111010000"; -- -0.12547851719440484
	pesos_i(2848) := b"1111111111111111_1111111111111111_1110010111101000_1001110101010011"; -- -0.10191933378234297
	pesos_i(2849) := b"0000000000000000_0000000000000000_0001111001001010_1110100011100001"; -- 0.11833053094031552
	pesos_i(2850) := b"1111111111111111_1111111111111111_1101001010011101_0100110010010011"; -- -0.1772873058893956
	pesos_i(2851) := b"0000000000000000_0000000000000000_0000001011110011_1100011110000000"; -- 0.011532276839623538
	pesos_i(2852) := b"0000000000000000_0000000000000000_0000001001010001_0100111111011100"; -- 0.009053221996426318
	pesos_i(2853) := b"0000000000000000_0000000000000000_0001010000011010_1001100110011000"; -- 0.07853088352552036
	pesos_i(2854) := b"1111111111111111_1111111111111111_1101100000011001_0001010010111110"; -- -0.15586729401864682
	pesos_i(2855) := b"1111111111111111_1111111111111111_1101000101001100_1100010000010001"; -- -0.18242239560607904
	pesos_i(2856) := b"0000000000000000_0000000000000000_0011001100100001_1101011100110100"; -- 0.1997351171346083
	pesos_i(2857) := b"0000000000000000_0000000000000000_0001011000111110_0111010010000100"; -- 0.0868904898594282
	pesos_i(2858) := b"1111111111111111_1111111111111111_1101011001010000_1000111101001100"; -- -0.16283325583146227
	pesos_i(2859) := b"0000000000000000_0000000000000000_0001100001001111_1100111101010010"; -- 0.09496780167158947
	pesos_i(2860) := b"1111111111111111_1111111111111111_1111011111000001_0001110010001000"; -- -0.03220960304075484
	pesos_i(2861) := b"0000000000000000_0000000000000000_0001101101101101_0110110100000011"; -- 0.10713845558526401
	pesos_i(2862) := b"0000000000000000_0000000000000000_0000001000100100_0010100001010101"; -- 0.008364220466048098
	pesos_i(2863) := b"0000000000000000_0000000000000000_0001011010000101_0001101110110010"; -- 0.0879685697105261
	pesos_i(2864) := b"0000000000000000_0000000000000000_0000001110000010_1000111010101111"; -- 0.01371089711668777
	pesos_i(2865) := b"1111111111111111_1111111111111111_1110100101001010_0101111000000100"; -- -0.08870899594582383
	pesos_i(2866) := b"0000000000000000_0000000000000000_0000111111100100_0110001110111010"; -- 0.06207869811537149
	pesos_i(2867) := b"0000000000000000_0000000000000000_0001000110011111_0000110000101000"; -- 0.06883312201093074
	pesos_i(2868) := b"0000000000000000_0000000000000000_0001010100000101_0111010000011110"; -- 0.08211446506987152
	pesos_i(2869) := b"0000000000000000_0000000000000000_0010001100001111_1100101111100000"; -- 0.13695978374317583
	pesos_i(2870) := b"1111111111111111_1111111111111111_1101110000001010_1111001100110101"; -- -0.14045791585414252
	pesos_i(2871) := b"1111111111111111_1111111111111111_1110011110001001_1001110000111111"; -- -0.09555648282411255
	pesos_i(2872) := b"1111111111111111_1111111111111111_1110011110101000_1000011001101000"; -- -0.09508476222387187
	pesos_i(2873) := b"1111111111111111_1111111111111111_1111111110011001_0000000011111010"; -- -0.0015715971806798236
	pesos_i(2874) := b"1111111111111111_1111111111111111_1100111110111001_1011000001110001"; -- -0.18857285726383471
	pesos_i(2875) := b"0000000000000000_0000000000000000_0001001001101110_0001011110101001"; -- 0.07199237698299911
	pesos_i(2876) := b"1111111111111111_1111111111111111_1101110010110010_1011100000101111"; -- -0.1378979572398379
	pesos_i(2877) := b"0000000000000000_0000000000000000_0011000011010000_0101000101010010"; -- 0.19067867520608908
	pesos_i(2878) := b"1111111111111111_1111111111111111_1110010001101001_0001110000101001"; -- -0.10777114873241969
	pesos_i(2879) := b"1111111111111111_1111111111111111_1110100101001101_1101011111101101"; -- -0.08865595297948108
	pesos_i(2880) := b"0000000000000000_0000000000000000_0001011000100001_0010101101110010"; -- 0.08644362950650447
	pesos_i(2881) := b"1111111111111111_1111111111111111_1111110000000110_1101101101101111"; -- -0.015520368031525423
	pesos_i(2882) := b"1111111111111111_1111111111111111_1101111110000100_1011100100000100"; -- -0.12688106209096495
	pesos_i(2883) := b"0000000000000000_0000000000000000_0000100111010100_0010101110101110"; -- 0.03839371680640593
	pesos_i(2884) := b"0000000000000000_0000000000000000_0001111100000000_1100111111110011"; -- 0.12110614464012484
	pesos_i(2885) := b"0000000000000000_0000000000000000_0001101000011001_1101110101010100"; -- 0.10195716182465188
	pesos_i(2886) := b"0000000000000000_0000000000000000_0010000011100110_0111010111010111"; -- 0.12851654530336706
	pesos_i(2887) := b"1111111111111111_1111111111111111_1110101100011011_0110010100000000"; -- -0.0816132425366824
	pesos_i(2888) := b"0000000000000000_0000000000000000_0001001111011010_1111000100000100"; -- 0.07755953158675986
	pesos_i(2889) := b"1111111111111111_1111111111111111_1101011011110101_1010001111101100"; -- -0.16031432616998578
	pesos_i(2890) := b"1111111111111111_1111111111111111_1111101010011100_0000011001011010"; -- -0.021056750330346576
	pesos_i(2891) := b"0000000000000000_0000000000000000_0001000110111000_1110000101110010"; -- 0.06922730485206488
	pesos_i(2892) := b"1111111111111111_1111111111111111_1111101001110010_0001011110000111"; -- -0.02169659559277894
	pesos_i(2893) := b"1111111111111111_1111111111111111_1111110100011101_1101111110000111"; -- -0.011262921753519997
	pesos_i(2894) := b"0000000000000000_0000000000000000_0001010011100111_1101111110001011"; -- 0.08166310441169455
	pesos_i(2895) := b"1111111111111111_1111111111111111_1111111100101110_0101011101100011"; -- -0.003199137138057768
	pesos_i(2896) := b"0000000000000000_0000000000000000_0001110111100001_0100111101101110"; -- 0.11671921196819346
	pesos_i(2897) := b"1111111111111111_1111111111111111_1111111011001111_1010001010101000"; -- -0.004644235562102
	pesos_i(2898) := b"1111111111111111_1111111111111111_1101110000000000_0110101100011111"; -- -0.14061861501862366
	pesos_i(2899) := b"1111111111111111_1111111111111111_1111111101100010_1001010001010001"; -- -0.002402048245717196
	pesos_i(2900) := b"0000000000000000_0000000000000000_0010001011011110_1001011101001011"; -- 0.13620896900850993
	pesos_i(2901) := b"0000000000000000_0000000000000000_0000011001101110_1001100001110010"; -- 0.025125053167924988
	pesos_i(2902) := b"0000000000000000_0000000000000000_0010000111101101_1010010101000100"; -- 0.13253243352949903
	pesos_i(2903) := b"0000000000000000_0000000000000000_0001011101000111_0101100111011101"; -- 0.09093248035628178
	pesos_i(2904) := b"1111111111111111_1111111111111111_1110010000000010_0000001110010011"; -- -0.10934426934960909
	pesos_i(2905) := b"0000000000000000_0000000000000000_0010010001101101_1111100100001111"; -- 0.14230305305466684
	pesos_i(2906) := b"1111111111111111_1111111111111111_1111011110000110_1111110011111000"; -- -0.03309649424582166
	pesos_i(2907) := b"0000000000000000_0000000000000000_0001011000001001_1101111000000011"; -- 0.08608806214096876
	pesos_i(2908) := b"1111111111111111_1111111111111111_1110001100110011_1111001111001000"; -- -0.1124885212192743
	pesos_i(2909) := b"1111111111111111_1111111111111111_1110111001100111_1100001000000000"; -- -0.06872928150743877
	pesos_i(2910) := b"1111111111111111_1111111111111111_1111100100000111_1010001111000000"; -- -0.027227178239161157
	pesos_i(2911) := b"1111111111111111_1111111111111111_1101100000001101_1101000101001111"; -- -0.15603916006279023
	pesos_i(2912) := b"1111111111111111_1111111111111111_1100110100110100_0100001001100000"; -- -0.19842133667277548
	pesos_i(2913) := b"0000000000000000_0000000000000000_0000100101101010_0111111110110101"; -- 0.03678129349373149
	pesos_i(2914) := b"1111111111111111_1111111111111111_1100110011110100_0101100001010011"; -- -0.19939659100281285
	pesos_i(2915) := b"1111111111111111_1111111111111111_1111100111101010_1010100101111101"; -- -0.023763091071886167
	pesos_i(2916) := b"1111111111111111_1111111111111111_1110011110010011_1100000100000001"; -- -0.09540170398197298
	pesos_i(2917) := b"1111111111111111_1111111111111111_1111111000011010_0010100001011101"; -- -0.007413365533509655
	pesos_i(2918) := b"0000000000000000_0000000000000000_0010000001001110_0101000011001101"; -- 0.12619500168332906
	pesos_i(2919) := b"1111111111111111_1111111111111111_1101010100011100_0010000110110111"; -- -0.16753949442937688
	pesos_i(2920) := b"1111111111111111_1111111111111111_1111010011101010_0001010000111000"; -- -0.04330323831019604
	pesos_i(2921) := b"1111111111111111_1111111111111111_1110101111111011_1000100100001111"; -- -0.07819312471154817
	pesos_i(2922) := b"0000000000000000_0000000000000000_0001011010111100_0111100000101101"; -- 0.08881331528257247
	pesos_i(2923) := b"0000000000000000_0000000000000000_0000110100110010_1000011100010010"; -- 0.05155224026268538
	pesos_i(2924) := b"0000000000000000_0000000000000000_0000000001001110_1101111101101110"; -- 0.0012035031036125346
	pesos_i(2925) := b"1111111111111111_1111111111111111_1111000110011010_1000001011111111"; -- -0.05623608854532452
	pesos_i(2926) := b"0000000000000000_0000000000000000_0000010111100001_1000111000100100"; -- 0.022972949740547772
	pesos_i(2927) := b"0000000000000000_0000000000000000_0010010001000100_0100100110000011"; -- 0.14166697925636737
	pesos_i(2928) := b"1111111111111111_1111111111111111_1100101101101111_0010011001110001"; -- -0.20533523311352983
	pesos_i(2929) := b"1111111111111111_1111111111111111_1111111000101001_1001011000101110"; -- -0.007177938206262583
	pesos_i(2930) := b"1111111111111111_1111111111111111_1111111111110110_0010001001111110"; -- -0.00015053201163642713
	pesos_i(2931) := b"0000000000000000_0000000000000000_0010011011111100_0000001011001100"; -- 0.15228288162559236
	pesos_i(2932) := b"1111111111111111_1111111111111111_1110011010011111_0000111001110111"; -- -0.09913549031105823
	pesos_i(2933) := b"0000000000000000_0000000000000000_0000001000010110_0101010000010000"; -- 0.008153203969805472
	pesos_i(2934) := b"1111111111111111_1111111111111111_1101100000010101_0010010100001110"; -- -0.15592735682530617
	pesos_i(2935) := b"1111111111111111_1111111111111111_1111111110010101_0110000001101101"; -- -0.0016269429389217185
	pesos_i(2936) := b"0000000000000000_0000000000000000_0000011011011001_0000000000100100"; -- 0.02674866557148989
	pesos_i(2937) := b"1111111111111111_1111111111111111_1111100011011010_0001110101101001"; -- -0.027921830894079985
	pesos_i(2938) := b"1111111111111111_1111111111111111_1110011100100010_0111100100100110"; -- -0.09713023018104419
	pesos_i(2939) := b"0000000000000000_0000000000000000_0010001111101001_0000110101111010"; -- 0.14027485117106403
	pesos_i(2940) := b"0000000000000000_0000000000000000_0010000010001001_0110101010111110"; -- 0.1270968164777769
	pesos_i(2941) := b"1111111111111111_1111111111111111_1110000001011111_1011110100101101"; -- -0.12353913920898545
	pesos_i(2942) := b"1111111111111111_1111111111111111_1101101000111110_1001010100000011"; -- -0.1474825732435096
	pesos_i(2943) := b"0000000000000000_0000000000000000_0000010010110101_0100101100110011"; -- 0.018391322995801346
	pesos_i(2944) := b"0000000000000000_0000000000000000_0010010110001101_0100010111111111"; -- 0.14668691124941344
	pesos_i(2945) := b"1111111111111111_1111111111111111_1110100101001111_1010001101101101"; -- -0.08862856474445767
	pesos_i(2946) := b"0000000000000000_0000000000000000_0001110001101110_0101101001110110"; -- 0.11105885861423556
	pesos_i(2947) := b"1111111111111111_1111111111111111_1111010011001010_1011101111110010"; -- -0.04378152209323649
	pesos_i(2948) := b"0000000000000000_0000000000000000_0001101010000100_0100011011110111"; -- 0.10358088989873383
	pesos_i(2949) := b"0000000000000000_0000000000000000_0001011111000011_1110000100101001"; -- 0.09283263442891712
	pesos_i(2950) := b"1111111111111111_1111111111111111_1111010001010001_1110011000111101"; -- -0.045625314811700096
	pesos_i(2951) := b"1111111111111111_1111111111111111_1110111001111011_1100101001101000"; -- -0.06842360465549793
	pesos_i(2952) := b"1111111111111111_1111111111111111_1111100101000010_1001010100010101"; -- -0.026327784040332716
	pesos_i(2953) := b"0000000000000000_0000000000000000_0001101110001000_1010001000010100"; -- 0.10755360586565035
	pesos_i(2954) := b"0000000000000000_0000000000000000_0011000010001110_1010111111000110"; -- 0.1896772248971534
	pesos_i(2955) := b"0000000000000000_0000000000000000_0001011111000001_1100011010111110"; -- 0.09280054232740406
	pesos_i(2956) := b"1111111111111111_1111111111111111_1110110001010010_0111110110111000"; -- -0.07686628592511884
	pesos_i(2957) := b"0000000000000000_0000000000000000_0010001000111001_1100010000001011"; -- 0.13369393612752167
	pesos_i(2958) := b"0000000000000000_0000000000000000_0010001101010100_0001011011010010"; -- 0.13800184846206054
	pesos_i(2959) := b"1111111111111111_1111111111111111_1101110111010011_0010001010101000"; -- -0.13349707989066992
	pesos_i(2960) := b"1111111111111111_1111111111111111_1101101011110000_0011011101110001"; -- -0.14477208605912603
	pesos_i(2961) := b"1111111111111111_1111111111111111_1111000010001001_1110011010100000"; -- -0.060395799561461815
	pesos_i(2962) := b"0000000000000000_0000000000000000_0001001111011101_1100011011101111"; -- 0.0776027997108893
	pesos_i(2963) := b"0000000000000000_0000000000000000_0000101111001100_1001000111001100"; -- 0.04609023316231135
	pesos_i(2964) := b"1111111111111111_1111111111111111_1100111010111110_0000000100111100"; -- -0.19241325659738995
	pesos_i(2965) := b"1111111111111111_1111111111111111_1111111011001000_1001110110101111"; -- -0.004751343492751068
	pesos_i(2966) := b"1111111111111111_1111111111111111_1110111011100010_1110001000011101"; -- -0.06685053636666514
	pesos_i(2967) := b"0000000000000000_0000000000000000_0000111110100001_1011001011000101"; -- 0.061061070508014376
	pesos_i(2968) := b"1111111111111111_1111111111111111_1111110110100111_1000000001110010"; -- -0.009162876209146822
	pesos_i(2969) := b"1111111111111111_1111111111111111_1111101000000011_0011101011100111"; -- -0.023388212838793592
	pesos_i(2970) := b"0000000000000000_0000000000000000_0000001101001000_1111100000000111"; -- 0.012832166415202031
	pesos_i(2971) := b"0000000000000000_0000000000000000_0001000000010111_1100111001101011"; -- 0.06286325568026273
	pesos_i(2972) := b"0000000000000000_0000000000000000_0010000001110010_0011001111011101"; -- 0.1267425933149827
	pesos_i(2973) := b"1111111111111111_1111111111111111_1111101001000000_0111110111001001"; -- -0.022453440170099672
	pesos_i(2974) := b"1111111111111111_1111111111111111_1101101010000101_0011110100011011"; -- -0.1464044389199879
	pesos_i(2975) := b"1111111111111111_1111111111111111_1110010000000011_0000111100101111"; -- -0.10932831871921164
	pesos_i(2976) := b"0000000000000000_0000000000000000_0001011111010111_1110110111111000"; -- 0.09313857361454042
	pesos_i(2977) := b"0000000000000000_0000000000000000_0000001001000111_1000010011000000"; -- 0.00890378645268014
	pesos_i(2978) := b"1111111111111111_1111111111111111_1101100011001101_0100001011011010"; -- -0.15311796346405918
	pesos_i(2979) := b"1111111111111111_1111111111111111_1101010101000010_0100001000101110"; -- -0.1669577251911105
	pesos_i(2980) := b"0000000000000000_0000000000000000_0010111011000110_0110100100110100"; -- 0.18271501082258565
	pesos_i(2981) := b"0000000000000000_0000000000000000_0000100010010111_0000000000100101"; -- 0.033554085836883345
	pesos_i(2982) := b"1111111111111111_1111111111111111_1100111100111001_0101101011001100"; -- -0.19053108707464814
	pesos_i(2983) := b"1111111111111111_1111111111111111_1101000010011100_0111011101100010"; -- -0.18511251309703247
	pesos_i(2984) := b"1111111111111111_1111111111111111_1101110101001011_0010001010001001"; -- -0.13557228226905457
	pesos_i(2985) := b"1111111111111111_1111111111111111_1110000101111101_0010100100010011"; -- -0.11918395308862582
	pesos_i(2986) := b"1111111111111111_1111111111111111_1110001100100101_1101100111101101"; -- -0.11270368534838507
	pesos_i(2987) := b"0000000000000000_0000000000000000_0000100010000000_1110101001101100"; -- 0.033217097604083194
	pesos_i(2988) := b"0000000000000000_0000000000000000_0010101011111011_1010101010110100"; -- 0.16790263081089754
	pesos_i(2989) := b"1111111111111111_1111111111111111_1101001101101001_1110111100001101"; -- -0.17416482867891236
	pesos_i(2990) := b"0000000000000000_0000000000000000_0010100000001100_0111010101000000"; -- 0.15644009421537716
	pesos_i(2991) := b"1111111111111111_1111111111111111_1111101011100100_1010001011111101"; -- -0.019948781242740965
	pesos_i(2992) := b"0000000000000000_0000000000000000_0010001101110011_1000100111110011"; -- 0.13848173305456266
	pesos_i(2993) := b"1111111111111111_1111111111111111_1110100110001110_1000001001110011"; -- -0.08766922651729059
	pesos_i(2994) := b"1111111111111111_1111111111111111_1101010101000011_1110010110110100"; -- -0.1669327198626351
	pesos_i(2995) := b"0000000000000000_0000000000000000_0000110001110100_0101000010001101"; -- 0.04864982081920885
	pesos_i(2996) := b"0000000000000000_0000000000000000_0001001110111011_0000010111001000"; -- 0.07707248821853324
	pesos_i(2997) := b"0000000000000000_0000000000000000_0010010111001100_1011010011000001"; -- 0.1476548167461194
	pesos_i(2998) := b"0000000000000000_0000000000000000_0001010111010001_0111000001101110"; -- 0.08522703820093007
	pesos_i(2999) := b"0000000000000000_0000000000000000_0000001011000000_1000101011000101"; -- 0.010750458788645658
	pesos_i(3000) := b"1111111111111111_1111111111111111_1110100010110001_1000101100011101"; -- -0.09104090244847768
	pesos_i(3001) := b"1111111111111111_1111111111111111_1110111000000010_1000110110101101"; -- -0.07027353796071303
	pesos_i(3002) := b"1111111111111111_1111111111111111_1110011111101101_1000000110001000"; -- -0.09403219624905179
	pesos_i(3003) := b"1111111111111111_1111111111111111_1101110101000011_1000101101001010"; -- -0.1356881087736303
	pesos_i(3004) := b"0000000000000000_0000000000000000_0000110111101001_0011101111110001"; -- 0.05434012060890517
	pesos_i(3005) := b"1111111111111111_1111111111111111_1111011110110100_0011001010011011"; -- -0.03240665155453403
	pesos_i(3006) := b"0000000000000000_0000000000000000_0000111011001010_0011110010111110"; -- 0.05777339579326889
	pesos_i(3007) := b"0000000000000000_0000000000000000_0001101001110111_1101000111111100"; -- 0.10339081205267346
	pesos_i(3008) := b"0000000000000000_0000000000000000_0000010100111010_1111011000010010"; -- 0.020430926770128883
	pesos_i(3009) := b"0000000000000000_0000000000000000_0001101110010010_0001000001101110"; -- 0.1076975124296193
	pesos_i(3010) := b"1111111111111111_1111111111111111_1101110010001111_0100011110101011"; -- -0.13843872148857797
	pesos_i(3011) := b"0000000000000000_0000000000000000_0000100000111001_1111111100010001"; -- 0.032134954015060474
	pesos_i(3012) := b"1111111111111111_1111111111111111_1101100111110011_1001110001000011"; -- -0.14862655025989593
	pesos_i(3013) := b"1111111111111111_1111111111111111_1101101101011110_1111101100110001"; -- -0.143081951604529
	pesos_i(3014) := b"1111111111111111_1111111111111111_1111101001001110_0001110011101101"; -- -0.022245590438736095
	pesos_i(3015) := b"1111111111111111_1111111111111111_1111001110101001_1110110110110011"; -- -0.048188346698679656
	pesos_i(3016) := b"0000000000000000_0000000000000000_0000001001010011_0110001011101100"; -- 0.009084875597741515
	pesos_i(3017) := b"1111111111111111_1111111111111111_1111011100110111_1010110011100100"; -- -0.03430671152067456
	pesos_i(3018) := b"1111111111111111_1111111111111111_1110011011011010_0001111011010101"; -- -0.09823424635760192
	pesos_i(3019) := b"1111111111111111_1111111111111111_1101000111111100_1011101000100101"; -- -0.17973744012771042
	pesos_i(3020) := b"0000000000000000_0000000000000000_0000111000011010_0010101010110001"; -- 0.055086773088752455
	pesos_i(3021) := b"0000000000000000_0000000000000000_0000000100111111_1001101010100011"; -- 0.004876770684409784
	pesos_i(3022) := b"1111111111111111_1111111111111111_1110110000110111_1000000010000110"; -- -0.0772781059050017
	pesos_i(3023) := b"1111111111111111_1111111111111111_1100100011100111_1010100001000110"; -- -0.2152151897869227
	pesos_i(3024) := b"1111111111111111_1111111111111111_1100110101101001_0110110011011100"; -- -0.1976100885984808
	pesos_i(3025) := b"0000000000000000_0000000000000000_0001001001001111_1010001001011011"; -- 0.07152762153165568
	pesos_i(3026) := b"1111111111111111_1111111111111111_1111111101100111_1010000000010111"; -- -0.0023250526555373342
	pesos_i(3027) := b"1111111111111111_1111111111111111_1110011101111100_0001011101010000"; -- -0.0957627706870017
	pesos_i(3028) := b"1111111111111111_1111111111111111_1100101111000110_1001100010000110"; -- -0.20400091866155726
	pesos_i(3029) := b"0000000000000000_0000000000000000_0010100110100100_0110100100011001"; -- 0.16266495566165562
	pesos_i(3030) := b"1111111111111111_1111111111111111_1110011111101101_1011111011000011"; -- -0.094028546684194
	pesos_i(3031) := b"0000000000000000_0000000000000000_0000110111111111_1010010110100010"; -- 0.054682113683158215
	pesos_i(3032) := b"1111111111111111_1111111111111111_1111000010101111_1111010011101100"; -- -0.05981511333511601
	pesos_i(3033) := b"1111111111111111_1111111111111111_1111000110101100_1111101110010100"; -- -0.05595424297401101
	pesos_i(3034) := b"1111111111111111_1111111111111111_1110000111110111_0011101000100101"; -- -0.117321363393707
	pesos_i(3035) := b"1111111111111111_1111111111111111_1110100111010001_0010010000000111"; -- -0.08665251564789717
	pesos_i(3036) := b"0000000000000000_0000000000000000_0001010000101101_0110000010111000"; -- 0.07881741049153242
	pesos_i(3037) := b"1111111111111111_1111111111111111_1111010111010100_1110101010010000"; -- -0.039719905621984464
	pesos_i(3038) := b"1111111111111111_1111111111111111_1110001110000010_1111110101100111"; -- -0.11128250358159919
	pesos_i(3039) := b"0000000000000000_0000000000000000_0010001010111101_0100100000010011"; -- 0.13570070713250584
	pesos_i(3040) := b"0000000000000000_0000000000000000_0001100001101100_0111011011000011"; -- 0.0954050278718722
	pesos_i(3041) := b"0000000000000000_0000000000000000_0001011010011110_0100111111001011"; -- 0.08835314472520428
	pesos_i(3042) := b"1111111111111111_1111111111111111_1111111101000111_0000100010110001"; -- -0.002822358037630285
	pesos_i(3043) := b"1111111111111111_1111111111111111_1111001111011111_1111010111101110"; -- -0.04736388154295762
	pesos_i(3044) := b"1111111111111111_1111111111111111_1101101100010010_0000000101001111"; -- -0.1442565138860796
	pesos_i(3045) := b"1111111111111111_1111111111111111_1111010110101011_0010000101001010"; -- -0.04035751284239821
	pesos_i(3046) := b"0000000000000000_0000000000000000_0001010011101010_0101001110100111"; -- 0.08170054262432247
	pesos_i(3047) := b"1111111111111111_1111111111111111_1110000011100000_1100111100011110"; -- -0.12156968605858759
	pesos_i(3048) := b"1111111111111111_1111111111111111_1110100000010011_1111011111111000"; -- -0.09344530284009331
	pesos_i(3049) := b"1111111111111111_1111111111111111_1111110111010001_0000111010001011"; -- -0.008528796173882462
	pesos_i(3050) := b"1111111111111111_1111111111111111_1110011001111000_1110100001011110"; -- -0.0997175951199468
	pesos_i(3051) := b"0000000000000000_0000000000000000_0001111000101111_0101100110011001"; -- 0.11791000352002255
	pesos_i(3052) := b"1111111111111111_1111111111111111_1111000000100111_1011100110100100"; -- -0.061893842296866945
	pesos_i(3053) := b"1111111111111111_1111111111111111_1110011101100101_1001001011110011"; -- -0.09610635345880222
	pesos_i(3054) := b"1111111111111111_1111111111111111_1111011111100101_1000010000110111"; -- -0.03165410666050925
	pesos_i(3055) := b"0000000000000000_0000000000000000_0001000111000110_1000011001110110"; -- 0.06943550466971819
	pesos_i(3056) := b"0000000000000000_0000000000000000_0001100101110101_1101111000101001"; -- 0.09945477017851065
	pesos_i(3057) := b"1111111111111111_1111111111111111_1111100100001101_0010100100000100"; -- -0.027142941020279147
	pesos_i(3058) := b"1111111111111111_1111111111111111_1110111001000111_1000100000100100"; -- -0.06922101135919767
	pesos_i(3059) := b"1111111111111111_1111111111111111_1111001010011101_1011110110110111"; -- -0.05228056221707408
	pesos_i(3060) := b"0000000000000000_0000000000000000_0000111011111000_1100101101010010"; -- 0.05848379841654759
	pesos_i(3061) := b"0000000000000000_0000000000000000_0000000011101000_0111110101111011"; -- 0.0035475182754967187
	pesos_i(3062) := b"0000000000000000_0000000000000000_0000001100011010_0111000111100000"; -- 0.012122266085014884
	pesos_i(3063) := b"0000000000000000_0000000000000000_0011011101001101_0110101000100010"; -- 0.2160250028294586
	pesos_i(3064) := b"0000000000000000_0000000000000000_0000100100110001_1111010011110001"; -- 0.03591853040910549
	pesos_i(3065) := b"0000000000000000_0000000000000000_0001000000000000_1110000111001110"; -- 0.06251345912285229
	pesos_i(3066) := b"0000000000000000_0000000000000000_0001101001010011_1011100100111011"; -- 0.10284002015315072
	pesos_i(3067) := b"1111111111111111_1111111111111111_1111111001111100_1110000110110000"; -- -0.005906958056715912
	pesos_i(3068) := b"0000000000000000_0000000000000000_0010000000001010_0110100111110101"; -- 0.12515890345384553
	pesos_i(3069) := b"0000000000000000_0000000000000000_0010111110001000_0000010000000101"; -- 0.18566918495760346
	pesos_i(3070) := b"1111111111111111_1111111111111111_1101110100111101_1100010110100100"; -- -0.1357761835758266
	pesos_i(3071) := b"0000000000000000_0000000000000000_0001100101001101_0111111000001000"; -- 0.0988386887907725
	pesos_i(3072) := b"1111111111111111_1111111111111111_1110000101111100_1111000001011010"; -- -0.11918733410734385
	pesos_i(3073) := b"1111111111111111_1111111111111111_1111100100101100_1111110001000101"; -- -0.02665732683686858
	pesos_i(3074) := b"0000000000000000_0000000000000000_0001101011101010_1101000110111000"; -- 0.10514555694211745
	pesos_i(3075) := b"1111111111111111_1111111111111111_1101100101100101_1110001100000110"; -- -0.15078908058656407
	pesos_i(3076) := b"0000000000000000_0000000000000000_0011010010110000_1111001100000011"; -- 0.20582503154366166
	pesos_i(3077) := b"0000000000000000_0000000000000000_0000011111011101_1100110110001110"; -- 0.030728194400195086
	pesos_i(3078) := b"1111111111111111_1111111111111111_1101010111011111_1010111100010010"; -- -0.1645556049252599
	pesos_i(3079) := b"1111111111111111_1111111111111111_1111010001101001_0001110101000101"; -- -0.04527108245293797
	pesos_i(3080) := b"1111111111111111_1111111111111111_1110100000111110_1111010011100010"; -- -0.09278935901017434
	pesos_i(3081) := b"0000000000000000_0000000000000000_0000111000110010_0001101010110010"; -- 0.05545203051864854
	pesos_i(3082) := b"0000000000000000_0000000000000000_0001000001000110_0110001100101100"; -- 0.06357402624768221
	pesos_i(3083) := b"1111111111111111_1111111111111111_1111110101101101_0111100100010110"; -- -0.01004832472013176
	pesos_i(3084) := b"0000000000000000_0000000000000000_0001001011101010_1001001010001011"; -- 0.07389179118396902
	pesos_i(3085) := b"1111111111111111_1111111111111111_1110111101011101_1110110010000100"; -- -0.06497308528398336
	pesos_i(3086) := b"1111111111111111_1111111111111111_1101111010011010_0000001110001000"; -- -0.13046243596332288
	pesos_i(3087) := b"0000000000000000_0000000000000000_0010000100010111_1100000111100111"; -- 0.1292687595937574
	pesos_i(3088) := b"1111111111111111_1111111111111111_1111111100011000_0000111101110001"; -- -0.0035391185856788413
	pesos_i(3089) := b"0000000000000000_0000000000000000_0000111100110000_0010101011101011"; -- 0.05932872988242293
	pesos_i(3090) := b"1111111111111111_1111111111111111_1101111110100100_0101100001010000"; -- -0.12639854483367383
	pesos_i(3091) := b"1111111111111111_1111111111111111_1111101111011000_0011100100011110"; -- -0.016231947144802694
	pesos_i(3092) := b"0000000000000000_0000000000000000_0001110111110101_1101000110011111"; -- 0.11703214776528152
	pesos_i(3093) := b"1111111111111111_1111111111111111_1110001101010110_1000011111010101"; -- -0.11196089784867352
	pesos_i(3094) := b"0000000000000000_0000000000000000_0000110111001010_1001111100110010"; -- 0.053873014268604746
	pesos_i(3095) := b"1111111111111111_1111111111111111_1110101111111001_0101101000010000"; -- -0.07822644327825805
	pesos_i(3096) := b"1111111111111111_1111111111111111_1110110100101001_0001011101101100"; -- -0.07359174359100429
	pesos_i(3097) := b"1111111111111111_1111111111111111_1101010001110101_1101011011000011"; -- -0.17007692084320675
	pesos_i(3098) := b"0000000000000000_0000000000000000_0001010010000001_0100000000101011"; -- 0.080097208452361
	pesos_i(3099) := b"1111111111111111_1111111111111111_1110100110110101_1110000101000100"; -- -0.08706848232312094
	pesos_i(3100) := b"0000000000000000_0000000000000000_0000001000001000_0000011100111011"; -- 0.007935001273025932
	pesos_i(3101) := b"0000000000000000_0000000000000000_0001000110111101_0101110001100110"; -- 0.06929566852500146
	pesos_i(3102) := b"0000000000000000_0000000000000000_0001100011010111_1011010010001110"; -- 0.0970414016196216
	pesos_i(3103) := b"1111111111111111_1111111111111111_1110011000110000_1101001000001010"; -- -0.10081755890127247
	pesos_i(3104) := b"0000000000000000_0000000000000000_0010011100010100_0010011010010001"; -- 0.15265122462239777
	pesos_i(3105) := b"1111111111111111_1111111111111111_1101100011001000_0100101011101111"; -- -0.15319377568123993
	pesos_i(3106) := b"1111111111111111_1111111111111111_1111110010101100_0100000000010110"; -- -0.012996668396032252
	pesos_i(3107) := b"0000000000000000_0000000000000000_0000110010011011_1000001001000110"; -- 0.049247877290259895
	pesos_i(3108) := b"0000000000000000_0000000000000000_0001100100111011_0000111010111010"; -- 0.0985573963011444
	pesos_i(3109) := b"0000000000000000_0000000000000000_0010001100100000_1001010100001101"; -- 0.13721591530630334
	pesos_i(3110) := b"1111111111111111_1111111111111111_1111000111100111_0101000001110110"; -- -0.05506417379884737
	pesos_i(3111) := b"0000000000000000_0000000000000000_0000001111111101_0101101011111101"; -- 0.01558464690470196
	pesos_i(3112) := b"1111111111111111_1111111111111111_1110011110110000_0000101001110011"; -- -0.09497008037516758
	pesos_i(3113) := b"0000000000000000_0000000000000000_0000101010010111_1101101100000010"; -- 0.04137963104717965
	pesos_i(3114) := b"1111111111111111_1111111111111111_1101001111110001_1001100010111111"; -- -0.17209477744922483
	pesos_i(3115) := b"1111111111111111_1111111111111111_1111100000101100_0101110011001001"; -- -0.030573082856652112
	pesos_i(3116) := b"0000000000000000_0000000000000000_0001010101111111_1100110001011001"; -- 0.08398129618209577
	pesos_i(3117) := b"0000000000000000_0000000000000000_0001011111110111_1010101111101001"; -- 0.09362291742796414
	pesos_i(3118) := b"1111111111111111_1111111111111111_1110111101001100_1101001111111011"; -- -0.06523394690576756
	pesos_i(3119) := b"0000000000000000_0000000000000000_0001110110111101_0111100001111001"; -- 0.1161723418381827
	pesos_i(3120) := b"1111111111111111_1111111111111111_1111111001100010_0001101011101110"; -- -0.006315533615220276
	pesos_i(3121) := b"0000000000000000_0000000000000000_0001100001011111_1100111011101001"; -- 0.09521191768034704
	pesos_i(3122) := b"0000000000000000_0000000000000000_0010011110011101_0001111011110111"; -- 0.15474122556344844
	pesos_i(3123) := b"0000000000000000_0000000000000000_0001100110110111_1010100111100100"; -- 0.1004587346229342
	pesos_i(3124) := b"1111111111111111_1111111111111111_1111111110110101_1101010101100111"; -- -0.0011316893027838448
	pesos_i(3125) := b"0000000000000000_0000000000000000_0001010011010100_1101011101010101"; -- 0.08137269801196823
	pesos_i(3126) := b"1111111111111111_1111111111111111_1111101011010100_0110100001101100"; -- -0.020196412590010454
	pesos_i(3127) := b"1111111111111111_1111111111111111_1101001100110001_1100111010001101"; -- -0.17502125786224576
	pesos_i(3128) := b"0000000000000000_0000000000000000_0000011100111100_0010100011110101"; -- 0.028261718574390693
	pesos_i(3129) := b"1111111111111111_1111111111111111_1111110000000101_0110000000010100"; -- -0.015542979453046502
	pesos_i(3130) := b"0000000000000000_0000000000000000_0010010100100010_1100101011100110"; -- 0.1450621424298441
	pesos_i(3131) := b"0000000000000000_0000000000000000_0010001101100011_1111111011100110"; -- 0.13824456313338113
	pesos_i(3132) := b"0000000000000000_0000000000000000_0000110110111101_1111101100000111"; -- 0.05368012348605666
	pesos_i(3133) := b"0000000000000000_0000000000000000_0010110100111100_0001011100000011"; -- 0.17669814898693892
	pesos_i(3134) := b"0000000000000000_0000000000000000_0001110010000110_1110110010101000"; -- 0.11143378349029276
	pesos_i(3135) := b"0000000000000000_0000000000000000_0001111110111101_1000110101011000"; -- 0.1239860858087597
	pesos_i(3136) := b"1111111111111111_1111111111111111_1111100100011001_1010100001001111"; -- -0.026952248291546382
	pesos_i(3137) := b"0000000000000000_0000000000000000_0010001010100100_1111001011000100"; -- 0.13532941130667325
	pesos_i(3138) := b"1111111111111111_1111111111111111_1110110110000111_0111010111001010"; -- -0.07215179274805933
	pesos_i(3139) := b"1111111111111111_1111111111111111_1111110110001000_0010100000110110"; -- -0.009641157882162327
	pesos_i(3140) := b"1111111111111111_1111111111111111_1111001111110101_0011110100111001"; -- -0.04703919763814629
	pesos_i(3141) := b"0000000000000000_0000000000000000_0010000010011100_1100001100111111"; -- 0.12739200869070533
	pesos_i(3142) := b"1111111111111111_1111111111111111_1110100101111100_1101100100001001"; -- -0.087938723816068
	pesos_i(3143) := b"0000000000000000_0000000000000000_0001011101011110_0010011011111101"; -- 0.0912804001328576
	pesos_i(3144) := b"1111111111111111_1111111111111111_1111001100110110_0111111100010001"; -- -0.04994970170354837
	pesos_i(3145) := b"0000000000000000_0000000000000000_0000100000111110_1001110111000000"; -- 0.032205447665053094
	pesos_i(3146) := b"1111111111111111_1111111111111111_1111010000010000_0100011011011110"; -- -0.04662663538104775
	pesos_i(3147) := b"0000000000000000_0000000000000000_0001011011110100_0101100001100000"; -- 0.08966591210901742
	pesos_i(3148) := b"1111111111111111_1111111111111111_1101001100011110_1011001010111001"; -- -0.17531283361749272
	pesos_i(3149) := b"1111111111111111_1111111111111111_1101101100001011_0000100110011111"; -- -0.14436282986036605
	pesos_i(3150) := b"1111111111111111_1111111111111111_1101001100101111_1101001001010010"; -- -0.17505155077826784
	pesos_i(3151) := b"1111111111111111_1111111111111111_1110111101001101_1111000110010111"; -- -0.06521692343754695
	pesos_i(3152) := b"0000000000000000_0000000000000000_0000000001110010_0010110101101111"; -- 0.0017422100862176937
	pesos_i(3153) := b"1111111111111111_1111111111111111_1101010010110010_0001010010110101"; -- -0.169157701244817
	pesos_i(3154) := b"0000000000000000_0000000000000000_0011000000000000_0010010010001010"; -- 0.18750217785015727
	pesos_i(3155) := b"1111111111111111_1111111111111111_1101011011100100_0110000010111100"; -- -0.16057773029136493
	pesos_i(3156) := b"1111111111111111_1111111111111111_1101110101110001_0011110001110010"; -- -0.13499090397914348
	pesos_i(3157) := b"1111111111111111_1111111111111111_1111111011101101_1000000101111000"; -- -0.004188449956780083
	pesos_i(3158) := b"1111111111111111_1111111111111111_1111100100001001_0101101010111010"; -- -0.027201013063964052
	pesos_i(3159) := b"1111111111111111_1111111111111111_1110010100100000_1010111010111000"; -- -0.10497005480939027
	pesos_i(3160) := b"0000000000000000_0000000000000000_0010110011010101_0101010001001010"; -- 0.1751301460802705
	pesos_i(3161) := b"0000000000000000_0000000000000000_0010100000100111_0011100010111110"; -- 0.15684847494928728
	pesos_i(3162) := b"1111111111111111_1111111111111111_1110011100010000_0110100110110111"; -- -0.09740580818192306
	pesos_i(3163) := b"1111111111111111_1111111111111111_1111101111001001_1110011001100101"; -- -0.016450500749311092
	pesos_i(3164) := b"0000000000000000_0000000000000000_0000111001001111_1000101000011011"; -- 0.055901176048224144
	pesos_i(3165) := b"0000000000000000_0000000000000000_0001100100100011_0111101010000111"; -- 0.09819761075309574
	pesos_i(3166) := b"1111111111111111_1111111111111111_1101001010111010_0011101000100011"; -- -0.17684589998907524
	pesos_i(3167) := b"0000000000000000_0000000000000000_0001000100011010_1111000101110100"; -- 0.06681737015352451
	pesos_i(3168) := b"1111111111111111_1111111111111111_1101011001101101_0000101110010010"; -- -0.16239860243018805
	pesos_i(3169) := b"1111111111111111_1111111111111111_1111010010110101_0101110000010100"; -- -0.04410767098099827
	pesos_i(3170) := b"1111111111111111_1111111111111111_1111000010010111_0100101111011000"; -- -0.06019140226390007
	pesos_i(3171) := b"0000000000000000_0000000000000000_0001100100101001_0000101011101001"; -- 0.0982825107515301
	pesos_i(3172) := b"1111111111111111_1111111111111111_1111011100000110_0000000010000111"; -- -0.03506466587733592
	pesos_i(3173) := b"1111111111111111_1111111111111111_1110111111001111_0111100000010111"; -- -0.06324052274715233
	pesos_i(3174) := b"0000000000000000_0000000000000000_0000000011010111_0100000000001111"; -- 0.0032844579105156257
	pesos_i(3175) := b"1111111111111111_1111111111111111_1111110010000001_0111011010110011"; -- -0.013649541180068225
	pesos_i(3176) := b"0000000000000000_0000000000000000_0001000110011011_0110100101100101"; -- 0.06877764435368855
	pesos_i(3177) := b"0000000000000000_0000000000000000_0001100010010101_1100111110001011"; -- 0.0960359300448671
	pesos_i(3178) := b"1111111111111111_1111111111111111_1111111111000001_0011010111010111"; -- -0.0009580945310152522
	pesos_i(3179) := b"0000000000000000_0000000000000000_0000100010011100_1010111101101100"; -- 0.0336408270235683
	pesos_i(3180) := b"0000000000000000_0000000000000000_0001011000001010_0110110111111100"; -- 0.0860966434020991
	pesos_i(3181) := b"1111111111111111_1111111111111111_1111101111010010_0001011001110001"; -- -0.01632556678494229
	pesos_i(3182) := b"1111111111111111_1111111111111111_1110100100011111_1100100001110111"; -- -0.089358778951373
	pesos_i(3183) := b"1111111111111111_1111111111111111_1110101100111001_1000011001010100"; -- -0.08115349249897343
	pesos_i(3184) := b"1111111111111111_1111111111111111_1111110011001011_1000101101000110"; -- -0.012519164498251911
	pesos_i(3185) := b"1111111111111111_1111111111111111_1110011101100110_0100010011000110"; -- -0.09609575433952375
	pesos_i(3186) := b"1111111111111111_1111111111111111_1111111011111111_0110111010001110"; -- -0.0039149191400768835
	pesos_i(3187) := b"0000000000000000_0000000000000000_0000010001010110_1000001101001100"; -- 0.016945081824626812
	pesos_i(3188) := b"0000000000000000_0000000000000000_0011000000110100_1010010000100000"; -- 0.18830323961309509
	pesos_i(3189) := b"1111111111111111_1111111111111111_1110000101000111_0000101111000001"; -- -0.12000967547506354
	pesos_i(3190) := b"0000000000000000_0000000000000000_0010011100010101_0101101001101101"; -- 0.15266957425950023
	pesos_i(3191) := b"1111111111111111_1111111111111111_1101010011100101_0101001100100100"; -- -0.168375781779599
	pesos_i(3192) := b"1111111111111111_1111111111111111_1110001010101110_0010111111110000"; -- -0.11452961335606208
	pesos_i(3193) := b"1111111111111111_1111111111111111_1101010101010001_0010101011111011"; -- -0.16673022621652514
	pesos_i(3194) := b"0000000000000000_0000000000000000_0010011000100000_0111001000101000"; -- 0.14893258541371895
	pesos_i(3195) := b"1111111111111111_1111111111111111_1101000010111110_0001001111110010"; -- -0.18459964127624814
	pesos_i(3196) := b"1111111111111111_1111111111111111_1110001101011111_0010010000101010"; -- -0.11182950954328402
	pesos_i(3197) := b"1111111111111111_1111111111111111_1111001100010010_1100000100110101"; -- -0.050495075688657826
	pesos_i(3198) := b"0000000000000000_0000000000000000_0000101111011000_1101110100111000"; -- 0.046277834030228365
	pesos_i(3199) := b"0000000000000000_0000000000000000_0010000011110010_1000100111110100"; -- 0.12870084960693168
	pesos_i(3200) := b"0000000000000000_0000000000000000_0001101001001011_1110100001010011"; -- 0.10272075680683285
	pesos_i(3201) := b"1111111111111111_1111111111111111_1101000001111101_0000101100001111"; -- -0.1855919922011502
	pesos_i(3202) := b"0000000000000000_0000000000000000_0000011110100010_1011111001010101"; -- 0.029827018551963375
	pesos_i(3203) := b"0000000000000000_0000000000000000_0001001111010000_0011111000101010"; -- 0.07739628342431953
	pesos_i(3204) := b"0000000000000000_0000000000000000_0001101110101100_1101011100110111"; -- 0.10810608949146117
	pesos_i(3205) := b"1111111111111111_1111111111111111_1110000100000001_1111011011101101"; -- -0.12106377332800183
	pesos_i(3206) := b"1111111111111111_1111111111111111_1101100110000111_1101101001111100"; -- -0.15027079072881036
	pesos_i(3207) := b"0000000000000000_0000000000000000_0010110001001001_1001111010011001"; -- 0.17299834483384924
	pesos_i(3208) := b"1111111111111111_1111111111111111_1110010100000100_0111101110100101"; -- -0.10540034496989426
	pesos_i(3209) := b"0000000000000000_0000000000000000_0000000110011111_0101101110010101"; -- 0.006337856099485978
	pesos_i(3210) := b"1111111111111111_1111111111111111_1101000001111011_0000111100100100"; -- -0.18562226649259778
	pesos_i(3211) := b"1111111111111111_1111111111111111_1111100010100001_1001001111111010"; -- -0.0287845149406028
	pesos_i(3212) := b"1111111111111111_1111111111111111_1111110101111100_1001001101010000"; -- -0.009817879615025504
	pesos_i(3213) := b"1111111111111111_1111111111111111_1110001001111101_1000100011111100"; -- -0.11527198637098607
	pesos_i(3214) := b"1111111111111111_1111111111111111_1111001101010000_0000011001000010"; -- -0.04956017395307283
	pesos_i(3215) := b"0000000000000000_0000000000000000_0001101011000110_1110101000000111"; -- 0.10459768939310399
	pesos_i(3216) := b"0000000000000000_0000000000000000_0000010010010100_0010000110000110"; -- 0.01788529886264459
	pesos_i(3217) := b"0000000000000000_0000000000000000_0000101000000111_0101001100000101"; -- 0.039174259825996344
	pesos_i(3218) := b"1111111111111111_1111111111111111_1110011011111010_0000101101110010"; -- -0.09774712057935725
	pesos_i(3219) := b"1111111111111111_1111111111111111_1110010010011010_1101100011100111"; -- -0.10701221798824423
	pesos_i(3220) := b"0000000000000000_0000000000000000_0001010010111100_0111111010100100"; -- 0.08100120071119188
	pesos_i(3221) := b"1111111111111111_1111111111111111_1110000100100010_1000000100100011"; -- -0.12056725408083142
	pesos_i(3222) := b"0000000000000000_0000000000000000_0010101100010110_0010100010101001"; -- 0.16830686690169
	pesos_i(3223) := b"1111111111111111_1111111111111111_1101000111100111_0000100100101000"; -- -0.18006842404465465
	pesos_i(3224) := b"0000000000000000_0000000000000000_0010000111001011_0001010010001010"; -- 0.1320050084416527
	pesos_i(3225) := b"1111111111111111_1111111111111111_1110100000101011_0001000111000001"; -- -0.09309281389633517
	pesos_i(3226) := b"1111111111111111_1111111111111111_1110011111001001_0111110001000010"; -- -0.09458182705217151
	pesos_i(3227) := b"0000000000000000_0000000000000000_0000011111101011_0101001010000111"; -- 0.030934484461651868
	pesos_i(3228) := b"0000000000000000_0000000000000000_0010001111100111_1110000010111111"; -- 0.14025692610281815
	pesos_i(3229) := b"0000000000000000_0000000000000000_0000011100110000_1000101110110010"; -- 0.028084498318643125
	pesos_i(3230) := b"1111111111111111_1111111111111111_1101000010000110_1111000101110111"; -- -0.1854409299468016
	pesos_i(3231) := b"1111111111111111_1111111111111111_1101100111011001_1110001101000111"; -- -0.14901904602473237
	pesos_i(3232) := b"1111111111111111_1111111111111111_1101110010001000_0100001110101100"; -- -0.13854577101835538
	pesos_i(3233) := b"1111111111111111_1111111111111111_1100111111010011_1111011011001111"; -- -0.18817193452383338
	pesos_i(3234) := b"0000000000000000_0000000000000000_0000101010011011_1011011110010100"; -- 0.04143855447044806
	pesos_i(3235) := b"0000000000000000_0000000000000000_0001100100100110_1010111100010110"; -- 0.09824651994966732
	pesos_i(3236) := b"0000000000000000_0000000000000000_0001111000000101_1000000000101011"; -- 0.11727143327754025
	pesos_i(3237) := b"1111111111111111_1111111111111111_1101110010101001_0010001110110110"; -- -0.13804413612933675
	pesos_i(3238) := b"0000000000000000_0000000000000000_0010111111100001_0000010111011010"; -- 0.1870273262505293
	pesos_i(3239) := b"1111111111111111_1111111111111111_1111000010111011_0110100101000110"; -- -0.05964033163949983
	pesos_i(3240) := b"0000000000000000_0000000000000000_0000011000000101_1010111110001100"; -- 0.02352425739871969
	pesos_i(3241) := b"1111111111111111_1111111111111111_1110110101110000_0111110101110101"; -- -0.07250228785565282
	pesos_i(3242) := b"1111111111111111_1111111111111111_1110001101110000_0011110110101100"; -- -0.11156858977701543
	pesos_i(3243) := b"1111111111111111_1111111111111111_1110110010011011_1000010001110110"; -- -0.07575199236154011
	pesos_i(3244) := b"1111111111111111_1111111111111111_1101000100011000_1100010110101000"; -- -0.18321575785199704
	pesos_i(3245) := b"1111111111111111_1111111111111111_1101101000111010_1110110010110011"; -- -0.14753838179991646
	pesos_i(3246) := b"1111111111111111_1111111111111111_1111111000011111_1110100101110011"; -- -0.007325562820416798
	pesos_i(3247) := b"1111111111111111_1111111111111111_1101110000011111_0110101000001010"; -- -0.14014565700843695
	pesos_i(3248) := b"1111111111111111_1111111111111111_1111000000100110_1110111111001101"; -- -0.061905872811453516
	pesos_i(3249) := b"1111111111111111_1111111111111111_1111111101011101_1110110010010010"; -- -0.002473082007371147
	pesos_i(3250) := b"0000000000000000_0000000000000000_0010001001110101_0101001000000011"; -- 0.13460266664253784
	pesos_i(3251) := b"1111111111111111_1111111111111111_1101101101101100_1100111001000110"; -- -0.14287100586345977
	pesos_i(3252) := b"1111111111111111_1111111111111111_1111011011001100_1000010111101101"; -- -0.035941724483311954
	pesos_i(3253) := b"0000000000000000_0000000000000000_0001010010011010_0110100011111101"; -- 0.08048111136540292
	pesos_i(3254) := b"1111111111111111_1111111111111111_1101101001000101_1001010110110110"; -- -0.14737572017426367
	pesos_i(3255) := b"1111111111111111_1111111111111111_1110100010101100_0101111110110100"; -- -0.09111978385952599
	pesos_i(3256) := b"1111111111111111_1111111111111111_1111011000110110_1111110100101001"; -- -0.03822343578223178
	pesos_i(3257) := b"1111111111111111_1111111111111111_1111000100000101_0111001110000000"; -- -0.058510571640065484
	pesos_i(3258) := b"0000000000000000_0000000000000000_0010001010100110_1001010110000101"; -- 0.1353543709849721
	pesos_i(3259) := b"0000000000000000_0000000000000000_0000101001101110_1010111110001101"; -- 0.040751430459447346
	pesos_i(3260) := b"1111111111111111_1111111111111111_1101100010100101_1000010001101011"; -- -0.15372440718884806
	pesos_i(3261) := b"1111111111111111_1111111111111111_1101100010101001_1100000100010101"; -- -0.15365975614865732
	pesos_i(3262) := b"0000000000000000_0000000000000000_0010101101000000_0011110101100110"; -- 0.168948972136436
	pesos_i(3263) := b"1111111111111111_1111111111111111_1111100011101000_0010111010011110"; -- -0.02770718223685706
	pesos_i(3264) := b"0000000000000000_0000000000000000_0000001011110111_0001100000001101"; -- 0.011582854439019102
	pesos_i(3265) := b"0000000000000000_0000000000000000_0010100101010000_0100001011101011"; -- 0.16138094165910521
	pesos_i(3266) := b"0000000000000000_0000000000000000_0001000001100010_1101101011000010"; -- 0.0640084002623576
	pesos_i(3267) := b"0000000000000000_0000000000000000_0010101100101010_1100011011110110"; -- 0.16862147803241967
	pesos_i(3268) := b"0000000000000000_0000000000000000_0001111100100101_0100101011010100"; -- 0.12166278527604063
	pesos_i(3269) := b"1111111111111111_1111111111111111_1101100100010001_0010010111000101"; -- -0.15208209936265898
	pesos_i(3270) := b"0000000000000000_0000000000000000_0000100010100110_1100010101010001"; -- 0.03379471984523599
	pesos_i(3271) := b"0000000000000000_0000000000000000_0010011010110110_1011100110100111"; -- 0.15122566541215826
	pesos_i(3272) := b"0000000000000000_0000000000000000_0000100000110111_0110011011000100"; -- 0.032095358810860036
	pesos_i(3273) := b"1111111111111111_1111111111111111_1110001001100000_1011001000001001"; -- -0.11571204442737103
	pesos_i(3274) := b"1111111111111111_1111111111111111_1101011001111010_0100100000101110"; -- -0.16219662560536366
	pesos_i(3275) := b"1111111111111111_1111111111111111_1110110000011000_1010111101000110"; -- -0.07774834196413402
	pesos_i(3276) := b"1111111111111111_1111111111111111_1110001000011000_0100001100000110"; -- -0.11681729417833334
	pesos_i(3277) := b"0000000000000000_0000000000000000_0010110111101101_0100101100100000"; -- 0.17940206082046006
	pesos_i(3278) := b"0000000000000000_0000000000000000_0010000101101101_0000001101101100"; -- 0.1305696619231661
	pesos_i(3279) := b"1111111111111111_1111111111111111_1111101101110001_0100000011110001"; -- -0.017803136114479423
	pesos_i(3280) := b"1111111111111111_1111111111111111_1111000110111010_1110111001110100"; -- -0.05574140236834446
	pesos_i(3281) := b"1111111111111111_1111111111111111_1101010111001010_0011001011001111"; -- -0.16488344617248862
	pesos_i(3282) := b"0000000000000000_0000000000000000_0000100010000100_1111110000000110"; -- 0.03327918187553633
	pesos_i(3283) := b"0000000000000000_0000000000000000_0010010001001000_1000011101110111"; -- 0.14173170704239563
	pesos_i(3284) := b"0000000000000000_0000000000000000_0010010000101011_1101001000111100"; -- 0.1412936588602139
	pesos_i(3285) := b"0000000000000000_0000000000000000_0010111000010010_0110000111001111"; -- 0.17996798799879404
	pesos_i(3286) := b"0000000000000000_0000000000000000_0010010110111001_1010010111010000"; -- 0.14736400920255183
	pesos_i(3287) := b"1111111111111111_1111111111111111_1101101010010000_1111000000100101"; -- -0.14622592062444678
	pesos_i(3288) := b"0000000000000000_0000000000000000_0010000101100101_0100100001000000"; -- 0.13045169418154912
	pesos_i(3289) := b"1111111111111111_1111111111111111_1110101011011111_1100101100000001"; -- -0.08252269005608343
	pesos_i(3290) := b"1111111111111111_1111111111111111_1110111100001000_0110111011010001"; -- -0.06627757457752213
	pesos_i(3291) := b"1111111111111111_1111111111111111_1111000110101011_0100101100011111"; -- -0.05598001940200917
	pesos_i(3292) := b"0000000000000000_0000000000000000_0010001010011010_0001001011111110"; -- 0.13516348548881196
	pesos_i(3293) := b"1111111111111111_1111111111111111_1110001001010001_0010001001010110"; -- -0.11594949148468126
	pesos_i(3294) := b"1111111111111111_1111111111111111_1111000011011111_1111001100100110"; -- -0.059082797216263444
	pesos_i(3295) := b"0000000000000000_0000000000000000_0001001100101111_1000110001111001"; -- 0.07494428594345282
	pesos_i(3296) := b"0000000000000000_0000000000000000_0001010011000000_1101110100000110"; -- 0.08106786163302843
	pesos_i(3297) := b"1111111111111111_1111111111111111_1101101010000010_1011100011100101"; -- -0.14644283684353449
	pesos_i(3298) := b"1111111111111111_1111111111111111_1110011111111110_0101111110000001"; -- -0.09377482519119691
	pesos_i(3299) := b"0000000000000000_0000000000000000_0001111110001010_1001001101101101"; -- 0.12320825017967285
	pesos_i(3300) := b"0000000000000000_0000000000000000_0000101011011010_1100010111000000"; -- 0.042400702815358016
	pesos_i(3301) := b"1111111111111111_1111111111111111_1110000111100101_0010000111000010"; -- -0.11759747524194052
	pesos_i(3302) := b"1111111111111111_1111111111111111_1110111010111111_1001011101100101"; -- -0.06738904738910115
	pesos_i(3303) := b"1111111111111111_1111111111111111_1110010101011111_0000000111011111"; -- -0.10401905360618684
	pesos_i(3304) := b"1111111111111111_1111111111111111_1111010001101000_0010001101010101"; -- -0.0452859800630424
	pesos_i(3305) := b"1111111111111111_1111111111111111_1111101111010010_1001100110010101"; -- -0.016317750185530645
	pesos_i(3306) := b"1111111111111111_1111111111111111_1110010110011101_1010110110110011"; -- -0.10306276681694228
	pesos_i(3307) := b"1111111111111111_1111111111111111_1110000000111110_1101111010001010"; -- -0.12404069060403995
	pesos_i(3308) := b"0000000000000000_0000000000000000_0000111101001111_1001101111001110"; -- 0.05980848094852901
	pesos_i(3309) := b"1111111111111111_1111111111111111_1111000001001010_1011011011101000"; -- -0.06135994764561588
	pesos_i(3310) := b"0000000000000000_0000000000000000_0000100000101111_1010010100111110"; -- 0.03197701233499085
	pesos_i(3311) := b"1111111111111111_1111111111111111_1111010101001000_1000101011010011"; -- -0.041861842642567815
	pesos_i(3312) := b"1111111111111111_1111111111111111_1101010110100010_1110000110001000"; -- -0.16548338356563222
	pesos_i(3313) := b"0000000000000000_0000000000000000_0010110001100111_1010111001001010"; -- 0.17345704382628413
	pesos_i(3314) := b"0000000000000000_0000000000000000_0000010010101001_1100111110011101"; -- 0.01821611005465727
	pesos_i(3315) := b"0000000000000000_0000000000000000_0010110011001111_0010111110111100"; -- 0.17503641451290664
	pesos_i(3316) := b"1111111111111111_1111111111111111_1110110100001101_1100110110111101"; -- -0.07400812275978866
	pesos_i(3317) := b"1111111111111111_1111111111111111_1110100100000001_0001001101010100"; -- -0.08982733922257206
	pesos_i(3318) := b"0000000000000000_0000000000000000_0000000110110110_0010100101111000"; -- 0.006685821324674202
	pesos_i(3319) := b"0000000000000000_0000000000000000_0001111111110010_1110101101101000"; -- 0.12480040827037588
	pesos_i(3320) := b"0000000000000000_0000000000000000_0001000011100100_0011001000101110"; -- 0.06598199482951453
	pesos_i(3321) := b"0000000000000000_0000000000000000_0000010110001100_1000000000111000"; -- 0.02167512281744032
	pesos_i(3322) := b"0000000000000000_0000000000000000_0000000010011100_1111010000010010"; -- 0.002394918889419395
	pesos_i(3323) := b"0000000000000000_0000000000000000_0000101100011001_1011110011110100"; -- 0.043361482154125296
	pesos_i(3324) := b"1111111111111111_1111111111111111_1110101101011100_0100000110101110"; -- -0.0806235265544107
	pesos_i(3325) := b"1111111111111111_1111111111111111_1100111011000101_0110011011110001"; -- -0.19230038269402697
	pesos_i(3326) := b"1111111111111111_1111111111111111_1110011101000110_1111001010011110"; -- -0.09657367358231865
	pesos_i(3327) := b"0000000000000000_0000000000000000_0000001101000111_1101101001110010"; -- 0.012815144274026108
	pesos_i(3328) := b"1111111111111111_1111111111111111_1110111100011110_1111010000111011"; -- -0.0659339289895544
	pesos_i(3329) := b"1111111111111111_1111111111111111_1101001010000111_1100000100101100"; -- -0.17761604964165192
	pesos_i(3330) := b"0000000000000000_0000000000000000_0000000100111100_1100001000000001"; -- 0.004833340865850296
	pesos_i(3331) := b"0000000000000000_0000000000000000_0001011010010100_0001110101000100"; -- 0.08819754516773866
	pesos_i(3332) := b"1111111111111111_1111111111111111_1101110110111000_0011001001000100"; -- -0.13390813665631587
	pesos_i(3333) := b"0000000000000000_0000000000000000_0000100111110101_0101011111110110"; -- 0.038899896159267804
	pesos_i(3334) := b"0000000000000000_0000000000000000_0010011000110100_0010111001101010"; -- 0.14923372356335915
	pesos_i(3335) := b"0000000000000000_0000000000000000_0001011010110111_1000100011011110"; -- 0.08873801630091632
	pesos_i(3336) := b"0000000000000000_0000000000000000_0000001001100110_1000110011111101"; -- 0.009377300153911283
	pesos_i(3337) := b"1111111111111111_1111111111111111_1111111111001101_1011000011101100"; -- -0.0007676529594972871
	pesos_i(3338) := b"1111111111111111_1111111111111111_1111000010100110_0111110010101101"; -- -0.05995960975320883
	pesos_i(3339) := b"1111111111111111_1111111111111111_1110100001111111_1101101110101101"; -- -0.09179904002317603
	pesos_i(3340) := b"0000000000000000_0000000000000000_0001000110111100_1011100000110010"; -- 0.06928588130216283
	pesos_i(3341) := b"0000000000000000_0000000000000000_0010010101011011_1011010111010111"; -- 0.14593063823050462
	pesos_i(3342) := b"1111111111111111_1111111111111111_1101111100100111_0110101111100101"; -- -0.12830472623333636
	pesos_i(3343) := b"1111111111111111_1111111111111111_1101101000001000_1101101011011110"; -- -0.14830238413369595
	pesos_i(3344) := b"1111111111111111_1111111111111111_1111111000011001_0101000000101010"; -- -0.007426252131610053
	pesos_i(3345) := b"0000000000000000_0000000000000000_0000011001001010_0000001001110101"; -- 0.024566796783148766
	pesos_i(3346) := b"0000000000000000_0000000000000000_0001111011001000_0000011111010000"; -- 0.12023972346263635
	pesos_i(3347) := b"0000000000000000_0000000000000000_0001111101110101_1011000011011000"; -- 0.12288956897043046
	pesos_i(3348) := b"0000000000000000_0000000000000000_0001110000111100_1000011010000100"; -- 0.11029854502506822
	pesos_i(3349) := b"0000000000000000_0000000000000000_0010011101011011_1101011000010001"; -- 0.1537450591588214
	pesos_i(3350) := b"0000000000000000_0000000000000000_0010111100110000_0100010011101100"; -- 0.18433027991542497
	pesos_i(3351) := b"0000000000000000_0000000000000000_0001100100000110_0010000101110001"; -- 0.0977497960395562
	pesos_i(3352) := b"1111111111111111_1111111111111111_1111111100100110_0111001101100110"; -- -0.0033195376458124946
	pesos_i(3353) := b"0000000000000000_0000000000000000_0010110001101001_0100010000000111"; -- 0.17348122753710016
	pesos_i(3354) := b"0000000000000000_0000000000000000_0000100100011010_0010100100010011"; -- 0.035555426653150785
	pesos_i(3355) := b"1111111111111111_1111111111111111_1111010111101110_0010100101101101"; -- -0.039334688955654264
	pesos_i(3356) := b"1111111111111111_1111111111111111_1110001000010000_1110111101100010"; -- -0.11692909102895775
	pesos_i(3357) := b"1111111111111111_1111111111111111_1110111001010111_1110001000001100"; -- -0.06897151190202842
	pesos_i(3358) := b"1111111111111111_1111111111111111_1111111000111000_0110011111000111"; -- -0.006951822093284992
	pesos_i(3359) := b"1111111111111111_1111111111111111_1110110100000000_0000100101101010"; -- -0.07421818880802823
	pesos_i(3360) := b"1111111111111111_1111111111111111_1101101101110101_0110001111010000"; -- -0.14274002237114783
	pesos_i(3361) := b"0000000000000000_0000000000000000_0011011100000111_0111111010011100"; -- 0.2149581079999505
	pesos_i(3362) := b"0000000000000000_0000000000000000_0001100111110100_1010111100000010"; -- 0.10138982571534756
	pesos_i(3363) := b"0000000000000000_0000000000000000_0010101000111100_1000000101110110"; -- 0.16498574385698117
	pesos_i(3364) := b"1111111111111111_1111111111111111_1101010101001011_1000101110111010"; -- -0.16681601235602095
	pesos_i(3365) := b"0000000000000000_0000000000000000_0011010011100100_0010010011101011"; -- 0.20660620449987946
	pesos_i(3366) := b"0000000000000000_0000000000000000_0000100001011100_1011110100011011"; -- 0.03266508005631935
	pesos_i(3367) := b"1111111111111111_1111111111111111_1110011100010010_0110011001000101"; -- -0.09737549617015691
	pesos_i(3368) := b"1111111111111111_1111111111111111_1111010100111010_0110000101111110"; -- -0.042077929178142466
	pesos_i(3369) := b"1111111111111111_1111111111111111_1111110101100000_1000001001011010"; -- -0.010246136791557593
	pesos_i(3370) := b"1111111111111111_1111111111111111_1101101011011011_1100110110000000"; -- -0.1450835764307962
	pesos_i(3371) := b"0000000000000000_0000000000000000_0000100110100101_1011111101101110"; -- 0.03768536029071435
	pesos_i(3372) := b"1111111111111111_1111111111111111_1110111110101001_0000011110110100"; -- -0.06382705541136562
	pesos_i(3373) := b"0000000000000000_0000000000000000_0010001000101100_1110100111011000"; -- 0.1334978249833165
	pesos_i(3374) := b"0000000000000000_0000000000000000_0001101011100010_1010110001000101"; -- 0.1050212543542035
	pesos_i(3375) := b"0000000000000000_0000000000000000_0011010010010000_0101111100001111"; -- 0.2053279316521809
	pesos_i(3376) := b"0000000000000000_0000000000000000_0000101111000100_1001001011011111"; -- 0.045968226764738954
	pesos_i(3377) := b"0000000000000000_0000000000000000_0011001110101011_0000101111100001"; -- 0.20182871088898094
	pesos_i(3378) := b"1111111111111111_1111111111111111_1110011101010101_1001011101100010"; -- -0.09635022979450215
	pesos_i(3379) := b"0000000000000000_0000000000000000_0000000100001101_0001101011001001"; -- 0.004106210875112187
	pesos_i(3380) := b"0000000000000000_0000000000000000_0000101000111101_0100010011001010"; -- 0.03999738634416884
	pesos_i(3381) := b"0000000000000000_0000000000000000_0000100000010101_1000101111000101"; -- 0.03157876548112654
	pesos_i(3382) := b"1111111111111111_1111111111111111_1100101001011100_0011110010010011"; -- -0.20953008081460764
	pesos_i(3383) := b"0000000000000000_0000000000000000_0000111110101111_0001111011000010"; -- 0.061265871414222725
	pesos_i(3384) := b"0000000000000000_0000000000000000_0000101010111000_1011100110111101"; -- 0.04188118814555177
	pesos_i(3385) := b"1111111111111111_1111111111111111_1111010011100110_0000101100001100"; -- -0.0433648200946446
	pesos_i(3386) := b"1111111111111111_1111111111111111_1101001000011001_1011000000000101"; -- -0.1792955386156467
	pesos_i(3387) := b"1111111111111111_1111111111111111_1111110100111111_1010110001111101"; -- -0.010747165273611518
	pesos_i(3388) := b"1111111111111111_1111111111111111_1110011101111010_1010010000000101"; -- -0.0957849013814513
	pesos_i(3389) := b"0000000000000000_0000000000000000_0001101101011010_1000100100011110"; -- 0.10685021391871935
	pesos_i(3390) := b"1111111111111111_1111111111111111_1101010101111000_0000100000110010"; -- -0.16613720683272645
	pesos_i(3391) := b"1111111111111111_1111111111111111_1111111011000010_1110010110011100"; -- -0.00483860923207349
	pesos_i(3392) := b"1111111111111111_1111111111111111_1111110101011100_0100010011010000"; -- -0.01031083987961907
	pesos_i(3393) := b"1111111111111111_1111111111111111_1110001000010000_0000101111010111"; -- -0.11694265366608002
	pesos_i(3394) := b"1111111111111111_1111111111111111_1111110010001000_1000000111010100"; -- -0.013542066356545812
	pesos_i(3395) := b"1111111111111111_1111111111111111_1111000001000011_1110000111010111"; -- -0.06146419998984728
	pesos_i(3396) := b"1111111111111111_1111111111111111_1101111010111101_1100101110011111"; -- -0.12991645216079234
	pesos_i(3397) := b"0000000000000000_0000000000000000_0000110000111110_1100011001110011"; -- 0.04783287339831732
	pesos_i(3398) := b"1111111111111111_1111111111111111_1111011100010000_1000111000011001"; -- -0.03490363978771352
	pesos_i(3399) := b"1111111111111111_1111111111111111_1111001111000100_0001110101101000"; -- -0.04778877463773726
	pesos_i(3400) := b"0000000000000000_0000000000000000_0000101111100011_1101100010001110"; -- 0.0464454027744629
	pesos_i(3401) := b"1111111111111111_1111111111111111_1110001011000110_0111000001100100"; -- -0.11415956076822391
	pesos_i(3402) := b"0000000000000000_0000000000000000_0000001000110010_1101111101001001"; -- 0.008588748269055277
	pesos_i(3403) := b"0000000000000000_0000000000000000_0010000111010001_0101100110101101"; -- 0.1321006820733249
	pesos_i(3404) := b"1111111111111111_1111111111111111_1111100001111110_0111001111001110"; -- -0.029320490027193304
	pesos_i(3405) := b"1111111111111111_1111111111111111_1110100100011110_0101000001001011"; -- -0.08938120043327799
	pesos_i(3406) := b"1111111111111111_1111111111111111_1101110011001010_0111001111111010"; -- -0.1375358117920989
	pesos_i(3407) := b"1111111111111111_1111111111111111_1110110000111101_1010000001000101"; -- -0.0771846610677057
	pesos_i(3408) := b"0000000000000000_0000000000000000_0001010101001010_0101111010101010"; -- 0.08316604276651424
	pesos_i(3409) := b"1111111111111111_1111111111111111_1111011101110011_0001101000011110"; -- -0.0333999325902543
	pesos_i(3410) := b"1111111111111111_1111111111111111_1101111100111000_1001000100000000"; -- -0.128043115146513
	pesos_i(3411) := b"1111111111111111_1111111111111111_1110100000001010_1100010000110100"; -- -0.09358571748513128
	pesos_i(3412) := b"1111111111111111_1111111111111111_1111001110001100_0010111011110111"; -- -0.048642220196499324
	pesos_i(3413) := b"0000000000000000_0000000000000000_0000000010100010_0011010011100101"; -- 0.002475076703011219
	pesos_i(3414) := b"1111111111111111_1111111111111111_1101011000010111_0100010100010101"; -- -0.163707430214229
	pesos_i(3415) := b"1111111111111111_1111111111111111_1111100111011110_0100000000000100"; -- -0.023952483113459946
	pesos_i(3416) := b"0000000000000000_0000000000000000_0000001110101000_0110100111010111"; -- 0.014288535180997526
	pesos_i(3417) := b"0000000000000000_0000000000000000_0010101100011011_1111111100100010"; -- 0.1683959443811298
	pesos_i(3418) := b"0000000000000000_0000000000000000_0001101101001100_0011011101001110"; -- 0.10663171431208342
	pesos_i(3419) := b"0000000000000000_0000000000000000_0010010110011011_1010110000111011"; -- 0.1469066279373098
	pesos_i(3420) := b"0000000000000000_0000000000000000_0001101010011110_1011110101001110"; -- 0.10398467208303121
	pesos_i(3421) := b"0000000000000000_0000000000000000_0000100101110010_1010001101001010"; -- 0.03690548467117264
	pesos_i(3422) := b"1111111111111111_1111111111111111_1111110011100011_1101010000010110"; -- -0.012148613536609426
	pesos_i(3423) := b"0000000000000000_0000000000000000_0000010000111001_0100100011001101"; -- 0.01649909026535501
	pesos_i(3424) := b"1111111111111111_1111111111111111_1101001011100101_0111111001001010"; -- -0.17618571000299035
	pesos_i(3425) := b"0000000000000000_0000000000000000_0000100100011101_0010001111001001"; -- 0.03560088790085628
	pesos_i(3426) := b"1111111111111111_1111111111111111_1111100001110010_0001101101110101"; -- -0.029508861369860417
	pesos_i(3427) := b"1111111111111111_1111111111111111_1111000110100001_0101011000110001"; -- -0.05613194745914039
	pesos_i(3428) := b"1111111111111111_1111111111111111_1110011001010111_1100100010111010"; -- -0.10022302116377278
	pesos_i(3429) := b"0000000000000000_0000000000000000_0010001110100101_0100000001100001"; -- 0.139240287417842
	pesos_i(3430) := b"0000000000000000_0000000000000000_0010001101000111_1101110001000101"; -- 0.13781525300902206
	pesos_i(3431) := b"1111111111111111_1111111111111111_1101010111101001_0110100000011010"; -- -0.16440724711866855
	pesos_i(3432) := b"1111111111111111_1111111111111111_1101010010101001_1010110001001100"; -- -0.16928599501910319
	pesos_i(3433) := b"0000000000000000_0000000000000000_0010100110111000_1110100110100010"; -- 0.1629777928202213
	pesos_i(3434) := b"1111111111111111_1111111111111111_1111110000000110_0000111100000111"; -- -0.015532551467055834
	pesos_i(3435) := b"0000000000000000_0000000000000000_0000000000010100_0011001101000001"; -- 0.0003082307128424847
	pesos_i(3436) := b"1111111111111111_1111111111111111_1101010111100110_0000000100011111"; -- -0.16445916160685572
	pesos_i(3437) := b"1111111111111111_1111111111111111_1110001101011000_0111111101100000"; -- -0.11193088432604066
	pesos_i(3438) := b"1111111111111111_1111111111111111_1111111001110001_0111011011000101"; -- -0.006081177542601919
	pesos_i(3439) := b"0000000000000000_0000000000000000_0001001001001010_0110101100011111"; -- 0.07144803521826684
	pesos_i(3440) := b"0000000000000000_0000000000000000_0001110111000000_0110101110010110"; -- 0.1162173500159347
	pesos_i(3441) := b"1111111111111111_1111111111111111_1101100100011000_0010100011110010"; -- -0.15197509860815006
	pesos_i(3442) := b"1111111111111111_1111111111111111_1101101010011110_0100011001101001"; -- -0.14602241444450909
	pesos_i(3443) := b"1111111111111111_1111111111111111_1100110010000000_0010101011011110"; -- -0.20116931995779694
	pesos_i(3444) := b"1111111111111111_1111111111111111_1110001111100110_0111101101111000"; -- -0.10976436913539289
	pesos_i(3445) := b"1111111111111111_1111111111111111_1110110101011011_1111000101000000"; -- -0.07281582050093631
	pesos_i(3446) := b"1111111111111111_1111111111111111_1111100010100101_0100001111011001"; -- -0.028728255673585577
	pesos_i(3447) := b"1111111111111111_1111111111111111_1110110101011101_0101110001110101"; -- -0.07279417165511969
	pesos_i(3448) := b"0000000000000000_0000000000000000_0001011101111111_0111101100001100"; -- 0.09178895047861019
	pesos_i(3449) := b"0000000000000000_0000000000000000_0001001111011111_1110101101010010"; -- 0.07763548605298282
	pesos_i(3450) := b"0000000000000000_0000000000000000_0011010001001100_0111011011010010"; -- 0.20429175028937446
	pesos_i(3451) := b"1111111111111111_1111111111111111_1100110110000010_0100000001111010"; -- -0.19723126422427242
	pesos_i(3452) := b"0000000000000000_0000000000000000_0011000110110101_0100110100101010"; -- 0.1941726902222552
	pesos_i(3453) := b"1111111111111111_1111111111111111_1111111110110100_1000010100001010"; -- -0.0011517382327283381
	pesos_i(3454) := b"1111111111111111_1111111111111111_1110011011001111_1010111100000010"; -- -0.09839349945881896
	pesos_i(3455) := b"1111111111111111_1111111111111111_1101101011010000_1100000100000101"; -- -0.1452521669919761
	pesos_i(3456) := b"0000000000000000_0000000000000000_0011100000011111_1100011011011001"; -- 0.21923487473816014
	pesos_i(3457) := b"0000000000000000_0000000000000000_0010001001011011_0101001011111001"; -- 0.13420599536983718
	pesos_i(3458) := b"1111111111111111_1111111111111111_1110100001000101_1100011100100100"; -- -0.09268527373255851
	pesos_i(3459) := b"0000000000000000_0000000000000000_0001110011000000_0100001001100100"; -- 0.11230864469767192
	pesos_i(3460) := b"0000000000000000_0000000000000000_0000000101011100_0100010101010011"; -- 0.00531419062472704
	pesos_i(3461) := b"0000000000000000_0000000000000000_0001000011101110_1000000101011111"; -- 0.06613930302989729
	pesos_i(3462) := b"1111111111111111_1111111111111111_1110101001111010_1010011000110001"; -- -0.08406602194266831
	pesos_i(3463) := b"1111111111111111_1111111111111111_1110110110010000_0101000111001101"; -- -0.07201660866904748
	pesos_i(3464) := b"1111111111111111_1111111111111111_1110110101001010_0010101100011110"; -- -0.07308702953900843
	pesos_i(3465) := b"1111111111111111_1111111111111111_1110100010011101_0111101010110111"; -- -0.09134705576699755
	pesos_i(3466) := b"0000000000000000_0000000000000000_0001010001101110_1010000100011010"; -- 0.07981306912586605
	pesos_i(3467) := b"1111111111111111_1111111111111111_1110111011110110_1101100100010101"; -- -0.06654589882631294
	pesos_i(3468) := b"0000000000000000_0000000000000000_0001111110000011_1011110100111101"; -- 0.12310393080786697
	pesos_i(3469) := b"1111111111111111_1111111111111111_1111000010110000_0010111111011000"; -- -0.05981160141408967
	pesos_i(3470) := b"0000000000000000_0000000000000000_0000010000100101_1000011000110011"; -- 0.016197574122402608
	pesos_i(3471) := b"0000000000000000_0000000000000000_0001101110011000_1100010011111110"; -- 0.10779982764010282
	pesos_i(3472) := b"0000000000000000_0000000000000000_0001001110010110_1110010111111101"; -- 0.07652127665493365
	pesos_i(3473) := b"1111111111111111_1111111111111111_1110000000010001_1010110010011100"; -- -0.12473031224096148
	pesos_i(3474) := b"0000000000000000_0000000000000000_0010011010011010_1101001010000100"; -- 0.15079990125620818
	pesos_i(3475) := b"0000000000000000_0000000000000000_0000110001111010_1100011100100010"; -- 0.04874844160994085
	pesos_i(3476) := b"1111111111111111_1111111111111111_1111100010011110_0110001111000100"; -- -0.028833164948174464
	pesos_i(3477) := b"0000000000000000_0000000000000000_0000100100111101_0010000000100011"; -- 0.03608895170736585
	pesos_i(3478) := b"1111111111111111_1111111111111111_1100111000111110_0011111000111011"; -- -0.19436274594272
	pesos_i(3479) := b"1111111111111111_1111111111111111_1111000100000011_1001111000000000"; -- -0.05853855602748089
	pesos_i(3480) := b"1111111111111111_1111111111111111_1111100001111001_1010101010010100"; -- -0.02939351930318758
	pesos_i(3481) := b"1111111111111111_1111111111111111_1101010111110100_1010000111100110"; -- -0.16423595558317733
	pesos_i(3482) := b"0000000000000000_0000000000000000_0010001101110110_1110001110011100"; -- 0.1385328536280414
	pesos_i(3483) := b"1111111111111111_1111111111111111_1111101111011001_1011001001111011"; -- -0.016209454570071048
	pesos_i(3484) := b"1111111111111111_1111111111111111_1111001011110100_0100001111001010"; -- -0.050960314975974835
	pesos_i(3485) := b"1111111111111111_1111111111111111_1111110101111010_1111100111100111"; -- -0.009842282469988554
	pesos_i(3486) := b"1111111111111111_1111111111111111_1111111101000011_0101101001001001"; -- -0.002878529778901932
	pesos_i(3487) := b"1111111111111111_1111111111111111_1111010011000101_1011111101101000"; -- -0.043857609795863964
	pesos_i(3488) := b"0000000000000000_0000000000000000_0001000111000001_1000110100001000"; -- 0.06935960246028369
	pesos_i(3489) := b"0000000000000000_0000000000000000_0001010101011000_1011111110011111"; -- 0.08338544495896093
	pesos_i(3490) := b"0000000000000000_0000000000000000_0000111010010000_0101111100000101"; -- 0.056890429146906125
	pesos_i(3491) := b"1111111111111111_1111111111111111_1110010110010001_0000100010110010"; -- -0.10325570740553247
	pesos_i(3492) := b"1111111111111111_1111111111111111_1110011011011111_1110100101000001"; -- -0.09814588705602967
	pesos_i(3493) := b"0000000000000000_0000000000000000_0001110010110000_0101100000000000"; -- 0.11206579209393693
	pesos_i(3494) := b"0000000000000000_0000000000000000_0000001011010011_0010110100111001"; -- 0.011034800034235653
	pesos_i(3495) := b"1111111111111111_1111111111111111_1101110111100010_0001101000110011"; -- -0.13326870202003285
	pesos_i(3496) := b"1111111111111111_1111111111111111_1110010111010100_0100011100100110"; -- -0.1022296458512943
	pesos_i(3497) := b"1111111111111111_1111111111111111_1110010011011000_1100001010000000"; -- -0.10606750850436851
	pesos_i(3498) := b"0000000000000000_0000000000000000_0001100000111111_0001101100110101"; -- 0.0947129254647969
	pesos_i(3499) := b"0000000000000000_0000000000000000_0001011000000110_0101010001101100"; -- 0.0860340845573271
	pesos_i(3500) := b"1111111111111111_1111111111111111_1110100110000100_1010100111010010"; -- -0.08781946786432046
	pesos_i(3501) := b"0000000000000000_0000000000000000_0001100111110000_1000111100101011"; -- 0.10132689275727326
	pesos_i(3502) := b"1111111111111111_1111111111111111_1110010100010001_1010010110100100"; -- -0.10519947758121433
	pesos_i(3503) := b"0000000000000000_0000000000000000_0010010001011010_1110111001011110"; -- 0.14201249887329198
	pesos_i(3504) := b"1111111111111111_1111111111111111_1101011001101101_1011100010011001"; -- -0.1623882891360663
	pesos_i(3505) := b"1111111111111111_1111111111111111_1111100000110011_0001000010010000"; -- -0.03047081455027229
	pesos_i(3506) := b"1111111111111111_1111111111111111_1111000001011000_1011111100001111"; -- -0.06114583864905227
	pesos_i(3507) := b"0000000000000000_0000000000000000_0001101000010000_0111011110110011"; -- 0.10181377529951442
	pesos_i(3508) := b"0000000000000000_0000000000000000_0010010000110101_1100111010001111"; -- 0.14144602777358553
	pesos_i(3509) := b"1111111111111111_1111111111111111_1110101010110100_0010001101101000"; -- -0.0831888076844928
	pesos_i(3510) := b"0000000000000000_0000000000000000_0001101011110111_0000010001110001"; -- 0.10533168563222109
	pesos_i(3511) := b"0000000000000000_0000000000000000_0001100011010110_1111110010101101"; -- 0.09703044154419893
	pesos_i(3512) := b"1111111111111111_1111111111111111_1110000000010010_1010000110001001"; -- -0.12471571356806627
	pesos_i(3513) := b"1111111111111111_1111111111111111_1110110111111011_0110111100001110"; -- -0.0703821746584517
	pesos_i(3514) := b"1111111111111111_1111111111111111_1111111010111100_1110110101101000"; -- -0.004929697191068113
	pesos_i(3515) := b"0000000000000000_0000000000000000_0000110001101001_1110100011110011"; -- 0.048491057630027416
	pesos_i(3516) := b"1111111111111111_1111111111111111_1110111010110010_0111011010100101"; -- -0.06758936383486489
	pesos_i(3517) := b"0000000000000000_0000000000000000_0010011110100010_0110101010010011"; -- 0.15482202621398877
	pesos_i(3518) := b"0000000000000000_0000000000000000_0010011100011111_0100100001100111"; -- 0.1528210879399091
	pesos_i(3519) := b"0000000000000000_0000000000000000_0000011001101101_0011100100101110"; -- 0.025104116178504672
	pesos_i(3520) := b"1111111111111111_1111111111111111_1101111100001111_0100011100001110"; -- -0.1286731329558849
	pesos_i(3521) := b"1111111111111111_1111111111111111_1101010100011000_0000001110101000"; -- -0.1676023210683052
	pesos_i(3522) := b"1111111111111111_1111111111111111_1111010111101110_0100101100000101"; -- -0.03933268672220966
	pesos_i(3523) := b"0000000000000000_0000000000000000_0010111001010011_1100010100011011"; -- 0.1809657278997008
	pesos_i(3524) := b"1111111111111111_1111111111111111_1111001111110110_0000101001101100"; -- -0.04702696662117074
	pesos_i(3525) := b"1111111111111111_1111111111111111_1101100001000111_1000010100111100"; -- -0.1551586846651718
	pesos_i(3526) := b"1111111111111111_1111111111111111_1111011101101011_0101100110000010"; -- -0.03351822449367355
	pesos_i(3527) := b"1111111111111111_1111111111111111_1111111110011010_1010000000001110"; -- -0.0015468563924446173
	pesos_i(3528) := b"0000000000000000_0000000000000000_0001010001010110_1010110110100001"; -- 0.07944760501319542
	pesos_i(3529) := b"1111111111111111_1111111111111111_1101101101011101_1101100001011111"; -- -0.14309928580569314
	pesos_i(3530) := b"0000000000000000_0000000000000000_0000000011000110_1101100101110101"; -- 0.0030342015678082885
	pesos_i(3531) := b"0000000000000000_0000000000000000_0010110010111001_0101110001001110"; -- 0.17470337783375298
	pesos_i(3532) := b"0000000000000000_0000000000000000_0010111001100101_0101100000110010"; -- 0.18123389449886035
	pesos_i(3533) := b"1111111111111111_1111111111111111_1111111000101101_1100010110010110"; -- -0.007114077530804067
	pesos_i(3534) := b"1111111111111111_1111111111111111_1110101100100110_0010010011100000"; -- -0.08144921813171015
	pesos_i(3535) := b"1111111111111111_1111111111111111_1111010000011101_1011110010010000"; -- -0.0464212559380333
	pesos_i(3536) := b"1111111111111111_1111111111111111_1111100111001101_0011111010000010"; -- -0.0242119724886451
	pesos_i(3537) := b"1111111111111111_1111111111111111_1110101101001101_0010001111010111"; -- -0.08085418706090863
	pesos_i(3538) := b"1111111111111111_1111111111111111_1111110000110100_1100000101101001"; -- -0.014820014854655983
	pesos_i(3539) := b"1111111111111111_1111111111111111_1111010000100000_0001011110101101"; -- -0.04638530752507927
	pesos_i(3540) := b"0000000000000000_0000000000000000_0010000001011111_1010111011100101"; -- 0.12646000941353489
	pesos_i(3541) := b"1111111111111111_1111111111111111_1101101011111100_1011001110111010"; -- -0.14458157266870322
	pesos_i(3542) := b"0000000000000000_0000000000000000_0010011101010010_1011101011010001"; -- 0.15360610591650325
	pesos_i(3543) := b"0000000000000000_0000000000000000_0001011111110010_0000110010111110"; -- 0.09353713648787622
	pesos_i(3544) := b"0000000000000000_0000000000000000_0001101011110111_0001111010000100"; -- 0.10533323969457123
	pesos_i(3545) := b"1111111111111111_1111111111111111_1111101011110111_0111110110011110"; -- -0.01966109179714031
	pesos_i(3546) := b"1111111111111111_1111111111111111_1101101101110011_0100110100000100"; -- -0.14277189885952968
	pesos_i(3547) := b"0000000000000000_0000000000000000_0001111101010001_1011101001111101"; -- 0.12234082759103039
	pesos_i(3548) := b"0000000000000000_0000000000000000_0000111000000001_1011001100010001"; -- 0.05471343199933659
	pesos_i(3549) := b"0000000000000000_0000000000000000_0001110011011011_1000010001110010"; -- 0.11272456913767168
	pesos_i(3550) := b"0000000000000000_0000000000000000_0000000100001100_0001100000000001"; -- 0.004090786214456345
	pesos_i(3551) := b"1111111111111111_1111111111111111_1101011010010001_1010111000101111"; -- -0.16183959345152266
	pesos_i(3552) := b"1111111111111111_1111111111111111_1101110001011110_1001010001110010"; -- -0.13918182582699543
	pesos_i(3553) := b"0000000000000000_0000000000000000_0000111100000101_1010111001100011"; -- 0.05868043810425908
	pesos_i(3554) := b"1111111111111111_1111111111111111_1110011001100111_0000010001010010"; -- -0.09999058714259705
	pesos_i(3555) := b"1111111111111111_1111111111111111_1110001000011010_1110111010100110"; -- -0.11677654683575041
	pesos_i(3556) := b"1111111111111111_1111111111111111_1110100101101001_1111111010011010"; -- -0.08822640163150988
	pesos_i(3557) := b"1111111111111111_1111111111111111_1101111001101000_1101100001110110"; -- -0.13121268388733695
	pesos_i(3558) := b"1111111111111111_1111111111111111_1111011101010110_1010010111010000"; -- -0.033834110942836046
	pesos_i(3559) := b"0000000000000000_0000000000000000_0000000010001010_1000111110011000"; -- 0.0021142717355516183
	pesos_i(3560) := b"1111111111111111_1111111111111111_1101110100100010_1100101110001000"; -- -0.13618781968562577
	pesos_i(3561) := b"1111111111111111_1111111111111111_1101101010100011_0000100011011011"; -- -0.1459497895012496
	pesos_i(3562) := b"0000000000000000_0000000000000000_0000101010111110_0101100010010100"; -- 0.041966949680957044
	pesos_i(3563) := b"0000000000000000_0000000000000000_0000000100001011_1100010100110001"; -- 0.004085850190826856
	pesos_i(3564) := b"1111111111111111_1111111111111111_1111110101011010_0000010111111110"; -- -0.010345101912571831
	pesos_i(3565) := b"1111111111111111_1111111111111111_1111010111010000_0010010100001011"; -- -0.03979271387966895
	pesos_i(3566) := b"1111111111111111_1111111111111111_1101001000101101_1001110011101110"; -- -0.17899150074936387
	pesos_i(3567) := b"0000000000000000_0000000000000000_0010110111100110_1000110010010101"; -- 0.17929915085802356
	pesos_i(3568) := b"0000000000000000_0000000000000000_0001111010011101_0100110010110101"; -- 0.11958770194710648
	pesos_i(3569) := b"0000000000000000_0000000000000000_0000011000100111_1101100110001011"; -- 0.024045559228608654
	pesos_i(3570) := b"0000000000000000_0000000000000000_0000110100011000_0000000010011010"; -- 0.051147496754867294
	pesos_i(3571) := b"1111111111111111_1111111111111111_1110110100010010_1001010001100001"; -- -0.07393524773264906
	pesos_i(3572) := b"0000000000000000_0000000000000000_0000101011110110_1010000110100011"; -- 0.0428257965081665
	pesos_i(3573) := b"0000000000000000_0000000000000000_0001101010001000_1101110000101011"; -- 0.10365081829233393
	pesos_i(3574) := b"0000000000000000_0000000000000000_0010000010000000_0110000011110100"; -- 0.12695890379432942
	pesos_i(3575) := b"1111111111111111_1111111111111111_1111001100111010_0110001010110111"; -- -0.04989035635346779
	pesos_i(3576) := b"0000000000000000_0000000000000000_0000101101000010_1100000001110101"; -- 0.04398730152155225
	pesos_i(3577) := b"0000000000000000_0000000000000000_0000001010100011_0101001000110001"; -- 0.01030458149875142
	pesos_i(3578) := b"0000000000000000_0000000000000000_0010000111111101_0101110110101110"; -- 0.13277230734119194
	pesos_i(3579) := b"0000000000000000_0000000000000000_0000111100111001_1001011001100000"; -- 0.05947246400059332
	pesos_i(3580) := b"1111111111111111_1111111111111111_1111011011000110_0001110001001101"; -- -0.036039572848820825
	pesos_i(3581) := b"0000000000000000_0000000000000000_0010000001011101_1100010000001100"; -- 0.1264307527382841
	pesos_i(3582) := b"1111111111111111_1111111111111111_1100101000100010_0110110001110001"; -- -0.21041223745882695
	pesos_i(3583) := b"0000000000000000_0000000000000000_0000010101011001_1100100000110000"; -- 0.02090121444671626
	pesos_i(3584) := b"1111111111111111_1111111111111111_1111001101110001_1101100101100110"; -- -0.04904404885750388
	pesos_i(3585) := b"1111111111111111_1111111111111111_1111111111101100_0000100001100101"; -- -0.00030467535656628173
	pesos_i(3586) := b"1111111111111111_1111111111111111_1101010101000110_1000100100101101"; -- -0.16689245838008002
	pesos_i(3587) := b"0000000000000000_0000000000000000_0000011110111111_0001101010010101"; -- 0.030259763152484343
	pesos_i(3588) := b"1111111111111111_1111111111111111_1111100000000011_1100010111001111"; -- -0.03119243324522975
	pesos_i(3589) := b"0000000000000000_0000000000000000_0010010011110111_1011100111011100"; -- 0.14440499898659
	pesos_i(3590) := b"1111111111111111_1111111111111111_1111111011110011_0011000011000010"; -- -0.00410170815811031
	pesos_i(3591) := b"0000000000000000_0000000000000000_0001101011110000_0101000011001011"; -- 0.1052294251213048
	pesos_i(3592) := b"0000000000000000_0000000000000000_0001011011100111_1000011011010101"; -- 0.08947031682930595
	pesos_i(3593) := b"0000000000000000_0000000000000000_0000100010101010_0001011011101000"; -- 0.033845359396559235
	pesos_i(3594) := b"1111111111111111_1111111111111111_1111110011100101_1001011111100001"; -- -0.01212168465939234
	pesos_i(3595) := b"0000000000000000_0000000000000000_0010001001101010_1111010110011110"; -- 0.13444457150967212
	pesos_i(3596) := b"1111111111111111_1111111111111111_1110111010010010_0110011110110011"; -- -0.06807853592694524
	pesos_i(3597) := b"1111111111111111_1111111111111111_1101010110010111_1001011111101000"; -- -0.16565561848694615
	pesos_i(3598) := b"0000000000000000_0000000000000000_0001010001010011_1010101001000101"; -- 0.0794016283634572
	pesos_i(3599) := b"1111111111111111_1111111111111111_1111011001101000_0011000000100010"; -- -0.03747271692253258
	pesos_i(3600) := b"1111111111111111_1111111111111111_1111101111110100_0001101011010001"; -- -0.015806507174590815
	pesos_i(3601) := b"1111111111111111_1111111111111111_1101000011001000_0000010001101111"; -- -0.18444797796921833
	pesos_i(3602) := b"0000000000000000_0000000000000000_0000111010011101_1011110000111001"; -- 0.05709434882902151
	pesos_i(3603) := b"1111111111111111_1111111111111111_1110011110101110_1010110111000111"; -- -0.09499086265485253
	pesos_i(3604) := b"1111111111111111_1111111111111111_1111011001100000_1010101111011111"; -- -0.03758741201729805
	pesos_i(3605) := b"0000000000000000_0000000000000000_0001100111011110_1110001101000011"; -- 0.10105724697293576
	pesos_i(3606) := b"1111111111111111_1111111111111111_1101111110110101_1100110101100010"; -- -0.1261321674431295
	pesos_i(3607) := b"1111111111111111_1111111111111111_1111101111001111_0000110010000001"; -- -0.016371935386708555
	pesos_i(3608) := b"0000000000000000_0000000000000000_0000000000011101_0011100001101001"; -- 0.0004458673063529026
	pesos_i(3609) := b"0000000000000000_0000000000000000_0000110100001101_1100011000000101"; -- 0.050991417252790584
	pesos_i(3610) := b"1111111111111111_1111111111111111_1101000111000101_1111001111001001"; -- -0.18057323779800424
	pesos_i(3611) := b"1111111111111111_1111111111111111_1101001100110000_0011110001001001"; -- -0.17504523485840284
	pesos_i(3612) := b"0000000000000000_0000000000000000_0010011110001101_0010000111001101"; -- 0.1544972538592703
	pesos_i(3613) := b"1111111111111111_1111111111111111_1110101011010101_0110000011101011"; -- -0.0826816012407704
	pesos_i(3614) := b"1111111111111111_1111111111111111_1111010110000010_1111111100111110"; -- -0.04096989370484214
	pesos_i(3615) := b"0000000000000000_0000000000000000_0010101011011111_0001001101100001"; -- 0.16746636514910374
	pesos_i(3616) := b"1111111111111111_1111111111111111_1111101101000101_1010000111100010"; -- -0.018468744648977835
	pesos_i(3617) := b"1111111111111111_1111111111111111_1110110111101111_0011001001001001"; -- -0.0705689021035829
	pesos_i(3618) := b"1111111111111111_1111111111111111_1110110111011111_0100100110110100"; -- -0.07081164699617555
	pesos_i(3619) := b"0000000000000000_0000000000000000_0000001000011001_0011010110101100"; -- 0.008197168858658415
	pesos_i(3620) := b"1111111111111111_1111111111111111_1101101010001000_1100001011110100"; -- -0.14635068451430555
	pesos_i(3621) := b"0000000000000000_0000000000000000_0010011011101101_0101101000010011"; -- 0.15205920195637126
	pesos_i(3622) := b"1111111111111111_1111111111111111_1101111101010101_1011111100100010"; -- -0.12759786052723926
	pesos_i(3623) := b"1111111111111111_1111111111111111_1101101001001110_0000001001100100"; -- -0.14724717198751158
	pesos_i(3624) := b"0000000000000000_0000000000000000_0001001001001100_0001010100110000"; -- 0.07147343075955807
	pesos_i(3625) := b"0000000000000000_0000000000000000_0000110001011110_0101000111100010"; -- 0.048314206719288044
	pesos_i(3626) := b"0000000000000000_0000000000000000_0001110001101001_0001110111110110"; -- 0.11097895868551327
	pesos_i(3627) := b"1111111111111111_1111111111111111_1110101011110111_0000000011101011"; -- -0.08216852449170282
	pesos_i(3628) := b"0000000000000000_0000000000000000_0000010101001101_0100011101000001"; -- 0.02071042381578597
	pesos_i(3629) := b"1111111111111111_1111111111111111_1111100010011110_1001101000010100"; -- -0.028829927472151635
	pesos_i(3630) := b"0000000000000000_0000000000000000_0000101100000110_0001111011011010"; -- 0.04306214167640674
	pesos_i(3631) := b"1111111111111111_1111111111111111_1111100011011001_1101010100101110"; -- -0.027926136359080995
	pesos_i(3632) := b"0000000000000000_0000000000000000_0000010110111110_0011010111010100"; -- 0.022433628425947108
	pesos_i(3633) := b"1111111111111111_1111111111111111_1110110111001000_1101011001001110"; -- -0.07115421856327701
	pesos_i(3634) := b"0000000000000000_0000000000000000_0010000001101101_1010101111011010"; -- 0.1266734510927807
	pesos_i(3635) := b"0000000000000000_0000000000000000_0000100111101111_0001000000000000"; -- 0.038804054178233585
	pesos_i(3636) := b"1111111111111111_1111111111111111_1101110001001101_1000011000011101"; -- -0.1394420795340578
	pesos_i(3637) := b"0000000000000000_0000000000000000_0000101000100110_1000001111011110"; -- 0.039650193937802156
	pesos_i(3638) := b"1111111111111111_1111111111111111_1110101010100100_1101101000000000"; -- -0.08342206481251685
	pesos_i(3639) := b"0000000000000000_0000000000000000_0001011000100010_1101100011101110"; -- 0.0864692289150526
	pesos_i(3640) := b"1111111111111111_1111111111111111_1110110110101001_1001100100010110"; -- -0.07163088990067856
	pesos_i(3641) := b"1111111111111111_1111111111111111_1101101110110110_1011100100011110"; -- -0.14174311659899227
	pesos_i(3642) := b"0000000000000000_0000000000000000_0000111010111101_1011110011010101"; -- 0.057582666429226714
	pesos_i(3643) := b"0000000000000000_0000000000000000_0000111100110111_1001001101101110"; -- 0.05944177094209063
	pesos_i(3644) := b"0000000000000000_0000000000000000_0001011110011101_0111001000000010"; -- 0.09224617521650869
	pesos_i(3645) := b"1111111111111111_1111111111111111_1111001011010011_0011001011101110"; -- -0.05146485990169354
	pesos_i(3646) := b"0000000000000000_0000000000000000_0001000111011000_1111101000010111"; -- 0.06971705494634944
	pesos_i(3647) := b"0000000000000000_0000000000000000_0010000010001011_0111111110011011"; -- 0.12712857746989598
	pesos_i(3648) := b"0000000000000000_0000000000000000_0000010110110001_1100111100000011"; -- 0.02224439446971757
	pesos_i(3649) := b"0000000000000000_0000000000000000_0000010001011111_1111000111110100"; -- 0.017089006383432345
	pesos_i(3650) := b"1111111111111111_1111111111111111_1111010100111111_1110010010010110"; -- -0.04199382147895063
	pesos_i(3651) := b"1111111111111111_1111111111111111_1110111000001111_1001111011010111"; -- -0.07007415054561551
	pesos_i(3652) := b"0000000000000000_0000000000000000_0000000110100100_0101101110110101"; -- 0.0064141576665490115
	pesos_i(3653) := b"1111111111111111_1111111111111111_1110101100111010_1011011111000101"; -- -0.08113528664740059
	pesos_i(3654) := b"1111111111111111_1111111111111111_1111000001000010_0000111110101001"; -- -0.06149198645563099
	pesos_i(3655) := b"0000000000000000_0000000000000000_0001101100011110_1001000010100110"; -- 0.10593513528035864
	pesos_i(3656) := b"0000000000000000_0000000000000000_0000010000010000_0001011111110100"; -- 0.01587056829341115
	pesos_i(3657) := b"1111111111111111_1111111111111111_1101111011110010_0000110110001111"; -- -0.12911906496924067
	pesos_i(3658) := b"1111111111111111_1111111111111111_1101000010001011_0010010001010111"; -- -0.185376862310842
	pesos_i(3659) := b"0000000000000000_0000000000000000_0001110100011111_0111000000011100"; -- 0.11376095464259953
	pesos_i(3660) := b"0000000000000000_0000000000000000_0001010000011011_1101101011100111"; -- 0.07855003497551434
	pesos_i(3661) := b"0000000000000000_0000000000000000_0000001010010101_0100110000111011"; -- 0.010090603312513971
	pesos_i(3662) := b"0000000000000000_0000000000000000_0000110100001001_1000110000110001"; -- 0.050926935047696756
	pesos_i(3663) := b"1111111111111111_1111111111111111_1101101100000100_0110001010110000"; -- -0.14446433267537548
	pesos_i(3664) := b"1111111111111111_1111111111111111_1110111011001010_0010010000110100"; -- -0.06722806662848833
	pesos_i(3665) := b"1111111111111111_1111111111111111_1101110111000010_0111011011110011"; -- -0.1337514549881362
	pesos_i(3666) := b"1111111111111111_1111111111111111_1101100000111000_1010100010110110"; -- -0.15538545191450065
	pesos_i(3667) := b"1111111111111111_1111111111111111_1110100000010000_1000110001110100"; -- -0.09349748780490177
	pesos_i(3668) := b"0000000000000000_0000000000000000_0010101000110100_0011000101000011"; -- 0.16485889315111993
	pesos_i(3669) := b"0000000000000000_0000000000000000_0000110010100010_0111111010100001"; -- 0.0493544714642472
	pesos_i(3670) := b"0000000000000000_0000000000000000_0010001111100001_1011111010000001"; -- 0.14016333236419481
	pesos_i(3671) := b"1111111111111111_1111111111111111_1110100100100010_0100110101010001"; -- -0.08932034277856278
	pesos_i(3672) := b"0000000000000000_0000000000000000_0010011011101110_0001001001010000"; -- 0.15207018334080674
	pesos_i(3673) := b"1111111111111111_1111111111111111_1110100000110000_1011110001101111"; -- -0.09300634656289247
	pesos_i(3674) := b"1111111111111111_1111111111111111_1101010010111001_1111001001010110"; -- -0.16903767965066974
	pesos_i(3675) := b"0000000000000000_0000000000000000_0000111100100000_0111101111101000"; -- 0.059089416700010076
	pesos_i(3676) := b"1111111111111111_1111111111111111_1111010000111011_0000011010010001"; -- -0.04597434016470644
	pesos_i(3677) := b"0000000000000000_0000000000000000_0011000011010011_0011011100010010"; -- 0.19072288690268735
	pesos_i(3678) := b"0000000000000000_0000000000000000_0000011001110100_0101010110011100"; -- 0.025212622241499574
	pesos_i(3679) := b"0000000000000000_0000000000000000_0000010000000001_0001110001000000"; -- 0.0156419426507992
	pesos_i(3680) := b"1111111111111111_1111111111111111_1110010101100001_1110110000000110"; -- -0.10397457935251549
	pesos_i(3681) := b"1111111111111111_1111111111111111_1101110110010000_0011100011110101"; -- -0.1345180895585957
	pesos_i(3682) := b"0000000000000000_0000000000000000_0000010001010001_1000111111111110"; -- 0.016869544620904342
	pesos_i(3683) := b"1111111111111111_1111111111111111_1111010111110011_1100111010101001"; -- -0.03924854624827644
	pesos_i(3684) := b"0000000000000000_0000000000000000_0001110010110011_1110101101001101"; -- 0.11212034825517084
	pesos_i(3685) := b"0000000000000000_0000000000000000_0010010010010010_1011100001100000"; -- 0.14286377274727066
	pesos_i(3686) := b"0000000000000000_0000000000000000_0001110010001101_0001111100100110"; -- 0.11152834574767347
	pesos_i(3687) := b"0000000000000000_0000000000000000_0010100010010101_1000110001000110"; -- 0.15853192041176264
	pesos_i(3688) := b"1111111111111111_1111111111111111_1110101011110101_0101100111010110"; -- -0.08219374199465686
	pesos_i(3689) := b"0000000000000000_0000000000000000_0010100111000000_0001001000100101"; -- 0.16308701898446604
	pesos_i(3690) := b"0000000000000000_0000000000000000_0000011000000000_0000000111110110"; -- 0.023437616867077963
	pesos_i(3691) := b"0000000000000000_0000000000000000_0010101011101010_0100111000101001"; -- 0.16763771535092334
	pesos_i(3692) := b"0000000000000000_0000000000000000_0010101111101000_0000010001110011"; -- 0.17150905427972105
	pesos_i(3693) := b"1111111111111111_1111111111111111_1110110101010001_0010011110001101"; -- -0.07298043062714793
	pesos_i(3694) := b"0000000000000000_0000000000000000_0010100100111011_0010000000110000"; -- 0.161058437020759
	pesos_i(3695) := b"1111111111111111_1111111111111111_1101100001100110_1000101100100111"; -- -0.1546853093528898
	pesos_i(3696) := b"1111111111111111_1111111111111111_1110111001010100_0011101010111001"; -- -0.06902726164744517
	pesos_i(3697) := b"0000000000000000_0000000000000000_0000010111011101_1101101101000110"; -- 0.022916512029733854
	pesos_i(3698) := b"1111111111111111_1111111111111111_1101111001100111_1101100010101100"; -- -0.13122793002187888
	pesos_i(3699) := b"1111111111111111_1111111111111111_1101100001111001_1010000000011011"; -- -0.15439414347993904
	pesos_i(3700) := b"1111111111111111_1111111111111111_1110001011001011_0011010010010010"; -- -0.11408683229946648
	pesos_i(3701) := b"1111111111111111_1111111111111111_1101001000110000_1101011100011010"; -- -0.17894225712745293
	pesos_i(3702) := b"1111111111111111_1111111111111111_1100110110010101_0111101001101000"; -- -0.1969378944706519
	pesos_i(3703) := b"0000000000000000_0000000000000000_0010010100011110_1010000100101101"; -- 0.1449986203870389
	pesos_i(3704) := b"1111111111111111_1111111111111111_1101101100100011_1001110110001010"; -- -0.1439878024386409
	pesos_i(3705) := b"1111111111111111_1111111111111111_1101101111111010_1101011100011000"; -- -0.14070373224819632
	pesos_i(3706) := b"0000000000000000_0000000000000000_0010011001101110_0011001011101101"; -- 0.15011900228453817
	pesos_i(3707) := b"0000000000000000_0000000000000000_0010000011010101_1101100010101110"; -- 0.12826303723079102
	pesos_i(3708) := b"1111111111111111_1111111111111111_1101110110100100_1001000100110000"; -- -0.13420765484531136
	pesos_i(3709) := b"1111111111111111_1111111111111111_1100101110000110_1001011010110101"; -- -0.20497758931443785
	pesos_i(3710) := b"0000000000000000_0000000000000000_0001111110000001_1010011111100000"; -- 0.12307213991971623
	pesos_i(3711) := b"0000000000000000_0000000000000000_0000001010101010_1101000101001011"; -- 0.010418969011717238
	pesos_i(3712) := b"1111111111111111_1111111111111111_1101000101001110_0101010010001000"; -- -0.18239852590372724
	pesos_i(3713) := b"1111111111111111_1111111111111111_1101001000010101_0101011001011011"; -- -0.17936191818361205
	pesos_i(3714) := b"1111111111111111_1111111111111111_1111001110011000_1001101110110011"; -- -0.0484526337088566
	pesos_i(3715) := b"1111111111111111_1111111111111111_1111101011111111_1011010010101000"; -- -0.019535740944382343
	pesos_i(3716) := b"1111111111111111_1111111111111111_1111101010011100_1101110101011000"; -- -0.021043935905343487
	pesos_i(3717) := b"1111111111111111_1111111111111111_1110110001011010_1110001010100010"; -- -0.07673820071790229
	pesos_i(3718) := b"1111111111111111_1111111111111111_1110101100000110_0101001101111100"; -- -0.08193472120980796
	pesos_i(3719) := b"0000000000000000_0000000000000000_0001100101011100_0011100001000100"; -- 0.09906341226341296
	pesos_i(3720) := b"0000000000000000_0000000000000000_0010010101001100_0010111100001010"; -- 0.1456937216483844
	pesos_i(3721) := b"1111111111111111_1111111111111111_1110110010000000_1100011011111011"; -- -0.07616001486124502
	pesos_i(3722) := b"1111111111111111_1111111111111111_1110001001001111_0000010110100110"; -- -0.1159817190691883
	pesos_i(3723) := b"1111111111111111_1111111111111111_1101101011001000_1000111101100001"; -- -0.14537719611183098
	pesos_i(3724) := b"0000000000000000_0000000000000000_0010010110000111_0101000011111000"; -- 0.1465960126394002
	pesos_i(3725) := b"0000000000000000_0000000000000000_0000100001000110_1001011100101111"; -- 0.032327126590351765
	pesos_i(3726) := b"1111111111111111_1111111111111111_1110001001011001_0011100000000000"; -- -0.11582612987215253
	pesos_i(3727) := b"1111111111111111_1111111111111111_1101101000101010_0100001010111010"; -- -0.14779265357110324
	pesos_i(3728) := b"1111111111111111_1111111111111111_1111000001010001_1101101111010110"; -- -0.06125093486354518
	pesos_i(3729) := b"0000000000000000_0000000000000000_0001010101111100_1100110010010001"; -- 0.0839355329198709
	pesos_i(3730) := b"0000000000000000_0000000000000000_0001101110100011_0011001010100100"; -- 0.10795895107716307
	pesos_i(3731) := b"0000000000000000_0000000000000000_0000110110011101_1110110111110010"; -- 0.05319106254066306
	pesos_i(3732) := b"1111111111111111_1111111111111111_1101111011110111_1100001000010010"; -- -0.12903201153188285
	pesos_i(3733) := b"0000000000000000_0000000000000000_0001001011000001_0010100110110001"; -- 0.07325993136310403
	pesos_i(3734) := b"0000000000000000_0000000000000000_0001101010000011_0101111110010110"; -- 0.10356709863629004
	pesos_i(3735) := b"0000000000000000_0000000000000000_0001011100110010_1100111111011101"; -- 0.09061907896340628
	pesos_i(3736) := b"1111111111111111_1111111111111111_1111100010011100_0111101010011111"; -- -0.028862320027131884
	pesos_i(3737) := b"1111111111111111_1111111111111111_1110001010011101_1110101011101110"; -- -0.11477786726274619
	pesos_i(3738) := b"0000000000000000_0000000000000000_0001000101111011_0010100101101011"; -- 0.06828554974162122
	pesos_i(3739) := b"1111111111111111_1111111111111111_1111100110101011_1001000000111001"; -- -0.024725900714847548
	pesos_i(3740) := b"1111111111111111_1111111111111111_1101100101111110_1101111111111011"; -- -0.15040779229679055
	pesos_i(3741) := b"1111111111111111_1111111111111111_1111000001001000_0001101101010100"; -- -0.06139973821461091
	pesos_i(3742) := b"0000000000000000_0000000000000000_0010111010011010_1011110100110011"; -- 0.18204863062129956
	pesos_i(3743) := b"1111111111111111_1111111111111111_1100011101100010_0000001101100000"; -- -0.2211606874535236
	pesos_i(3744) := b"1111111111111111_1111111111111111_1111011101101101_0010100000010011"; -- -0.03349065328829993
	pesos_i(3745) := b"1111111111111111_1111111111111111_1100111010100101_0111011100110000"; -- -0.1927876955879099
	pesos_i(3746) := b"0000000000000000_0000000000000000_0000000000001111_0011111101011000"; -- 0.00023265730430443697
	pesos_i(3747) := b"0000000000000000_0000000000000000_0001110010110101_1110100001110001"; -- 0.1121506954155773
	pesos_i(3748) := b"1111111111111111_1111111111111111_1111111110001111_0110101100000100"; -- -0.0017178644657421653
	pesos_i(3749) := b"1111111111111111_1111111111111111_1101110100000010_1001011101100000"; -- -0.13667920980423764
	pesos_i(3750) := b"0000000000000000_0000000000000000_0010111001101100_0000101010100010"; -- 0.18133608293925876
	pesos_i(3751) := b"0000000000000000_0000000000000000_0010100011101010_0101101101101100"; -- 0.15982600572674116
	pesos_i(3752) := b"0000000000000000_0000000000000000_0001000001001101_0011111000101100"; -- 0.06367863254176503
	pesos_i(3753) := b"0000000000000000_0000000000000000_0001011100111110_0000100000001001"; -- 0.09079027384498284
	pesos_i(3754) := b"0000000000000000_0000000000000000_0000010101101011_1011010001001000"; -- 0.02117468605668331
	pesos_i(3755) := b"0000000000000000_0000000000000000_0000001001110011_0100110010011011"; -- 0.009571826827935611
	pesos_i(3756) := b"1111111111111111_1111111111111111_1101110001110110_0011110001011010"; -- -0.13882086575424718
	pesos_i(3757) := b"0000000000000000_0000000000000000_0000001101001011_1111010000111001"; -- 0.012877716033040441
	pesos_i(3758) := b"0000000000000000_0000000000000000_0000010100001101_1101010000010110"; -- 0.019742255671398277
	pesos_i(3759) := b"1111111111111111_1111111111111111_1101101000110110_0101011011001010"; -- -0.14760835242519105
	pesos_i(3760) := b"1111111111111111_1111111111111111_1110010101101000_1011001111010010"; -- -0.10387111771693243
	pesos_i(3761) := b"0000000000000000_0000000000000000_0000001111011110_1011110001010110"; -- 0.01511742684915654
	pesos_i(3762) := b"1111111111111111_1111111111111111_1111010111110000_1101000110110100"; -- -0.03929414128167459
	pesos_i(3763) := b"0000000000000000_0000000000000000_0000100001101010_1001011001100110"; -- 0.03287639611218606
	pesos_i(3764) := b"1111111111111111_1111111111111111_1110011000101001_0000010001000101"; -- -0.10093663523379585
	pesos_i(3765) := b"0000000000000000_0000000000000000_0001000100001100_0111110110110110"; -- 0.06659684845512755
	pesos_i(3766) := b"0000000000000000_0000000000000000_0010011111101010_0011001001101101"; -- 0.15591731214008947
	pesos_i(3767) := b"1111111111111111_1111111111111111_1110110000100011_0010100011000010"; -- -0.07758851303956148
	pesos_i(3768) := b"0000000000000000_0000000000000000_0010000001001100_0010110100000111"; -- 0.12616235169221024
	pesos_i(3769) := b"0000000000000000_0000000000000000_0001110000101111_0101010110000011"; -- 0.11009726008452084
	pesos_i(3770) := b"1111111111111111_1111111111111111_1111000011011111_0010000011011000"; -- -0.05909533244048994
	pesos_i(3771) := b"0000000000000000_0000000000000000_0010101011110101_1100111110010110"; -- 0.1678132764167976
	pesos_i(3772) := b"1111111111111111_1111111111111111_1111001111001110_0111010010110001"; -- -0.04763098405616692
	pesos_i(3773) := b"0000000000000000_0000000000000000_0010000000100110_1011010010010010"; -- 0.12559059680596987
	pesos_i(3774) := b"0000000000000000_0000000000000000_0000010111111001_0010000110001001"; -- 0.023332687373480994
	pesos_i(3775) := b"1111111111111111_1111111111111111_1111100001110101_1000000010000110"; -- -0.029457061154937455
	pesos_i(3776) := b"1111111111111111_1111111111111111_1111000101101011_1001110000010110"; -- -0.05695175621017285
	pesos_i(3777) := b"0000000000000000_0000000000000000_0001010001001011_0001101111110101"; -- 0.0792710756206698
	pesos_i(3778) := b"0000000000000000_0000000000000000_0010000110101110_1111010100111110"; -- 0.13157589693350646
	pesos_i(3779) := b"0000000000000000_0000000000000000_0000101110111101_1101001001101100"; -- 0.04586520319788321
	pesos_i(3780) := b"0000000000000000_0000000000000000_0001101010001101_1111011101101101"; -- 0.10372873704603688
	pesos_i(3781) := b"0000000000000000_0000000000000000_0010101000100110_0010010001101111"; -- 0.16464450556491222
	pesos_i(3782) := b"0000000000000000_0000000000000000_0010010100100100_0101000100010100"; -- 0.1450853990062742
	pesos_i(3783) := b"0000000000000000_0000000000000000_0001011011101101_1010110101011011"; -- 0.08956416587591336
	pesos_i(3784) := b"0000000000000000_0000000000000000_0000000101101001_1110000101011111"; -- 0.0055218559521879014
	pesos_i(3785) := b"0000000000000000_0000000000000000_0000000001110001_0110110101000000"; -- 0.0017307549474060685
	pesos_i(3786) := b"0000000000000000_0000000000000000_0000000011110001_0111101001001011"; -- 0.0036846573629484578
	pesos_i(3787) := b"0000000000000000_0000000000000000_0000111101101001_1010011100100010"; -- 0.06020588476211893
	pesos_i(3788) := b"0000000000000000_0000000000000000_0000110000000001_0100010101001111"; -- 0.04689438990959837
	pesos_i(3789) := b"1111111111111111_1111111111111111_1111100110100101_1100100010100000"; -- -0.0248140916609417
	pesos_i(3790) := b"1111111111111111_1111111111111111_1111000001000111_0110101010000100"; -- -0.061410277246802224
	pesos_i(3791) := b"1111111111111111_1111111111111111_1111110011010100_1010100100100001"; -- -0.012380055917713774
	pesos_i(3792) := b"1111111111111111_1111111111111111_1111000101000100_1110101100001011"; -- -0.05754214276971146
	pesos_i(3793) := b"0000000000000000_0000000000000000_0001110100100001_1110101101100001"; -- 0.1137988197631072
	pesos_i(3794) := b"1111111111111111_1111111111111111_1110000000010101_1100110011011111"; -- -0.12466735415888804
	pesos_i(3795) := b"1111111111111111_1111111111111111_1110001010101000_1101110111110110"; -- -0.1146107934971946
	pesos_i(3796) := b"0000000000000000_0000000000000000_0000011001101110_1111001111100110"; -- 0.02513050417056545
	pesos_i(3797) := b"0000000000000000_0000000000000000_0001000010000011_0001001001100011"; -- 0.06449999720169614
	pesos_i(3798) := b"1111111111111111_1111111111111111_1110111011101101_0111100110001101"; -- -0.06668892207407091
	pesos_i(3799) := b"0000000000000000_0000000000000000_0000110100110110_0000001000011100"; -- 0.05160535044670357
	pesos_i(3800) := b"0000000000000000_0000000000000000_0010100010101001_1010110110110011"; -- 0.15883908854705844
	pesos_i(3801) := b"1111111111111111_1111111111111111_1110001111010101_1100010011100101"; -- -0.11001939212655017
	pesos_i(3802) := b"1111111111111111_1111111111111111_1111110000001011_1100110000101011"; -- -0.015444983881890724
	pesos_i(3803) := b"0000000000000000_0000000000000000_0010010101001000_0001101001011111"; -- 0.14563145454817158
	pesos_i(3804) := b"1111111111111111_1111111111111111_1101101001011101_0101110010110101"; -- -0.14701290675259426
	pesos_i(3805) := b"0000000000000000_0000000000000000_0010001111010001_0011101010101011"; -- 0.13991133389231972
	pesos_i(3806) := b"1111111111111111_1111111111111111_1110100100111010_0100000100000101"; -- -0.0889548647164688
	pesos_i(3807) := b"0000000000000000_0000000000000000_0000111001000000_0111011100011001"; -- 0.05567116134311721
	pesos_i(3808) := b"1111111111111111_1111111111111111_1101111101110010_1001001101010111"; -- -0.12715796595993414
	pesos_i(3809) := b"0000000000000000_0000000000000000_0010101111010000_0000111000111010"; -- 0.1711434260139787
	pesos_i(3810) := b"0000000000000000_0000000000000000_0000110000011010_0010010110000110"; -- 0.04727396508953837
	pesos_i(3811) := b"1111111111111111_1111111111111111_1110110110001010_0110010000001100"; -- -0.07210707382303072
	pesos_i(3812) := b"1111111111111111_1111111111111111_1101101110000011_1110100111110100"; -- -0.14251840401341204
	pesos_i(3813) := b"1111111111111111_1111111111111111_1111000101100101_1101100000110011"; -- -0.05703972585028547
	pesos_i(3814) := b"1111111111111111_1111111111111111_1101001111101011_0010011011010000"; -- -0.17219312119501648
	pesos_i(3815) := b"0000000000000000_0000000000000000_0000001001000001_0100101000110100"; -- 0.008808744254184125
	pesos_i(3816) := b"0000000000000000_0000000000000000_0001011010110111_0010110000100111"; -- 0.08873249019034636
	pesos_i(3817) := b"1111111111111111_1111111111111111_1110000110010111_0011100101110111"; -- -0.1187862477291313
	pesos_i(3818) := b"1111111111111111_1111111111111111_1110100110010000_1101001101110000"; -- -0.08763388176142088
	pesos_i(3819) := b"1111111111111111_1111111111111111_1100111110110110_1110011111001100"; -- -0.18861533414032128
	pesos_i(3820) := b"0000000000000000_0000000000000000_0000001011001010_1100010111110001"; -- 0.010906573690752607
	pesos_i(3821) := b"1111111111111111_1111111111111111_1110100000001111_1000101101110011"; -- -0.09351280645866468
	pesos_i(3822) := b"0000000000000000_0000000000000000_0000000111101001_0111011100101011"; -- 0.007468650810093319
	pesos_i(3823) := b"1111111111111111_1111111111111111_1101100110111100_1010110101011000"; -- -0.14946476555138324
	pesos_i(3824) := b"1111111111111111_1111111111111111_1110011001011000_0111101101011011"; -- -0.10021237399617247
	pesos_i(3825) := b"0000000000000000_0000000000000000_0001001010011111_1110111100111101"; -- 0.072752907153055
	pesos_i(3826) := b"1111111111111111_1111111111111111_1110010011011000_0110110010011001"; -- -0.10607262865286526
	pesos_i(3827) := b"0000000000000000_0000000000000000_0001010101001001_0101001011100010"; -- 0.08315008171851586
	pesos_i(3828) := b"1111111111111111_1111111111111111_1100110010100111_0010110110100100"; -- -0.20057406180220194
	pesos_i(3829) := b"1111111111111111_1111111111111111_1101011011101000_1011100001111101"; -- -0.16051146455146342
	pesos_i(3830) := b"1111111111111111_1111111111111111_1110000110000000_1000111111110100"; -- -0.11913204472245893
	pesos_i(3831) := b"1111111111111111_1111111111111111_1111110011010110_0001000111000001"; -- -0.01235856083466541
	pesos_i(3832) := b"1111111111111111_1111111111111111_1111011110111110_1001100000110001"; -- -0.032248008830832085
	pesos_i(3833) := b"0000000000000000_0000000000000000_0010100101101110_1111001101110000"; -- 0.1618492267799121
	pesos_i(3834) := b"0000000000000000_0000000000000000_0000011100011110_1010100011001011"; -- 0.027811574595822047
	pesos_i(3835) := b"1111111111111111_1111111111111111_1111011000101101_1110010000011001"; -- -0.038362258698988565
	pesos_i(3836) := b"1111111111111111_1111111111111111_1111011101111011_0100101100001111"; -- -0.033274945109204056
	pesos_i(3837) := b"0000000000000000_0000000000000000_0000011111100101_1001011111111010"; -- 0.03084707126063283
	pesos_i(3838) := b"1111111111111111_1111111111111111_1110101101000000_0000100111111101"; -- -0.08105409217510885
	pesos_i(3839) := b"1111111111111111_1111111111111111_1110100001111110_0101001101100010"; -- -0.09182242253695926
	pesos_i(3840) := b"1111111111111111_1111111111111111_1110001011100010_1111110111001001"; -- -0.11372388701051345
	pesos_i(3841) := b"0000000000000000_0000000000000000_0000111001110001_0011111001000010"; -- 0.056415454063389915
	pesos_i(3842) := b"1111111111111111_1111111111111111_1110010001101011_0110110011110001"; -- -0.10773581609698073
	pesos_i(3843) := b"1111111111111111_1111111111111111_1101100010111100_1000011001011101"; -- -0.15337333898329653
	pesos_i(3844) := b"1111111111111111_1111111111111111_1111111000110101_1001001111110101"; -- -0.006994965269090835
	pesos_i(3845) := b"1111111111111111_1111111111111111_1110000100010101_0010010000011100"; -- -0.12077116307742405
	pesos_i(3846) := b"0000000000000000_0000000000000000_0000000010010011_0111001001001001"; -- 0.0022498538951066954
	pesos_i(3847) := b"0000000000000000_0000000000000000_0010010010101111_1010101101011111"; -- 0.1433055027035309
	pesos_i(3848) := b"1111111111111111_1111111111111111_1110010000011001_0011011100101000"; -- -0.10899024273744343
	pesos_i(3849) := b"0000000000000000_0000000000000000_0010111100110010_0110011000110101"; -- 0.18436278153654415
	pesos_i(3850) := b"1111111111111111_1111111111111111_1110111101010000_0101110101111001"; -- -0.06517997537074421
	pesos_i(3851) := b"0000000000000000_0000000000000000_0001011110101110_1110001101011110"; -- 0.09251233138483388
	pesos_i(3852) := b"1111111111111111_1111111111111111_1110100011110010_1110010111011100"; -- -0.09004367245828786
	pesos_i(3853) := b"0000000000000000_0000000000000000_0000101100011011_0111011001010011"; -- 0.043387790054602506
	pesos_i(3854) := b"1111111111111111_1111111111111111_1110001101011100_0110010110100000"; -- -0.11187138399249091
	pesos_i(3855) := b"0000000000000000_0000000000000000_0000101010011010_1000111110100011"; -- 0.04142091502247705
	pesos_i(3856) := b"0000000000000000_0000000000000000_0000010101100001_1110100100101110"; -- 0.02102525118397614
	pesos_i(3857) := b"0000000000000000_0000000000000000_0000000011110010_0001001001100010"; -- 0.0036937226146937724
	pesos_i(3858) := b"1111111111111111_1111111111111111_1110011010000110_1111110011110010"; -- -0.09950274545161533
	pesos_i(3859) := b"1111111111111111_1111111111111111_1110110100100111_1010111001001011"; -- -0.07361326849533133
	pesos_i(3860) := b"0000000000000000_0000000000000000_0001001110100010_1110100000011001"; -- 0.07670450799731089
	pesos_i(3861) := b"0000000000000000_0000000000000000_0010101010100000_0011110001011011"; -- 0.1665075038183203
	pesos_i(3862) := b"1111111111111111_1111111111111111_1111011101101100_0000101101001001"; -- -0.033507628168014364
	pesos_i(3863) := b"0000000000000000_0000000000000000_0000111110011111_0100110100111110"; -- 0.061024501451314175
	pesos_i(3864) := b"1111111111111111_1111111111111111_1101010011100100_0011010000110101"; -- -0.1683928842395496
	pesos_i(3865) := b"0000000000000000_0000000000000000_0000101011010011_0000110110110100"; -- 0.04228292125586335
	pesos_i(3866) := b"1111111111111111_1111111111111111_1111100010110110_0111110110100110"; -- -0.028465411196698775
	pesos_i(3867) := b"1111111111111111_1111111111111111_1110011010101101_1110010111101010"; -- -0.09890902548950141
	pesos_i(3868) := b"1111111111111111_1111111111111111_1111111111101011_0100111000110100"; -- -0.0003157733736876413
	pesos_i(3869) := b"1111111111111111_1111111111111111_1111000110100111_1011110001110001"; -- -0.056034300255185444
	pesos_i(3870) := b"0000000000000000_0000000000000000_0000000001000000_1101101111100010"; -- 0.0009896686012755879
	pesos_i(3871) := b"1111111111111111_1111111111111111_1111110011110000_1010111100111100"; -- -0.011952445783127012
	pesos_i(3872) := b"1111111111111111_1111111111111111_1111111101110000_0000101011110110"; -- -0.0021966123331554482
	pesos_i(3873) := b"0000000000000000_0000000000000000_0000001000111100_1111111111001100"; -- 0.008743274063331473
	pesos_i(3874) := b"0000000000000000_0000000000000000_0001111100001110_0000101000100011"; -- 0.12130797721348835
	pesos_i(3875) := b"1111111111111111_1111111111111111_1101000101001001_0110100111010110"; -- -0.18247355017229944
	pesos_i(3876) := b"1111111111111111_1111111111111111_1110100110100100_1011111111111011"; -- -0.0873298655838913
	pesos_i(3877) := b"0000000000000000_0000000000000000_0000010111011100_1111100001011100"; -- 0.02290298704306998
	pesos_i(3878) := b"0000000000000000_0000000000000000_0001010110010001_1010011110001011"; -- 0.08425376078749976
	pesos_i(3879) := b"0000000000000000_0000000000000000_0011001100111100_1010111111110101"; -- 0.20014476523021893
	pesos_i(3880) := b"1111111111111111_1111111111111111_1110001110010001_1101111010000100"; -- -0.11105546253723071
	pesos_i(3881) := b"0000000000000000_0000000000000000_0001100001100110_1011100010100011"; -- 0.09531740180675757
	pesos_i(3882) := b"1111111111111111_1111111111111111_1111100001011110_1010110001101001"; -- -0.02980539730582394
	pesos_i(3883) := b"0000000000000000_0000000000000000_0000101000110110_0010001000100001"; -- 0.039888508896464815
	pesos_i(3884) := b"1111111111111111_1111111111111111_1101100110001011_0100100110010111"; -- -0.15021839201517453
	pesos_i(3885) := b"1111111111111111_1111111111111111_1101000001011011_1011100000110101"; -- -0.18610047062544327
	pesos_i(3886) := b"1111111111111111_1111111111111111_1111001000111000_0101001001111100"; -- -0.05382809135995447
	pesos_i(3887) := b"0000000000000000_0000000000000000_0000001111011111_1001000100100000"; -- 0.015130110062705792
	pesos_i(3888) := b"1111111111111111_1111111111111111_1111110000101100_1100101000110010"; -- -0.01494156150804428
	pesos_i(3889) := b"0000000000000000_0000000000000000_0001010011011001_1111101110001010"; -- 0.08145115018579788
	pesos_i(3890) := b"0000000000000000_0000000000000000_0001000111001100_0101110001010111"; -- 0.06952454695703905
	pesos_i(3891) := b"0000000000000000_0000000000000000_0000011000000101_1001101100001101"; -- 0.023523035805138186
	pesos_i(3892) := b"0000000000000000_0000000000000000_0000000100010011_0001111110100010"; -- 0.004198052494823889
	pesos_i(3893) := b"0000000000000000_0000000000000000_0010100100001000_1011010100000010"; -- 0.1602891093054218
	pesos_i(3894) := b"1111111111111111_1111111111111111_1101000011101100_0111101101100010"; -- -0.18389157159247707
	pesos_i(3895) := b"1111111111111111_1111111111111111_1111100010001100_0000101000000011"; -- -0.029113172851744758
	pesos_i(3896) := b"1111111111111111_1111111111111111_1110010110101101_1000101000010111"; -- -0.1028207487169791
	pesos_i(3897) := b"0000000000000000_0000000000000000_0000011000011001_1111000011110101"; -- 0.02383333179136335
	pesos_i(3898) := b"0000000000000000_0000000000000000_0001000111101100_1001100010111010"; -- 0.07001642747578678
	pesos_i(3899) := b"1111111111111111_1111111111111111_1110110101001100_1001000100110101"; -- -0.07305042705134969
	pesos_i(3900) := b"1111111111111111_1111111111111111_1110100011001110_1101001100001110"; -- -0.09059410966618284
	pesos_i(3901) := b"0000000000000000_0000000000000000_0010110110011101_0110101011001110"; -- 0.17818324588332868
	pesos_i(3902) := b"1111111111111111_1111111111111111_1110111000111100_0100100101011011"; -- -0.0693926003074623
	pesos_i(3903) := b"1111111111111111_1111111111111111_1111011000100000_0000010101010110"; -- -0.03857390073130415
	pesos_i(3904) := b"0000000000000000_0000000000000000_0000100100110111_0111000101000010"; -- 0.036002234180623094
	pesos_i(3905) := b"0000000000000000_0000000000000000_0001111011000110_1111101100111100"; -- 0.12022371505523893
	pesos_i(3906) := b"1111111111111111_1111111111111111_1111011110001010_0000101000101100"; -- -0.03304993093341532
	pesos_i(3907) := b"0000000000000000_0000000000000000_0010000111010010_1000110101111001"; -- 0.13211902805648107
	pesos_i(3908) := b"0000000000000000_0000000000000000_0001111111100010_0111101110000101"; -- 0.12454959877639654
	pesos_i(3909) := b"1111111111111111_1111111111111111_1111010011001001_0101100011100111"; -- -0.043802684290834726
	pesos_i(3910) := b"1111111111111111_1111111111111111_1101001001101000_1100101001111000"; -- -0.17808851779674778
	pesos_i(3911) := b"1111111111111111_1111111111111111_1111101010011111_0100111011111000"; -- -0.021006645686554887
	pesos_i(3912) := b"0000000000000000_0000000000000000_0001101001001110_1011111101111011"; -- 0.10276409869929531
	pesos_i(3913) := b"0000000000000000_0000000000000000_0000001110100101_0110011110010100"; -- 0.014242623901566276
	pesos_i(3914) := b"0000000000000000_0000000000000000_0010010011101001_0100100111111101"; -- 0.14418470800357897
	pesos_i(3915) := b"1111111111111111_1111111111111111_1101110010110000_0111001011000100"; -- -0.13793261249331173
	pesos_i(3916) := b"1111111111111111_1111111111111111_1100111101000100_1010101101110111"; -- -0.19035843218961002
	pesos_i(3917) := b"0000000000000000_0000000000000000_0001101111011011_0010010011010101"; -- 0.10881262016185683
	pesos_i(3918) := b"1111111111111111_1111111111111111_1111110110010000_1011100101101101"; -- -0.009510432080213016
	pesos_i(3919) := b"0000000000000000_0000000000000000_0001100011100000_0001010110111101"; -- 0.09716926455104574
	pesos_i(3920) := b"1111111111111111_1111111111111111_1110101100010111_1010101010000010"; -- -0.08167013476422377
	pesos_i(3921) := b"1111111111111111_1111111111111111_1101110010101000_1000001011101100"; -- -0.13805371985086726
	pesos_i(3922) := b"0000000000000000_0000000000000000_0000011101010110_1010010000110110"; -- 0.028665793598629252
	pesos_i(3923) := b"0000000000000000_0000000000000000_0001101101111100_1111111110111100"; -- 0.10737608270550619
	pesos_i(3924) := b"1111111111111111_1111111111111111_1101110111111010_1000111100101110"; -- -0.13289551854655038
	pesos_i(3925) := b"1111111111111111_1111111111111111_1100111101010101_0110001001011001"; -- -0.19010339085920816
	pesos_i(3926) := b"0000000000000000_0000000000000000_0000011000101010_1001001011110000"; -- 0.024087127404474634
	pesos_i(3927) := b"0000000000000000_0000000000000000_0000111001000100_1100000101110001"; -- 0.055736627740955696
	pesos_i(3928) := b"1111111111111111_1111111111111111_1111000111000111_1000001111011001"; -- -0.05554939226350042
	pesos_i(3929) := b"0000000000000000_0000000000000000_0000000010110011_1101011111000111"; -- 0.0027441845905543383
	pesos_i(3930) := b"1111111111111111_1111111111111111_1110101100100111_0111111110110100"; -- -0.08142854560910369
	pesos_i(3931) := b"1111111111111111_1111111111111111_1110110100000110_1011000010111011"; -- -0.07411666330840123
	pesos_i(3932) := b"1111111111111111_1111111111111111_1110010000101100_1010100001011011"; -- -0.10869357861117081
	pesos_i(3933) := b"0000000000000000_0000000000000000_0000011101000100_0101101110011011"; -- 0.02838680773395358
	pesos_i(3934) := b"1111111111111111_1111111111111111_1111010000101001_0010111010111101"; -- -0.046246603754040244
	pesos_i(3935) := b"0000000000000000_0000000000000000_0001010000011011_0100000110000001"; -- 0.07854089157362448
	pesos_i(3936) := b"1111111111111111_1111111111111111_1110011001101011_1000101011011111"; -- -0.09992153217100294
	pesos_i(3937) := b"0000000000000000_0000000000000000_0001000010010010_1001001000100111"; -- 0.06473649461507963
	pesos_i(3938) := b"0000000000000000_0000000000000000_0001010101110010_1011001010000100"; -- 0.0837813922582556
	pesos_i(3939) := b"1111111111111111_1111111111111111_1110001101000101_1111101010100001"; -- -0.11221345493641618
	pesos_i(3940) := b"0000000000000000_0000000000000000_0001111111111101_1100111110011001"; -- 0.12496659734247234
	pesos_i(3941) := b"1111111111111111_1111111111111111_1101111101100001_1101111100001110"; -- -0.12741285236181005
	pesos_i(3942) := b"1111111111111111_1111111111111111_1111111011010011_1010010000110111"; -- -0.004583107546610704
	pesos_i(3943) := b"0000000000000000_0000000000000000_0001101100001101_1101001000100010"; -- 0.10567963912150397
	pesos_i(3944) := b"1111111111111111_1111111111111111_1101111100111100_0101011000010100"; -- -0.12798559205522486
	pesos_i(3945) := b"0000000000000000_0000000000000000_0010100010000010_1100101000010100"; -- 0.15824568746393264
	pesos_i(3946) := b"0000000000000000_0000000000000000_0000011000001101_0000100111101110"; -- 0.023636456213182694
	pesos_i(3947) := b"1111111111111111_1111111111111111_1111100001101011_0111101010000110"; -- -0.02961000654974752
	pesos_i(3948) := b"1111111111111111_1111111111111111_1110010000010100_1110010011100000"; -- -0.1090561821308297
	pesos_i(3949) := b"1111111111111111_1111111111111111_1101100101010010_1110011010111110"; -- -0.15107877605515613
	pesos_i(3950) := b"0000000000000000_0000000000000000_0000000111111000_1101000111000011"; -- 0.007702932401773832
	pesos_i(3951) := b"1111111111111111_1111111111111111_1111100000111101_0110101011101000"; -- -0.030312841642366
	pesos_i(3952) := b"0000000000000000_0000000000000000_0001111100001011_0010001010110111"; -- 0.12126366581245396
	pesos_i(3953) := b"0000000000000000_0000000000000000_0001100110010100_0100101110100100"; -- 0.09991905937637369
	pesos_i(3954) := b"0000000000000000_0000000000000000_0010101101001010_0011010110001110"; -- 0.1691010924289954
	pesos_i(3955) := b"0000000000000000_0000000000000000_0001111100110100_1110010011111101"; -- 0.1219008559027061
	pesos_i(3956) := b"1111111111111111_1111111111111111_1110111111101001_1001001111000111"; -- -0.06284214389137335
	pesos_i(3957) := b"1111111111111111_1111111111111111_1101001111011010_1001011001001101"; -- -0.17244587542709489
	pesos_i(3958) := b"1111111111111111_1111111111111111_1110110101100110_0011001000111110"; -- -0.07265935891418346
	pesos_i(3959) := b"1111111111111111_1111111111111111_1101001110110101_1111000110111011"; -- -0.17300500083135284
	pesos_i(3960) := b"1111111111111111_1111111111111111_1111011011101100_0111111001110001"; -- -0.03545388929998919
	pesos_i(3961) := b"1111111111111111_1111111111111111_1110110110011010_1011001111011100"; -- -0.07185817601453211
	pesos_i(3962) := b"1111111111111111_1111111111111111_1110111010100110_0101001101000101"; -- -0.0677745778627129
	pesos_i(3963) := b"1111111111111111_1111111111111111_1101011100011010_1111100100110101"; -- -0.1597446675107606
	pesos_i(3964) := b"1111111111111111_1111111111111111_1101101010110001_0000000110110101"; -- -0.1457365924788884
	pesos_i(3965) := b"1111111111111111_1111111111111111_1101100100000001_1010011011111111"; -- -0.1523185373634895
	pesos_i(3966) := b"0000000000000000_0000000000000000_0011000001010010_0111010110100111"; -- 0.1887582333828282
	pesos_i(3967) := b"0000000000000000_0000000000000000_0001100101110100_1000000101101001"; -- 0.09943398303187478
	pesos_i(3968) := b"0000000000000000_0000000000000000_0010101111111101_1000011010000101"; -- 0.17183724155836738
	pesos_i(3969) := b"1111111111111111_1111111111111111_1111111101101111_1010011110100110"; -- -0.00220253185811331
	pesos_i(3970) := b"0000000000000000_0000000000000000_0001011111011010_1110111101110101"; -- 0.09318443877338545
	pesos_i(3971) := b"1111111111111111_1111111111111111_1101010100111111_0001011011110001"; -- -0.16700607875990067
	pesos_i(3972) := b"0000000000000000_0000000000000000_0001001110110011_0110111001110111"; -- 0.07695665735368129
	pesos_i(3973) := b"0000000000000000_0000000000000000_0001001110001011_0100100101110010"; -- 0.07634409934322467
	pesos_i(3974) := b"1111111111111111_1111111111111111_1101000110111001_0000100000011111"; -- -0.18077038999911182
	pesos_i(3975) := b"1111111111111111_1111111111111111_1111111011100100_0111011111001100"; -- -0.004326355564558709
	pesos_i(3976) := b"1111111111111111_1111111111111111_1100111100001100_1101000010111101"; -- -0.19121070269829177
	pesos_i(3977) := b"1111111111111111_1111111111111111_1111101111111010_0101111010010010"; -- -0.015710915924631363
	pesos_i(3978) := b"1111111111111111_1111111111111111_1111011110001010_1111001000000000"; -- -0.033036112685965874
	pesos_i(3979) := b"1111111111111111_1111111111111111_1100111100010010_0000001100111010"; -- -0.19113139936313112
	pesos_i(3980) := b"1111111111111111_1111111111111111_1111101011111001_1101100101010100"; -- -0.019625107816296644
	pesos_i(3981) := b"1111111111111111_1111111111111111_1111011101010010_0010001011011100"; -- -0.03390295149189404
	pesos_i(3982) := b"1111111111111111_1111111111111111_1101000100011010_1101101100001001"; -- -0.18318396598252268
	pesos_i(3983) := b"0000000000000000_0000000000000000_0000110011100111_0011101001100111"; -- 0.0504032613085193
	pesos_i(3984) := b"1111111111111111_1111111111111111_1110100000001011_1001100101100100"; -- -0.0935730104321495
	pesos_i(3985) := b"1111111111111111_1111111111111111_1101011100111111_1110010001011001"; -- -0.15918133571846976
	pesos_i(3986) := b"1111111111111111_1111111111111111_1101101011010001_0101000000101000"; -- -0.1452436355019232
	pesos_i(3987) := b"0000000000000000_0000000000000000_0010010100000000_1010111010111100"; -- 0.1445416649204414
	pesos_i(3988) := b"0000000000000000_0000000000000000_0010011001100101_1110100000001100"; -- 0.14999246877225414
	pesos_i(3989) := b"1111111111111111_1111111111111111_1111110011101011_1110110001001100"; -- -0.01202510023843642
	pesos_i(3990) := b"1111111111111111_1111111111111111_1101001100110011_1000110111000101"; -- -0.17499460168360625
	pesos_i(3991) := b"0000000000000000_0000000000000000_0001000110100000_1111010000110000"; -- 0.06886221088467082
	pesos_i(3992) := b"0000000000000000_0000000000000000_0010100100101011_1000111101010110"; -- 0.16082092130767378
	pesos_i(3993) := b"1111111111111111_1111111111111111_1110011011101011_0111100101011100"; -- -0.0979694510417026
	pesos_i(3994) := b"1111111111111111_1111111111111111_1110101101000011_1000100011010011"; -- -0.08100075587849849
	pesos_i(3995) := b"0000000000000000_0000000000000000_0010010001110011_0010010100101100"; -- 0.14238197630029575
	pesos_i(3996) := b"0000000000000000_0000000000000000_0010111011010111_0010000100100000"; -- 0.182970114062473
	pesos_i(3997) := b"1111111111111111_1111111111111111_1110000010000101_1010111001000100"; -- -0.1229601939039028
	pesos_i(3998) := b"1111111111111111_1111111111111111_1100111101001010_1110110011100001"; -- -0.19026298050853294
	pesos_i(3999) := b"0000000000000000_0000000000000000_0000111000011111_1111001110010110"; -- 0.05517504121638114
	pesos_i(4000) := b"0000000000000000_0000000000000000_0000111011100101_1001000101001111"; -- 0.05819042378686298
	pesos_i(4001) := b"0000000000000000_0000000000000000_0001010100101010_0001000101011111"; -- 0.08267315444234502
	pesos_i(4002) := b"0000000000000000_0000000000000000_0000000011111011_1101011101010101"; -- 0.0038427907848495313
	pesos_i(4003) := b"1111111111111111_1111111111111111_1110011111011000_0100001001011111"; -- -0.09435639563997146
	pesos_i(4004) := b"0000000000000000_0000000000000000_0000101111100000_0010011010101011"; -- 0.046389023546428404
	pesos_i(4005) := b"0000000000000000_0000000000000000_0010001100010100_0000101001101100"; -- 0.13702454705959477
	pesos_i(4006) := b"0000000000000000_0000000000000000_0010001001000010_1101110010111001"; -- 0.1338327362684697
	pesos_i(4007) := b"1111111111111111_1111111111111111_1111011111101011_0000111011110100"; -- -0.03156954332801276
	pesos_i(4008) := b"1111111111111111_1111111111111111_1111101001011010_0001000010110111"; -- -0.022063212763686224
	pesos_i(4009) := b"1111111111111111_1111111111111111_1111111111100111_0101101001001001"; -- -0.000376088195546076
	pesos_i(4010) := b"0000000000000000_0000000000000000_0001101100001100_0110110100011010"; -- 0.10565835844839788
	pesos_i(4011) := b"1111111111111111_1111111111111111_1110011010010011_0100110010001101"; -- -0.09931489526300472
	pesos_i(4012) := b"1111111111111111_1111111111111111_1101111011001111_0010001111000001"; -- -0.1296517995001708
	pesos_i(4013) := b"1111111111111111_1111111111111111_1101001001111001_0011010001101110"; -- -0.17783806135955016
	pesos_i(4014) := b"1111111111111111_1111111111111111_1101010011011000_1110101100011111"; -- -0.16856508728624114
	pesos_i(4015) := b"0000000000000000_0000000000000000_0001100111100011_0011000111011100"; -- 0.10112296700613677
	pesos_i(4016) := b"0000000000000000_0000000000000000_0010000000000111_1001100110111011"; -- 0.12511597468735713
	pesos_i(4017) := b"1111111111111111_1111111111111111_1110100000111010_0010100111001000"; -- -0.09286249979530048
	pesos_i(4018) := b"1111111111111111_1111111111111111_1101001110000010_0001011001110100"; -- -0.17379626917977645
	pesos_i(4019) := b"0000000000000000_0000000000000000_0001110000100111_0110000011110101"; -- 0.10997587190127267
	pesos_i(4020) := b"1111111111111111_1111111111111111_1111100101110011_1101101100001000"; -- -0.025575934079760054
	pesos_i(4021) := b"0000000000000000_0000000000000000_0000111110011000_1011111010110000"; -- 0.060924451754025055
	pesos_i(4022) := b"1111111111111111_1111111111111111_1101001101100010_1000001011010111"; -- -0.17427808997255845
	pesos_i(4023) := b"0000000000000000_0000000000000000_0000101001110100_1011000101100011"; -- 0.040843092591899194
	pesos_i(4024) := b"0000000000000000_0000000000000000_0001111111011101_0001011010010111"; -- 0.1244672888930235
	pesos_i(4025) := b"0000000000000000_0000000000000000_0010000011000001_0010011001110000"; -- 0.12794723738248043
	pesos_i(4026) := b"1111111111111111_1111111111111111_1110011001001001_1101001101010100"; -- -0.10043601223742164
	pesos_i(4027) := b"0000000000000000_0000000000000000_0000100111100010_0010001100011111"; -- 0.03860682972931981
	pesos_i(4028) := b"0000000000000000_0000000000000000_0010110111100101_0001000000101011"; -- 0.17927647629242072
	pesos_i(4029) := b"0000000000000000_0000000000000000_0000010011001011_1010101101011101"; -- 0.018732748260641946
	pesos_i(4030) := b"0000000000000000_0000000000000000_0001011000101100_0000000010100000"; -- 0.08660892395684677
	pesos_i(4031) := b"1111111111111111_1111111111111111_1101101000101100_1011100011101010"; -- -0.14775509164495618
	pesos_i(4032) := b"1111111111111111_1111111111111111_1111101111110100_1110101010101100"; -- -0.015794117900900878
	pesos_i(4033) := b"1111111111111111_1111111111111111_1111000101010011_0001001101000111"; -- -0.05732612154241329
	pesos_i(4034) := b"0000000000000000_0000000000000000_0000101011010100_1110111000101100"; -- 0.04231155949037396
	pesos_i(4035) := b"0000000000000000_0000000000000000_0001101010011010_0001001011111001"; -- 0.10391348434234182
	pesos_i(4036) := b"0000000000000000_0000000000000000_0010111100011110_1010001000101101"; -- 0.18406118007484717
	pesos_i(4037) := b"0000000000000000_0000000000000000_0001010011110111_0010001110111111"; -- 0.08189605145095791
	pesos_i(4038) := b"0000000000000000_0000000000000000_0010110000011101_1101101100000110"; -- 0.17233055972063138
	pesos_i(4039) := b"1111111111111111_1111111111111111_1111111000111001_1000000000000011"; -- -0.006935118935583295
	pesos_i(4040) := b"1111111111111111_1111111111111111_1101011101111111_1101101100111101"; -- -0.15820531627693069
	pesos_i(4041) := b"0000000000000000_0000000000000000_0000001011010001_1101100001100011"; -- 0.011014484669869123
	pesos_i(4042) := b"0000000000000000_0000000000000000_0000010101010010_0010001011011100"; -- 0.020784548582696932
	pesos_i(4043) := b"0000000000000000_0000000000000000_0010010010111001_0111111000111000"; -- 0.1434553992248369
	pesos_i(4044) := b"1111111111111111_1111111111111111_1110100011001111_0100010101000101"; -- -0.09058730188656672
	pesos_i(4045) := b"1111111111111111_1111111111111111_1101100011000001_0100000110011000"; -- -0.15330114407177173
	pesos_i(4046) := b"0000000000000000_0000000000000000_0001000010011010_1001011010011111"; -- 0.06485883125680825
	pesos_i(4047) := b"0000000000000000_0000000000000000_0001011110101010_1101011000010011"; -- 0.09245050392485904
	pesos_i(4048) := b"0000000000000000_0000000000000000_0001101101011010_0001001111111110"; -- 0.10684323265613876
	pesos_i(4049) := b"1111111111111111_1111111111111111_1110010101000100_1000101000010110"; -- -0.1044229216873268
	pesos_i(4050) := b"0000000000000000_0000000000000000_0001011001011011_0010001110011011"; -- 0.0873281719993172
	pesos_i(4051) := b"0000000000000000_0000000000000000_0010100110100001_0100010111111000"; -- 0.16261708545633746
	pesos_i(4052) := b"1111111111111111_1111111111111111_1101000110101100_1011111000010111"; -- -0.18095790807172907
	pesos_i(4053) := b"1111111111111111_1111111111111111_1101011010110010_1010101001111010"; -- -0.16133627444104212
	pesos_i(4054) := b"0000000000000000_0000000000000000_0010000011111001_0111011111010001"; -- 0.12880658013206348
	pesos_i(4055) := b"1111111111111111_1111111111111111_1101101101111110_0101100001101001"; -- -0.14260337286886615
	pesos_i(4056) := b"0000000000000000_0000000000000000_0001010010001000_0000110011010011"; -- 0.08020095979396602
	pesos_i(4057) := b"1111111111111111_1111111111111111_1111000111100101_1111100100011010"; -- -0.05508463973524813
	pesos_i(4058) := b"1111111111111111_1111111111111111_1110101110100111_0111111100001000"; -- -0.07947546060186039
	pesos_i(4059) := b"0000000000000000_0000000000000000_0000111010010010_1000011010010011"; -- 0.0569233044499724
	pesos_i(4060) := b"1111111111111111_1111111111111111_1101101111000110_0101100110001011"; -- -0.14150467257591698
	pesos_i(4061) := b"1111111111111111_1111111111111111_1101110111001010_0100000100001101"; -- -0.13363259717420903
	pesos_i(4062) := b"0000000000000000_0000000000000000_0010111110111000_0000000101110000"; -- 0.1864014528872866
	pesos_i(4063) := b"1111111111111111_1111111111111111_1110100100101010_1100000001001100"; -- -0.0891914189654516
	pesos_i(4064) := b"0000000000000000_0000000000000000_0000111100110101_0100101000011010"; -- 0.059406882593553645
	pesos_i(4065) := b"0000000000000000_0000000000000000_0010101110101101_0001111000000000"; -- 0.1706103085631493
	pesos_i(4066) := b"0000000000000000_0000000000000000_0000011111110100_1110111100101111"; -- 0.031081150994528572
	pesos_i(4067) := b"1111111111111111_1111111111111111_1110110100110110_1111010110011100"; -- -0.07338013583823783
	pesos_i(4068) := b"0000000000000000_0000000000000000_0001010110011101_1011101011101110"; -- 0.08443802174551318
	pesos_i(4069) := b"1111111111111111_1111111111111111_1111010000001011_0111010110001101"; -- -0.046700146860794184
	pesos_i(4070) := b"0000000000000000_0000000000000000_0010010110011101_0110100001111001"; -- 0.14693310691205885
	pesos_i(4071) := b"1111111111111111_1111111111111111_1101010001010000_1100010001010111"; -- -0.1706425940128287
	pesos_i(4072) := b"1111111111111111_1111111111111111_1111001011000011_1101000100110011"; -- -0.05169956677232562
	pesos_i(4073) := b"0000000000000000_0000000000000000_0001011011011111_0010100110101001"; -- 0.089342693026013
	pesos_i(4074) := b"1111111111111111_1111111111111111_1111100100110000_1101101000000001"; -- -0.02659833405447054
	pesos_i(4075) := b"1111111111111111_1111111111111111_1111000010110110_1000110100100101"; -- -0.05971448743449953
	pesos_i(4076) := b"0000000000000000_0000000000000000_0000011110001010_0100011001111111"; -- 0.029453664801525725
	pesos_i(4077) := b"0000000000000000_0000000000000000_0010101010110000_1001011111101010"; -- 0.1667571015516774
	pesos_i(4078) := b"1111111111111111_1111111111111111_1111001011100100_1111010111011111"; -- -0.051193840975747806
	pesos_i(4079) := b"1111111111111111_1111111111111111_1111111111101101_0100011100101101"; -- -0.00028567451734953786
	pesos_i(4080) := b"0000000000000000_0000000000000000_0001110000000101_0110010111110111"; -- 0.1094573714381053
	pesos_i(4081) := b"0000000000000000_0000000000000000_0001010000100111_0011010101001100"; -- 0.07872326959363773
	pesos_i(4082) := b"0000000000000000_0000000000000000_0001100011111111_0010010111111111"; -- 0.09764325600716928
	pesos_i(4083) := b"1111111111111111_1111111111111111_1101010001100111_0101011010000111"; -- -0.17029818729042753
	pesos_i(4084) := b"1111111111111111_1111111111111111_1110101010000110_1110111010001100"; -- -0.08387860387263893
	pesos_i(4085) := b"0000000000000000_0000000000000000_0001001110011000_1011011011010010"; -- 0.07654898292888856
	pesos_i(4086) := b"0000000000000000_0000000000000000_0010100010110001_0001110001101000"; -- 0.15895249874131218
	pesos_i(4087) := b"0000000000000000_0000000000000000_0011000000110101_0101100110111100"; -- 0.18831406448250992
	pesos_i(4088) := b"0000000000000000_0000000000000000_0000011110011010_1110011110101001"; -- 0.029707411422800423
	pesos_i(4089) := b"1111111111111111_1111111111111111_1111001000000110_1001001111010100"; -- -0.054587136097236616
	pesos_i(4090) := b"0000000000000000_0000000000000000_0001101001001111_0110100001111110"; -- 0.1027741725801804
	pesos_i(4091) := b"1111111111111111_1111111111111111_1101010110011100_0000011110001001"; -- -0.16558792967194794
	pesos_i(4092) := b"1111111111111111_1111111111111111_1111111001011111_0001100001011001"; -- -0.006361463858227584
	pesos_i(4093) := b"0000000000000000_0000000000000000_0010001000011101_1010100011010110"; -- 0.13326506835660146
	pesos_i(4094) := b"1111111111111111_1111111111111111_1101100001010010_0010101000011000"; -- -0.15499627032107646
	pesos_i(4095) := b"1111111111111111_1111111111111111_1111110001111111_1100011110011100"; -- -0.013675236154224113
	pesos_i(4096) := b"1111111111111111_1111111111111111_1111110101001100_1001110010000110"; -- -0.01054975240759004
	pesos_i(4097) := b"1111111111111111_1111111111111111_1110011000110011_1101110111010100"; -- -0.1007710797944256
	pesos_i(4098) := b"0000000000000000_0000000000000000_0001010011110101_1101110110111111"; -- 0.08187662048938976
	pesos_i(4099) := b"0000000000000000_0000000000000000_0010010000101001_1101110010001111"; -- 0.14126375659209145
	pesos_i(4100) := b"0000000000000000_0000000000000000_0000110000010011_1111010000010110"; -- 0.047179465687129
	pesos_i(4101) := b"1111111111111111_1111111111111111_1101101010000101_0100001011101101"; -- -0.14640409194318152
	pesos_i(4102) := b"1111111111111111_1111111111111111_1110001000010111_0111100101110110"; -- -0.11682930811126555
	pesos_i(4103) := b"1111111111111111_1111111111111111_1111011111001100_0110101001001111"; -- -0.03203712056593108
	pesos_i(4104) := b"1111111111111111_1111111111111111_1101001010001111_1001100001100101"; -- -0.17749640964544502
	pesos_i(4105) := b"1111111111111111_1111111111111111_1111110101000111_1011110100001011"; -- -0.01062410820424252
	pesos_i(4106) := b"1111111111111111_1111111111111111_1110111001001000_0011010101111010"; -- -0.06921067981667604
	pesos_i(4107) := b"1111111111111111_1111111111111111_1110101110000111_0101100100011010"; -- -0.0799660025151487
	pesos_i(4108) := b"1111111111111111_1111111111111111_1101100010011001_1001010000011101"; -- -0.15390657707182628
	pesos_i(4109) := b"1111111111111111_1111111111111111_1111100111110100_0101010000001000"; -- -0.02361559686783602
	pesos_i(4110) := b"0000000000000000_0000000000000000_0010111101010110_1011111101000001"; -- 0.18491740558513362
	pesos_i(4111) := b"1111111111111111_1111111111111111_1100111110111000_0111000010011011"; -- -0.18859192100139266
	pesos_i(4112) := b"0000000000000000_0000000000000000_0001011111000001_1111101100000101"; -- 0.09280365827845777
	pesos_i(4113) := b"1111111111111111_1111111111111111_1110111110000111_1000100001101000"; -- -0.06433818310540804
	pesos_i(4114) := b"0000000000000000_0000000000000000_0000111010000101_0100010011101110"; -- 0.056721027460757904
	pesos_i(4115) := b"0000000000000000_0000000000000000_0001100101001001_0111001011100010"; -- 0.09877698924104113
	pesos_i(4116) := b"0000000000000000_0000000000000000_0010001010011111_1000010000000100"; -- 0.13524651610940377
	pesos_i(4117) := b"1111111111111111_1111111111111111_1101101111000011_0010110101101110"; -- -0.14155307824382807
	pesos_i(4118) := b"1111111111111111_1111111111111111_1101000101101000_0000101000111101"; -- -0.18200622575724867
	pesos_i(4119) := b"0000000000000000_0000000000000000_0000110111001000_0111001000101110"; -- 0.053839813545332925
	pesos_i(4120) := b"1111111111111111_1111111111111111_1111010000111110_1001101100000011"; -- -0.04591971555113834
	pesos_i(4121) := b"1111111111111111_1111111111111111_1110010011011001_0110010011011100"; -- -0.10605783112560646
	pesos_i(4122) := b"1111111111111111_1111111111111111_1111011000110111_0101010000110001"; -- -0.03821824846085797
	pesos_i(4123) := b"0000000000000000_0000000000000000_0000011010011000_0011111111001000"; -- 0.025760637560358204
	pesos_i(4124) := b"1111111111111111_1111111111111111_1101001100001010_1111001000110011"; -- -0.17561422586430203
	pesos_i(4125) := b"1111111111111111_1111111111111111_1101000000101101_0000000000100010"; -- -0.18681334657398888
	pesos_i(4126) := b"1111111111111111_1111111111111111_1110001110001111_0000010100101101"; -- -0.11109893458964895
	pesos_i(4127) := b"1111111111111111_1111111111111111_1110101011000001_1111000000000010"; -- -0.08297824803467284
	pesos_i(4128) := b"1111111111111111_1111111111111111_1111010100010111_1001001111101100"; -- -0.04260898107538493
	pesos_i(4129) := b"1111111111111111_1111111111111111_1101111011010100_1111110111110110"; -- -0.1295624994299086
	pesos_i(4130) := b"1111111111111111_1111111111111111_1111100100110101_0110100100101101"; -- -0.026528765305936047
	pesos_i(4131) := b"0000000000000000_0000000000000000_0001110101100100_0001101100110000"; -- 0.11480874934650868
	pesos_i(4132) := b"0000000000000000_0000000000000000_0000000110010010_1100111111010110"; -- 0.006146421176449496
	pesos_i(4133) := b"0000000000000000_0000000000000000_0001111101100111_0100101011111000"; -- 0.1226698738479301
	pesos_i(4134) := b"0000000000000000_0000000000000000_0010001111110101_1010100101011000"; -- 0.14046724694973464
	pesos_i(4135) := b"1111111111111111_1111111111111111_1110111010100100_1000000110100001"; -- -0.06780233213955941
	pesos_i(4136) := b"1111111111111111_1111111111111111_1110111011011111_0110001001011011"; -- -0.06690392760297936
	pesos_i(4137) := b"0000000000000000_0000000000000000_0001101010001110_1010000111111110"; -- 0.10373890357254757
	pesos_i(4138) := b"0000000000000000_0000000000000000_0000100010001000_0001010100101001"; -- 0.033326456619458524
	pesos_i(4139) := b"1111111111111111_1111111111111111_1101010011100110_0011001111010010"; -- -0.16836238969083853
	pesos_i(4140) := b"1111111111111111_1111111111111111_1111010111011100_0101010010011010"; -- -0.039606773713908874
	pesos_i(4141) := b"1111111111111111_1111111111111111_1101001001111000_1000011111110100"; -- -0.17784834195975907
	pesos_i(4142) := b"0000000000000000_0000000000000000_0010101101100001_1101110111100011"; -- 0.16946207801064278
	pesos_i(4143) := b"1111111111111111_1111111111111111_1110101101011101_0011110111101010"; -- -0.08060849221177707
	pesos_i(4144) := b"0000000000000000_0000000000000000_0001101011111111_1010100100100101"; -- 0.105463573005612
	pesos_i(4145) := b"1111111111111111_1111111111111111_1111010100100011_1101000111111011"; -- -0.042422176648569884
	pesos_i(4146) := b"0000000000000000_0000000000000000_0000110111010001_1110011010101101"; -- 0.05398408622499053
	pesos_i(4147) := b"0000000000000000_0000000000000000_0000101100110111_0010111001011101"; -- 0.04381074694769693
	pesos_i(4148) := b"0000000000000000_0000000000000000_0010000101101101_1001100111111010"; -- 0.13057863562285557
	pesos_i(4149) := b"1111111111111111_1111111111111111_1111100110010111_0010010110111001"; -- -0.025037424326144104
	pesos_i(4150) := b"0000000000000000_0000000000000000_0001011000100001_1110010011000101"; -- 0.08645467584392146
	pesos_i(4151) := b"1111111111111111_1111111111111111_1110111101000001_0100010110111101"; -- -0.06541027192083018
	pesos_i(4152) := b"0000000000000000_0000000000000000_0001011000011101_1000011110110010"; -- 0.08638809301890696
	pesos_i(4153) := b"1111111111111111_1111111111111111_1101111111111100_1111101110100101"; -- -0.125046035991521
	pesos_i(4154) := b"0000000000000000_0000000000000000_0000010100101011_0001111011000001"; -- 0.020189211053752244
	pesos_i(4155) := b"0000000000000000_0000000000000000_0010100111100001_0010011011010000"; -- 0.16359179092575674
	pesos_i(4156) := b"1111111111111111_1111111111111111_1100010100001010_1100111001010100"; -- -0.2303038640994807
	pesos_i(4157) := b"0000000000000000_0000000000000000_0011010001000000_1000011011101000"; -- 0.2041096035894619
	pesos_i(4158) := b"1111111111111111_1111111111111111_1100101110000011_1010110110001001"; -- -0.20502200522106195
	pesos_i(4159) := b"1111111111111111_1111111111111111_1110100010101111_0001011111010011"; -- -0.09107829183807281
	pesos_i(4160) := b"0000000000000000_0000000000000000_0010101011000110_1100100010000100"; -- 0.1670956918361955
	pesos_i(4161) := b"0000000000000000_0000000000000000_0000100111100101_0110001011000111"; -- 0.03865640027759805
	pesos_i(4162) := b"0000000000000000_0000000000000000_0001111001001110_1100010000010000"; -- 0.11838937179491373
	pesos_i(4163) := b"0000000000000000_0000000000000000_0001110101111101_0110110101000001"; -- 0.11519511069509937
	pesos_i(4164) := b"0000000000000000_0000000000000000_0000000011001110_0100110000001111"; -- 0.0031478439087519166
	pesos_i(4165) := b"1111111111111111_1111111111111111_1110001011001110_0111100000111100"; -- -0.11403702288301087
	pesos_i(4166) := b"0000000000000000_0000000000000000_0010011000001111_1110001101111011"; -- 0.14867994076112115
	pesos_i(4167) := b"0000000000000000_0000000000000000_0000011011100101_1010001111011011"; -- 0.026941529139592378
	pesos_i(4168) := b"1111111111111111_1111111111111111_1110110111011011_0111110101111100"; -- -0.07086959581345943
	pesos_i(4169) := b"0000000000000000_0000000000000000_0010010000111110_0101111101101110"; -- 0.14157673301215795
	pesos_i(4170) := b"0000000000000000_0000000000000000_0000011110001000_0010010011101110"; -- 0.029421146485262326
	pesos_i(4171) := b"1111111111111111_1111111111111111_1111011010101000_1100011001011111"; -- -0.03648719960561564
	pesos_i(4172) := b"0000000000000000_0000000000000000_0010110111100110_0000111100000110"; -- 0.1792916669522627
	pesos_i(4173) := b"0000000000000000_0000000000000000_0001110001111100_0011001101100001"; -- 0.11127015234980764
	pesos_i(4174) := b"0000000000000000_0000000000000000_0001111010100001_0001000000011001"; -- 0.11964512453215165
	pesos_i(4175) := b"1111111111111111_1111111111111111_1101111101111111_1101101110111110"; -- -0.12695528607145176
	pesos_i(4176) := b"0000000000000000_0000000000000000_0000000011011011_0011000101001111"; -- 0.003344613853378597
	pesos_i(4177) := b"0000000000000000_0000000000000000_0000101011101011_0110111111010010"; -- 0.04265498054595734
	pesos_i(4178) := b"1111111111111111_1111111111111111_1111000000000110_0101001100010111"; -- -0.062403494744722704
	pesos_i(4179) := b"1111111111111111_1111111111111111_1110001000010100_0101110010010100"; -- -0.11687680620056305
	pesos_i(4180) := b"1111111111111111_1111111111111111_1111001110001101_0110111100111110"; -- -0.04862313029938407
	pesos_i(4181) := b"0000000000000000_0000000000000000_0001011100000110_0010101101111101"; -- 0.08993789494253758
	pesos_i(4182) := b"1111111111111111_1111111111111111_1111011001000101_1100100010010001"; -- -0.037997688922919354
	pesos_i(4183) := b"0000000000000000_0000000000000000_0000110010011101_0101111011111101"; -- 0.049276291601395836
	pesos_i(4184) := b"1111111111111111_1111111111111111_1101111001110000_1000110001000111"; -- -0.13109515441863087
	pesos_i(4185) := b"0000000000000000_0000000000000000_0000000100111111_0111111001001010"; -- 0.004875081033248067
	pesos_i(4186) := b"0000000000000000_0000000000000000_0000110101011110_1010011010010110"; -- 0.052225505407409445
	pesos_i(4187) := b"0000000000000000_0000000000000000_0001001101110001_0101111110000011"; -- 0.07594868612331111
	pesos_i(4188) := b"0000000000000000_0000000000000000_0001100010111010_1110011101001110"; -- 0.09660192170673869
	pesos_i(4189) := b"1111111111111111_1111111111111111_1101110011011011_0111111000111110"; -- -0.13727580050576813
	pesos_i(4190) := b"0000000000000000_0000000000000000_0010000101001101_0111010001010000"; -- 0.13008810959717862
	pesos_i(4191) := b"0000000000000000_0000000000000000_0000000000000010_1010010001011100"; -- 4.0314162671155396e-05
	pesos_i(4192) := b"0000000000000000_0000000000000000_0001011000101011_0100100111101000"; -- 0.08659803315279556
	pesos_i(4193) := b"0000000000000000_0000000000000000_0010000100101001_0111101111110000"; -- 0.12953924765883035
	pesos_i(4194) := b"1111111111111111_1111111111111111_1110111011110001_1001010000000010"; -- -0.06662630987195522
	pesos_i(4195) := b"0000000000000000_0000000000000000_0010111110100110_0001111001000010"; -- 0.18612851252146195
	pesos_i(4196) := b"1111111111111111_1111111111111111_1110001100101001_0000011011100100"; -- -0.11265522899934996
	pesos_i(4197) := b"0000000000000000_0000000000000000_0000101011010011_1001000010011001"; -- 0.04229072325353084
	pesos_i(4198) := b"0000000000000000_0000000000000000_0010100101001111_0001101100001010"; -- 0.16136330607606397
	pesos_i(4199) := b"1111111111111111_1111111111111111_1101011010010100_0000011011100101"; -- -0.16180378823416547
	pesos_i(4200) := b"0000000000000000_0000000000000000_0001100011110110_1000001010101101"; -- 0.09751145110199494
	pesos_i(4201) := b"0000000000000000_0000000000000000_0010000100010101_1110011001110111"; -- 0.1292404213490937
	pesos_i(4202) := b"1111111111111111_1111111111111111_1101100001100111_1101101111001001"; -- -0.1546652445153304
	pesos_i(4203) := b"0000000000000000_0000000000000000_0010100110111111_1110100110010101"; -- 0.1630846013300858
	pesos_i(4204) := b"1111111111111111_1111111111111111_1110011010101110_0100100101100110"; -- -0.09890309581546834
	pesos_i(4205) := b"0000000000000000_0000000000000000_0000010101101001_1010010011101011"; -- 0.021143252633061323
	pesos_i(4206) := b"1111111111111111_1111111111111111_1111000110101100_0101000010111101"; -- -0.05596442590743792
	pesos_i(4207) := b"0000000000000000_0000000000000000_0001011111011111_0101110011000100"; -- 0.0932519891978492
	pesos_i(4208) := b"1111111111111111_1111111111111111_1111111000011100_0010100111011101"; -- -0.0073827585782372225
	pesos_i(4209) := b"1111111111111111_1111111111111111_1101111000100101_0111001101111000"; -- -0.1322410424278484
	pesos_i(4210) := b"1111111111111111_1111111111111111_1111110101111110_1000101010101000"; -- -0.009787878069863174
	pesos_i(4211) := b"1111111111111111_1111111111111111_1111101011011000_1101101111010001"; -- -0.020128499505613212
	pesos_i(4212) := b"1111111111111111_1111111111111111_1110010100110000_1101100011000100"; -- -0.10472340793113438
	pesos_i(4213) := b"1111111111111111_1111111111111111_1110110010001001_1011000111010111"; -- -0.0760239457908687
	pesos_i(4214) := b"1111111111111111_1111111111111111_1110101100110010_0110011011101101"; -- -0.08126217569257173
	pesos_i(4215) := b"0000000000000000_0000000000000000_0000011110110010_0110111011010011"; -- 0.0300664200650492
	pesos_i(4216) := b"1111111111111111_1111111111111111_1111001110010000_0001000010001111"; -- -0.0485829973281118
	pesos_i(4217) := b"0000000000000000_0000000000000000_0000101001010010_1001010010100111"; -- 0.0403225811384328
	pesos_i(4218) := b"1111111111111111_1111111111111111_1100111011101011_1001110010000011"; -- -0.19171735578827948
	pesos_i(4219) := b"1111111111111111_1111111111111111_1111000011000000_0100010110110100"; -- -0.05956615776572489
	pesos_i(4220) := b"1111111111111111_1111111111111111_1111101011111111_1110000001101101"; -- -0.019533131975098404
	pesos_i(4221) := b"1111111111111111_1111111111111111_1111101010010011_1001001001100100"; -- -0.02118573238154267
	pesos_i(4222) := b"1111111111111111_1111111111111111_1111011001001110_0110011100011000"; -- -0.03786616954195682
	pesos_i(4223) := b"1111111111111111_1111111111111111_1100101101000010_0111011101100100"; -- -0.20601705378370144
	pesos_i(4224) := b"1111111111111111_1111111111111111_1110000111001110_0001001100100100"; -- -0.11794929861320429
	pesos_i(4225) := b"1111111111111111_1111111111111111_1110111101001010_0011110011011011"; -- -0.06527347233873147
	pesos_i(4226) := b"1111111111111111_1111111111111111_1111110110101100_1100110011010001"; -- -0.009082030174169382
	pesos_i(4227) := b"0000000000000000_0000000000000000_0000100011110101_1000010001011001"; -- 0.034996291766208935
	pesos_i(4228) := b"0000000000000000_0000000000000000_0010000011001010_0110011111010001"; -- 0.12808846327799306
	pesos_i(4229) := b"1111111111111111_1111111111111111_1101101100001010_1101111110110000"; -- -0.14436532922571768
	pesos_i(4230) := b"0000000000000000_0000000000000000_0000010111010111_0110001001000000"; -- 0.022817745811395528
	pesos_i(4231) := b"1111111111111111_1111111111111111_1111101100101101_1011100111111110"; -- -0.018833518588218627
	pesos_i(4232) := b"1111111111111111_1111111111111111_1110001110111000_0000110010000111"; -- -0.11047288619754925
	pesos_i(4233) := b"1111111111111111_1111111111111111_1111100010010111_0010001000100110"; -- -0.02894388755572871
	pesos_i(4234) := b"0000000000000000_0000000000000000_0000110011110011_0000100001110011"; -- 0.05058338933821452
	pesos_i(4235) := b"0000000000000000_0000000000000000_0000110101011101_0000011011110110"; -- 0.0522007322743144
	pesos_i(4236) := b"1111111111111111_1111111111111111_1111111011111111_1111011010110011"; -- -0.003906804282219646
	pesos_i(4237) := b"1111111111111111_1111111111111111_1111100011001000_1111101100110110"; -- -0.028183268798149187
	pesos_i(4238) := b"1111111111111111_1111111111111111_1111101110001010_1010001011010100"; -- -0.01741583173214558
	pesos_i(4239) := b"0000000000000000_0000000000000000_0000111111011010_0000000011000110"; -- 0.06192021215593582
	pesos_i(4240) := b"0000000000000000_0000000000000000_0000111010110010_0100010111011000"; -- 0.057407727497091235
	pesos_i(4241) := b"1111111111111111_1111111111111111_1110010110000000_1110001110101111"; -- -0.10350205405155931
	pesos_i(4242) := b"1111111111111111_1111111111111111_1101001001011101_0110011110010111"; -- -0.17826225808165308
	pesos_i(4243) := b"1111111111111111_1111111111111111_1110011110100100_1101101000110010"; -- -0.09514080325262678
	pesos_i(4244) := b"1111111111111111_1111111111111111_1110011010000110_1011101010100000"; -- -0.09950669855516667
	pesos_i(4245) := b"1111111111111111_1111111111111111_1101011110111110_0010111011011100"; -- -0.1572542869940466
	pesos_i(4246) := b"0000000000000000_0000000000000000_0001100000010010_0011010111000111"; -- 0.09402786347444164
	pesos_i(4247) := b"1111111111111111_1111111111111111_1110010111011011_1010101100001010"; -- -0.1021168804345603
	pesos_i(4248) := b"1111111111111111_1111111111111111_1111000100010111_0001111011100011"; -- -0.058240956946962734
	pesos_i(4249) := b"0000000000000000_0000000000000000_0000101010011101_1110011010010100"; -- 0.041471873325464224
	pesos_i(4250) := b"1111111111111111_1111111111111111_1110101000100111_1111111001100111"; -- -0.08532724356820719
	pesos_i(4251) := b"1111111111111111_1111111111111111_1110101111111101_1111110100100101"; -- -0.07815568785679834
	pesos_i(4252) := b"1111111111111111_1111111111111111_1111011110100110_0011101111000001"; -- -0.032619729343861675
	pesos_i(4253) := b"0000000000000000_0000000000000000_0001111011100110_1100110010101010"; -- 0.12070922029860838
	pesos_i(4254) := b"0000000000000000_0000000000000000_0000000111001110_0000011111000101"; -- 0.0070500236074491456
	pesos_i(4255) := b"0000000000000000_0000000000000000_0001010101110010_1101110110010110"; -- 0.08378395961644738
	pesos_i(4256) := b"0000000000000000_0000000000000000_0010100010111101_0111111000011011"; -- 0.15914142761568467
	pesos_i(4257) := b"1111111111111111_1111111111111111_1111011010101100_1011101100000011"; -- -0.03642684160845918
	pesos_i(4258) := b"1111111111111111_1111111111111111_1110001100110100_1100100101010101"; -- -0.11247579257678617
	pesos_i(4259) := b"0000000000000000_0000000000000000_0001010101000001_1101111001011110"; -- 0.08303632536845447
	pesos_i(4260) := b"1111111111111111_1111111111111111_1110100100100001_0110101000011010"; -- -0.08933388571926841
	pesos_i(4261) := b"0000000000000000_0000000000000000_0001010110111110_0100010111010000"; -- 0.0849345811313614
	pesos_i(4262) := b"0000000000000000_0000000000000000_0001011001100110_1010011011011001"; -- 0.0875038413366664
	pesos_i(4263) := b"0000000000000000_0000000000000000_0000110001110010_0010001111010001"; -- 0.04861663671110902
	pesos_i(4264) := b"1111111111111111_1111111111111111_1110011011111010_0010001111110101"; -- -0.0977456594658094
	pesos_i(4265) := b"1111111111111111_1111111111111111_1110011011000010_0100101101111001"; -- -0.09859779631424744
	pesos_i(4266) := b"1111111111111111_1111111111111111_1111100001000100_1000001101000110"; -- -0.030204577742409987
	pesos_i(4267) := b"0000000000000000_0000000000000000_0010001010111101_1001110001011110"; -- 0.13570573126426982
	pesos_i(4268) := b"0000000000000000_0000000000000000_0000011101001111_0000100001010000"; -- 0.028549689892161542
	pesos_i(4269) := b"0000000000000000_0000000000000000_0000110011011010_0010011100000100"; -- 0.050203741432890255
	pesos_i(4270) := b"0000000000000000_0000000000000000_0001010000001100_0011111110001011"; -- 0.07831189293307708
	pesos_i(4271) := b"1111111111111111_1111111111111111_1100111011111101_1100100110011000"; -- -0.19144001055581678
	pesos_i(4272) := b"1111111111111111_1111111111111111_1110000110100011_0011110110110110"; -- -0.11860288905848003
	pesos_i(4273) := b"0000000000000000_0000000000000000_0010101001000011_1000011111101110"; -- 0.1650929409222367
	pesos_i(4274) := b"1111111111111111_1111111111111111_1110101100100001_0110100000111111"; -- -0.08152149638158665
	pesos_i(4275) := b"1111111111111111_1111111111111111_1110110111001111_0101011010111000"; -- -0.07105501178001314
	pesos_i(4276) := b"1111111111111111_1111111111111111_1101100110101010_1010011111001110"; -- -0.14973975392223443
	pesos_i(4277) := b"0000000000000000_0000000000000000_0000100110111000_1000011110101001"; -- 0.03797195308095201
	pesos_i(4278) := b"1111111111111111_1111111111111111_1101100101011010_0000000100101101"; -- -0.15097038896850296
	pesos_i(4279) := b"0000000000000000_0000000000000000_0010101010111010_0000100011111000"; -- 0.1669011693842669
	pesos_i(4280) := b"1111111111111111_1111111111111111_1101100101101010_0101010000000010"; -- -0.15072131107729653
	pesos_i(4281) := b"0000000000000000_0000000000000000_0010011000011101_1100111111000110"; -- 0.14889238922354497
	pesos_i(4282) := b"1111111111111111_1111111111111111_1111100111100111_0100000010000100"; -- -0.02381512427268607
	pesos_i(4283) := b"1111111111111111_1111111111111111_1101010000011001_1000000110110111"; -- -0.17148579876761028
	pesos_i(4284) := b"0000000000000000_0000000000000000_0001110111011111_0001000011010100"; -- 0.11668496297350342
	pesos_i(4285) := b"1111111111111111_1111111111111111_1111000010111001_1111010110011110"; -- -0.059662483985099345
	pesos_i(4286) := b"1111111111111111_1111111111111111_1101001001001110_1011010011000111"; -- -0.17848653918957977
	pesos_i(4287) := b"1111111111111111_1111111111111111_1110110010110000_1111111011101000"; -- -0.0754242595773444
	pesos_i(4288) := b"1111111111111111_1111111111111111_1110000010101101_1100110111100110"; -- -0.1223479570430953
	pesos_i(4289) := b"0000000000000000_0000000000000000_0000100111100011_0101111010110110"; -- 0.03862564030011298
	pesos_i(4290) := b"1111111111111111_1111111111111111_1111000110100111_1011001110101001"; -- -0.05603482369782532
	pesos_i(4291) := b"1111111111111111_1111111111111111_1101101010010011_1110000001000001"; -- -0.14618109148506386
	pesos_i(4292) := b"0000000000000000_0000000000000000_0000010110111111_0001100110110001"; -- 0.022447210145147025
	pesos_i(4293) := b"0000000000000000_0000000000000000_0000001100001011_0010100101001010"; -- 0.011889057595488604
	pesos_i(4294) := b"0000000000000000_0000000000000000_0000000010100010_0110111110100000"; -- 0.0024785771415966606
	pesos_i(4295) := b"0000000000000000_0000000000000000_0001000111000111_1101010011111100"; -- 0.06945544383582992
	pesos_i(4296) := b"1111111111111111_1111111111111111_1101111001100101_0000111010100100"; -- -0.13127048972005373
	pesos_i(4297) := b"1111111111111111_1111111111111111_1111100101000101_1110110000110111"; -- -0.02627681396655726
	pesos_i(4298) := b"1111111111111111_1111111111111111_1101101010011001_1011111001010001"; -- -0.14609156150304844
	pesos_i(4299) := b"0000000000000000_0000000000000000_0001100001100101_1010000101111110"; -- 0.09530076336538604
	pesos_i(4300) := b"0000000000000000_0000000000000000_0000001011000101_1111001101111111"; -- 0.010832995020785885
	pesos_i(4301) := b"1111111111111111_1111111111111111_1101000011101101_0110101000010100"; -- -0.18387734414779522
	pesos_i(4302) := b"0000000000000000_0000000000000000_0010001000001011_1001011111110001"; -- 0.13298940310307703
	pesos_i(4303) := b"1111111111111111_1111111111111111_1111111001100101_0010111010011000"; -- -0.0062685850952936
	pesos_i(4304) := b"1111111111111111_1111111111111111_1111000000101100_0100111111010000"; -- -0.06182385603720586
	pesos_i(4305) := b"0000000000000000_0000000000000000_0010000010100000_0010100110100000"; -- 0.12744388725378747
	pesos_i(4306) := b"1111111111111111_1111111111111111_1110011001101011_1010011100010001"; -- -0.09991985152721239
	pesos_i(4307) := b"0000000000000000_0000000000000000_0001101101001101_1001110010101110"; -- 0.10665301566707973
	pesos_i(4308) := b"0000000000000000_0000000000000000_0001001111001100_1010101101100111"; -- 0.07734175943733443
	pesos_i(4309) := b"1111111111111111_1111111111111111_1110110010010011_1111111010011111"; -- -0.07586678131541434
	pesos_i(4310) := b"1111111111111111_1111111111111111_1110011010101100_1010111110110100"; -- -0.09892751548890516
	pesos_i(4311) := b"0000000000000000_0000000000000000_0001100000111101_1101001100010010"; -- 0.09469336682216573
	pesos_i(4312) := b"1111111111111111_1111111111111111_1111011111010110_1110010010001001"; -- -0.03187724739909758
	pesos_i(4313) := b"1111111111111111_1111111111111111_1111101010010001_1111010110001111"; -- -0.021210339212159098
	pesos_i(4314) := b"0000000000000000_0000000000000000_0001000111011010_0101010011110101"; -- 0.06973772991122282
	pesos_i(4315) := b"1111111111111111_1111111111111111_1110010100010011_1111111000110100"; -- -0.10516368122203372
	pesos_i(4316) := b"0000000000000000_0000000000000000_0001011110000010_1110010110000011"; -- 0.09184107245172164
	pesos_i(4317) := b"1111111111111111_1111111111111111_1111111110101001_1010000110001001"; -- -0.0013178863943840947
	pesos_i(4318) := b"0000000000000000_0000000000000000_0001000001001101_0110011010011100"; -- 0.06368104280766831
	pesos_i(4319) := b"1111111111111111_1111111111111111_1101100101011111_0110100010111001"; -- -0.15088792302654103
	pesos_i(4320) := b"0000000000000000_0000000000000000_0001010010111010_0110101000000000"; -- 0.08096945280149202
	pesos_i(4321) := b"0000000000000000_0000000000000000_0000111011000110_1010001110111001"; -- 0.05771849885895994
	pesos_i(4322) := b"1111111111111111_1111111111111111_1111100001101000_1000111000011011"; -- -0.029654615778082816
	pesos_i(4323) := b"0000000000000000_0000000000000000_0010011010101110_1000001111010011"; -- 0.15110038673997886
	pesos_i(4324) := b"1111111111111111_1111111111111111_1100101110010100_1011010100011001"; -- -0.20476215499720485
	pesos_i(4325) := b"1111111111111111_1111111111111111_1111000111110110_1110011010001000"; -- -0.054826347243024445
	pesos_i(4326) := b"1111111111111111_1111111111111111_1101111100001000_1101000110111100"; -- -0.12877167851318483
	pesos_i(4327) := b"1111111111111111_1111111111111111_1111010110110111_0010101010111111"; -- -0.04017384375282694
	pesos_i(4328) := b"1111111111111111_1111111111111111_1101101110110100_0001001000100010"; -- -0.14178358721980047
	pesos_i(4329) := b"0000000000000000_0000000000000000_0010011110100110_0000011000110110"; -- 0.15487707906994133
	pesos_i(4330) := b"0000000000000000_0000000000000000_0000001100011011_0011110110100100"; -- 0.01213441128405248
	pesos_i(4331) := b"1111111111111111_1111111111111111_1111111110010110_0100100000010110"; -- -0.0016131350736859594
	pesos_i(4332) := b"0000000000000000_0000000000000000_0000010010110111_0011000000011111"; -- 0.018420226662893415
	pesos_i(4333) := b"1111111111111111_1111111111111111_1110000110110001_1110000111010100"; -- -0.11837948395588073
	pesos_i(4334) := b"0000000000000000_0000000000000000_0000000100010011_0111001110110101"; -- 0.0042030636648662315
	pesos_i(4335) := b"1111111111111111_1111111111111111_1111110111100011_1000111101100001"; -- -0.008246458815552221
	pesos_i(4336) := b"1111111111111111_1111111111111111_1101001111100000_1110110010110100"; -- -0.17234917268127767
	pesos_i(4337) := b"0000000000000000_0000000000000000_0001000011100001_0100010000110011"; -- 0.06593729253195031
	pesos_i(4338) := b"0000000000000000_0000000000000000_0000110011110101_0101010010101111"; -- 0.05061845090293969
	pesos_i(4339) := b"0000000000000000_0000000000000000_0010010011010111_0011011001111000"; -- 0.14390888633360782
	pesos_i(4340) := b"1111111111111111_1111111111111111_1110111010000011_0000100111001100"; -- -0.06831301473338888
	pesos_i(4341) := b"0000000000000000_0000000000000000_0010001100001111_0111100101101100"; -- 0.13695486911335672
	pesos_i(4342) := b"1111111111111111_1111111111111111_1111110111111001_0101011100001010"; -- -0.007914123606588414
	pesos_i(4343) := b"0000000000000000_0000000000000000_0010011010011000_1111101101000010"; -- 0.15077181207102988
	pesos_i(4344) := b"0000000000000000_0000000000000000_0000001111000010_1011011001101101"; -- 0.014689828487704176
	pesos_i(4345) := b"1111111111111111_1111111111111111_1110000111100100_1001101101111100"; -- -0.1176054784848433
	pesos_i(4346) := b"0000000000000000_0000000000000000_0001010111011101_0110100011000010"; -- 0.08540968649796386
	pesos_i(4347) := b"1111111111111111_1111111111111111_1101001010010010_0100000101011110"; -- -0.17745582057278164
	pesos_i(4348) := b"1111111111111111_1111111111111111_1110110001000001_1011011110001001"; -- -0.07712223904752805
	pesos_i(4349) := b"0000000000000000_0000000000000000_0000000101110101_0111110001111101"; -- 0.005698948509495896
	pesos_i(4350) := b"1111111111111111_1111111111111111_1110000101010000_0001111100111111"; -- -0.11987118437667646
	pesos_i(4351) := b"1111111111111111_1111111111111111_1111101101100101_0001110001100011"; -- -0.017988420211763785
	pesos_i(4352) := b"1111111111111111_1111111111111111_1101110100011010_1110000111101010"; -- -0.1363085559533882
	pesos_i(4353) := b"1111111111111111_1111111111111111_1110110101111100_1011111101101111"; -- -0.07231524981894535
	pesos_i(4354) := b"1111111111111111_1111111111111111_1110011111011001_0010100100100001"; -- -0.09434264121024576
	pesos_i(4355) := b"1111111111111111_1111111111111111_1110100011010000_0101010110001001"; -- -0.09057107366296854
	pesos_i(4356) := b"0000000000000000_0000000000000000_0000101000110011_1101110001100000"; -- 0.03985383361725974
	pesos_i(4357) := b"0000000000000000_0000000000000000_0010010111110010_1011100100101101"; -- 0.1482349143810144
	pesos_i(4358) := b"0000000000000000_0000000000000000_0001101011111001_0111100100110000"; -- 0.10536916186733328
	pesos_i(4359) := b"0000000000000000_0000000000000000_0010000011111111_0011011100100110"; -- 0.1288942782047755
	pesos_i(4360) := b"0000000000000000_0000000000000000_0010000101101100_1010010000100110"; -- 0.13056398327873325
	pesos_i(4361) := b"0000000000000000_0000000000000000_0000100011010011_0001101000001100"; -- 0.03447115709887318
	pesos_i(4362) := b"1111111111111111_1111111111111111_1111000111001100_0111101101100100"; -- -0.05547360226905979
	pesos_i(4363) := b"0000000000000000_0000000000000000_0000100011100010_1101110100110010"; -- 0.03471167068794603
	pesos_i(4364) := b"0000000000000000_0000000000000000_0000101101111010_0010010101100001"; -- 0.04483255030575521
	pesos_i(4365) := b"0000000000000000_0000000000000000_0001110110011100_1010100110010100"; -- 0.11567172866723707
	pesos_i(4366) := b"1111111111111111_1111111111111111_1110001001001010_1000010000001100"; -- -0.11605047896031992
	pesos_i(4367) := b"0000000000000000_0000000000000000_0000010100000101_0101111100001110"; -- 0.01961320970575205
	pesos_i(4368) := b"1111111111111111_1111111111111111_1110111000111100_0100000100000010"; -- -0.069393097881813
	pesos_i(4369) := b"0000000000000000_0000000000000000_0001100111011111_1100001101000000"; -- 0.10107059771061637
	pesos_i(4370) := b"1111111111111111_1111111111111111_1101111101001000_1000101100100110"; -- -0.12779932339639033
	pesos_i(4371) := b"0000000000000000_0000000000000000_0000000110001011_0010001100101100"; -- 0.006029318003649787
	pesos_i(4372) := b"0000000000000000_0000000000000000_0000100100001101_0010111010010001"; -- 0.03535738992136795
	pesos_i(4373) := b"1111111111111111_1111111111111111_1110010010000110_0010101000111000"; -- -0.10732780593314024
	pesos_i(4374) := b"1111111111111111_1111111111111111_1100111110001111_1111000100001101"; -- -0.18920987547684248
	pesos_i(4375) := b"1111111111111111_1111111111111111_1101000000110101_0111101010101101"; -- -0.18668397218110427
	pesos_i(4376) := b"1111111111111111_1111111111111111_1101100000110100_0011100010110110"; -- -0.155453162622005
	pesos_i(4377) := b"0000000000000000_0000000000000000_0001100000110000_1010000011001011"; -- 0.09449200595508402
	pesos_i(4378) := b"1111111111111111_1111111111111111_1110110100000010_1011101000101000"; -- -0.07417713663908254
	pesos_i(4379) := b"0000000000000000_0000000000000000_0001101011111011_0010100100000010"; -- 0.10539490035498912
	pesos_i(4380) := b"0000000000000000_0000000000000000_0000100101001111_0000110110110111"; -- 0.036362511772098045
	pesos_i(4381) := b"1111111111111111_1111111111111111_1101011111110011_0010100111011010"; -- -0.15644586963088555
	pesos_i(4382) := b"0000000000000000_0000000000000000_0000001101101110_0111110001000011"; -- 0.013404623359249345
	pesos_i(4383) := b"0000000000000000_0000000000000000_0010000000010100_0110001000000000"; -- 0.12531101693881527
	pesos_i(4384) := b"1111111111111111_1111111111111111_1111001111111100_1110001110011100"; -- -0.04692246854425063
	pesos_i(4385) := b"1111111111111111_1111111111111111_1110011010100000_0000001110111111"; -- -0.0991208704404842
	pesos_i(4386) := b"1111111111111111_1111111111111111_1101110001011100_0110010001110011"; -- -0.13921520409502244
	pesos_i(4387) := b"0000000000000000_0000000000000000_0001111000010111_0000110110110011"; -- 0.11753926873220724
	pesos_i(4388) := b"1111111111111111_1111111111111111_1111000010001110_1011000011100110"; -- -0.06032270809571263
	pesos_i(4389) := b"0000000000000000_0000000000000000_0001110011110010_1111100011111011"; -- 0.11308246743229507
	pesos_i(4390) := b"0000000000000000_0000000000000000_0000111111000110_0001100110011010"; -- 0.06161651610245946
	pesos_i(4391) := b"1111111111111111_1111111111111111_1100110001101101_0100100010001011"; -- -0.20145746813515444
	pesos_i(4392) := b"0000000000000000_0000000000000000_0001011101010100_1011100001111100"; -- 0.09113648433301638
	pesos_i(4393) := b"1111111111111111_1111111111111111_1101100011111110_1100010000011001"; -- -0.15236257929741684
	pesos_i(4394) := b"0000000000000000_0000000000000000_0000001100110111_0110101111011001"; -- 0.012564411610641757
	pesos_i(4395) := b"1111111111111111_1111111111111111_1110000001100101_1011110111001001"; -- -0.12344755032156085
	pesos_i(4396) := b"1111111111111111_1111111111111111_1111111100000000_0011000101001011"; -- -0.003903312014137378
	pesos_i(4397) := b"0000000000000000_0000000000000000_0000010011111101_1001110111011110"; -- 0.01949488327386989
	pesos_i(4398) := b"1111111111111111_1111111111111111_1101100010110111_0111110100001110"; -- -0.15345018785143683
	pesos_i(4399) := b"1111111111111111_1111111111111111_1110101011000011_0000000011001000"; -- -0.08296198952926827
	pesos_i(4400) := b"0000000000000000_0000000000000000_0000011110010010_0000000101110100"; -- 0.029571619825005287
	pesos_i(4401) := b"0000000000000000_0000000000000000_0000110001010111_0010001011111000"; -- 0.04820459891081524
	pesos_i(4402) := b"1111111111111111_1111111111111111_1101010000110001_1011010101001111"; -- -0.17111651254724058
	pesos_i(4403) := b"0000000000000000_0000000000000000_0010110010000001_0000011110011010"; -- 0.1738438368068042
	pesos_i(4404) := b"1111111111111111_1111111111111111_1111111010010011_0101111000111101"; -- -0.005563841004723794
	pesos_i(4405) := b"1111111111111111_1111111111111111_1110001000011100_0001001001100100"; -- -0.11675915772509414
	pesos_i(4406) := b"0000000000000000_0000000000000000_0011000101100110_0100011001011010"; -- 0.1929668397182854
	pesos_i(4407) := b"0000000000000000_0000000000000000_0000011101100101_1000100000011101"; -- 0.028893000641439466
	pesos_i(4408) := b"1111111111111111_1111111111111111_1100101100011011_0110011110110110"; -- -0.20661308114645152
	pesos_i(4409) := b"0000000000000000_0000000000000000_0010001111001100_0001110000000010"; -- 0.1398332122797792
	pesos_i(4410) := b"1111111111111111_1111111111111111_1101100000110100_1100111101101001"; -- -0.15544418033416177
	pesos_i(4411) := b"1111111111111111_1111111111111111_1111111111001110_1110100101100000"; -- -0.0007490292218547412
	pesos_i(4412) := b"0000000000000000_0000000000000000_0001000000011110_0010100011000011"; -- 0.06296019335864733
	pesos_i(4413) := b"1111111111111111_1111111111111111_1110100100010000_1000010011000100"; -- -0.08959169583944064
	pesos_i(4414) := b"0000000000000000_0000000000000000_0010100101011000_1000110101101010"; -- 0.16150745243647832
	pesos_i(4415) := b"1111111111111111_1111111111111111_1101110001101000_0100011100111000"; -- -0.13903384089739765
	pesos_i(4416) := b"1111111111111111_1111111111111111_1110000101001010_1110011011011111"; -- -0.11995083869770098
	pesos_i(4417) := b"0000000000000000_0000000000000000_0001101101011101_0111101000100010"; -- 0.10689509709001088
	pesos_i(4418) := b"0000000000000000_0000000000000000_0010000100101101_1010011110000001"; -- 0.12960287945742793
	pesos_i(4419) := b"0000000000000000_0000000000000000_0010110110111110_1101010110100000"; -- 0.17869315303532138
	pesos_i(4420) := b"0000000000000000_0000000000000000_0011100111000010_0001001110010010"; -- 0.22561762153298787
	pesos_i(4421) := b"0000000000000000_0000000000000000_0001101110010010_1111111100001000"; -- 0.10771173423202189
	pesos_i(4422) := b"1111111111111111_1111111111111111_1110101000101001_0101010011101111"; -- -0.08530682715603437
	pesos_i(4423) := b"1111111111111111_1111111111111111_1101110111011001_1100001011011111"; -- -0.13339597762612068
	pesos_i(4424) := b"1111111111111111_1111111111111111_1111010101101100_1010110001011010"; -- -0.04131052786993935
	pesos_i(4425) := b"1111111111111111_1111111111111111_1100110111111000_0101010001011111"; -- -0.19542954148335012
	pesos_i(4426) := b"0000000000000000_0000000000000000_0000101000010010_1000001101001100"; -- 0.03934498401535236
	pesos_i(4427) := b"1111111111111111_1111111111111111_1111010010101010_1110110000100111"; -- -0.044266930072193005
	pesos_i(4428) := b"0000000000000000_0000000000000000_0000110001100010_0000100111110011"; -- 0.048370954323001994
	pesos_i(4429) := b"0000000000000000_0000000000000000_0000000111000000_0100000010010011"; -- 0.006839786491030592
	pesos_i(4430) := b"0000000000000000_0000000000000000_0001110100000000_0011101100001101"; -- 0.11328476960238967
	pesos_i(4431) := b"0000000000000000_0000000000000000_0000111000110111_0100000000101111"; -- 0.05553055908613598
	pesos_i(4432) := b"0000000000000000_0000000000000000_0010001101111110_1100101011011010"; -- 0.13865344840223603
	pesos_i(4433) := b"0000000000000000_0000000000000000_0010100011110000_0010010111100110"; -- 0.1599143682894022
	pesos_i(4434) := b"0000000000000000_0000000000000000_0001101001111000_0101101010110100"; -- 0.10339896094614046
	pesos_i(4435) := b"1111111111111111_1111111111111111_1110111111010011_1100000001010111"; -- -0.06317518114374467
	pesos_i(4436) := b"1111111111111111_1111111111111111_1111100100010101_1000011011111010"; -- -0.027015270137021097
	pesos_i(4437) := b"1111111111111111_1111111111111111_1110100101101100_1010001111100010"; -- -0.08818603266420508
	pesos_i(4438) := b"1111111111111111_1111111111111111_1111101001010011_1110100111100111"; -- -0.0221570788165442
	pesos_i(4439) := b"1111111111111111_1111111111111111_1110011001100101_1111101011011000"; -- -0.10000641085253394
	pesos_i(4440) := b"0000000000000000_0000000000000000_0000100100101101_0001011100001110"; -- 0.035844269686272065
	pesos_i(4441) := b"0000000000000000_0000000000000000_0010100011111111_0011001010100001"; -- 0.16014400885835148
	pesos_i(4442) := b"1111111111111111_1111111111111111_1110111101010011_0101011001100000"; -- -0.06513462209118692
	pesos_i(4443) := b"0000000000000000_0000000000000000_0010100010110010_1101001011011101"; -- 0.15897863278293822
	pesos_i(4444) := b"0000000000000000_0000000000000000_0001101001001001_0100101000101000"; -- 0.10268081167095723
	pesos_i(4445) := b"0000000000000000_0000000000000000_0010000011110110_0101010110101001"; -- 0.12875876777529893
	pesos_i(4446) := b"1111111111111111_1111111111111111_1111011001000010_0101101000110000"; -- -0.038050044307637754
	pesos_i(4447) := b"1111111111111111_1111111111111111_1111000101101000_1010000101000010"; -- -0.05699722420072335
	pesos_i(4448) := b"1111111111111111_1111111111111111_1110110111101010_0001010100010011"; -- -0.07064693723664867
	pesos_i(4449) := b"0000000000000000_0000000000000000_0001111100011101_1011011110011000"; -- 0.12154719786378215
	pesos_i(4450) := b"0000000000000000_0000000000000000_0010111101001000_1100010101001001"; -- 0.18470414191118653
	pesos_i(4451) := b"0000000000000000_0000000000000000_0000010111000100_1110101100000001"; -- 0.022535979961610605
	pesos_i(4452) := b"0000000000000000_0000000000000000_0011100001111000_1110110001001011"; -- 0.22059513877079018
	pesos_i(4453) := b"1111111111111111_1111111111111111_1101001111110101_1010000001011110"; -- -0.17203328815814647
	pesos_i(4454) := b"0000000000000000_0000000000000000_0001010001101011_0010110000011110"; -- 0.07976032007325878
	pesos_i(4455) := b"1111111111111111_1111111111111111_1101100111100000_1010000001010101"; -- -0.14891622473819646
	pesos_i(4456) := b"1111111111111111_1111111111111111_1101111000011011_0101101101000100"; -- -0.13239507274019366
	pesos_i(4457) := b"1111111111111111_1111111111111111_1111110101100110_1000000111001000"; -- -0.010154617883803079
	pesos_i(4458) := b"1111111111111111_1111111111111111_1101100000001001_0001111000101100"; -- -0.1561108725103323
	pesos_i(4459) := b"1111111111111111_1111111111111111_1111101111110110_1100011100111001"; -- -0.01576571329388231
	pesos_i(4460) := b"1111111111111111_1111111111111111_1111101000000110_1010110000001101"; -- -0.023335692167054507
	pesos_i(4461) := b"1111111111111111_1111111111111111_1110101000000110_0111111011100001"; -- -0.08583838478138074
	pesos_i(4462) := b"1111111111111111_1111111111111111_1110111000000110_0101010000011110"; -- -0.07021593360358985
	pesos_i(4463) := b"0000000000000000_0000000000000000_0001001001010001_0000110111111000"; -- 0.0715492945388134
	pesos_i(4464) := b"1111111111111111_1111111111111111_1110000100100000_0000000100100101"; -- -0.1206054004912823
	pesos_i(4465) := b"0000000000000000_0000000000000000_0000111100101011_1000110000101100"; -- 0.05925823273526743
	pesos_i(4466) := b"1111111111111111_1111111111111111_1111000111101111_0010111110110100"; -- -0.054944056076100097
	pesos_i(4467) := b"1111111111111111_1111111111111111_1101101001100011_0010001100100001"; -- -0.14692478596725772
	pesos_i(4468) := b"1111111111111111_1111111111111111_1111111000001110_0110010010100110"; -- -0.007592877758892823
	pesos_i(4469) := b"1111111111111111_1111111111111111_1111111010011010_0100100100110011"; -- -0.005458283585496817
	pesos_i(4470) := b"1111111111111111_1111111111111111_1110110100011000_0010101001100001"; -- -0.07385001305929707
	pesos_i(4471) := b"1111111111111111_1111111111111111_1101010111111101_1111011010000110"; -- -0.16409358234047025
	pesos_i(4472) := b"1111111111111111_1111111111111111_1110100111100110_0111011000111111"; -- -0.08632718042219127
	pesos_i(4473) := b"1111111111111111_1111111111111111_1110110111000000_1011010101001000"; -- -0.07127825734915993
	pesos_i(4474) := b"1111111111111111_1111111111111111_1111101001010011_0011000011110111"; -- -0.022168102016570542
	pesos_i(4475) := b"1111111111111111_1111111111111111_1111011010001000_1101010101111001"; -- -0.03697458068840239
	pesos_i(4476) := b"1111111111111111_1111111111111111_1110101110001101_1001011110000001"; -- -0.07987073051710926
	pesos_i(4477) := b"1111111111111111_1111111111111111_1101010110111001_0110110000101100"; -- -0.16513942659002248
	pesos_i(4478) := b"1111111111111111_1111111111111111_1110100101001111_0001101111101111"; -- -0.08863664057706004
	pesos_i(4479) := b"0000000000000000_0000000000000000_0000000011100100_0001110111001001"; -- 0.003480779210182029
	pesos_i(4480) := b"0000000000000000_0000000000000000_0000000011100000_0100010011011000"; -- 0.0034220721152894897
	pesos_i(4481) := b"0000000000000000_0000000000000000_0000001110011101_1110000110000001"; -- 0.014127820966814812
	pesos_i(4482) := b"1111111111111111_1111111111111111_1111000000001101_0110011101001000"; -- -0.06229547962508385
	pesos_i(4483) := b"0000000000000000_0000000000000000_0010100101000100_1000011110101010"; -- 0.16120193387728748
	pesos_i(4484) := b"0000000000000000_0000000000000000_0000100110001110_1101101010010110"; -- 0.037336026858632694
	pesos_i(4485) := b"0000000000000000_0000000000000000_0000111000010000_1111100100001101"; -- 0.054946485125028206
	pesos_i(4486) := b"1111111111111111_1111111111111111_1101111011110101_0001010011001011"; -- -0.1290728572296823
	pesos_i(4487) := b"0000000000000000_0000000000000000_0000001101000000_1101111101001111"; -- 0.012708622647015114
	pesos_i(4488) := b"0000000000000000_0000000000000000_0001000100011111_0100100100001101"; -- 0.06688362657693996
	pesos_i(4489) := b"0000000000000000_0000000000000000_0001000000100110_0101001100110111"; -- 0.06308479403413429
	pesos_i(4490) := b"0000000000000000_0000000000000000_0010011000101011_1000010110001100"; -- 0.1491015879400422
	pesos_i(4491) := b"0000000000000000_0000000000000000_0000000100000101_1011111011101101"; -- 0.003993924061475948
	pesos_i(4492) := b"0000000000000000_0000000000000000_0000100001100011_0001001000001011"; -- 0.03276169559775854
	pesos_i(4493) := b"0000000000000000_0000000000000000_0010011001110000_0011010001011011"; -- 0.15014960501135796
	pesos_i(4494) := b"0000000000000000_0000000000000000_0010010110111011_0011101000010100"; -- 0.1473881053535862
	pesos_i(4495) := b"1111111111111111_1111111111111111_1110000000111011_1011101110000101"; -- -0.12408855440335598
	pesos_i(4496) := b"1111111111111111_1111111111111111_1111110110101010_1011011110001011"; -- -0.009113815880195358
	pesos_i(4497) := b"1111111111111111_1111111111111111_1101001011111100_0110000110000010"; -- -0.17583647312932657
	pesos_i(4498) := b"0000000000000000_0000000000000000_0000111010001100_1001011111010101"; -- 0.05683278030127613
	pesos_i(4499) := b"1111111111111111_1111111111111111_1110100101011100_0000001000000010"; -- -0.08843982170894822
	pesos_i(4500) := b"0000000000000000_0000000000000000_0001100111100101_0001011000001111"; -- 0.10115182745375569
	pesos_i(4501) := b"1111111111111111_1111111111111111_1101110110011111_0000001010111110"; -- -0.13429243910692712
	pesos_i(4502) := b"0000000000000000_0000000000000000_0000000000110011_1010110001110010"; -- 0.0007884767629022835
	pesos_i(4503) := b"1111111111111111_1111111111111111_1110110111001010_0010001010100111"; -- -0.0711344091117524
	pesos_i(4504) := b"1111111111111111_1111111111111111_1110000111111100_1101101010110111"; -- -0.11723549873761897
	pesos_i(4505) := b"1111111111111111_1111111111111111_1101100010010110_0101111100111111"; -- -0.15395550461865123
	pesos_i(4506) := b"1111111111111111_1111111111111111_1111100000000101_0100111100011101"; -- -0.03116899043414446
	pesos_i(4507) := b"1111111111111111_1111111111111111_1110000001110001_1000011000000111"; -- -0.12326776822164115
	pesos_i(4508) := b"1111111111111111_1111111111111111_1100111010001110_0000011100011011"; -- -0.19314532842426277
	pesos_i(4509) := b"1111111111111111_1111111111111111_1100110011000011_0010011110010010"; -- -0.20014717751548589
	pesos_i(4510) := b"1111111111111111_1111111111111111_1110011001100001_0000011001100111"; -- -0.10008201588738297
	pesos_i(4511) := b"1111111111111111_1111111111111111_1101110110010110_0100100100011101"; -- -0.1344255736726233
	pesos_i(4512) := b"1111111111111111_1111111111111111_1101110101110110_0111001100101110"; -- -0.13491134762601578
	pesos_i(4513) := b"1111111111111111_1111111111111111_1111111010110100_0010111001000111"; -- -0.005063159632090148
	pesos_i(4514) := b"1111111111111111_1111111111111111_1101101111000101_1111111111101100"; -- -0.14151001435617033
	pesos_i(4515) := b"1111111111111111_1111111111111111_1110010100110100_0110011110110001"; -- -0.10466911237087184
	pesos_i(4516) := b"0000000000000000_0000000000000000_0011001101101100_0001001100001010"; -- 0.2008678340200044
	pesos_i(4517) := b"1111111111111111_1111111111111111_1101111110000101_0010011111111010"; -- -0.12687444817562868
	pesos_i(4518) := b"1111111111111111_1111111111111111_1101001000110000_1000001000111100"; -- -0.17894731558844756
	pesos_i(4519) := b"0000000000000000_0000000000000000_0001010101001101_1010001011111111"; -- 0.08321589206059744
	pesos_i(4520) := b"1111111111111111_1111111111111111_1111010100100100_1010001001001101"; -- -0.042409759789434974
	pesos_i(4521) := b"0000000000000000_0000000000000000_0000101011011011_1100100110100111"; -- 0.04241619422105291
	pesos_i(4522) := b"0000000000000000_0000000000000000_0001000110011111_0011011110110100"; -- 0.0688357176397218
	pesos_i(4523) := b"0000000000000000_0000000000000000_0010001111000111_0101101010100001"; -- 0.1397606508774957
	pesos_i(4524) := b"0000000000000000_0000000000000000_0001111000000110_1001011100000111"; -- 0.11728805472955285
	pesos_i(4525) := b"1111111111111111_1111111111111111_1111110010101001_1101111101011110"; -- -0.013032950813325749
	pesos_i(4526) := b"0000000000000000_0000000000000000_0001110011000000_0001011110010100"; -- 0.11230609276769893
	pesos_i(4527) := b"1111111111111111_1111111111111111_1101101101111101_0001001011010111"; -- -0.14262277842080948
	pesos_i(4528) := b"1111111111111111_1111111111111111_1101001001111111_1010110010110101"; -- -0.17773933953143692
	pesos_i(4529) := b"0000000000000000_0000000000000000_0000101100110011_0000111100110100"; -- 0.04374785447428861
	pesos_i(4530) := b"0000000000000000_0000000000000000_0000010111111110_1110000001001011"; -- 0.02342035142719337
	pesos_i(4531) := b"0000000000000000_0000000000000000_0000011101111110_1110110101110010"; -- 0.029280510353726308
	pesos_i(4532) := b"0000000000000000_0000000000000000_0001011010100101_1101100011011100"; -- 0.08846812600773674
	pesos_i(4533) := b"0000000000000000_0000000000000000_0010000010011110_1001010101100101"; -- 0.12741979329238617
	pesos_i(4534) := b"1111111111111111_1111111111111111_1101111111000010_0010001100101000"; -- -0.12594394937742928
	pesos_i(4535) := b"1111111111111111_1111111111111111_1101101001011011_0000100110100001"; -- -0.14704837621953779
	pesos_i(4536) := b"1111111111111111_1111111111111111_1101110110101010_0111100110001101"; -- -0.1341175109757484
	pesos_i(4537) := b"1111111111111111_1111111111111111_1100110100110110_0001100111011101"; -- -0.19839323381815308
	pesos_i(4538) := b"0000000000000000_0000000000000000_0001100011100111_0100000100110101"; -- 0.09727866702908693
	pesos_i(4539) := b"0000000000000000_0000000000000000_0000111111101100_0110110010100000"; -- 0.06220129880633124
	pesos_i(4540) := b"1111111111111111_1111111111111111_1101010000100100_0110111111001110"; -- -0.17131901953223164
	pesos_i(4541) := b"0000000000000000_0000000000000000_0000011001010010_0110011011001111"; -- 0.02469484853751236
	pesos_i(4542) := b"1111111111111111_1111111111111111_1101001010010110_1100101101011100"; -- -0.1773865605292213
	pesos_i(4543) := b"1111111111111111_1111111111111111_1101010111011110_0000010011101010"; -- -0.16458100596558528
	pesos_i(4544) := b"0000000000000000_0000000000000000_0000000111101111_1100001101110000"; -- 0.007564749629211194
	pesos_i(4545) := b"1111111111111111_1111111111111111_1101111100010101_0000111011110011"; -- -0.12858492447996808
	pesos_i(4546) := b"0000000000000000_0000000000000000_0010101110010110_0010111011000100"; -- 0.1702603556981381
	pesos_i(4547) := b"1111111111111111_1111111111111111_1101100000001000_0101110010100001"; -- -0.15612240853687073
	pesos_i(4548) := b"1111111111111111_1111111111111111_1101101011110011_1110000111001000"; -- -0.14471615665006074
	pesos_i(4549) := b"0000000000000000_0000000000000000_0000100111001101_1001000010111100"; -- 0.03829292865623203
	pesos_i(4550) := b"1111111111111111_1111111111111111_1110001111001101_1001011001011000"; -- -0.11014423698131579
	pesos_i(4551) := b"0000000000000000_0000000000000000_0001101000110011_0101111011011110"; -- 0.10234635277204282
	pesos_i(4552) := b"1111111111111111_1111111111111111_1101000011100101_0101000001111000"; -- -0.1840009409647417
	pesos_i(4553) := b"0000000000000000_0000000000000000_0001101011000111_0101101111111100"; -- 0.10460448167748719
	pesos_i(4554) := b"1111111111111111_1111111111111111_1110011111001111_0111010111100000"; -- -0.09449065476907274
	pesos_i(4555) := b"0000000000000000_0000000000000000_0000011101011001_1010111011010000"; -- 0.028712201914698386
	pesos_i(4556) := b"0000000000000000_0000000000000000_0001001110111111_1011000111001100"; -- 0.07714377624817194
	pesos_i(4557) := b"0000000000000000_0000000000000000_0001101100100000_0100001000101001"; -- 0.10596097471121353
	pesos_i(4558) := b"1111111111111111_1111111111111111_1101111011000000_1111110011010111"; -- -0.12986774214383845
	pesos_i(4559) := b"1111111111111111_1111111111111111_1110100110110001_1101101100110000"; -- -0.08712987980593973
	pesos_i(4560) := b"0000000000000000_0000000000000000_0010100101000111_0100010001101010"; -- 0.1612437018433722
	pesos_i(4561) := b"0000000000000000_0000000000000000_0000001111001110_1110111111001110"; -- 0.014876353955218634
	pesos_i(4562) := b"0000000000000000_0000000000000000_0010100101000001_0011100000110110"; -- 0.16115142181845707
	pesos_i(4563) := b"0000000000000000_0000000000000000_0010001111110110_0010011101011111"; -- 0.14047475890536892
	pesos_i(4564) := b"1111111111111111_1111111111111111_1111101111111100_1111100111011000"; -- -0.015671143395458862
	pesos_i(4565) := b"0000000000000000_0000000000000000_0010110000101100_0101000101101110"; -- 0.17255124033692637
	pesos_i(4566) := b"1111111111111111_1111111111111111_1101101101110001_0011111111000101"; -- -0.14280320594599494
	pesos_i(4567) := b"1111111111111111_1111111111111111_1111000000101000_1101000001001000"; -- -0.06187723396048131
	pesos_i(4568) := b"0000000000000000_0000000000000000_0010101010110100_0001101110111110"; -- 0.1668107355257308
	pesos_i(4569) := b"1111111111111111_1111111111111111_1100110111001101_1100001111111101"; -- -0.19607901651952048
	pesos_i(4570) := b"0000000000000000_0000000000000000_0000101101111100_1111101010000001"; -- 0.04487577092920185
	pesos_i(4571) := b"1111111111111111_1111111111111111_1111010011101101_0000000011101111"; -- -0.04325861137187705
	pesos_i(4572) := b"1111111111111111_1111111111111111_1110011011111111_0111011110001111"; -- -0.09766438251719105
	pesos_i(4573) := b"0000000000000000_0000000000000000_0000000110110100_1000110011111010"; -- 0.006661234819331608
	pesos_i(4574) := b"0000000000000000_0000000000000000_0001010101110101_1011010101110101"; -- 0.0838273439430556
	pesos_i(4575) := b"1111111111111111_1111111111111111_1111110001001101_0010111100001000"; -- -0.014447269861842658
	pesos_i(4576) := b"1111111111111111_1111111111111111_1110011111101101_1000011001111101"; -- -0.09403190075570743
	pesos_i(4577) := b"0000000000000000_0000000000000000_0000101101110011_0101001000101110"; -- 0.044728409055954134
	pesos_i(4578) := b"0000000000000000_0000000000000000_0000100010000010_0010011000011101"; -- 0.033235914306038714
	pesos_i(4579) := b"1111111111111111_1111111111111111_1110010001111010_1110101010101000"; -- -0.10749944119039427
	pesos_i(4580) := b"0000000000000000_0000000000000000_0001001111010010_1111011110001001"; -- 0.07743784993766369
	pesos_i(4581) := b"1111111111111111_1111111111111111_1111110000101010_0110011011110001"; -- -0.014977994966433983
	pesos_i(4582) := b"1111111111111111_1111111111111111_1110110000111100_1110101000110001"; -- -0.07719551368423008
	pesos_i(4583) := b"0000000000000000_0000000000000000_0001110111100110_1110000111001011"; -- 0.11680422978325747
	pesos_i(4584) := b"1111111111111111_1111111111111111_1101000000101000_1111011011001010"; -- -0.18687493868508206
	pesos_i(4585) := b"0000000000000000_0000000000000000_0000000000010010_1101011101111100"; -- 0.00028750196086432014
	pesos_i(4586) := b"1111111111111111_1111111111111111_1101100010110110_1110111010010000"; -- -0.15345868097746124
	pesos_i(4587) := b"1111111111111111_1111111111111111_1111101101001111_1111101101011111"; -- -0.018310822794183324
	pesos_i(4588) := b"0000000000000000_0000000000000000_0001010110000000_1101000000000001"; -- 0.08399677308474984
	pesos_i(4589) := b"1111111111111111_1111111111111111_1101110011111111_0000111011000001"; -- -0.136733129462913
	pesos_i(4590) := b"0000000000000000_0000000000000000_0000111111011000_1010111111110111"; -- 0.06190013667439965
	pesos_i(4591) := b"0000000000000000_0000000000000000_0001001111101110_0010110001000010"; -- 0.07785297974582148
	pesos_i(4592) := b"0000000000000000_0000000000000000_0011000001010100_1010000001010110"; -- 0.18879129498074365
	pesos_i(4593) := b"0000000000000000_0000000000000000_0000111101010111_0111011111001000"; -- 0.059928404168730486
	pesos_i(4594) := b"0000000000000000_0000000000000000_0000110111111010_0000000010011001"; -- 0.05459598280817682
	pesos_i(4595) := b"1111111111111111_1111111111111111_1111110011010010_0011110011100001"; -- -0.012417025569219807
	pesos_i(4596) := b"1111111111111111_1111111111111111_1101110100101011_0110101011001111"; -- -0.1360562557923951
	pesos_i(4597) := b"0000000000000000_0000000000000000_0001101010101010_1100000011111111"; -- 0.10416799759728834
	pesos_i(4598) := b"1111111111111111_1111111111111111_1100111011110111_1000100111110110"; -- -0.19153535594863952
	pesos_i(4599) := b"0000000000000000_0000000000000000_0001110110101011_1111111110000100"; -- 0.11590573291035094
	pesos_i(4600) := b"0000000000000000_0000000000000000_0010110100100010_0011101101010000"; -- 0.1763035842247648
	pesos_i(4601) := b"0000000000000000_0000000000000000_0001111000111001_0101000001101001"; -- 0.11806204372662366
	pesos_i(4602) := b"1111111111111111_1111111111111111_1101110001011111_1000000100011001"; -- -0.13916772025254295
	pesos_i(4603) := b"0000000000000000_0000000000000000_0001101001101011_1010101011010001"; -- 0.1032053717732896
	pesos_i(4604) := b"0000000000000000_0000000000000000_0010011111000000_0001001100101110"; -- 0.15527458070352398
	pesos_i(4605) := b"1111111111111111_1111111111111111_1101111001001110_1101101000000010"; -- -0.13160932007159593
	pesos_i(4606) := b"1111111111111111_1111111111111111_1110010001010010_1111000010111101"; -- -0.10810943023628113
	pesos_i(4607) := b"1111111111111111_1111111111111111_1110110010010100_1010010000000111"; -- -0.07585692237129299
	pesos_i(4608) := b"1111111111111111_1111111111111111_1111010010111111_0100010110000001"; -- -0.043956428492805996
	pesos_i(4609) := b"1111111111111111_1111111111111111_1110000110101011_0010101010111111"; -- -0.11848194916789212
	pesos_i(4610) := b"0000000000000000_0000000000000000_0010010110111000_1111001010110111"; -- 0.14735333406296772
	pesos_i(4611) := b"1111111111111111_1111111111111111_1110000111101100_1000010010011001"; -- -0.11748477245413533
	pesos_i(4612) := b"1111111111111111_1111111111111111_1101010100000001_1001011101011000"; -- -0.16794447045968008
	pesos_i(4613) := b"1111111111111111_1111111111111111_1111011010000011_0100100011010000"; -- -0.03705925864999722
	pesos_i(4614) := b"0000000000000000_0000000000000000_0000100000000111_1110101000000001"; -- 0.031370759164718175
	pesos_i(4615) := b"0000000000000000_0000000000000000_0000011101100011_1010001101101101"; -- 0.02886411101963474
	pesos_i(4616) := b"1111111111111111_1111111111111111_1110111000001010_1111100101101010"; -- -0.07014504579740816
	pesos_i(4617) := b"0000000000000000_0000000000000000_0010010000000101_1101101010000110"; -- 0.14071431890748007
	pesos_i(4618) := b"0000000000000000_0000000000000000_0001011101011011_0111110100100100"; -- 0.09123975868321174
	pesos_i(4619) := b"1111111111111111_1111111111111111_1110010111001100_0010010111100011"; -- -0.10235369879094124
	pesos_i(4620) := b"1111111111111111_1111111111111111_1110101110010011_0100111010010001"; -- -0.07978352506295855
	pesos_i(4621) := b"1111111111111111_1111111111111111_1101000111101001_1011101011101101"; -- -0.18002731051294746
	pesos_i(4622) := b"1111111111111111_1111111111111111_1110010101011111_1111110101111001"; -- -0.10400405694479392
	pesos_i(4623) := b"1111111111111111_1111111111111111_1110000011101001_1001100011010010"; -- -0.12143559327147799
	pesos_i(4624) := b"1111111111111111_1111111111111111_1100111110011110_1101010001001001"; -- -0.1889827080759928
	pesos_i(4625) := b"1111111111111111_1111111111111111_1110000011000000_1000001000110111"; -- -0.12206255103436017
	pesos_i(4626) := b"1111111111111111_1111111111111111_1111101101010100_0100101100110011"; -- -0.018245029425154012
	pesos_i(4627) := b"1111111111111111_1111111111111111_1111111011100011_1101111110100010"; -- -0.0043354253543651826
	pesos_i(4628) := b"1111111111111111_1111111111111111_1111101011010111_0011011100101000"; -- -0.020153572848166892
	pesos_i(4629) := b"0000000000000000_0000000000000000_0000010110110100_1010110110011110"; -- 0.022288180402142487
	pesos_i(4630) := b"1111111111111111_1111111111111111_1111011100100010_0011110000011100"; -- -0.03463386827377467
	pesos_i(4631) := b"0000000000000000_0000000000000000_0000011010101111_1001101111000101"; -- 0.026117072668575266
	pesos_i(4632) := b"0000000000000000_0000000000000000_0001011000010111_0101010111001010"; -- 0.0862935656756867
	pesos_i(4633) := b"1111111111111111_1111111111111111_1110011110111101_1111010100100100"; -- -0.09475772744775823
	pesos_i(4634) := b"1111111111111111_1111111111111111_1110100110001001_0100101111100100"; -- -0.08774877237283946
	pesos_i(4635) := b"0000000000000000_0000000000000000_0000011000010111_1001000001110001"; -- 0.023797061523380958
	pesos_i(4636) := b"0000000000000000_0000000000000000_0000101010100111_1100000010011011"; -- 0.041622197952811996
	pesos_i(4637) := b"0000000000000000_0000000000000000_0011100100101101_1010100100100000"; -- 0.2233529762420373
	pesos_i(4638) := b"0000000000000000_0000000000000000_0001001111001100_0000011000101111"; -- 0.07733191153523963
	pesos_i(4639) := b"1111111111111111_1111111111111111_1111111111110100_0010101100000011"; -- -0.00018054185726047495
	pesos_i(4640) := b"1111111111111111_1111111111111111_1101001101100000_0000110111010111"; -- -0.17431558134648223
	pesos_i(4641) := b"1111111111111111_1111111111111111_1111100110111100_1010010001101010"; -- -0.024465297754467333
	pesos_i(4642) := b"1111111111111111_1111111111111111_1110111111001001_1101111001011110"; -- -0.06332597916943405
	pesos_i(4643) := b"0000000000000000_0000000000000000_0001001001100000_1010100100111001"; -- 0.07178743018657296
	pesos_i(4644) := b"0000000000000000_0000000000000000_0011111101101001_1001011011000001"; -- 0.24770490857470207
	pesos_i(4645) := b"1111111111111111_1111111111111111_1111100110100011_1100101011111001"; -- -0.024844469239952566
	pesos_i(4646) := b"1111111111111111_1111111111111111_1110011100001111_1101100011010101"; -- -0.0974144438983965
	pesos_i(4647) := b"1111111111111111_1111111111111111_1110110010010000_0001010100011111"; -- -0.07592647550098945
	pesos_i(4648) := b"1111111111111111_1111111111111111_1111000100110111_1001010001110010"; -- -0.05774566868158359
	pesos_i(4649) := b"0000000000000000_0000000000000000_0000111111011011_1100101101000100"; -- 0.061947540341178144
	pesos_i(4650) := b"0000000000000000_0000000000000000_0010010000011011_1001010010100101"; -- 0.14104584724638064
	pesos_i(4651) := b"1111111111111111_1111111111111111_1110000000111010_1010001001111100"; -- -0.12410530543607415
	pesos_i(4652) := b"0000000000000000_0000000000000000_0000000001110001_0010001000110101"; -- 0.0017262819667674854
	pesos_i(4653) := b"0000000000000000_0000000000000000_0010001101111111_1100110000010001"; -- 0.1386687796252221
	pesos_i(4654) := b"1111111111111111_1111111111111111_1110000000101110_1010100011111100"; -- -0.12428802350998983
	pesos_i(4655) := b"1111111111111111_1111111111111111_1110111010110000_1001001001111010"; -- -0.06761822237446424
	pesos_i(4656) := b"0000000000000000_0000000000000000_0010110100011111_1101110000000011"; -- 0.17626738617147933
	pesos_i(4657) := b"0000000000000000_0000000000000000_0010001000001110_0100011110110011"; -- 0.1330303965809804
	pesos_i(4658) := b"1111111111111111_1111111111111111_1111000111100001_1000110100011110"; -- -0.05515211131077011
	pesos_i(4659) := b"0000000000000000_0000000000000000_0000000000100010_1001110011111010"; -- 0.0005281552983525391
	pesos_i(4660) := b"0000000000000000_0000000000000000_0000101101101111_0000100010011011"; -- 0.04466298841861547
	pesos_i(4661) := b"0000000000000000_0000000000000000_0010001101001011_1101100110111111"; -- 0.13787613784398592
	pesos_i(4662) := b"1111111111111111_1111111111111111_1101010000010000_1101001001101101"; -- -0.17161831697453475
	pesos_i(4663) := b"1111111111111111_1111111111111111_1101111010100101_1010010000011111"; -- -0.13028501746373303
	pesos_i(4664) := b"1111111111111111_1111111111111111_1110010101100101_1101010000111101"; -- -0.10391496182703416
	pesos_i(4665) := b"1111111111111111_1111111111111111_1101001010101010_0111101000010111"; -- -0.17708622863005916
	pesos_i(4666) := b"1111111111111111_1111111111111111_1101111010010111_0011101001001001"; -- -0.1305049487407306
	pesos_i(4667) := b"1111111111111111_1111111111111111_1110011100000111_1100101110110101"; -- -0.09753729661050094
	pesos_i(4668) := b"0000000000000000_0000000000000000_0010010011000110_1011111101011101"; -- 0.14365764628785607
	pesos_i(4669) := b"0000000000000000_0000000000000000_0000111111101110_1101110101001100"; -- 0.06223853223153679
	pesos_i(4670) := b"1111111111111111_1111111111111111_1101101000101001_1011000100001110"; -- -0.14780133626935446
	pesos_i(4671) := b"0000000000000000_0000000000000000_0001010000001100_0100100000011001"; -- 0.07831240281673378
	pesos_i(4672) := b"0000000000000000_0000000000000000_0001101000011011_0100001111000001"; -- 0.10197852580442536
	pesos_i(4673) := b"1111111111111111_1111111111111111_1101101010100000_1001011111010001"; -- -0.14598704480903404
	pesos_i(4674) := b"0000000000000000_0000000000000000_0001100100011101_1001011111000000"; -- 0.0981077999028647
	pesos_i(4675) := b"0000000000000000_0000000000000000_0000100010101110_0000100001101001"; -- 0.03390553068985579
	pesos_i(4676) := b"1111111111111111_1111111111111111_1101100011111000_0101100010001011"; -- -0.1524605426950976
	pesos_i(4677) := b"0000000000000000_0000000000000000_0001110011110010_1010100000110001"; -- 0.11307765193889299
	pesos_i(4678) := b"1111111111111111_1111111111111111_1110011010101001_1101111001100010"; -- -0.09897050953808219
	pesos_i(4679) := b"1111111111111111_1111111111111111_1111000011000100_1010101001000111"; -- -0.05949912799148953
	pesos_i(4680) := b"0000000000000000_0000000000000000_0001010010001010_0001111100011100"; -- 0.08023256719492866
	pesos_i(4681) := b"0000000000000000_0000000000000000_0001001101010001_1100101011101110"; -- 0.07546680757002477
	pesos_i(4682) := b"0000000000000000_0000000000000000_0010000111001111_0010111101100100"; -- 0.13206764409477023
	pesos_i(4683) := b"0000000000000000_0000000000000000_0000000110110000_0010100100001111"; -- 0.006594244263612281
	pesos_i(4684) := b"1111111111111111_1111111111111111_1110001110010111_1100010110100111"; -- -0.11096539183157349
	pesos_i(4685) := b"0000000000000000_0000000000000000_0000110101100100_0000100001011111"; -- 0.052307627932532005
	pesos_i(4686) := b"0000000000000000_0000000000000000_0000111111100111_0111110000110100"; -- 0.06212593326448615
	pesos_i(4687) := b"0000000000000000_0000000000000000_0001110110000011_0001110001011001"; -- 0.11528184090851534
	pesos_i(4688) := b"0000000000000000_0000000000000000_0010100101100101_0110101011111101"; -- 0.16170376474847853
	pesos_i(4689) := b"1111111111111111_1111111111111111_1111010000000101_1010000011001100"; -- -0.04678912173638495
	pesos_i(4690) := b"1111111111111111_1111111111111111_1111010101011111_1011110110010001"; -- -0.04150786611082193
	pesos_i(4691) := b"1111111111111111_1111111111111111_1111000011111111_0100010000111000"; -- -0.05860494265029926
	pesos_i(4692) := b"1111111111111111_1111111111111111_1111010001100111_0101100110010000"; -- -0.04529800644100728
	pesos_i(4693) := b"1111111111111111_1111111111111111_1101110110011101_0100001111111001"; -- -0.13431906867008994
	pesos_i(4694) := b"0000000000000000_0000000000000000_0000001010000101_1010100010011000"; -- 0.009851967849832333
	pesos_i(4695) := b"1111111111111111_1111111111111111_1110111111111010_1001001101001100"; -- -0.06258277327271011
	pesos_i(4696) := b"1111111111111111_1111111111111111_1101011111010010_0011101101010111"; -- -0.156948367467656
	pesos_i(4697) := b"0000000000000000_0000000000000000_0010110101010011_0010010110011011"; -- 0.17704997094515984
	pesos_i(4698) := b"1111111111111111_1111111111111111_1111011101111101_1010010010001111"; -- -0.03323909279665169
	pesos_i(4699) := b"0000000000000000_0000000000000000_0010110101111000_0001010011010111"; -- 0.1776135469404805
	pesos_i(4700) := b"1111111111111111_1111111111111111_1110000011011010_1000101001010111"; -- -0.12166533829473732
	pesos_i(4701) := b"0000000000000000_0000000000000000_0010111100001011_1111011101011101"; -- 0.18377634060599052
	pesos_i(4702) := b"1111111111111111_1111111111111111_1101111001011111_1011111100101010"; -- -0.1313515207019971
	pesos_i(4703) := b"1111111111111111_1111111111111111_1111111011111110_0000110010100110"; -- -0.0039360137593039005
	pesos_i(4704) := b"1111111111111111_1111111111111111_1101011000011110_1011011101111111"; -- -0.1635937991931531
	pesos_i(4705) := b"1111111111111111_1111111111111111_1101100001010000_0100000011010001"; -- -0.15502543353417508
	pesos_i(4706) := b"0000000000000000_0000000000000000_0010000000000101_0101110100101100"; -- 0.12508184735867173
	pesos_i(4707) := b"1111111111111111_1111111111111111_1111101101001000_1010010001011001"; -- -0.01842282136213028
	pesos_i(4708) := b"1111111111111111_1111111111111111_1110010011110000_0110110000000101"; -- -0.10570645209085278
	pesos_i(4709) := b"0000000000000000_0000000000000000_0000110001100101_0001000101101000"; -- 0.04841717524177644
	pesos_i(4710) := b"1111111111111111_1111111111111111_1111011000111011_1110101011000011"; -- -0.0381482386678232
	pesos_i(4711) := b"0000000000000000_0000000000000000_0010000000010010_0111001000000101"; -- 0.12528145437278781
	pesos_i(4712) := b"1111111111111111_1111111111111111_1111100111011010_1001011011100101"; -- -0.024008340066077688
	pesos_i(4713) := b"1111111111111111_1111111111111111_1111000101001101_0010101010011000"; -- -0.05741628449355593
	pesos_i(4714) := b"1111111111111111_1111111111111111_1111001001010011_1001010100101101"; -- -0.05341212892571079
	pesos_i(4715) := b"1111111111111111_1111111111111111_1101001110110010_1110111101100111"; -- -0.1730509161262473
	pesos_i(4716) := b"1111111111111111_1111111111111111_1110101100010000_0111111001101010"; -- -0.08177957451841647
	pesos_i(4717) := b"1111111111111111_1111111111111111_1110111010011001_0010101111101011"; -- -0.06797528756679135
	pesos_i(4718) := b"0000000000000000_0000000000000000_0010110101011100_1100100110001100"; -- 0.17719707163754359
	pesos_i(4719) := b"1111111111111111_1111111111111111_1111101101100111_0010000010100000"; -- -0.017957650111666126
	pesos_i(4720) := b"1111111111111111_1111111111111111_1110100010111110_1011001110110000"; -- -0.09084011987865086
	pesos_i(4721) := b"0000000000000000_0000000000000000_0000101111010010_0001101011001011"; -- 0.04617469260754506
	pesos_i(4722) := b"0000000000000000_0000000000000000_0010000011011001_1101010011100010"; -- 0.12832384599530866
	pesos_i(4723) := b"0000000000000000_0000000000000000_0011000001010001_1101111110111011"; -- 0.18874929719432848
	pesos_i(4724) := b"0000000000000000_0000000000000000_0001011110010110_0000010001100001"; -- 0.09213282926816052
	pesos_i(4725) := b"0000000000000000_0000000000000000_0001000110101010_1111011110010100"; -- 0.06901500095624415
	pesos_i(4726) := b"1111111111111111_1111111111111111_1101110000000001_0000001101110001"; -- -0.14060953601073756
	pesos_i(4727) := b"1111111111111111_1111111111111111_1110111000111000_0010101111001010"; -- -0.06945539789109938
	pesos_i(4728) := b"0000000000000000_0000000000000000_0001010011101010_0100111010001100"; -- 0.0817002384004647
	pesos_i(4729) := b"1111111111111111_1111111111111111_1110100010001111_0001101001100101"; -- -0.09156641995715836
	pesos_i(4730) := b"0000000000000000_0000000000000000_0010110000010000_0001100000111100"; -- 0.17212058510872477
	pesos_i(4731) := b"0000000000000000_0000000000000000_0001101010010111_1010110110111100"; -- 0.1038769325433585
	pesos_i(4732) := b"1111111111111111_1111111111111111_1111001101010111_0010110001101111"; -- -0.049451086794856686
	pesos_i(4733) := b"1111111111111111_1111111111111111_1011101111110000_0000010111110000"; -- -0.2658687866375512
	pesos_i(4734) := b"0000000000000000_0000000000000000_0001110000011101_0111000100001000"; -- 0.10982424201747433
	pesos_i(4735) := b"1111111111111111_1111111111111111_1101101011011011_1000011001011011"; -- -0.14508781691856784
	pesos_i(4736) := b"1111111111111111_1111111111111111_1110010110100100_1100101010110100"; -- -0.10295422665241308
	pesos_i(4737) := b"0000000000000000_0000000000000000_0000001010011011_1011011001110110"; -- 0.0101884877828477
	pesos_i(4738) := b"0000000000000000_0000000000000000_0000001100100011_1110100011010110"; -- 0.01226668579392809
	pesos_i(4739) := b"1111111111111111_1111111111111111_1111110101000100_0011001010110011"; -- -0.010678130487730093
	pesos_i(4740) := b"1111111111111111_1111111111111111_1101101001101001_0000001000010011"; -- -0.14683520346984974
	pesos_i(4741) := b"0000000000000000_0000000000000000_0000110101111100_1100111101110001"; -- 0.052685704299811016
	pesos_i(4742) := b"1111111111111111_1111111111111111_1110111101010010_0100011110100011"; -- -0.06515075943359355
	pesos_i(4743) := b"0000000000000000_0000000000000000_0000011001010000_0011100010101000"; -- 0.02466158017533857
	pesos_i(4744) := b"0000000000000000_0000000000000000_0101001101001110_0110111111001011"; -- 0.3254155988276059
	pesos_i(4745) := b"1111111111111111_1111111111111111_1111111011011001_0011000101110001"; -- -0.004498395768820206
	pesos_i(4746) := b"1111111111111111_1111111111111111_1111101110000100_0101011000011110"; -- -0.01751195683800433
	pesos_i(4747) := b"0000000000000000_0000000000000000_0000001010101011_1011000000110000"; -- 0.010432254460442547
	pesos_i(4748) := b"1111111111111111_1111111111111111_1011011100011111_1110011010001110"; -- -0.284669485375416
	pesos_i(4749) := b"0000000000000000_0000000000000000_0010010101110011_1110111111111000"; -- 0.14630031394883655
	pesos_i(4750) := b"1111111111111111_1111111111111111_1101000000011110_0010010111011101"; -- -0.18703997948507306
	pesos_i(4751) := b"1111111111111111_1111111111111111_1111001101110010_1011111101011001"; -- -0.049030342837195
	pesos_i(4752) := b"1111111111111111_1111111111111111_1111101011111001_1011101010101011"; -- -0.0196269351822639
	pesos_i(4753) := b"1111111111111111_1111111111111111_1111100111101100_0000011001100000"; -- -0.023742295735434987
	pesos_i(4754) := b"1111111111111111_1111111111111111_1101111011111111_1101101011000000"; -- -0.12890847038860637
	pesos_i(4755) := b"0000000000000000_0000000000000000_0010111011111110_0011011111110000"; -- 0.1835665666485824
	pesos_i(4756) := b"1111111111111111_1111111111111111_1110100000100101_0001100111000000"; -- -0.09318388997352225
	pesos_i(4757) := b"1111111111111111_1111111111111111_1110000011000110_0100000011011101"; -- -0.12197489369548598
	pesos_i(4758) := b"0000000000000000_0000000000000000_0010101010001000_0000110110100111"; -- 0.16613850904482824
	pesos_i(4759) := b"0000000000000000_0000000000000000_0010001011110101_0100101110101010"; -- 0.13655541328413137
	pesos_i(4760) := b"0000000000000000_0000000000000000_0001111101001011_0010111001111000"; -- 0.12224092893973054
	pesos_i(4761) := b"0000000000000000_0000000000000000_0000000001101010_0000110111110011"; -- 0.0016182631489991568
	pesos_i(4762) := b"0000000000000000_0000000000000000_0011001000010001_0000000100000001"; -- 0.19557195921232992
	pesos_i(4763) := b"1111111111111111_1111111111111111_1101011001001111_0110011000111110"; -- -0.16285096163059845
	pesos_i(4764) := b"1111111111111111_1111111111111111_1110000000011010_0010011100101001"; -- -0.1246009372974633
	pesos_i(4765) := b"1111111111111111_1111111111111111_1111011111111110_0101110001101011"; -- -0.031275008964426476
	pesos_i(4766) := b"1111111111111111_1111111111111111_1111010111000100_1000010010010100"; -- -0.039970125017921465
	pesos_i(4767) := b"0000000000000000_0000000000000000_0000011010000101_0110110101101000"; -- 0.025473440164902217
	pesos_i(4768) := b"1111111111111111_1111111111111111_1101011101011110_1011101011100111"; -- -0.1587107836747184
	pesos_i(4769) := b"1111111111111111_1111111111111111_1110010111111010_0111010100100110"; -- -0.10164707003790048
	pesos_i(4770) := b"0000000000000000_0000000000000000_0000001111001010_1011111111011010"; -- 0.014812460605800187
	pesos_i(4771) := b"1111111111111111_1111111111111111_1101011110001100_0101101100110010"; -- -0.15801458380217942
	pesos_i(4772) := b"1111111111111111_1111111111111111_1110100101111111_0011101111010100"; -- -0.08790231777438406
	pesos_i(4773) := b"1111111111111111_1111111111111111_1110010000011101_0001010001110100"; -- -0.10893127603438575
	pesos_i(4774) := b"1111111111111111_1111111111111111_1110001110111001_1111001001100011"; -- -0.11044392657569074
	pesos_i(4775) := b"0000000000000000_0000000000000000_0010010100101101_0011001000010111"; -- 0.14522088108056994
	pesos_i(4776) := b"0000000000000000_0000000000000000_0010100000100010_1100111000000000"; -- 0.15678107733659802
	pesos_i(4777) := b"1111111111111111_1111111111111111_1111001111110101_0010111010110111"; -- -0.04704006221510968
	pesos_i(4778) := b"0000000000000000_0000000000000000_0001000000101111_0001111101111010"; -- 0.06321903919571897
	pesos_i(4779) := b"0000000000000000_0000000000000000_0000100010010101_1011110100111110"; -- 0.03353483929260313
	pesos_i(4780) := b"1111111111111111_1111111111111111_1100011010101101_1111110111000101"; -- -0.22390760362448736
	pesos_i(4781) := b"1111111111111111_1111111111111111_1101100111000011_0001101111001000"; -- -0.14936663033356068
	pesos_i(4782) := b"0000000000000000_0000000000000000_0000101010111110_1001101011011110"; -- 0.041970900742221984
	pesos_i(4783) := b"0000000000000000_0000000000000000_0001100001101011_1100100111110011"; -- 0.0953947276038891
	pesos_i(4784) := b"0000000000000000_0000000000000000_0010101010110100_0000101001100010"; -- 0.1668097008481142
	pesos_i(4785) := b"1111111111111111_1111111111111111_1110001000000110_1011010110011110"; -- -0.11708512197610907
	pesos_i(4786) := b"1111111111111111_1111111111111111_1110111111010001_1000000101111010"; -- -0.06320944560265598
	pesos_i(4787) := b"1111111111111111_1111111111111111_1010101101110101_1001110000101000"; -- -0.3302366641045879
	pesos_i(4788) := b"1111111111111111_1111111111111111_1101101000001011_0000010111001110"; -- -0.14826930739152622
	pesos_i(4789) := b"0000000000000000_0000000000000000_0001111010111111_1100001010000110"; -- 0.1201135231058156
	pesos_i(4790) := b"1111111111111111_1111111111111111_1100100011110000_0101101000101110"; -- -0.21508251557704833
	pesos_i(4791) := b"0000000000000000_0000000000000000_0000011110011111_0111010000101010"; -- 0.029776821300777273
	pesos_i(4792) := b"1111111111111111_1111111111111111_1101001010101011_0000111010000111"; -- -0.17707738118071636
	pesos_i(4793) := b"1111111111111111_1111111111111111_1111011101111100_1111110101110111"; -- -0.033249052565991935
	pesos_i(4794) := b"1111111111111111_1111111111111111_1110100111001011_1001100111111010"; -- -0.08673703813940449
	pesos_i(4795) := b"1111111111111111_1111111111111111_1111111100010101_1010101110111111"; -- -0.0035755784507086608
	pesos_i(4796) := b"0000000000000000_0000000000000000_0000011001011111_1100010111010111"; -- 0.024898877145337478
	pesos_i(4797) := b"0000000000000000_0000000000000000_0001101011100011_0100100011101101"; -- 0.10503059188329888
	pesos_i(4798) := b"0000000000000000_0000000000000000_0001100010111111_1100111101010001"; -- 0.0966767858423332
	pesos_i(4799) := b"0000000000000000_0000000000000000_0011011000100001_0100101000000110"; -- 0.21144545222833255
	pesos_i(4800) := b"1111111111111111_1111111111111111_1101110101101011_0110000000110011"; -- -0.13508032558145144
	pesos_i(4801) := b"0000000000000000_0000000000000000_0000000011100101_0101010000001011"; -- 0.0034992720398038524
	pesos_i(4802) := b"1111111111111111_1111111111111111_1111011001000110_0111001001011011"; -- -0.0379875686202745
	pesos_i(4803) := b"1111111111111111_1111111111111111_1110101100101110_0111001100110010"; -- -0.08132247945191629
	pesos_i(4804) := b"1111111111111111_1111111111111111_1110000101011100_1010100011100010"; -- -0.11967987520186021
	pesos_i(4805) := b"0000000000000000_0000000000000000_0000001100000011_1010001011010010"; -- 0.011774231245666567
	pesos_i(4806) := b"1111111111111111_1111111111111111_1110000110001101_0001000110101001"; -- -0.11894120807639479
	pesos_i(4807) := b"1111111111111111_1111111111111111_1110111110001100_0110001011010001"; -- -0.0642641296963464
	pesos_i(4808) := b"0000000000000000_0000000000000000_0010100110100001_0101010100100100"; -- 0.1626179898797681
	pesos_i(4809) := b"0000000000000000_0000000000000000_0001101101101101_0110010100101100"; -- 0.10713798841989014
	pesos_i(4810) := b"0000000000000000_0000000000000000_0010010101110010_1001001011101111"; -- 0.14627950977317128
	pesos_i(4811) := b"0000000000000000_0000000000000000_0001101001001001_0110001011110000"; -- 0.10268228868277768
	pesos_i(4812) := b"1111111111111111_1111111111111111_1111111110101010_0011000101000010"; -- -0.0013093198208705692
	pesos_i(4813) := b"0000000000000000_0000000000000000_0000111100000001_1010000101100010"; -- 0.05861862791667696
	pesos_i(4814) := b"1111111111111111_1111111111111111_1101110110000100_0000000010000100"; -- -0.13470455915644125
	pesos_i(4815) := b"0000000000000000_0000000000000000_0000101001101000_1100111111111110"; -- 0.04066181134814814
	pesos_i(4816) := b"0000000000000000_0000000000000000_0010111100110001_0011001011100111"; -- 0.18434446465559395
	pesos_i(4817) := b"1111111111111111_1111111111111111_1110011010111000_0101010011111101"; -- -0.09874981713011237
	pesos_i(4818) := b"0000000000000000_0000000000000000_0001000011011010_0111101110100111"; -- 0.06583378628024261
	pesos_i(4819) := b"1111111111111111_1111111111111111_1101100110100111_1111000011001010"; -- -0.14978117998264454
	pesos_i(4820) := b"0000000000000000_0000000000000000_0001101011100100_1110010010100000"; -- 0.10505513100261954
	pesos_i(4821) := b"0000000000000000_0000000000000000_0001100100001000_1110001110001011"; -- 0.09779188282388102
	pesos_i(4822) := b"1111111111111111_1111111111111111_1101010110000110_0100000110000000"; -- -0.1659201682432452
	pesos_i(4823) := b"1111111111111111_1111111111111111_1110111100100100_1110100011011001"; -- -0.06584305468157978
	pesos_i(4824) := b"1111111111111111_1111111111111111_1101000011000111_1010100100011011"; -- -0.18445342160107606
	pesos_i(4825) := b"0000000000000000_0000000000000000_0010100011001111_0110111011010100"; -- 0.15941517529694688
	pesos_i(4826) := b"0000000000000000_0000000000000000_0000011010110011_0101111000011011"; -- 0.026174432305897083
	pesos_i(4827) := b"0000000000000000_0000000000000000_0001100000110000_0100000010101000"; -- 0.09448627575836477
	pesos_i(4828) := b"0000000000000000_0000000000000000_0000001001101101_1010011010101011"; -- 0.0094856421106565
	pesos_i(4829) := b"1111111111111111_1111111111111111_1110100011000000_1110011000100100"; -- -0.09080659512635474
	pesos_i(4830) := b"1111111111111111_1111111111111111_1110011000010100_0011011111111010"; -- -0.10125398786727564
	pesos_i(4831) := b"1111111111111111_1111111111111111_1111111100001000_1000101111111111"; -- -0.0037758351977999483
	pesos_i(4832) := b"0000000000000000_0000000000000000_0001111010110111_0101011110100111"; -- 0.11998508277531572
	pesos_i(4833) := b"1111111111111111_1111111111111111_1110100011101111_0010110000001101"; -- -0.09010052372880885
	pesos_i(4834) := b"0000000000000000_0000000000000000_0001100101100100_1000111111101110"; -- 0.09919070774843342
	pesos_i(4835) := b"0000000000000000_0000000000000000_0000010101001101_0010110010001000"; -- 0.020708831091811597
	pesos_i(4836) := b"0000000000000000_0000000000000000_0010101111110101_0011011101010101"; -- 0.17171045138783353
	pesos_i(4837) := b"0000000000000000_0000000000000000_0000000000111101_1001010100110110"; -- 0.0009396798533060913
	pesos_i(4838) := b"0000000000000000_0000000000000000_0000011110100111_0010111100111001"; -- 0.02989478245605326
	pesos_i(4839) := b"1111111111111111_1111111111111111_1111100010000110_1010110010011110"; -- -0.029195033372757667
	pesos_i(4840) := b"1111111111111111_1111111111111111_1110111010111010_0100100111001011"; -- -0.06746996690410947
	pesos_i(4841) := b"0000000000000000_0000000000000000_0000001100010111_0110001110000111"; -- 0.012075634507839578
	pesos_i(4842) := b"0000000000000000_0000000000000000_0001001111000011_1110001000110111"; -- 0.07720769727748622
	pesos_i(4843) := b"1111111111111111_1111111111111111_1101010101101011_1001000001111001"; -- -0.166327448392247
	pesos_i(4844) := b"0000000000000000_0000000000000000_0001111001100010_1011110101010101"; -- 0.11869414628912722
	pesos_i(4845) := b"1111111111111111_1111111111111111_1101100111000011_0011111110001000"; -- -0.14936449932153
	pesos_i(4846) := b"0000000000000000_0000000000000000_0010011100111101_0101101110101101"; -- 0.1532800004773957
	pesos_i(4847) := b"0000000000000000_0000000000000000_0010001101111100_1000001011101010"; -- 0.1386186429544955
	pesos_i(4848) := b"1111111111111111_1111111111111111_1110010011110000_1010001010001011"; -- -0.10570320239384604
	pesos_i(4849) := b"0000000000000000_0000000000000000_0010111111011101_1000000001100111"; -- 0.18697359574367922
	pesos_i(4850) := b"0000000000000000_0000000000000000_0010011111000000_1000011000100011"; -- 0.15528143267409145
	pesos_i(4851) := b"0000000000000000_0000000000000000_0001100011111111_1111001111011101"; -- 0.09765552664491522
	pesos_i(4852) := b"0000000000000000_0000000000000000_0000010000110011_0011000010001100"; -- 0.016406091772037612
	pesos_i(4853) := b"1111111111111111_1111111111111111_1110001000010101_1011000111101100"; -- -0.11685646042329773
	pesos_i(4854) := b"0000000000000000_0000000000000000_0001101010000000_1011011010011011"; -- 0.10352650903558319
	pesos_i(4855) := b"0000000000000000_0000000000000000_0010111011100111_0001100011110011"; -- 0.1832137672834248
	pesos_i(4856) := b"0000000000000000_0000000000000000_0001011110010010_0010001010110001"; -- 0.09207360090164984
	pesos_i(4857) := b"1111111111111111_1111111111111111_1111010011000011_0101011001001111"; -- -0.04389439184684077
	pesos_i(4858) := b"1111111111111111_1111111111111111_1111110101100000_1011010110111011"; -- -0.010243074295960913
	pesos_i(4859) := b"1111111111111111_1111111111111111_1100111100100111_1011011100100010"; -- -0.1908002416140575
	pesos_i(4860) := b"0000000000000000_0000000000000000_0000000000101111_1001010000011011"; -- 0.0007259907872942672
	pesos_i(4861) := b"1111111111111111_1111111111111111_1101111011101011_1110101100011011"; -- -0.12921267130265332
	pesos_i(4862) := b"0000000000000000_0000000000000000_0001000101110110_0110011001100011"; -- 0.06821288991228236
	pesos_i(4863) := b"1111111111111111_1111111111111111_1101101111100100_0100111001010010"; -- -0.14104757786225494
	pesos_i(4864) := b"1111111111111111_1111111111111111_1101100000110101_1110001000010111"; -- -0.15542780822040436
	pesos_i(4865) := b"1111111111111111_1111111111111111_1111000000111011_0001001001111110"; -- -0.06159862913898334
	pesos_i(4866) := b"1111111111111111_1111111111111111_1111001100110110_0010111000100110"; -- -0.04995452483371185
	pesos_i(4867) := b"1111111111111111_1111111111111111_1110100100100110_0001000001101100"; -- -0.08926293719652757
	pesos_i(4868) := b"1111111111111111_1111111111111111_1101101100110001_1011101001101100"; -- -0.14377245774942032
	pesos_i(4869) := b"0000000000000000_0000000000000000_0000000010010110_0010010101000100"; -- 0.002291039678513379
	pesos_i(4870) := b"0000000000000000_0000000000000000_0010000010110110_0010011100001110"; -- 0.12777942734544578
	pesos_i(4871) := b"1111111111111111_1111111111111111_1101000110000100_1000000110111110"; -- -0.18157185671437692
	pesos_i(4872) := b"1111111111111111_1111111111111111_1111101000010001_0001100100011010"; -- -0.023176604418336216
	pesos_i(4873) := b"1111111111111111_1111111111111111_1101011110110101_0111000011100110"; -- -0.1573876798635902
	pesos_i(4874) := b"0000000000000000_0000000000000000_0010010011001010_0011001100101101"; -- 0.14371032571655812
	pesos_i(4875) := b"0000000000000000_0000000000000000_0010010111010110_0001100001100101"; -- 0.14779808484724616
	pesos_i(4876) := b"1111111111111111_1111111111111111_1101001110001110_0011110101011000"; -- -0.17361084554442566
	pesos_i(4877) := b"0000000000000000_0000000000000000_0011000010110111_1010101110111011"; -- 0.19030259433427127
	pesos_i(4878) := b"0000000000000000_0000000000000000_0010110001100001_0110001000100111"; -- 0.1733609527793889
	pesos_i(4879) := b"1111111111111111_1111111111111111_1111000000110100_1001001110001100"; -- -0.06169774837832773
	pesos_i(4880) := b"0000000000000000_0000000000000000_0001101100010110_0111000000100011"; -- 0.10581112731591136
	pesos_i(4881) := b"0000000000000000_0000000000000000_0001111111111110_1111111010100111"; -- 0.12498466094424415
	pesos_i(4882) := b"0000000000000000_0000000000000000_0000110001111110_0110000101001111"; -- 0.04880340737398889
	pesos_i(4883) := b"1111111111111111_1111111111111111_1101111001100011_1100100011100111"; -- -0.13128990513295835
	pesos_i(4884) := b"1111111111111111_1111111111111111_1110000101010011_0001010011001101"; -- -0.119826030607514
	pesos_i(4885) := b"1111111111111111_1111111111111111_1111111011111011_0010001010010010"; -- -0.003980483363293069
	pesos_i(4886) := b"0000000000000000_0000000000000000_0010000111100010_0111011011111110"; -- 0.13236182874326086
	pesos_i(4887) := b"1111111111111111_1111111111111111_1110100000100010_1011110011001000"; -- -0.09321994888356544
	pesos_i(4888) := b"0000000000000000_0000000000000000_0001110010101010_1111100111000000"; -- 0.11198388047528973
	pesos_i(4889) := b"1111111111111111_1111111111111111_1101110110100010_0000110111111111"; -- -0.13424599188914302
	pesos_i(4890) := b"0000000000000000_0000000000000000_0000011011010110_1001011110111101"; -- 0.026711925218040194
	pesos_i(4891) := b"1111111111111111_1111111111111111_1101101010100101_0010111101001100"; -- -0.14591698073919385
	pesos_i(4892) := b"1111111111111111_1111111111111111_1111011101110011_0001100010001011"; -- -0.033400026278383205
	pesos_i(4893) := b"1111111111111111_1111111111111111_1111100100001000_0000011111001001"; -- -0.0272212155541518
	pesos_i(4894) := b"1111111111111111_1111111111111111_1110110000001001_0100011111100010"; -- -0.07798338625547868
	pesos_i(4895) := b"0000000000000000_0000000000000000_0000000111111101_0100111101111101"; -- 0.007771461571552785
	pesos_i(4896) := b"1111111111111111_1111111111111111_1111100100111100_1110001101000100"; -- -0.02641467656693275
	pesos_i(4897) := b"1111111111111111_1111111111111111_1101101001101001_0001000011101101"; -- -0.146834318229932
	pesos_i(4898) := b"0000000000000000_0000000000000000_0010101101001100_0100100010010000"; -- 0.16913274311872256
	pesos_i(4899) := b"1111111111111111_1111111111111111_1110111000110100_1101101001011010"; -- -0.0695060282912734
	pesos_i(4900) := b"0000000000000000_0000000000000000_0001100111010111_1101110001110100"; -- 0.10095002961403918
	pesos_i(4901) := b"1111111111111111_1111111111111111_1101010100010110_1111010011101101"; -- -0.16761845785524973
	pesos_i(4902) := b"0000000000000000_0000000000000000_0001101101000101_0100100011000011"; -- 0.10652594344396893
	pesos_i(4903) := b"1111111111111111_1111111111111111_1110100100001100_0000011110010101"; -- -0.08966019271608318
	pesos_i(4904) := b"1111111111111111_1111111111111111_1111010100101011_1011110010111101"; -- -0.04230137250719672
	pesos_i(4905) := b"0000000000000000_0000000000000000_0001110100000101_0100010111001101"; -- 0.11336170446815187
	pesos_i(4906) := b"1111111111111111_1111111111111111_1111010011010011_0101110110011100"; -- -0.04364981599087284
	pesos_i(4907) := b"1111111111111111_1111111111111111_1101110100111001_1100101000001111"; -- -0.13583695541310786
	pesos_i(4908) := b"1111111111111111_1111111111111111_1110111110110110_0000000001000110"; -- -0.06362913416277792
	pesos_i(4909) := b"1111111111111111_1111111111111111_1110101010100110_1100011011101010"; -- -0.08339268482118817
	pesos_i(4910) := b"1111111111111111_1111111111111111_1110100010110101_0010010101001011"; -- -0.09098593632647113
	pesos_i(4911) := b"0000000000000000_0000000000000000_0001011111001001_1100011010001001"; -- 0.09292260028481314
	pesos_i(4912) := b"1111111111111111_1111111111111111_1111011001110110_0011110011000101"; -- -0.0372583406493353
	pesos_i(4913) := b"1111111111111111_1111111111111111_1111101001110010_1000110111011010"; -- -0.021689543015132318
	pesos_i(4914) := b"1111111111111111_1111111111111111_1101110100000001_1000111100111111"; -- -0.13669495298295958
	pesos_i(4915) := b"1111111111111111_1111111111111111_1111001010110110_1111010000011010"; -- -0.05189585076539352
	pesos_i(4916) := b"0000000000000000_0000000000000000_0000010000110001_0011000011110011"; -- 0.0163755983079985
	pesos_i(4917) := b"1111111111111111_1111111111111111_1101011011110100_1100001111011111"; -- -0.16032768054238175
	pesos_i(4918) := b"1111111111111111_1111111111111111_1100100011010011_0101100110100010"; -- -0.2155250530572933
	pesos_i(4919) := b"1111111111111111_1111111111111111_1110111111010100_1000011001001000"; -- -0.06316338290882334
	pesos_i(4920) := b"0000000000000000_0000000000000000_0000101001101011_1000010011011111"; -- 0.040703110108559336
	pesos_i(4921) := b"1111111111111111_1111111111111111_1101111010001110_1111110111100111"; -- -0.13063061811373455
	pesos_i(4922) := b"1111111111111111_1111111111111111_1101111000001000_1011001001110000"; -- -0.13267979399043775
	pesos_i(4923) := b"1111111111111111_1111111111111111_1110101000110111_0001111101101011"; -- -0.08509639394303496
	pesos_i(4924) := b"0000000000000000_0000000000000000_0001110011111111_0011000101100110"; -- 0.1132689355465572
	pesos_i(4925) := b"1111111111111111_1111111111111111_1101000011110000_0110001000001000"; -- -0.18383204743337622
	pesos_i(4926) := b"0000000000000000_0000000000000000_0010000001111110_1000011011011000"; -- 0.12693064475580185
	pesos_i(4927) := b"0000000000000000_0000000000000000_0010111100111100_0001000000111101"; -- 0.1845102453059512
	pesos_i(4928) := b"1111111111111111_1111111111111111_1101100011000010_1100111111111111"; -- -0.15327739730810583
	pesos_i(4929) := b"1111111111111111_1111111111111111_1111001000000110_0001011011001010"; -- -0.05459458884098666
	pesos_i(4930) := b"1111111111111111_1111111111111111_1111011110111010_0011101111110111"; -- -0.03231454094017232
	pesos_i(4931) := b"1111111111111111_1111111111111111_1101011111110000_0010000100000111"; -- -0.1564921720207809
	pesos_i(4932) := b"0000000000000000_0000000000000000_0000111000101010_0011101101001111"; -- 0.05533190411197943
	pesos_i(4933) := b"0000000000000000_0000000000000000_0010001110000010_1111101010000000"; -- 0.13871732357002048
	pesos_i(4934) := b"0000000000000000_0000000000000000_0010111000110100_1000011011010100"; -- 0.18048899337866994
	pesos_i(4935) := b"0000000000000000_0000000000000000_0010101000110101_0011011010101100"; -- 0.16487447447374678
	pesos_i(4936) := b"1111111111111111_1111111111111111_1110111001100000_0110000011001011"; -- -0.0688418868795674
	pesos_i(4937) := b"1111111111111111_1111111111111111_1110010111001011_0010011111011011"; -- -0.10236884026563463
	pesos_i(4938) := b"0000000000000000_0000000000000000_0010001111010011_1000110011001101"; -- 0.13994674689850228
	pesos_i(4939) := b"1111111111111111_1111111111111111_1111100101010000_0000100000100101"; -- -0.026122561487121197
	pesos_i(4940) := b"1111111111111111_1111111111111111_1110110000011100_0111110110010001"; -- -0.07769026951419862
	pesos_i(4941) := b"0000000000000000_0000000000000000_0000010010001111_0000011110001111"; -- 0.01780745731199869
	pesos_i(4942) := b"1111111111111111_1111111111111111_1111011001111011_1000101010000001"; -- -0.03717741347972675
	pesos_i(4943) := b"0000000000000000_0000000000000000_0001001010111000_0110110011110101"; -- 0.07312661154324494
	pesos_i(4944) := b"0000000000000000_0000000000000000_0010100101100010_1010100100110110"; -- 0.1616616970062664
	pesos_i(4945) := b"1111111111111111_1111111111111111_1101000001000110_0110100000101010"; -- -0.18642567612056146
	pesos_i(4946) := b"0000000000000000_0000000000000000_0000001000111100_0010100011001101"; -- 0.008730459357839037
	pesos_i(4947) := b"1111111111111111_1111111111111111_1110010001001010_0110110101100111"; -- -0.10823932866591385
	pesos_i(4948) := b"1111111111111111_1111111111111111_1111001001101011_0010100100010001"; -- -0.05305236184553913
	pesos_i(4949) := b"0000000000000000_0000000000000000_0000111100000001_1000110111000001"; -- 0.05861745804064165
	pesos_i(4950) := b"1111111111111111_1111111111111111_1111001110101110_1011100111001111"; -- -0.048115145589193636
	pesos_i(4951) := b"1111111111111111_1111111111111111_1110100101001101_1110101010110110"; -- -0.08865483331782532
	pesos_i(4952) := b"0000000000000000_0000000000000000_0000011100111101_1001000110111001"; -- 0.02828322199357177
	pesos_i(4953) := b"1111111111111111_1111111111111111_1100110111001010_1001011011000011"; -- -0.196127488472281
	pesos_i(4954) := b"1111111111111111_1111111111111111_1101110110110101_1110010011110101"; -- -0.13394326226677564
	pesos_i(4955) := b"0000000000000000_0000000000000000_0000001111101101_1001100100001100"; -- 0.01534420541758788
	pesos_i(4956) := b"0000000000000000_0000000000000000_0001001011000001_0110000010010100"; -- 0.07326320269579026
	pesos_i(4957) := b"0000000000000000_0000000000000000_0001101001111110_0010100001111110"; -- 0.1034875209935705
	pesos_i(4958) := b"0000000000000000_0000000000000000_0000000110111111_0000100110001110"; -- 0.006821248104253907
	pesos_i(4959) := b"1111111111111111_1111111111111111_1111111001010000_0000111100110100"; -- -0.006590890766090941
	pesos_i(4960) := b"1111111111111111_1111111111111111_1111001111100000_1110000001010001"; -- -0.0473499108534281
	pesos_i(4961) := b"1111111111111111_1111111111111111_1110111111000111_0111011001000000"; -- -0.06336270261636667
	pesos_i(4962) := b"1111111111111111_1111111111111111_1111010010000010_1000111011100101"; -- -0.04488284017321168
	pesos_i(4963) := b"0000000000000000_0000000000000000_0001000110011011_1011001110001011"; -- 0.06878206395109386
	pesos_i(4964) := b"1111111111111111_1111111111111111_1101101100101001_0101101111110000"; -- -0.14390015967760225
	pesos_i(4965) := b"0000000000000000_0000000000000000_0010111110011010_0010110100111001"; -- 0.18594629890394557
	pesos_i(4966) := b"0000000000000000_0000000000000000_0010000100011000_1011000000000000"; -- 0.1292829514177243
	pesos_i(4967) := b"0000000000000000_0000000000000000_0000000011100101_0111100100111001"; -- 0.003501488129135164
	pesos_i(4968) := b"1111111111111111_1111111111111111_1111101010111011_1101110001100010"; -- -0.020570970720787538
	pesos_i(4969) := b"1111111111111111_1111111111111111_1111101011111011_1111000011000001"; -- -0.019593193808435917
	pesos_i(4970) := b"1111111111111111_1111111111111111_1101010110110100_0010101100011101"; -- -0.16521959829417723
	pesos_i(4971) := b"1111111111111111_1111111111111111_1111100011011010_1100000010100110"; -- -0.02791210114673656
	pesos_i(4972) := b"1111111111111111_1111111111111111_1101010101000011_1110010000011000"; -- -0.16693281575944627
	pesos_i(4973) := b"1111111111111111_1111111111111111_1111000011101000_1011101111110010"; -- -0.05894875851757463
	pesos_i(4974) := b"1111111111111111_1111111111111111_1110100110001010_1101101001110100"; -- -0.08772501633434426
	pesos_i(4975) := b"0000000000000000_0000000000000000_0001011101100111_1110001011000000"; -- 0.09142892064719464
	pesos_i(4976) := b"0000000000000000_0000000000000000_0000101000000110_1111001000000111"; -- 0.039168478762013605
	pesos_i(4977) := b"1111111111111111_1111111111111111_1111111100100010_0100000010100000"; -- -0.0033835991243207717
	pesos_i(4978) := b"1111111111111111_1111111111111111_1111110100111010_1011000111100110"; -- -0.01082313664043581
	pesos_i(4979) := b"1111111111111111_1111111111111111_1110110110000110_1011001100001100"; -- -0.07216340015574109
	pesos_i(4980) := b"0000000000000000_0000000000000000_0000111010001001_0100010111101110"; -- 0.056782122121816214
	pesos_i(4981) := b"1111111111111111_1111111111111111_1100111110000011_1101001001111100"; -- -0.1893948028254341
	pesos_i(4982) := b"1111111111111111_1111111111111111_1111011110000101_1111111111101100"; -- -0.03311157684102615
	pesos_i(4983) := b"0000000000000000_0000000000000000_0001000101001110_1010111100110011"; -- 0.0676068781609095
	pesos_i(4984) := b"1111111111111111_1111111111111111_1110010111010011_1110001110000110"; -- -0.1022355841309118
	pesos_i(4985) := b"0000000000000000_0000000000000000_0000000000000100_1001010000111010"; -- 6.987007023602254e-05
	pesos_i(4986) := b"0000000000000000_0000000000000000_0000100001100111_0001100111000000"; -- 0.032823190119129445
	pesos_i(4987) := b"1111111111111111_1111111111111111_1110011011000100_1000100111011000"; -- -0.09856356118310838
	pesos_i(4988) := b"1111111111111111_1111111111111111_1111110001010011_0010101001011011"; -- -0.014355995904853973
	pesos_i(4989) := b"1111111111111111_1111111111111111_1101000110100111_1011010010001110"; -- -0.18103477038674312
	pesos_i(4990) := b"1111111111111111_1111111111111111_1110010000010101_1010000111011100"; -- -0.10904491795864413
	pesos_i(4991) := b"0000000000000000_0000000000000000_0100010000100011_1011010100101001"; -- 0.2661698555953491
	pesos_i(4992) := b"1111111111111111_1111111111111111_1110111111001111_1100111011001100"; -- -0.06323535465288445
	pesos_i(4993) := b"1111111111111111_1111111111111111_1100111000101010_1100011111011000"; -- -0.19465971917589836
	pesos_i(4994) := b"0000000000000000_0000000000000000_0000110110110001_0011010110111000"; -- 0.05348525747906485
	pesos_i(4995) := b"0000000000000000_0000000000000000_0001010010111100_1011000111001100"; -- 0.08100424989121631
	pesos_i(4996) := b"1111111111111111_1111111111111111_1101110001100111_1110110100110011"; -- -0.13903920655408603
	pesos_i(4997) := b"1111111111111111_1111111111111111_1110101100011110_1010001001000110"; -- -0.08156381405519875
	pesos_i(4998) := b"1111111111111111_1111111111111111_1110011011000110_1011111100100011"; -- -0.09852986712956747
	pesos_i(4999) := b"1111111111111111_1111111111111111_1101101101100001_1000000010100100"; -- -0.143043479822933
	pesos_i(5000) := b"0000000000000000_0000000000000000_0001000101001110_0000100101000100"; -- 0.067596987837238
	pesos_i(5001) := b"1111111111111111_1111111111111111_1111001000001101_0011001110110000"; -- -0.05448605494478489
	pesos_i(5002) := b"1111111111111111_1111111111111111_1110110010000100_0000110011001011"; -- -0.07611007742471336
	pesos_i(5003) := b"1111111111111111_1111111111111111_1101000100101101_0101010100110110"; -- -0.1829020255572864
	pesos_i(5004) := b"1111111111111111_1111111111111111_1110010001100010_1100101101001100"; -- -0.10786752124677873
	pesos_i(5005) := b"1111111111111111_1111111111111111_1110011110101011_1101110011000100"; -- -0.09503383830865501
	pesos_i(5006) := b"1111111111111111_1111111111111111_1111100111001111_0000111111110001"; -- -0.024184230565759923
	pesos_i(5007) := b"0000000000000000_0000000000000000_0000010001011011_0011111011001000"; -- 0.017017291838580004
	pesos_i(5008) := b"1111111111111111_1111111111111111_1110010110011011_1100100111001101"; -- -0.1030916094611483
	pesos_i(5009) := b"0000000000000000_0000000000000000_0000011000010100_0101100100000100"; -- 0.023747981440852325
	pesos_i(5010) := b"1111111111111111_1111111111111111_1101101101000110_0110101111001001"; -- -0.1434567101967363
	pesos_i(5011) := b"0000000000000000_0000000000000000_0001100010101001_0011110011100101"; -- 0.09633236486256941
	pesos_i(5012) := b"1111111111111111_1111111111111111_1101011000110110_0111010011011001"; -- -0.16323156073239165
	pesos_i(5013) := b"0000000000000000_0000000000000000_0001001001101101_0011011110001100"; -- 0.07197901877960655
	pesos_i(5014) := b"0000000000000000_0000000000000000_0001011010000010_1011011111011111"; -- 0.08793210216255258
	pesos_i(5015) := b"0000000000000000_0000000000000000_0000101001010110_1010000101100010"; -- 0.040384375041044876
	pesos_i(5016) := b"0000000000000000_0000000000000000_0000001010010111_1001010100100100"; -- 0.010125466719915065
	pesos_i(5017) := b"1111111111111111_1111111111111111_1111110011110110_0100110010011010"; -- -0.011866772026643005
	pesos_i(5018) := b"0000000000000000_0000000000000000_0010010100100100_0111100111000010"; -- 0.14508782363649902
	pesos_i(5019) := b"0000000000000000_0000000000000000_0000100010011111_1011111100110001"; -- 0.03368754338908504
	pesos_i(5020) := b"1111111111111111_1111111111111111_1111110010100110_0101101110000111"; -- -0.013086585600642377
	pesos_i(5021) := b"1111111111111111_1111111111111111_1110011101010111_0100010011001110"; -- -0.09632463417612323
	pesos_i(5022) := b"0000000000000000_0000000000000000_0010100100110110_1110100101110111"; -- 0.16099414011535462
	pesos_i(5023) := b"0000000000000000_0000000000000000_0000100101010001_1001110110010100"; -- 0.03640160420628479
	pesos_i(5024) := b"1111111111111111_1111111111111111_1111101011100011_0010111001100011"; -- -0.019970989917579538
	pesos_i(5025) := b"1111111111111111_1111111111111111_1101001011001111_0111110001101010"; -- -0.17652151494251442
	pesos_i(5026) := b"1111111111111111_1111111111111111_1101111101101011_0100001100000110"; -- -0.12726956463819641
	pesos_i(5027) := b"0000000000000000_0000000000000000_0000110010110111_0000111111100110"; -- 0.049668306118456004
	pesos_i(5028) := b"0000000000000000_0000000000000000_0001001000011110_0100010101100001"; -- 0.07077439889107388
	pesos_i(5029) := b"0000000000000000_0000000000000000_0000010100111001_0011001010011011"; -- 0.020404017242134816
	pesos_i(5030) := b"1111111111111111_1111111111111111_1111101100101101_1111111011001111"; -- -0.018829416773825693
	pesos_i(5031) := b"1111111111111111_1111111111111111_1110110111010101_0100010111111000"; -- -0.07096445757239808
	pesos_i(5032) := b"1111111111111111_1111111111111111_1110101111000100_0000001111110011"; -- -0.07904029187980123
	pesos_i(5033) := b"1111111111111111_1111111111111111_1111011011011010_0100110111001101"; -- -0.035731446584694404
	pesos_i(5034) := b"1111111111111111_1111111111111111_1101000101101101_1111001010110001"; -- -0.18191607655126116
	pesos_i(5035) := b"0000000000000000_0000000000000000_0000111000101011_0010111001000101"; -- 0.055346385907669146
	pesos_i(5036) := b"1111111111111111_1111111111111111_1110000111100011_0101010101000110"; -- -0.11762492229877095
	pesos_i(5037) := b"0000000000000000_0000000000000000_0010010100001010_0000111000001011"; -- 0.14468467488935516
	pesos_i(5038) := b"1111111111111111_1111111111111111_1110000100001110_0010100000010111"; -- -0.12087773734647339
	pesos_i(5039) := b"1111111111111111_1111111111111111_1111110111101010_0100111000111010"; -- -0.00814353076212635
	pesos_i(5040) := b"1111111111111111_1111111111111111_1111011000100100_0110110100010010"; -- -0.03850668241878843
	pesos_i(5041) := b"1111111111111111_1111111111111111_1111011101000101_1000001000011001"; -- -0.03409563902700452
	pesos_i(5042) := b"1111111111111111_1111111111111111_1101111010100011_1111001001000010"; -- -0.1303108777891625
	pesos_i(5043) := b"0000000000000000_0000000000000000_0000000101001101_1001010100101011"; -- 0.005090067849481315
	pesos_i(5044) := b"0000000000000000_0000000000000000_0001000110100011_1001110110100001"; -- 0.06890282799381434
	pesos_i(5045) := b"0000000000000000_0000000000000000_0010000110010110_0110001011001100"; -- 0.13120095700852125
	pesos_i(5046) := b"0000000000000000_0000000000000000_0001110010000110_0110010110010100"; -- 0.11142573231870675
	pesos_i(5047) := b"1111111111111111_1111111111111111_1101000100000100_0100110010011010"; -- -0.18352814893138428
	pesos_i(5048) := b"1111111111111111_1111111111111111_1110111010101101_0010110110111001"; -- -0.06767000416710509
	pesos_i(5049) := b"1111111111111111_1111111111111111_1111010010111101_0000111101101001"; -- -0.043990170372087696
	pesos_i(5050) := b"0000000000000000_0000000000000000_0000101010000110_1011000111100011"; -- 0.0411177805239905
	pesos_i(5051) := b"0000000000000000_0000000000000000_0001111010100111_0010001010001111"; -- 0.11973777759607794
	pesos_i(5052) := b"1111111111111111_1111111111111111_1101101001011011_1101011011011110"; -- -0.14703614321614597
	pesos_i(5053) := b"0000000000000000_0000000000000000_0000100100111011_1100000011100101"; -- 0.03606801597507841
	pesos_i(5054) := b"1111111111111111_1111111111111111_1110100001011011_1010111000100011"; -- -0.09235107076906302
	pesos_i(5055) := b"0000000000000000_0000000000000000_0001100010011011_0111011101001011"; -- 0.09612222275199866
	pesos_i(5056) := b"0000000000000000_0000000000000000_0000000000011010_0101010001100001"; -- 0.00040175786953740896
	pesos_i(5057) := b"0000000000000000_0000000000000000_0001110000100000_0110100111110100"; -- 0.10986959648753758
	pesos_i(5058) := b"0000000000000000_0000000000000000_0010100001100110_1011101101110100"; -- 0.15781756946496311
	pesos_i(5059) := b"0000000000000000_0000000000000000_0010001100000110_1001110100011000"; -- 0.13681966620225566
	pesos_i(5060) := b"0000000000000000_0000000000000000_0010001110101110_1011000101111000"; -- 0.13938435731718285
	pesos_i(5061) := b"0000000000000000_0000000000000000_0010010111101101_1001101010000100"; -- 0.1481567929504748
	pesos_i(5062) := b"0000000000000000_0000000000000000_0000100001100001_0001100110011101"; -- 0.0327316293153818
	pesos_i(5063) := b"1111111111111111_1111111111111111_1100110010101010_0100111111110000"; -- -0.20052624124826093
	pesos_i(5064) := b"0000000000000000_0000000000000000_0000100101111110_1011101000010100"; -- 0.037089948457726035
	pesos_i(5065) := b"1111111111111111_1111111111111111_1101010111001101_0101010100011000"; -- -0.16483562637195737
	pesos_i(5066) := b"1111111111111111_1111111111111111_1101011000100010_1000111101001011"; -- -0.16353516013135866
	pesos_i(5067) := b"1111111111111111_1111111111111111_1101100000010010_1111001000101100"; -- -0.1559609072800233
	pesos_i(5068) := b"0000000000000000_0000000000000000_0000000100010010_1110000010110110"; -- 0.004194302089482239
	pesos_i(5069) := b"0000000000000000_0000000000000000_0001001110100001_1001001011010000"; -- 0.07668416569486172
	pesos_i(5070) := b"0000000000000000_0000000000000000_0010100110100110_0001010001010001"; -- 0.16269041987186322
	pesos_i(5071) := b"1111111111111111_1111111111111111_1110000011010101_0001000011111110"; -- -0.12174886516258848
	pesos_i(5072) := b"1111111111111111_1111111111111111_1111011010111111_0010001000110000"; -- -0.03614603353596573
	pesos_i(5073) := b"0000000000000000_0000000000000000_0001110011000011_1110011000011101"; -- 0.11236417960548221
	pesos_i(5074) := b"1111111111111111_1111111111111111_1110011010100100_1111010100000000"; -- -0.09904545539148148
	pesos_i(5075) := b"0000000000000000_0000000000000000_0001101010010011_0011011011111100"; -- 0.10380881932212088
	pesos_i(5076) := b"1111111111111111_1111111111111111_1111111010101101_1111111010001111"; -- -0.005157556505431607
	pesos_i(5077) := b"0000000000000000_0000000000000000_0001110111110101_0110111000010001"; -- 0.1170262138439987
	pesos_i(5078) := b"1111111111111111_1111111111111111_1101001000000010_0101111101101011"; -- -0.17965129517789016
	pesos_i(5079) := b"1111111111111111_1111111111111111_1111001101010101_1000010111100011"; -- -0.04947627270498862
	pesos_i(5080) := b"0000000000000000_0000000000000000_0010000101100101_0110110110110011"; -- 0.13045392620666202
	pesos_i(5081) := b"0000000000000000_0000000000000000_0000111011010110_1001110101101110"; -- 0.05796226431984245
	pesos_i(5082) := b"0000000000000000_0000000000000000_0001110011010010_1001011110101100"; -- 0.11258838596688144
	pesos_i(5083) := b"1111111111111111_1111111111111111_1111001010000101_1001101111111111"; -- -0.05264878303518953
	pesos_i(5084) := b"1111111111111111_1111111111111111_1110001001110111_1100100101010011"; -- -0.11535970423297864
	pesos_i(5085) := b"0000000000000000_0000000000000000_0010010110001110_1101010110101011"; -- 0.14671073367432877
	pesos_i(5086) := b"0000000000000000_0000000000000000_0000101010101010_0110111010110111"; -- 0.04166309317079702
	pesos_i(5087) := b"1111111111111111_1111111111111111_1111010011101110_1011110111010110"; -- -0.043232092987123105
	pesos_i(5088) := b"0000000000000000_0000000000000000_0010011010101111_1110000100000011"; -- 0.15112119982117223
	pesos_i(5089) := b"1111111111111111_1111111111111111_1110110110101011_1010101110010000"; -- -0.07159927116278987
	pesos_i(5090) := b"1111111111111111_1111111111111111_1111110010010110_0100001101010001"; -- -0.013332169358755046
	pesos_i(5091) := b"1111111111111111_1111111111111111_1111101000111000_1111100110010110"; -- -0.022568131438849736
	pesos_i(5092) := b"1111111111111111_1111111111111111_1110111010010000_0011011010100001"; -- -0.06811197827932267
	pesos_i(5093) := b"0000000000000000_0000000000000000_0010111000010110_0011111100001100"; -- 0.18002695118224007
	pesos_i(5094) := b"0000000000000000_0000000000000000_0010010110000000_1110101110000110"; -- 0.1464984132691881
	pesos_i(5095) := b"0000000000000000_0000000000000000_0010000010001011_0000101011110101"; -- 0.1271216246598611
	pesos_i(5096) := b"0000000000000000_0000000000000000_0000000111010111_0000011101101110"; -- 0.007187332542214597
	pesos_i(5097) := b"1111111111111111_1111111111111111_1101110111100101_0111101000010010"; -- -0.13321721131877468
	pesos_i(5098) := b"0000000000000000_0000000000000000_0000110110110011_0110000110011110"; -- 0.0535183916822551
	pesos_i(5099) := b"0000000000000000_0000000000000000_0001101001110000_1100100010101010"; -- 0.10328344484163567
	pesos_i(5100) := b"1111111111111111_1111111111111111_1110001011011110_0111010010100100"; -- -0.1137930963910143
	pesos_i(5101) := b"0000000000000000_0000000000000000_0010001100110000_1001100001110111"; -- 0.13746025953138458
	pesos_i(5102) := b"0000000000000000_0000000000000000_0000011001111001_0000011001011011"; -- 0.02528419232775412
	pesos_i(5103) := b"1111111111111111_1111111111111111_1111110000111100_0001001010101110"; -- -0.014708359332374783
	pesos_i(5104) := b"0000000000000000_0000000000000000_0001010000101000_1110110101000011"; -- 0.07874949338070154
	pesos_i(5105) := b"0000000000000000_0000000000000000_0010101010001111_0100101111010000"; -- 0.16624902559117036
	pesos_i(5106) := b"1111111111111111_1111111111111111_1100100011000101_0100101010101001"; -- -0.21573956834871352
	pesos_i(5107) := b"0000000000000000_0000000000000000_0001011100100010_0100100010010011"; -- 0.09036687460839324
	pesos_i(5108) := b"0000000000000000_0000000000000000_0010110000001000_1011100101010000"; -- 0.17200811589921036
	pesos_i(5109) := b"0000000000000000_0000000000000000_0000101000010111_0011000101011011"; -- 0.039416393878220046
	pesos_i(5110) := b"0000000000000000_0000000000000000_0000111101000001_1011001010001101"; -- 0.0595962138012512
	pesos_i(5111) := b"1111111111111111_1111111111111111_1110111001110110_0000001110011001"; -- -0.06851174845597517
	pesos_i(5112) := b"0000000000000000_0000000000000000_0000001101010110_1111101101111011"; -- 0.013045995192254724
	pesos_i(5113) := b"0000000000000000_0000000000000000_0000110101101011_1011100001110101"; -- 0.052424934865605385
	pesos_i(5114) := b"0000000000000000_0000000000000000_0010101111101101_0101111111110111"; -- 0.17159080300548213
	pesos_i(5115) := b"0000000000000000_0000000000000000_0001100001111011_0000010010101110"; -- 0.09562710991873122
	pesos_i(5116) := b"0000000000000000_0000000000000000_0000010101111001_1101100010111100"; -- 0.021390481917043326
	pesos_i(5117) := b"1111111111111111_1111111111111111_1111101101001010_1100111100101100"; -- -0.018389751130116417
	pesos_i(5118) := b"1111111111111111_1111111111111111_1111101110110110_0111111011010010"; -- -0.016746591369960585
	pesos_i(5119) := b"0000000000000000_0000000000000000_0000101001100101_0001010101101010"; -- 0.0406049139800319
	pesos_i(5120) := b"1111111111111111_1111111111111111_1110110100000110_0010110101011100"; -- -0.07412449367695571
	pesos_i(5121) := b"1111111111111111_1111111111111111_1100101111100101_0001010111100010"; -- -0.20353568302490238
	pesos_i(5122) := b"0000000000000000_0000000000000000_0010010101111000_0001100011001111"; -- 0.14636378348920626
	pesos_i(5123) := b"1111111111111111_1111111111111111_1110100001010011_1111011000100111"; -- -0.09246884857475383
	pesos_i(5124) := b"0000000000000000_0000000000000000_0000000001010110_1110101001010100"; -- 0.0013262229955778935
	pesos_i(5125) := b"0000000000000000_0000000000000000_0010100111101010_0110011000100011"; -- 0.16373289445642766
	pesos_i(5126) := b"0000000000000000_0000000000000000_0001101111111101_1111101101010001"; -- 0.10934420331670003
	pesos_i(5127) := b"1111111111111111_1111111111111111_1101001000111101_0010100111110001"; -- -0.17875421387899645
	pesos_i(5128) := b"1111111111111111_1111111111111111_1101001000111101_1000001001000111"; -- -0.1787489487279073
	pesos_i(5129) := b"1111111111111111_1111111111111111_1100110111100010_0000101001010111"; -- -0.19576964730890042
	pesos_i(5130) := b"1111111111111111_1111111111111111_1111100001110010_0111011110000011"; -- -0.02950337470379554
	pesos_i(5131) := b"0000000000000000_0000000000000000_0001010100010010_0010110101100001"; -- 0.08230861297753649
	pesos_i(5132) := b"1111111111111111_1111111111111111_1111011001100111_1000001101100000"; -- -0.03748301424132228
	pesos_i(5133) := b"0000000000000000_0000000000000000_0010101000100100_1101101010111111"; -- 0.16462485474882232
	pesos_i(5134) := b"0000000000000000_0000000000000000_0010101100001010_1011110100000111"; -- 0.16813260487706258
	pesos_i(5135) := b"1111111111111111_1111111111111111_1100111100011000_1111100001001000"; -- -0.1910252402693316
	pesos_i(5136) := b"0000000000000000_0000000000000000_0001110011110110_1110011100111010"; -- 0.11314244427817441
	pesos_i(5137) := b"1111111111111111_1111111111111111_1110001000110001_1100001111000011"; -- -0.1164281509783173
	pesos_i(5138) := b"0000000000000000_0000000000000000_0000100101101000_0000101010000011"; -- 0.036743790524522216
	pesos_i(5139) := b"0000000000000000_0000000000000000_0000111100100001_1111011010111011"; -- 0.05911199637058031
	pesos_i(5140) := b"0000000000000000_0000000000000000_0001110111000110_0011011010011011"; -- 0.11630574495758714
	pesos_i(5141) := b"0000000000000000_0000000000000000_0000010011100010_1011011100001101"; -- 0.019084396910956727
	pesos_i(5142) := b"1111111111111111_1111111111111111_1110110011100111_1110000111001101"; -- -0.07458676104144871
	pesos_i(5143) := b"1111111111111111_1111111111111111_1111010100001110_0110010000001010"; -- -0.04274916426844409
	pesos_i(5144) := b"1111111111111111_1111111111111111_1111000100110110_0110011001000011"; -- -0.05776368015586206
	pesos_i(5145) := b"0000000000000000_0000000000000000_0010001001001101_0101000111011111"; -- 0.1339923066060874
	pesos_i(5146) := b"1111111111111111_1111111111111111_1111100001011011_0100101111100011"; -- -0.029856927006579305
	pesos_i(5147) := b"1111111111111111_1111111111111111_1111100110010111_1111001001111001"; -- -0.025025220246883143
	pesos_i(5148) := b"1111111111111111_1111111111111111_1111000000101101_1101110111000110"; -- -0.061800135821508374
	pesos_i(5149) := b"0000000000000000_0000000000000000_0010000011010010_1100010010101010"; -- 0.12821606779688577
	pesos_i(5150) := b"0000000000000000_0000000000000000_0000101101101010_0101001100100110"; -- 0.04459113767787046
	pesos_i(5151) := b"0000000000000000_0000000000000000_0010011001000111_1011100100101101"; -- 0.14953191134727803
	pesos_i(5152) := b"0000000000000000_0000000000000000_0001100001101011_1001111011000110"; -- 0.09539215400753666
	pesos_i(5153) := b"0000000000000000_0000000000000000_0001011101111111_1001110000101001"; -- 0.09179092415495689
	pesos_i(5154) := b"0000000000000000_0000000000000000_0000111011101001_1010100111011100"; -- 0.05825292235090945
	pesos_i(5155) := b"1111111111111111_1111111111111111_1111010011100010_1011001100101111"; -- -0.043415833511484085
	pesos_i(5156) := b"0000000000000000_0000000000000000_0001111100001000_1000011100101101"; -- 0.12122387742032525
	pesos_i(5157) := b"0000000000000000_0000000000000000_0000000101101111_1001100101000011"; -- 0.005609110585488193
	pesos_i(5158) := b"0000000000000000_0000000000000000_0000111010011010_0111111010011100"; -- 0.05704489993379133
	pesos_i(5159) := b"0000000000000000_0000000000000000_0000110110000001_1010111011000100"; -- 0.05276005056146986
	pesos_i(5160) := b"1111111111111111_1111111111111111_1101111110100010_1111000001101111"; -- -0.12641999513559
	pesos_i(5161) := b"1111111111111111_1111111111111111_1101111001010011_0100000100101010"; -- -0.13154213647361063
	pesos_i(5162) := b"1111111111111111_1111111111111111_1110100100000000_0010000100000110"; -- -0.08984178167176801
	pesos_i(5163) := b"1111111111111111_1111111111111111_1110100000100111_0011111010011011"; -- -0.09315117572636618
	pesos_i(5164) := b"1111111111111111_1111111111111111_1101111111111110_1001011111111001"; -- -0.12502145941184642
	pesos_i(5165) := b"1111111111111111_1111111111111111_1110100100001100_0100101011001101"; -- -0.08965618600142984
	pesos_i(5166) := b"1111111111111111_1111111111111111_1110001111101001_0011010101100111"; -- -0.10972276922132132
	pesos_i(5167) := b"1111111111111111_1111111111111111_1110110111000110_1010101110100010"; -- -0.07118727961200091
	pesos_i(5168) := b"1111111111111111_1111111111111111_1111001000011101_1111101100110101"; -- -0.05423002212232581
	pesos_i(5169) := b"0000000000000000_0000000000000000_0001000100110111_0101011001010011"; -- 0.06725062882738679
	pesos_i(5170) := b"0000000000000000_0000000000000000_0001110000111101_1100110001010100"; -- 0.11031796509419155
	pesos_i(5171) := b"0000000000000000_0000000000000000_0000100110100110_1101100101100011"; -- 0.037702166225599056
	pesos_i(5172) := b"0000000000000000_0000000000000000_0000110111110111_1011000011100001"; -- 0.05456071365383534
	pesos_i(5173) := b"1111111111111111_1111111111111111_1101011001101000_0101010001001111"; -- -0.16247056081860733
	pesos_i(5174) := b"0000000000000000_0000000000000000_0010001111001110_0001000000111000"; -- 0.13986302716932622
	pesos_i(5175) := b"0000000000000000_0000000000000000_0010010101101001_1001011011110010"; -- 0.1461424198836482
	pesos_i(5176) := b"0000000000000000_0000000000000000_0000001111110101_0010100011011001"; -- 0.015459588002461812
	pesos_i(5177) := b"1111111111111111_1111111111111111_1111100001001000_0110010110001101"; -- -0.03014531423329925
	pesos_i(5178) := b"1111111111111111_1111111111111111_1111110111100101_1010000000010000"; -- -0.008214946821440637
	pesos_i(5179) := b"1111111111111111_1111111111111111_1111010101001101_1011101010001111"; -- -0.04178270352257775
	pesos_i(5180) := b"1111111111111111_1111111111111111_1110010001110100_0100000100100101"; -- -0.10760109756514613
	pesos_i(5181) := b"1111111111111111_1111111111111111_1101010001100100_0011110000001000"; -- -0.17034554291797024
	pesos_i(5182) := b"0000000000000000_0000000000000000_0000010010000001_1011101000000000"; -- 0.017604470231147674
	pesos_i(5183) := b"0000000000000000_0000000000000000_0001111010101111_0010110010101011"; -- 0.1198604504680377
	pesos_i(5184) := b"1111111111111111_1111111111111111_1110111010111100_1000011000010011"; -- -0.06743585620125986
	pesos_i(5185) := b"1111111111111111_1111111111111111_1101010000010100_0011100000101010"; -- -0.1715664766103991
	pesos_i(5186) := b"1111111111111111_1111111111111111_1111011001101111_0111000011100101"; -- -0.03736204545047004
	pesos_i(5187) := b"0000000000000000_0000000000000000_0001000110101100_0010101011111110"; -- 0.0690333242424979
	pesos_i(5188) := b"1111111111111111_1111111111111111_1101111010100001_1011100110001101"; -- -0.13034477531608904
	pesos_i(5189) := b"0000000000000000_0000000000000000_0001010001011110_1010101100111110"; -- 0.07956953289459143
	pesos_i(5190) := b"0000000000000000_0000000000000000_0000110100001110_1101000010010110"; -- 0.05100730569724211
	pesos_i(5191) := b"0000000000000000_0000000000000000_0010011110011011_1001100000010000"; -- 0.1547179258708444
	pesos_i(5192) := b"0000000000000000_0000000000000000_0000101010111000_0111101111100111"; -- 0.04187750225951357
	pesos_i(5193) := b"0000000000000000_0000000000000000_0010011100110010_0010101000000000"; -- 0.15310919295580466
	pesos_i(5194) := b"0000000000000000_0000000000000000_0001001110111111_0111111000100010"; -- 0.07714069688336711
	pesos_i(5195) := b"0000000000000000_0000000000000000_0000100011010101_1001000000001010"; -- 0.03450870738567752
	pesos_i(5196) := b"0000000000000000_0000000000000000_0001101010000100_1011101101100111"; -- 0.10358783010185008
	pesos_i(5197) := b"1111111111111111_1111111111111111_1110101101000101_0010011100000000"; -- -0.08097606904628198
	pesos_i(5198) := b"1111111111111111_1111111111111111_1101011001001000_0000101101000011"; -- -0.16296319590589975
	pesos_i(5199) := b"0000000000000000_0000000000000000_0010110010010000_0010000010010111"; -- 0.17407420812517496
	pesos_i(5200) := b"0000000000000000_0000000000000000_0000111111101111_0101100110100101"; -- 0.062245943904167086
	pesos_i(5201) := b"1111111111111111_1111111111111111_1110011110000011_0011001001111100"; -- -0.09565433959196232
	pesos_i(5202) := b"0000000000000000_0000000000000000_0010001100001000_0111110101011001"; -- 0.13684829171825388
	pesos_i(5203) := b"0000000000000000_0000000000000000_0001100011100010_0000110001111001"; -- 0.09719922975750357
	pesos_i(5204) := b"1111111111111111_1111111111111111_1101111011110011_1011011001100111"; -- -0.1290937421225862
	pesos_i(5205) := b"1111111111111111_1111111111111111_1111011110000011_1100011000010110"; -- -0.033145541740736605
	pesos_i(5206) := b"1111111111111111_1111111111111111_1111100011101000_0110110001101101"; -- -0.027703498281794286
	pesos_i(5207) := b"0000000000000000_0000000000000000_0000101000111010_1000010101001111"; -- 0.039955455657921864
	pesos_i(5208) := b"1111111111111111_1111111111111111_1111101111011101_0000001100111010"; -- -0.016158865312029296
	pesos_i(5209) := b"0000000000000000_0000000000000000_0000001000001010_0000101110111110"; -- 0.007965787833378075
	pesos_i(5210) := b"1111111111111111_1111111111111111_1110100000011000_0100111001100001"; -- -0.09337911735561807
	pesos_i(5211) := b"1111111111111111_1111111111111111_1111011111111101_1101011000100001"; -- -0.03128301322288829
	pesos_i(5212) := b"1111111111111111_1111111111111111_1111100110010000_0000110011001011"; -- -0.02514572185146328
	pesos_i(5213) := b"0000000000000000_0000000000000000_0000001101110010_1110111001110110"; -- 0.013472465364145179
	pesos_i(5214) := b"1111111111111111_1111111111111111_1110101000100001_0000000001001011"; -- -0.08543394253999502
	pesos_i(5215) := b"0000000000000000_0000000000000000_0010101010010011_0111111111010101"; -- 0.16631316133323115
	pesos_i(5216) := b"0000000000000000_0000000000000000_0010001100111111_1111001010010111"; -- 0.1376945132492879
	pesos_i(5217) := b"0000000000000000_0000000000000000_0001011101111000_1110110011001010"; -- 0.09168891845369502
	pesos_i(5218) := b"1111111111111111_1111111111111111_1101111111010001_0011110001100010"; -- -0.12571356400870518
	pesos_i(5219) := b"1111111111111111_1111111111111111_1101001101001101_0001101111000101"; -- -0.17460466796192978
	pesos_i(5220) := b"1111111111111111_1111111111111111_1111001000001100_1001111101100110"; -- -0.05449489362376698
	pesos_i(5221) := b"0000000000000000_0000000000000000_0001011011111001_0111011110110001"; -- 0.08974407262998486
	pesos_i(5222) := b"1111111111111111_1111111111111111_1101010110011010_1110000110010010"; -- -0.16560545151472295
	pesos_i(5223) := b"1111111111111111_1111111111111111_1110011100110110_1110000111111100"; -- -0.0968188056837253
	pesos_i(5224) := b"1111111111111111_1111111111111111_1111110101001100_0000001101010111"; -- -0.010558882870812544
	pesos_i(5225) := b"1111111111111111_1111111111111111_1101000011100111_1010100000111110"; -- -0.18396519167739128
	pesos_i(5226) := b"0000000000000000_0000000000000000_0001101001001100_1101111000011111"; -- 0.10273540735149553
	pesos_i(5227) := b"0000000000000000_0000000000000000_0000100010011010_1011101100001101"; -- 0.03361100256615906
	pesos_i(5228) := b"0000000000000000_0000000000000000_0010011111001101_1110010010100111"; -- 0.15548543058460607
	pesos_i(5229) := b"0000000000000000_0000000000000000_0001110001100010_0100100110011011"; -- 0.11087474865867067
	pesos_i(5230) := b"0000000000000000_0000000000000000_0000110001011001_0000010011110101"; -- 0.04823332761879364
	pesos_i(5231) := b"1111111111111111_1111111111111111_1111010000110001_0110011000111111"; -- -0.04612122493039848
	pesos_i(5232) := b"1111111111111111_1111111111111111_1101111010000100_1101110101010000"; -- -0.13078514863647459
	pesos_i(5233) := b"0000000000000000_0000000000000000_0001101000110010_0010100111001011"; -- 0.10232793059911037
	pesos_i(5234) := b"0000000000000000_0000000000000000_0000101010111111_0000100101011110"; -- 0.041977486951820506
	pesos_i(5235) := b"1111111111111111_1111111111111111_1101101011110110_1011000011110001"; -- -0.14467329130663614
	pesos_i(5236) := b"1111111111111111_1111111111111111_1110100101011010_1010101011000110"; -- -0.08846028011508286
	pesos_i(5237) := b"1111111111111111_1111111111111111_1111010001101110_1011110110001111"; -- -0.045185234733788694
	pesos_i(5238) := b"0000000000000000_0000000000000000_0010010010101000_1011011111110111"; -- 0.14319944178202668
	pesos_i(5239) := b"0000000000000000_0000000000000000_0010100110000111_0010100111001000"; -- 0.16221867686156594
	pesos_i(5240) := b"1111111111111111_1111111111111111_1111101001111000_0001110000111001"; -- -0.021604763038116283
	pesos_i(5241) := b"1111111111111111_1111111111111111_1111101010100011_0111011100110100"; -- -0.020943212269478647
	pesos_i(5242) := b"1111111111111111_1111111111111111_1111001010111111_1001011010110010"; -- -0.051764089110487854
	pesos_i(5243) := b"1111111111111111_1111111111111111_1111110010101010_0000110011010110"; -- -0.013030240883185475
	pesos_i(5244) := b"0000000000000000_0000000000000000_0001100111011110_0101011011000101"; -- 0.10104887310391601
	pesos_i(5245) := b"0000000000000000_0000000000000000_0010001100010110_0001111100010001"; -- 0.13705629500390606
	pesos_i(5246) := b"0000000000000000_0000000000000000_0000011111011110_1011010011011100"; -- 0.030741981332248522
	pesos_i(5247) := b"1111111111111111_1111111111111111_1110001100001001_1100111011011101"; -- -0.11313159079412206
	pesos_i(5248) := b"1111111111111111_1111111111111111_1101101010001101_0001101010100001"; -- -0.14628442342150536
	pesos_i(5249) := b"0000000000000000_0000000000000000_0001010010011111_0010100001111110"; -- 0.08055356098167792
	pesos_i(5250) := b"0000000000000000_0000000000000000_0010100101101110_0110001010110010"; -- 0.16184059943674495
	pesos_i(5251) := b"1111111111111111_1111111111111111_1101000000001101_0110101100010001"; -- -0.18729525403526892
	pesos_i(5252) := b"1111111111111111_1111111111111111_1101001001001110_0100111010101010"; -- -0.17849262560232645
	pesos_i(5253) := b"0000000000000000_0000000000000000_0000000010111001_1011010100111000"; -- 0.0028336775281048525
	pesos_i(5254) := b"0000000000000000_0000000000000000_0000001111101010_0000100001101101"; -- 0.01528980895513308
	pesos_i(5255) := b"0000000000000000_0000000000000000_0001111010000111_1000110000011011"; -- 0.1192557874858942
	pesos_i(5256) := b"0000000000000000_0000000000000000_0001000011111000_0010100111000001"; -- 0.06628666831401718
	pesos_i(5257) := b"1111111111111111_1111111111111111_1110101101111001_0000001101111000"; -- -0.08018472973161751
	pesos_i(5258) := b"0000000000000000_0000000000000000_0010101101101010_0001110010010001"; -- 0.16958788428959284
	pesos_i(5259) := b"0000000000000000_0000000000000000_0000101000101100_1010010010010111"; -- 0.039743697065041446
	pesos_i(5260) := b"0000000000000000_0000000000000000_0000111001001011_1110011011111100"; -- 0.055845677006025655
	pesos_i(5261) := b"1111111111111111_1111111111111111_1101110101010001_0100001111100111"; -- -0.13547874087416822
	pesos_i(5262) := b"0000000000000000_0000000000000000_0010100000000001_1000001000110100"; -- 0.156273019489455
	pesos_i(5263) := b"0000000000000000_0000000000000000_0010000000111110_0100111001100011"; -- 0.12595071714793962
	pesos_i(5264) := b"0000000000000000_0000000000000000_0010010101010000_0100010111000011"; -- 0.14575611117183573
	pesos_i(5265) := b"1111111111111111_1111111111111111_1111011101001101_0110010111110001"; -- -0.03397524714143875
	pesos_i(5266) := b"0000000000000000_0000000000000000_0001010000011100_0000011010100000"; -- 0.07855264108528393
	pesos_i(5267) := b"1111111111111111_1111111111111111_1110101101000011_0000101001110101"; -- -0.08100828783727577
	pesos_i(5268) := b"1111111111111111_1111111111111111_1111111110110101_1011101111010000"; -- -0.0011332146769359064
	pesos_i(5269) := b"1111111111111111_1111111111111111_1110101011011100_1011101001011110"; -- -0.08256945797401553
	pesos_i(5270) := b"0000000000000000_0000000000000000_0001001110010010_0011011011100001"; -- 0.07644980425652924
	pesos_i(5271) := b"0000000000000000_0000000000000000_0001100111101001_1100100111011100"; -- 0.10122357967564667
	pesos_i(5272) := b"1111111111111111_1111111111111111_1110101011000011_0111000010100100"; -- -0.08295532215266631
	pesos_i(5273) := b"0000000000000000_0000000000000000_0001001110000011_1011010110111001"; -- 0.07622848289896982
	pesos_i(5274) := b"0000000000000000_0000000000000000_0001011111000000_1010110010100111"; -- 0.09278372830712069
	pesos_i(5275) := b"0000000000000000_0000000000000000_0001011001001101_0111101110111100"; -- 0.0871198018195907
	pesos_i(5276) := b"0000000000000000_0000000000000000_0000110110011111_0100001001101000"; -- 0.053211355625094006
	pesos_i(5277) := b"1111111111111111_1111111111111111_1110011110110101_0110111001011000"; -- -0.09488783211731992
	pesos_i(5278) := b"0000000000000000_0000000000000000_0001011010111001_1100100001011110"; -- 0.08877231886420937
	pesos_i(5279) := b"0000000000000000_0000000000000000_0001001101011111_0111111010000011"; -- 0.07567587571062373
	pesos_i(5280) := b"0000000000000000_0000000000000000_0010100001111110_0110001011110100"; -- 0.1581785055519236
	pesos_i(5281) := b"0000000000000000_0000000000000000_0010011111000010_0001001110001110"; -- 0.15530512070086422
	pesos_i(5282) := b"1111111111111111_1111111111111111_1101111010011111_1010011101111111"; -- -0.13037636909414643
	pesos_i(5283) := b"0000000000000000_0000000000000000_0000110010100011_1000110101100010"; -- 0.04937060965782838
	pesos_i(5284) := b"1111111111111111_1111111111111111_1101001001001101_0000011010110000"; -- -0.1785121747059696
	pesos_i(5285) := b"1111111111111111_1111111111111111_1110100100011000_1111010101111010"; -- -0.08946290750208437
	pesos_i(5286) := b"1111111111111111_1111111111111111_1111011000000100_1001100001111111"; -- -0.0389923753232067
	pesos_i(5287) := b"0000000000000000_0000000000000000_0010001011001100_0100111111010001"; -- 0.13593005036379366
	pesos_i(5288) := b"1111111111111111_1111111111111111_1111001001010010_0000111010111101"; -- -0.0534354007771005
	pesos_i(5289) := b"1111111111111111_1111111111111111_1111000110111001_0111010001101100"; -- -0.055763934759156836
	pesos_i(5290) := b"0000000000000000_0000000000000000_0001011011111001_1100100110011001"; -- 0.08974895462557889
	pesos_i(5291) := b"1111111111111111_1111111111111111_1110000111000001_1010010111100111"; -- -0.11813891516676354
	pesos_i(5292) := b"0000000000000000_0000000000000000_0000001100110100_1100111110110011"; -- 0.012524586869046846
	pesos_i(5293) := b"0000000000000000_0000000000000000_0010011001101001_1101100001111110"; -- 0.15005257673020972
	pesos_i(5294) := b"1111111111111111_1111111111111111_1111010101001110_0000110001100101"; -- -0.04177782564907037
	pesos_i(5295) := b"1111111111111111_1111111111111111_1100110111001111_0000110000110001"; -- -0.19605945401289243
	pesos_i(5296) := b"1111111111111111_1111111111111111_1101000111000011_0011110111001100"; -- -0.18061460266626356
	pesos_i(5297) := b"0000000000000000_0000000000000000_0011000001111001_0000111011000111"; -- 0.18934719431400926
	pesos_i(5298) := b"1111111111111111_1111111111111111_1101010101010110_0001011110101101"; -- -0.16665508305089813
	pesos_i(5299) := b"0000000000000000_0000000000000000_0000000101110100_1010011011011101"; -- 0.005686215437815317
	pesos_i(5300) := b"0000000000000000_0000000000000000_0001001001001110_1100011010111000"; -- 0.07151453011603141
	pesos_i(5301) := b"0000000000000000_0000000000000000_0000110011010110_1010001111010011"; -- 0.05015014558292377
	pesos_i(5302) := b"0000000000000000_0000000000000000_0001010110111001_1010011100110000"; -- 0.08486409102485397
	pesos_i(5303) := b"1111111111111111_1111111111111111_1111111010100010_1001101001110110"; -- -0.005331369610066765
	pesos_i(5304) := b"0000000000000000_0000000000000000_0001100001110100_0100001111111111"; -- 0.09552407235762718
	pesos_i(5305) := b"1111111111111111_1111111111111111_1110011111011001_0101100110000100"; -- -0.09433975728838358
	pesos_i(5306) := b"1111111111111111_1111111111111111_1111111000001010_0111100100011110"; -- -0.007652692975685992
	pesos_i(5307) := b"1111111111111111_1111111111111111_1101101011000010_1111100010110011"; -- -0.1454624712462787
	pesos_i(5308) := b"0000000000000000_0000000000000000_0010101010110100_0111101110111110"; -- 0.16681645768921002
	pesos_i(5309) := b"0000000000000000_0000000000000000_0000010000010110_0101011101010001"; -- 0.015965897753575927
	pesos_i(5310) := b"1111111111111111_1111111111111111_1110000000110111_0001001111011100"; -- -0.12415958289700295
	pesos_i(5311) := b"1111111111111111_1111111111111111_1101100010110100_1010011111011010"; -- -0.15349341319154966
	pesos_i(5312) := b"0000000000000000_0000000000000000_0000001111101000_1101101011010101"; -- 0.015271832427573637
	pesos_i(5313) := b"0000000000000000_0000000000000000_0010000000001101_0010011010001000"; -- 0.12520066096450663
	pesos_i(5314) := b"0000000000000000_0000000000000000_0010110000101110_0110001111010001"; -- 0.1725828538942457
	pesos_i(5315) := b"1111111111111111_1111111111111111_1111010000010110_1110110011011111"; -- -0.046525187988408996
	pesos_i(5316) := b"1111111111111111_1111111111111111_1111110001111111_1110011010101101"; -- -0.01367338449404857
	pesos_i(5317) := b"0000000000000000_0000000000000000_0001100010010110_0000111010001010"; -- 0.09603968503014629
	pesos_i(5318) := b"1111111111111111_1111111111111111_1111010011101001_1111100001001001"; -- -0.043304903098018765
	pesos_i(5319) := b"1111111111111111_1111111111111111_1110111111110100_0101101001110001"; -- -0.0626777147019161
	pesos_i(5320) := b"1111111111111111_1111111111111111_1110010110001000_0001000100100001"; -- -0.1033925337907445
	pesos_i(5321) := b"1111111111111111_1111111111111111_1101100000100000_0100000011011010"; -- -0.1557578532484234
	pesos_i(5322) := b"1111111111111111_1111111111111111_1101001000000000_0011110111110110"; -- -0.1796838068218011
	pesos_i(5323) := b"1111111111111111_1111111111111111_1110010100011111_0100110000110100"; -- -0.10499118549580715
	pesos_i(5324) := b"0000000000000000_0000000000000000_0010101000101100_0000011001000001"; -- 0.16473425952494308
	pesos_i(5325) := b"0000000000000000_0000000000000000_0000010011001001_0101000100001010"; -- 0.018696846934110646
	pesos_i(5326) := b"1111111111111111_1111111111111111_1110101000111111_0001100101010101"; -- -0.0849746863082757
	pesos_i(5327) := b"1111111111111111_1111111111111111_1111101001011001_0101010011001000"; -- -0.02207441430168161
	pesos_i(5328) := b"1111111111111111_1111111111111111_1101001100010001_1100101110001111"; -- -0.1755097175529024
	pesos_i(5329) := b"1111111111111111_1111111111111111_1110000011001011_1111000001110010"; -- -0.12188813412371048
	pesos_i(5330) := b"1111111111111111_1111111111111111_1111101110111100_0001010111000111"; -- -0.016661299689379648
	pesos_i(5331) := b"1111111111111111_1111111111111111_1111101110000110_1100011111001101"; -- -0.01747466311888744
	pesos_i(5332) := b"1111111111111111_1111111111111111_1100111010010110_1000000111011111"; -- -0.19301594061900074
	pesos_i(5333) := b"0000000000000000_0000000000000000_0001110010010011_1110001001111011"; -- 0.11163154121764794
	pesos_i(5334) := b"1111111111111111_1111111111111111_1110011110010101_1101101001000100"; -- -0.09536968071262357
	pesos_i(5335) := b"0000000000000000_0000000000000000_0001000101100000_0100110101011001"; -- 0.06787570411287032
	pesos_i(5336) := b"0000000000000000_0000000000000000_0000010000000010_1111001100000101"; -- 0.01567000274332719
	pesos_i(5337) := b"0000000000000000_0000000000000000_0010111000100101_0000001001110011"; -- 0.180252221165115
	pesos_i(5338) := b"0000000000000000_0000000000000000_0000010001101100_0010010100001010"; -- 0.017275156926024444
	pesos_i(5339) := b"1111111111111111_1111111111111111_1101111000111010_1100001011101010"; -- -0.13191587252040501
	pesos_i(5340) := b"0000000000000000_0000000000000000_0000110111011100_0100110001000111"; -- 0.054142730061897355
	pesos_i(5341) := b"1111111111111111_1111111111111111_1101000110001110_1111010011010000"; -- -0.18141241001322267
	pesos_i(5342) := b"1111111111111111_1111111111111111_1101100101101110_1100011000111010"; -- -0.1506534679114699
	pesos_i(5343) := b"0000000000000000_0000000000000000_0011011100111101_0111100011100100"; -- 0.21578174180547818
	pesos_i(5344) := b"1111111111111111_1111111111111111_1110110000000011_1010010111010110"; -- -0.07806933908328412
	pesos_i(5345) := b"0000000000000000_0000000000000000_0010011100000011_0000001010110100"; -- 0.1523896874999761
	pesos_i(5346) := b"1111111111111111_1111111111111111_1110100000001001_0100101111100110"; -- -0.09360814708551349
	pesos_i(5347) := b"1111111111111111_1111111111111111_1111001000110111_0101010110110010"; -- -0.05384315887747385
	pesos_i(5348) := b"0000000000000000_0000000000000000_0001010001100101_1011110000100011"; -- 0.07967735142092922
	pesos_i(5349) := b"0000000000000000_0000000000000000_0000101110110101_1100000001100100"; -- 0.04574205823233556
	pesos_i(5350) := b"0000000000000000_0000000000000000_0000001110100111_1001001111101111"; -- 0.014275785246569033
	pesos_i(5351) := b"0000000000000000_0000000000000000_0001100011101111_1101000010011110"; -- 0.09740928523018073
	pesos_i(5352) := b"1111111111111111_1111111111111111_1110011010011000_0110000010011101"; -- -0.09923740547549159
	pesos_i(5353) := b"1111111111111111_1111111111111111_1110100010110001_1101011100111000"; -- -0.09103636622834213
	pesos_i(5354) := b"1111111111111111_1111111111111111_1111100011100101_0100101111111010"; -- -0.027751208638956696
	pesos_i(5355) := b"0000000000000000_0000000000000000_0001001100101111_0001011011011000"; -- 0.07493727477690827
	pesos_i(5356) := b"1111111111111111_1111111111111111_1100001001111001_0110011101111111"; -- -0.24033501772164023
	pesos_i(5357) := b"1111111111111111_1111111111111111_1111111010001110_0001000001101010"; -- -0.005644773551550894
	pesos_i(5358) := b"1111111111111111_1111111111111111_1110101010101101_0101100101010101"; -- -0.08329240492837552
	pesos_i(5359) := b"0000000000000000_0000000000000000_0010000101111101_1001010111011111"; -- 0.13082253158232213
	pesos_i(5360) := b"0000000000000000_0000000000000000_0010100110100001_1111100101111000"; -- 0.16262778464673552
	pesos_i(5361) := b"1111111111111111_1111111111111111_1111111010101100_0111101001101010"; -- -0.005180691919580226
	pesos_i(5362) := b"0000000000000000_0000000000000000_0001110010111010_1101100011010000"; -- 0.11222605779616622
	pesos_i(5363) := b"0000000000000000_0000000000000000_0001001111010110_1111111111100000"; -- 0.0774993821727162
	pesos_i(5364) := b"0000000000000000_0000000000000000_0001100011111000_1010100011011110"; -- 0.09754424483985004
	pesos_i(5365) := b"1111111111111111_1111111111111111_1111100101111111_0111111001111000"; -- -0.025398345575518656
	pesos_i(5366) := b"0000000000000000_0000000000000000_0001101100001000_0010010011001110"; -- 0.10559301414575954
	pesos_i(5367) := b"0000000000000000_0000000000000000_0001001010101111_1111111100111000"; -- 0.07299800021656346
	pesos_i(5368) := b"1111111111111111_1111111111111111_1111110001100101_0011010111100101"; -- -0.014080649864287706
	pesos_i(5369) := b"0000000000000000_0000000000000000_0001111111001100_1111001100000000"; -- 0.12422102696493371
	pesos_i(5370) := b"0000000000000000_0000000000000000_0000101011101101_0010101011110000"; -- 0.04268139235477545
	pesos_i(5371) := b"1111111111111111_1111111111111111_1100010111001111_0101011001111001"; -- -0.22730502657639398
	pesos_i(5372) := b"1111111111111111_1111111111111111_1101010100000111_1000111001101101"; -- -0.16785344921737114
	pesos_i(5373) := b"1111111111111111_1111111111111111_1110110000101000_0101001011101010"; -- -0.07750970627910128
	pesos_i(5374) := b"1111111111111111_1111111111111111_1101101101011111_1011111101111110"; -- -0.143070251222391
	pesos_i(5375) := b"0000000000000000_0000000000000000_0001100111110001_1111011110011001"; -- 0.10134837603857952
	pesos_i(5376) := b"1111111111111111_1111111111111111_1111110000110011_0101100000100000"; -- -0.014841549071466693
	pesos_i(5377) := b"0000000000000000_0000000000000000_0001110011001001_0101110000011100"; -- 0.11244750665260908
	pesos_i(5378) := b"1111111111111111_1111111111111111_1110000101011010_1101001011000011"; -- -0.11970789656427885
	pesos_i(5379) := b"0000000000000000_0000000000000000_0010110000101001_0011111000011011"; -- 0.17250431216278153
	pesos_i(5380) := b"1111111111111111_1111111111111111_1111000010001101_1011110000011111"; -- -0.0603372978294946
	pesos_i(5381) := b"0000000000000000_0000000000000000_0010100010100111_0000110100000101"; -- 0.15879899380674825
	pesos_i(5382) := b"1111111111111111_1111111111111111_1101111110110001_0111101101010001"; -- -0.1261980941176103
	pesos_i(5383) := b"1111111111111111_1111111111111111_1111000111000111_1001100010110101"; -- -0.055548148882628344
	pesos_i(5384) := b"1111111111111111_1111111111111111_1101110011100111_0101001011111001"; -- -0.1370952742580415
	pesos_i(5385) := b"0000000000000000_0000000000000000_0001001010000110_1111100110010000"; -- 0.07237205271272062
	pesos_i(5386) := b"1111111111111111_1111111111111111_1101101000001101_0001001110101101"; -- -0.14823796302007464
	pesos_i(5387) := b"0000000000000000_0000000000000000_0001010101011010_0001111100001010"; -- 0.08340639104252666
	pesos_i(5388) := b"1111111111111111_1111111111111111_1111001110001011_0001000101001001"; -- -0.04865924805733139
	pesos_i(5389) := b"0000000000000000_0000000000000000_0000111100000001_1010010101100010"; -- 0.05861886638177873
	pesos_i(5390) := b"1111111111111111_1111111111111111_1110001110011000_1101000001101010"; -- -0.11094949152800514
	pesos_i(5391) := b"0000000000000000_0000000000000000_0001010100100000_0011001001000111"; -- 0.08252252811199477
	pesos_i(5392) := b"0000000000000000_0000000000000000_0000111011000011_1110011011011010"; -- 0.05767672371981465
	pesos_i(5393) := b"1111111111111111_1111111111111111_1110011100101000_1100000111001101"; -- -0.09703434709024368
	pesos_i(5394) := b"1111111111111111_1111111111111111_1110111010110101_0100100011001111"; -- -0.0675463193977045
	pesos_i(5395) := b"1111111111111111_1111111111111111_1111111011110101_1110011100110100"; -- -0.004060315855107572
	pesos_i(5396) := b"0000000000000000_0000000000000000_0000101000111111_0001100111110100"; -- 0.04002535052303621
	pesos_i(5397) := b"1111111111111111_1111111111111111_1111110010100000_0101111111011010"; -- -0.013177880665355246
	pesos_i(5398) := b"0000000000000000_0000000000000000_0010011010010110_1001100011101000"; -- 0.15073543220187485
	pesos_i(5399) := b"1111111111111111_1111111111111111_1101101011011011_0000010101001011"; -- -0.14509550973246063
	pesos_i(5400) := b"0000000000000000_0000000000000000_0010010001001010_0010100010011111"; -- 0.14175657163168245
	pesos_i(5401) := b"1111111111111111_1111111111111111_1111000011000110_0011101110000101"; -- -0.05947521218328065
	pesos_i(5402) := b"0000000000000000_0000000000000000_0010011000011101_0000010010101100"; -- 0.14888028334738485
	pesos_i(5403) := b"1111111111111111_1111111111111111_1111010001000011_1110000011101100"; -- -0.04583925483372338
	pesos_i(5404) := b"1111111111111111_1111111111111111_1110001111101010_0010111011110110"; -- -0.10970789419386694
	pesos_i(5405) := b"0000000000000000_0000000000000000_0000011111001001_0100001101000001"; -- 0.030414775158853293
	pesos_i(5406) := b"0000000000000000_0000000000000000_0001010010100010_0110001011011000"; -- 0.08060281548676773
	pesos_i(5407) := b"0000000000000000_0000000000000000_0000010011010000_0011111011100101"; -- 0.01880257688585472
	pesos_i(5408) := b"0000000000000000_0000000000000000_0000111100100111_1010000101001111"; -- 0.0591984574380379
	pesos_i(5409) := b"1111111111111111_1111111111111111_1110110000110101_1011010011101011"; -- -0.07730550057775466
	pesos_i(5410) := b"0000000000000000_0000000000000000_0001010111100011_0010000000100010"; -- 0.08549691036314595
	pesos_i(5411) := b"1111111111111111_1111111111111111_1111010111111100_0101001111100101"; -- -0.039118534750848616
	pesos_i(5412) := b"0000000000000000_0000000000000000_0010110111000011_1000110101101100"; -- 0.1787651433582595
	pesos_i(5413) := b"0000000000000000_0000000000000000_0001100001101110_1111110011111100"; -- 0.09544354588832896
	pesos_i(5414) := b"0000000000000000_0000000000000000_0000001110100001_1001001100101011"; -- 0.014184186896401881
	pesos_i(5415) := b"1111111111111111_1111111111111111_1110110011010000_1110111000001011"; -- -0.07493698333669056
	pesos_i(5416) := b"1111111111111111_1111111111111111_1111001100110111_1011101101101011"; -- -0.04993084573340438
	pesos_i(5417) := b"0000000000000000_0000000000000000_0000001111111011_1011101000010101"; -- 0.015559797354185131
	pesos_i(5418) := b"0000000000000000_0000000000000000_0001001011000111_1100001101101111"; -- 0.07336064772212804
	pesos_i(5419) := b"0000000000000000_0000000000000000_0010101001011101_1010001101000000"; -- 0.16549129788160022
	pesos_i(5420) := b"0000000000000000_0000000000000000_0010111111110101_1011011011011010"; -- 0.18734305212217542
	pesos_i(5421) := b"1111111111111111_1111111111111111_1101110011001010_0111110000010110"; -- -0.13753532856204892
	pesos_i(5422) := b"1111111111111111_1111111111111111_1110010101011010_1000101010010101"; -- -0.10408719887224513
	pesos_i(5423) := b"1111111111111111_1111111111111111_1101111110100111_0000011010101110"; -- -0.12635763410748918
	pesos_i(5424) := b"0000000000000000_0000000000000000_0000011010110100_0100101110011100"; -- 0.026188588781369305
	pesos_i(5425) := b"1111111111111111_1111111111111111_1111011100010000_1111100011001111"; -- -0.034897279223860385
	pesos_i(5426) := b"0000000000000000_0000000000000000_0010011101010001_0110000011011111"; -- 0.1535854859591268
	pesos_i(5427) := b"0000000000000000_0000000000000000_0000110101000101_0011110000111100"; -- 0.051837696629984935
	pesos_i(5428) := b"0000000000000000_0000000000000000_0001101000111000_1111000101001011"; -- 0.10243137434337851
	pesos_i(5429) := b"0000000000000000_0000000000000000_0010010001111110_1111110111001100"; -- 0.14256273493451366
	pesos_i(5430) := b"1111111111111111_1111111111111111_1101100110011111_0011011000000011"; -- -0.149914383281781
	pesos_i(5431) := b"1111111111111111_1111111111111111_1101111101110001_0110000001101001"; -- -0.12717626044498445
	pesos_i(5432) := b"0000000000000000_0000000000000000_0000111111100000_1000110101100010"; -- 0.06202014588189844
	pesos_i(5433) := b"1111111111111111_1111111111111111_1111001001011010_1100101100001001"; -- -0.05330210710440015
	pesos_i(5434) := b"0000000000000000_0000000000000000_0010000000010001_0100000000001011"; -- 0.12526321677623456
	pesos_i(5435) := b"0000000000000000_0000000000000000_0001101101010000_1010110001011110"; -- 0.10669972694847782
	pesos_i(5436) := b"0000000000000000_0000000000000000_0001111111010110_1100010110101010"; -- 0.12437091263579496
	pesos_i(5437) := b"0000000000000000_0000000000000000_0001111100111001_1101101001001100"; -- 0.12197651243198938
	pesos_i(5438) := b"0000000000000000_0000000000000000_0001100000011010_0101101001001001"; -- 0.09415210994931825
	pesos_i(5439) := b"1111111111111111_1111111111111111_1101101101100001_1011001101111000"; -- -0.14304045028836082
	pesos_i(5440) := b"1111111111111111_1111111111111111_1101111000100101_1111001101100001"; -- -0.13223341832026744
	pesos_i(5441) := b"1111111111111111_1111111111111111_1101111100111101_0110110111101011"; -- -0.127968912228063
	pesos_i(5442) := b"1111111111111111_1111111111111111_1101010010111000_0111001110010101"; -- -0.16906049350406585
	pesos_i(5443) := b"0000000000000000_0000000000000000_0010101110101000_1100111001000011"; -- 0.17054452082361865
	pesos_i(5444) := b"0000000000000000_0000000000000000_0000100110100100_1111010110110101"; -- 0.03767333674820276
	pesos_i(5445) := b"0000000000000000_0000000000000000_0000100011100000_0110001101100110"; -- 0.03467389332629277
	pesos_i(5446) := b"1111111111111111_1111111111111111_1111100100001111_0011001111100001"; -- -0.02711177599339898
	pesos_i(5447) := b"1111111111111111_1111111111111111_1110111001100110_1101010110110101"; -- -0.06874336555970835
	pesos_i(5448) := b"0000000000000000_0000000000000000_0010100111011000_1001010100000000"; -- 0.16346102957065084
	pesos_i(5449) := b"0000000000000000_0000000000000000_0000101100000010_0110100011100101"; -- 0.04300551979970625
	pesos_i(5450) := b"1111111111111111_1111111111111111_1100111111111100_0101100010001111"; -- -0.18755575656828327
	pesos_i(5451) := b"0000000000000000_0000000000000000_0001010010010010_0000101110001101"; -- 0.08035347164490238
	pesos_i(5452) := b"0000000000000000_0000000000000000_0001111110111100_1000011110001000"; -- 0.12397048053452792
	pesos_i(5453) := b"1111111111111111_1111111111111111_1110110011100111_0101111010011001"; -- -0.07459458130655512
	pesos_i(5454) := b"1111111111111111_1111111111111111_1111001001001111_1010110000011001"; -- -0.053471797837178654
	pesos_i(5455) := b"1111111111111111_1111111111111111_1100111111000011_1100111000110001"; -- -0.18841849614439388
	pesos_i(5456) := b"1111111111111111_1111111111111111_1110100011100001_1111110010100001"; -- -0.09030171464072638
	pesos_i(5457) := b"1111111111111111_1111111111111111_1110100011110110_1000001111110101"; -- -0.08998847268393664
	pesos_i(5458) := b"1111111111111111_1111111111111111_1100111011000010_0110100010111010"; -- -0.1923460526774853
	pesos_i(5459) := b"1111111111111111_1111111111111111_1100110100110111_0111001011011000"; -- -0.19837267149345317
	pesos_i(5460) := b"0000000000000000_0000000000000000_0001100010011011_0100111011000100"; -- 0.09611980711471066
	pesos_i(5461) := b"1111111111111111_1111111111111111_1111101100010111_1001111100100110"; -- -0.01917081182051257
	pesos_i(5462) := b"0000000000000000_0000000000000000_0001111111101111_1011110000011000"; -- 0.1247518119358777
	pesos_i(5463) := b"0000000000000000_0000000000000000_0010000110010010_0010001110001000"; -- 0.1311361510434442
	pesos_i(5464) := b"0000000000000000_0000000000000000_0010001011101100_0010111101111111"; -- 0.13641640531902413
	pesos_i(5465) := b"1111111111111111_1111111111111111_1110111010011010_1111100010101011"; -- -0.06794782471202807
	pesos_i(5466) := b"1111111111111111_1111111111111111_1100110011001001_1010010101000111"; -- -0.20004813207579628
	pesos_i(5467) := b"1111111111111111_1111111111111111_1100101110010110_0101110010111110"; -- -0.20473690375396486
	pesos_i(5468) := b"0000000000000000_0000000000000000_0000101001100001_0000010001101011"; -- 0.04054286590196195
	pesos_i(5469) := b"1111111111111111_1111111111111111_1111101101100011_1011001010110010"; -- -0.018009978900655747
	pesos_i(5470) := b"0000000000000000_0000000000000000_0010101100111110_0100101100110111"; -- 0.16891927815517657
	pesos_i(5471) := b"0000000000000000_0000000000000000_0000111101110010_1111000110111010"; -- 0.060347660067724976
	pesos_i(5472) := b"1111111111111111_1111111111111111_1111110110011010_1011110001100110"; -- -0.009357667147455626
	pesos_i(5473) := b"1111111111111111_1111111111111111_1101000110000000_0001001000111100"; -- -0.18163953805995045
	pesos_i(5474) := b"1111111111111111_1111111111111111_1111100001100001_0001111100000010"; -- -0.029768049259019685
	pesos_i(5475) := b"0000000000000000_0000000000000000_0001111100001111_0001111000000001"; -- 0.1213244201747856
	pesos_i(5476) := b"0000000000000000_0000000000000000_0000101001001101_1001011010011110"; -- 0.04024640430801526
	pesos_i(5477) := b"0000000000000000_0000000000000000_0001000001000010_1010011001111011"; -- 0.06351700313500978
	pesos_i(5478) := b"1111111111111111_1111111111111111_1110100110000001_0111111001100111"; -- -0.08786783193324753
	pesos_i(5479) := b"0000000000000000_0000000000000000_0001110101100011_1000011011001010"; -- 0.11479990406328892
	pesos_i(5480) := b"1111111111111111_1111111111111111_1101111010000000_0001011010000101"; -- -0.13085803266147208
	pesos_i(5481) := b"1111111111111111_1111111111111111_1111101010101110_0111011001010110"; -- -0.02077541735710177
	pesos_i(5482) := b"1111111111111111_1111111111111111_1100111000011110_0100100110000010"; -- -0.19485035498546746
	pesos_i(5483) := b"1111111111111111_1111111111111111_1110110000011011_0110000001111110"; -- -0.07770726138083728
	pesos_i(5484) := b"1111111111111111_1111111111111111_1111000100110011_0110111001011100"; -- -0.057808973843892573
	pesos_i(5485) := b"1111111111111111_1111111111111111_1101100010010110_1101011010100000"; -- -0.15394838909023417
	pesos_i(5486) := b"1111111111111111_1111111111111111_1111101011001010_0010110100110010"; -- -0.020352530775957934
	pesos_i(5487) := b"1111111111111111_1111111111111111_1111111101110100_1111111100010011"; -- -0.0021210269269275033
	pesos_i(5488) := b"1111111111111111_1111111111111111_1110000110110001_1101000110111000"; -- -0.11838044403755292
	pesos_i(5489) := b"0000000000000000_0000000000000000_0011010001111001_1010101100111011"; -- 0.2049815195090906
	pesos_i(5490) := b"1111111111111111_1111111111111111_1111001010001000_0001110110111110"; -- -0.052610532022643666
	pesos_i(5491) := b"0000000000000000_0000000000000000_0000101011100101_0011100101101111"; -- 0.04256018591735503
	pesos_i(5492) := b"0000000000000000_0000000000000000_0000010000000011_0010110000111010"; -- 0.015673412562971632
	pesos_i(5493) := b"1111111111111111_1111111111111111_1110101011001001_0011011110010010"; -- -0.08286717116291996
	pesos_i(5494) := b"1111111111111111_1111111111111111_1110011000001001_0110010100000111"; -- -0.1014191491718629
	pesos_i(5495) := b"1111111111111111_1111111111111111_1101000101001100_1000101011010010"; -- -0.1824258076674026
	pesos_i(5496) := b"1111111111111111_1111111111111111_1111111000111111_0101001110100000"; -- -0.006846211818952147
	pesos_i(5497) := b"0000000000000000_0000000000000000_0000011010000110_0010000110000100"; -- 0.02548417530725236
	pesos_i(5498) := b"0000000000000000_0000000000000000_0010000011000111_1101110111110001"; -- 0.12804972766327832
	pesos_i(5499) := b"1111111111111111_1111111111111111_1111001111101000_0001101100001010"; -- -0.04723959938476065
	pesos_i(5500) := b"0000000000000000_0000000000000000_0000001010011000_1110011100111011"; -- 0.010145618254681254
	pesos_i(5501) := b"0000000000000000_0000000000000000_0001100110010100_0110011011100101"; -- 0.09992068369137652
	pesos_i(5502) := b"0000000000000000_0000000000000000_0001110010001100_0000010111001000"; -- 0.11151157504119003
	pesos_i(5503) := b"1111111111111111_1111111111111111_1110001111101011_1100010011001011"; -- -0.10968370469611853
	pesos_i(5504) := b"1111111111111111_1111111111111111_1111000000000010_1111001100010010"; -- -0.06245499437725834
	pesos_i(5505) := b"1111111111111111_1111111111111111_1110000011010111_0100100100101010"; -- -0.12171499950516158
	pesos_i(5506) := b"1111111111111111_1111111111111111_1101100010111010_0101100011111101"; -- -0.15340656121689625
	pesos_i(5507) := b"1111111111111111_1111111111111111_1100101011101111_0100110001011110"; -- -0.2072860976233616
	pesos_i(5508) := b"0000000000000000_0000000000000000_0010101110010101_0101100100101000"; -- 0.17024762360497925
	pesos_i(5509) := b"0000000000000000_0000000000000000_0001111001001100_1101011010011100"; -- 0.11835995975582397
	pesos_i(5510) := b"0000000000000000_0000000000000000_0000010001100010_0111111000100010"; -- 0.017127879480669315
	pesos_i(5511) := b"0000000000000000_0000000000000000_0010001011011111_1110111001110111"; -- 0.13622942354724638
	pesos_i(5512) := b"1111111111111111_1111111111111111_1110010001100101_1101000011011010"; -- -0.10782141369913331
	pesos_i(5513) := b"0000000000000000_0000000000000000_0001010101010001_0011000000011001"; -- 0.08327007870475416
	pesos_i(5514) := b"1111111111111111_1111111111111111_1111001101101010_0111011111100111"; -- -0.04915667165267341
	pesos_i(5515) := b"1111111111111111_1111111111111111_1101001011111010_1000111101111111"; -- -0.17586424958612398
	pesos_i(5516) := b"1111111111111111_1111111111111111_1111111110111000_0010110011101011"; -- -0.0010959554706297396
	pesos_i(5517) := b"0000000000000000_0000000000000000_0000001101101101_0000110000111010"; -- 0.013382686861497697
	pesos_i(5518) := b"1111111111111111_1111111111111111_1111111010101100_1100110111000001"; -- -0.005175724432171438
	pesos_i(5519) := b"1111111111111111_1111111111111111_1111010101101101_0111000111001100"; -- -0.041298759094781284
	pesos_i(5520) := b"0000000000000000_0000000000000000_0011010001000001_0000110000101001"; -- 0.20411754604432686
	pesos_i(5521) := b"1111111111111111_1111111111111111_1110101001100000_0010111001001101"; -- -0.08446989659278362
	pesos_i(5522) := b"1111111111111111_1111111111111111_1110011010001101_1000010011101101"; -- -0.09940308773574295
	pesos_i(5523) := b"0000000000000000_0000000000000000_0001100101111100_1010100100001010"; -- 0.09955841541396337
	pesos_i(5524) := b"0000000000000000_0000000000000000_0000100000111100_1110110101110111"; -- 0.03217968133702223
	pesos_i(5525) := b"1111111111111111_1111111111111111_1110101011000110_1101101110110110"; -- -0.0829031640169939
	pesos_i(5526) := b"0000000000000000_0000000000000000_0000101101010001_1100010110011111"; -- 0.04421649108039695
	pesos_i(5527) := b"1111111111111111_1111111111111111_1110000011011010_0111000111110101"; -- -0.12166679170631214
	pesos_i(5528) := b"1111111111111111_1111111111111111_1111101110110100_1000101010101001"; -- -0.016776403255394083
	pesos_i(5529) := b"0000000000000000_0000000000000000_0000011010011100_0010000100011010"; -- 0.02581984414361166
	pesos_i(5530) := b"0000000000000000_0000000000000000_0000011001001111_1000001011110110"; -- 0.024650750292560454
	pesos_i(5531) := b"0000000000000000_0000000000000000_0001111101101010_0110111000110011"; -- 0.12271774998575141
	pesos_i(5532) := b"0000000000000000_0000000000000000_0000011010101011_1101101111110010"; -- 0.0260598627777636
	pesos_i(5533) := b"1111111111111111_1111111111111111_1101010011001000_1001000111010001"; -- -0.16881455088557457
	pesos_i(5534) := b"1111111111111111_1111111111111111_1110001011101111_0000010110101100"; -- -0.11354031140876239
	pesos_i(5535) := b"1111111111111111_1111111111111111_1101101111000111_0010011110111100"; -- -0.14149238261843594
	pesos_i(5536) := b"0000000000000000_0000000000000000_0001001010100111_0111000011110000"; -- 0.07286744944919207
	pesos_i(5537) := b"1111111111111111_1111111111111111_1111111000110010_0010010111010011"; -- -0.007047306136950064
	pesos_i(5538) := b"1111111111111111_1111111111111111_1110011100111110_0011100110111110"; -- -0.09670676340100244
	pesos_i(5539) := b"1111111111111111_1111111111111111_1101000001111000_0010100110101101"; -- -0.18566646113951385
	pesos_i(5540) := b"1111111111111111_1111111111111111_1111111001011011_1000010100011011"; -- -0.006416016511568451
	pesos_i(5541) := b"1111111111111111_1111111111111111_1101100110100110_1001100000001101"; -- -0.14980172819750484
	pesos_i(5542) := b"1111111111111111_1111111111111111_1111001110001111_0000010010001111"; -- -0.04859897154503051
	pesos_i(5543) := b"0000000000000000_0000000000000000_0001100100110010_1110001011111110"; -- 0.09843271924441212
	pesos_i(5544) := b"1111111111111111_1111111111111111_1100000110011111_0011101101000101"; -- -0.24366406975199165
	pesos_i(5545) := b"1111111111111111_1111111111111111_1111011110010000_0001101000010100"; -- -0.03295743005979476
	pesos_i(5546) := b"0000000000000000_0000000000000000_0001101000110110_1110010000000001"; -- 0.10240006460847942
	pesos_i(5547) := b"0000000000000000_0000000000000000_0001100110000111_0100010011010010"; -- 0.09972028861410243
	pesos_i(5548) := b"1111111111111111_1111111111111111_1111001101110001_1000100110001110"; -- -0.04904880798292539
	pesos_i(5549) := b"1111111111111111_1111111111111111_1111100011101001_1110001101001001"; -- -0.027681154955980065
	pesos_i(5550) := b"1111111111111111_1111111111111111_1101101010010010_1000001111011010"; -- -0.14620185780355696
	pesos_i(5551) := b"1111111111111111_1111111111111111_1100110000011111_0111011011011101"; -- -0.20264489267637897
	pesos_i(5552) := b"0000000000000000_0000000000000000_0000101011110000_0100010010011111"; -- 0.04272869953423663
	pesos_i(5553) := b"0000000000000000_0000000000000000_0000011111001110_0100111110010010"; -- 0.03049180322842152
	pesos_i(5554) := b"1111111111111111_1111111111111111_1101110111101111_0011010101101010"; -- -0.13306871574823495
	pesos_i(5555) := b"0000000000000000_0000000000000000_0010000100111001_0100100010011001"; -- 0.12978032808178538
	pesos_i(5556) := b"0000000000000000_0000000000000000_0011011110100100_0101000010101111"; -- 0.21735100042361352
	pesos_i(5557) := b"1111111111111111_1111111111111111_1101111111100001_0000011011010110"; -- -0.12547261490961475
	pesos_i(5558) := b"0000000000000000_0000000000000000_0010001000111011_0010100101011101"; -- 0.13371523398566154
	pesos_i(5559) := b"1111111111111111_1111111111111111_1111101110100100_1001100011011001"; -- -0.017019698225634323
	pesos_i(5560) := b"0000000000000000_0000000000000000_0010101010110100_0000100100100000"; -- 0.16680962592481066
	pesos_i(5561) := b"0000000000000000_0000000000000000_0001110000100001_1111000111100010"; -- 0.10989295727501396
	pesos_i(5562) := b"1111111111111111_1111111111111111_1111101011111111_1111110011000110"; -- -0.019531442219371708
	pesos_i(5563) := b"1111111111111111_1111111111111111_1110000010000100_1010010000110110"; -- -0.12297605222164493
	pesos_i(5564) := b"1111111111111111_1111111111111111_1101110000101100_1101100100111011"; -- -0.13994066543761496
	pesos_i(5565) := b"1111111111111111_1111111111111111_1111001001101101_1101001101001101"; -- -0.053011697473081626
	pesos_i(5566) := b"0000000000000000_0000000000000000_0001001100011000_1001011110110000"; -- 0.07459400212206416
	pesos_i(5567) := b"1111111111111111_1111111111111111_1110110001011011_1001010000101001"; -- -0.07672761918557422
	pesos_i(5568) := b"0000000000000000_0000000000000000_0000101011101111_0010110011110111"; -- 0.04271203076310034
	pesos_i(5569) := b"1111111111111111_1111111111111111_1110001101100010_0001010101010011"; -- -0.11178461757802305
	pesos_i(5570) := b"1111111111111111_1111111111111111_1110100110101111_0101111110101100"; -- -0.08716775943810424
	pesos_i(5571) := b"1111111111111111_1111111111111111_1111110111010100_1111000001101001"; -- -0.00846955721222757
	pesos_i(5572) := b"0000000000000000_0000000000000000_0000101111010010_1001010100000101"; -- 0.04618197803929669
	pesos_i(5573) := b"0000000000000000_0000000000000000_0010101010010111_1100111101110010"; -- 0.1663789417702297
	pesos_i(5574) := b"0000000000000000_0000000000000000_0010010001101110_1001110011000010"; -- 0.14231281038148663
	pesos_i(5575) := b"1111111111111111_1111111111111111_1110100101011100_0010111010011110"; -- -0.08843716286118636
	pesos_i(5576) := b"0000000000000000_0000000000000000_0000001000000101_1011011000001011"; -- 0.007899644487932657
	pesos_i(5577) := b"1111111111111111_1111111111111111_1101111000100010_1101101011000110"; -- -0.13228066123652615
	pesos_i(5578) := b"0000000000000000_0000000000000000_0001010101111100_0001011110001101"; -- 0.08392474361435154
	pesos_i(5579) := b"1111111111111111_1111111111111111_1110101010111010_1001010001000100"; -- -0.08309052782618044
	pesos_i(5580) := b"0000000000000000_0000000000000000_0001101000110010_0111110100001011"; -- 0.102332892554435
	pesos_i(5581) := b"0000000000000000_0000000000000000_0000101111000100_1001101100001111"; -- 0.04596871477655002
	pesos_i(5582) := b"1111111111111111_1111111111111111_1101011000010000_0101001000000010"; -- -0.16381347128882823
	pesos_i(5583) := b"1111111111111111_1111111111111111_1110110111001001_1011111100000101"; -- -0.07114034768455024
	pesos_i(5584) := b"0000000000000000_0000000000000000_0001010000101001_0111010010010101"; -- 0.07875755918500049
	pesos_i(5585) := b"1111111111111111_1111111111111111_1101110111100001_1110100101001001"; -- -0.1332716176347154
	pesos_i(5586) := b"0000000000000000_0000000000000000_0001010001011101_0111111111011110"; -- 0.07955168889999133
	pesos_i(5587) := b"1111111111111111_1111111111111111_1111010111010011_1001001101100101"; -- -0.03974036001918426
	pesos_i(5588) := b"1111111111111111_1111111111111111_1110110101001000_0000011010110100"; -- -0.07311971770871617
	pesos_i(5589) := b"1111111111111111_1111111111111111_1101101000110100_0000001100001101"; -- -0.14764386106661076
	pesos_i(5590) := b"1111111111111111_1111111111111111_1110011011110101_0010110110011101"; -- -0.0978213778896217
	pesos_i(5591) := b"0000000000000000_0000000000000000_0001101111111111_1110011100111110"; -- 0.109373524428854
	pesos_i(5592) := b"0000000000000000_0000000000000000_0000001111010000_1010000110001110"; -- 0.014902207586255248
	pesos_i(5593) := b"0000000000000000_0000000000000000_0011110110011111_1100111111110101"; -- 0.2407197927017107
	pesos_i(5594) := b"0000000000000000_0000000000000000_0011000001100001_0000110000000100"; -- 0.18898081865826682
	pesos_i(5595) := b"0000000000000000_0000000000000000_0000101000101111_1010011010111001"; -- 0.0397896004239304
	pesos_i(5596) := b"1111111111111111_1111111111111111_1110100100010010_0001000101110001"; -- -0.08956805226913157
	pesos_i(5597) := b"0000000000000000_0000000000000000_0010000110010011_0110101100100100"; -- 0.13115567813034434
	pesos_i(5598) := b"1111111111111111_1111111111111111_1101111000101100_1111001011100000"; -- -0.13212663687656426
	pesos_i(5599) := b"1111111111111111_1111111111111111_1111001110010010_0010100001011101"; -- -0.048551060885089585
	pesos_i(5600) := b"0000000000000000_0000000000000000_0000010011011110_1111000110111100"; -- 0.019026859609323127
	pesos_i(5601) := b"0000000000000000_0000000000000000_0000100111001101_1000000001011100"; -- 0.03829195249044487
	pesos_i(5602) := b"0000000000000000_0000000000000000_0000000110101111_0011111000101111"; -- 0.0065802444963253826
	pesos_i(5603) := b"1111111111111111_1111111111111111_1110000010110010_0010010011001110"; -- -0.12228174187682787
	pesos_i(5604) := b"1111111111111111_1111111111111111_1101000101101101_0000001101110100"; -- -0.18193033616401405
	pesos_i(5605) := b"0000000000000000_0000000000000000_0010011111001011_0101011011010111"; -- 0.15544646019699693
	pesos_i(5606) := b"0000000000000000_0000000000000000_0000100000001111_0011101110110000"; -- 0.03148243938564507
	pesos_i(5607) := b"0000000000000000_0000000000000000_0010111110100011_1100010010010100"; -- 0.1860926496526018
	pesos_i(5608) := b"1111111111111111_1111111111111111_1110111011101000_1110001110000101"; -- -0.06675889961670764
	pesos_i(5609) := b"1111111111111111_1111111111111111_1101000011011100_1101010000100110"; -- -0.1841304214601543
	pesos_i(5610) := b"0000000000000000_0000000000000000_0010111010001101_1000010001101110"; -- 0.1818468827802322
	pesos_i(5611) := b"1111111111111111_1111111111111111_1110101011100011_1000000101011110"; -- -0.08246604400118518
	pesos_i(5612) := b"0000000000000000_0000000000000000_0001001010111001_1011000011001101"; -- 0.07314591420192323
	pesos_i(5613) := b"0000000000000000_0000000000000000_0001100110001011_0000111100010000"; -- 0.09977811946531401
	pesos_i(5614) := b"1111111111111111_1111111111111111_1101001001000001_0100010001100010"; -- -0.17869160269293954
	pesos_i(5615) := b"1111111111111111_1111111111111111_1111000001110101_1110010110111010"; -- -0.06070102901482735
	pesos_i(5616) := b"0000000000000000_0000000000000000_0001000111110110_1111000110101100"; -- 0.0701743168688872
	pesos_i(5617) := b"0000000000000000_0000000000000000_0001100001110111_0100000100100101"; -- 0.09556967881322742
	pesos_i(5618) := b"0000000000000000_0000000000000000_0010111101101011_0100010110100101"; -- 0.18523059162657407
	pesos_i(5619) := b"0000000000000000_0000000000000000_0010011111001100_0111101101100101"; -- 0.1554638977759375
	pesos_i(5620) := b"1111111111111111_1111111111111111_1111010111000001_1010101100110110"; -- -0.04001359879381247
	pesos_i(5621) := b"0000000000000000_0000000000000000_0010001001111110_1011101100000101"; -- 0.13474625469395368
	pesos_i(5622) := b"1111111111111111_1111111111111111_1101101101011011_0011101001101010"; -- -0.143139218553188
	pesos_i(5623) := b"1111111111111111_1111111111111111_1110001001011111_0000001111010011"; -- -0.11573768710221242
	pesos_i(5624) := b"1111111111111111_1111111111111111_1101001000010100_0001011100011111"; -- -0.17938094602712495
	pesos_i(5625) := b"0000000000000000_0000000000000000_0001010110100100_1101111111010000"; -- 0.0845470315801673
	pesos_i(5626) := b"0000000000000000_0000000000000000_0010001001110000_0001100001110011"; -- 0.1345229415705243
	pesos_i(5627) := b"1111111111111111_1111111111111111_1111010110101111_1001111001011101"; -- -0.04028902268467777
	pesos_i(5628) := b"0000000000000000_0000000000000000_0001000011100111_0100011000000010"; -- 0.0660289530584261
	pesos_i(5629) := b"0000000000000000_0000000000000000_0001001010000001_1110011011111010"; -- 0.07229465115337586
	pesos_i(5630) := b"1111111111111111_1111111111111111_1110111001110111_1111001010001110"; -- -0.06848224663108846
	pesos_i(5631) := b"0000000000000000_0000000000000000_0010100010100001_0100010010100110"; -- 0.15871075688571923
	pesos_i(5632) := b"1111111111111111_1111111111111111_1110100110011100_1100010111001111"; -- -0.08745158848574495
	pesos_i(5633) := b"1111111111111111_1111111111111111_1110111110000101_0111110100100110"; -- -0.06436937171493748
	pesos_i(5634) := b"1111111111111111_1111111111111111_1101111100010101_1000011001111000"; -- -0.12857780038081046
	pesos_i(5635) := b"1111111111111111_1111111111111111_1110011100010011_1111100001010001"; -- -0.0973515322910615
	pesos_i(5636) := b"0000000000000000_0000000000000000_0001101101110100_1101001100100011"; -- 0.10725135433784155
	pesos_i(5637) := b"0000000000000000_0000000000000000_0001011010101010_0111010101000010"; -- 0.08853848320467461
	pesos_i(5638) := b"0000000000000000_0000000000000000_0000101011111010_0001010010110001"; -- 0.04287843061298677
	pesos_i(5639) := b"1111111111111111_1111111111111111_1101000110111001_1010101011101010"; -- -0.18076068674279663
	pesos_i(5640) := b"0000000000000000_0000000000000000_0001011101111000_0010001011100101"; -- 0.09167688455582129
	pesos_i(5641) := b"0000000000000000_0000000000000000_0010011100001010_0000000100110011"; -- 0.152496409355099
	pesos_i(5642) := b"1111111111111111_1111111111111111_1101100111010010_0000001110111101"; -- -0.14913918152123437
	pesos_i(5643) := b"0000000000000000_0000000000000000_0000101010100110_0001110000000000"; -- 0.04159712802270327
	pesos_i(5644) := b"0000000000000000_0000000000000000_0000110011011010_1101110101110001"; -- 0.050214614885783576
	pesos_i(5645) := b"0000000000000000_0000000000000000_0000000010111011_1001000111000100"; -- 0.002862081901372965
	pesos_i(5646) := b"0000000000000000_0000000000000000_0000100000001101_1110111100011110"; -- 0.03146261670354708
	pesos_i(5647) := b"1111111111111111_1111111111111111_1101010010010011_0000110001100011"; -- -0.16963121961861688
	pesos_i(5648) := b"0000000000000000_0000000000000000_0000111110100011_1011101110010111"; -- 0.0610921138440611
	pesos_i(5649) := b"0000000000000000_0000000000000000_0010110110110010_0110000111111000"; -- 0.17850315390184857
	pesos_i(5650) := b"0000000000000000_0000000000000000_0001110100100001_0011110001111101"; -- 0.1137883955061662
	pesos_i(5651) := b"1111111111111111_1111111111111111_1111100001010000_0100001000110111"; -- -0.030025350122610123
	pesos_i(5652) := b"0000000000000000_0000000000000000_0010101000100011_1100100010101101"; -- 0.16460851885805972
	pesos_i(5653) := b"0000000000000000_0000000000000000_0000001110110010_1011010010100011"; -- 0.014445581134766822
	pesos_i(5654) := b"1111111111111111_1111111111111111_1111010011101110_1110010100011000"; -- -0.043229753201162485
	pesos_i(5655) := b"0000000000000000_0000000000000000_0000000101101000_0000000110111110"; -- 0.005493267946148822
	pesos_i(5656) := b"0000000000000000_0000000000000000_0010011010000001_0100001100010010"; -- 0.15040988155669188
	pesos_i(5657) := b"0000000000000000_0000000000000000_0001111000011110_0001101101010110"; -- 0.11764689302544712
	pesos_i(5658) := b"0000000000000000_0000000000000000_0010001001000100_1110010011110111"; -- 0.13386374510968346
	pesos_i(5659) := b"0000000000000000_0000000000000000_0010000111001101_0100100000100010"; -- 0.13203860117163813
	pesos_i(5660) := b"0000000000000000_0000000000000000_0010000100011011_1011111100101001"; -- 0.12932963127445596
	pesos_i(5661) := b"1111111111111111_1111111111111111_1110101011010110_1001100011101001"; -- -0.0826630050947023
	pesos_i(5662) := b"0000000000000000_0000000000000000_0000001110001101_1101000010100000"; -- 0.013882674185747207
	pesos_i(5663) := b"1111111111111111_1111111111111111_1110010110110100_0110100001100100"; -- -0.10271594575510191
	pesos_i(5664) := b"0000000000000000_0000000000000000_0001100000111101_0101111111010001"; -- 0.09468649728568507
	pesos_i(5665) := b"0000000000000000_0000000000000000_0001010010010110_0100000011110010"; -- 0.08041768941075272
	pesos_i(5666) := b"0000000000000000_0000000000000000_0001100101111110_1000101000100110"; -- 0.09958709163580981
	pesos_i(5667) := b"0000000000000000_0000000000000000_0010111101100010_1100110010101000"; -- 0.18510130985708712
	pesos_i(5668) := b"1111111111111111_1111111111111111_1101110010111101_0001101011011011"; -- -0.1377394882515827
	pesos_i(5669) := b"0000000000000000_0000000000000000_0001101000111100_0010000111010100"; -- 0.1024800436847143
	pesos_i(5670) := b"1111111111111111_1111111111111111_1101011000000110_1100100111011000"; -- -0.16395891645800564
	pesos_i(5671) := b"1111111111111111_1111111111111111_1111110000001100_1011001011111010"; -- -0.01543122665811622
	pesos_i(5672) := b"0000000000000000_0000000000000000_0001000111001001_0011100111000100"; -- 0.06947670972709741
	pesos_i(5673) := b"1111111111111111_1111111111111111_1110111101111101_0110001101110101"; -- -0.0644929733587847
	pesos_i(5674) := b"0000000000000000_0000000000000000_0001010001001110_0100011000111011"; -- 0.07931937159542518
	pesos_i(5675) := b"1111111111111111_1111111111111111_1110110000010101_1010010000110011"; -- -0.07779477828653414
	pesos_i(5676) := b"1111111111111111_1111111111111111_1110010001100000_0011000010000011"; -- -0.1079072646166664
	pesos_i(5677) := b"0000000000000000_0000000000000000_0010100010100010_0010011000101010"; -- 0.15872419868803833
	pesos_i(5678) := b"1111111111111111_1111111111111111_1111111101001001_1001110010001111"; -- -0.0027830268104963307
	pesos_i(5679) := b"0000000000000000_0000000000000000_0000001111110010_0000111010001101"; -- 0.01541224417882639
	pesos_i(5680) := b"1111111111111111_1111111111111111_1111010010010010_1111001101000001"; -- -0.04463271764192281
	pesos_i(5681) := b"1111111111111111_1111111111111111_1101011101011111_1110100001110000"; -- -0.15869281060758467
	pesos_i(5682) := b"1111111111111111_1111111111111111_1101101010010011_0011101001100001"; -- -0.1461909782374598
	pesos_i(5683) := b"1111111111111111_1111111111111111_1101001010101101_1101110010100101"; -- -0.17703457810119347
	pesos_i(5684) := b"1111111111111111_1111111111111111_1101111110011101_1000110100001000"; -- -0.12650221409129725
	pesos_i(5685) := b"0000000000000000_0000000000000000_0010010101101000_1100101000100111"; -- 0.14613021338998894
	pesos_i(5686) := b"1111111111111111_1111111111111111_1110010101101011_0100000101101101"; -- -0.1038321598183871
	pesos_i(5687) := b"0000000000000000_0000000000000000_0001010010001101_1010100100000011"; -- 0.08028656320261407
	pesos_i(5688) := b"1111111111111111_1111111111111111_1101000000010101_1100000011110100"; -- -0.18716806462474259
	pesos_i(5689) := b"1111111111111111_1111111111111111_1110011110100110_1011000110001001"; -- -0.09511270898624923
	pesos_i(5690) := b"1111111111111111_1111111111111111_1111001001111011_1101010101111000"; -- -0.052797945144056196
	pesos_i(5691) := b"0000000000000000_0000000000000000_0001111010100000_1100110001010000"; -- 0.11964108431892256
	pesos_i(5692) := b"1111111111111111_1111111111111111_1110110110000101_1110101101110000"; -- -0.07217529783908778
	pesos_i(5693) := b"0000000000000000_0000000000000000_0000110010011000_1101001011010010"; -- 0.04920690181172907
	pesos_i(5694) := b"1111111111111111_1111111111111111_1101110011001001_0010000000111010"; -- -0.1375560624510557
	pesos_i(5695) := b"0000000000000000_0000000000000000_0000010010111100_1001000001000111"; -- 0.018502252023582216
	pesos_i(5696) := b"1111111111111111_1111111111111111_1111111111000101_1000110011000101"; -- -0.0008918781206572746
	pesos_i(5697) := b"1111111111111111_1111111111111111_1101100000101011_0001011100111100"; -- -0.15559248727055588
	pesos_i(5698) := b"1111111111111111_1111111111111111_1101100111100101_1110000001010000"; -- -0.14883611715780937
	pesos_i(5699) := b"1111111111111111_1111111111111111_1101101000100110_0110010010010001"; -- -0.14785167169026484
	pesos_i(5700) := b"1111111111111111_1111111111111111_1111111011010010_0101011100011011"; -- -0.0046029622988766426
	pesos_i(5701) := b"0000000000000000_0000000000000000_0000011001000111_1011001101011011"; -- 0.024531564385372406
	pesos_i(5702) := b"0000000000000000_0000000000000000_0001110110000101_0011111110101111"; -- 0.1153144648976764
	pesos_i(5703) := b"1111111111111111_1111111111111111_1110101000010000_0111100001101110"; -- -0.08568618129621378
	pesos_i(5704) := b"1111111111111111_1111111111111111_1101100101101101_1001100001011011"; -- -0.15067146096694828
	pesos_i(5705) := b"1111111111111111_1111111111111111_1100111001100010_0010111000010111"; -- -0.19381439154316266
	pesos_i(5706) := b"0000000000000000_0000000000000000_0001010100111111_1100110101111001"; -- 0.08300480074215408
	pesos_i(5707) := b"1111111111111111_1111111111111111_1110110001011010_1010100011101001"; -- -0.07674164111363732
	pesos_i(5708) := b"1111111111111111_1111111111111111_1101010011011001_1001110100101110"; -- -0.16855447419207514
	pesos_i(5709) := b"0000000000000000_0000000000000000_0010000111101101_0111000000001011"; -- 0.13252926135834184
	pesos_i(5710) := b"0000000000000000_0000000000000000_0000011011100011_0111101101001110"; -- 0.02690859473392732
	pesos_i(5711) := b"1111111111111111_1111111111111111_1101100010100111_1110010111110110"; -- -0.15368807541275226
	pesos_i(5712) := b"0000000000000000_0000000000000000_0000001100100101_1000111101110111"; -- 0.012291876453292373
	pesos_i(5713) := b"0000000000000000_0000000000000000_0001110101000111_1101101100011110"; -- 0.11437768431989792
	pesos_i(5714) := b"0000000000000000_0000000000000000_0000001001101011_0100010110011100"; -- 0.009449339547165552
	pesos_i(5715) := b"0000000000000000_0000000000000000_0000000010010000_1011001100110101"; -- 0.002207947120777375
	pesos_i(5716) := b"0000000000000000_0000000000000000_0010100001100111_0111111101010000"; -- 0.1578292437631727
	pesos_i(5717) := b"0000000000000000_0000000000000000_0001010010001101_0000101010111111"; -- 0.08027712981089781
	pesos_i(5718) := b"0000000000000000_0000000000000000_0001011000000100_0100101100000011"; -- 0.0860030061791474
	pesos_i(5719) := b"0000000000000000_0000000000000000_0001001110011110_0010001111000010"; -- 0.07663176996906113
	pesos_i(5720) := b"0000000000000000_0000000000000000_0001011011100000_0110011111111100"; -- 0.08936166668642942
	pesos_i(5721) := b"1111111111111111_1111111111111111_1111000011101110_0100001100010101"; -- -0.0588644097696491
	pesos_i(5722) := b"1111111111111111_1111111111111111_1110000010111111_0000011111010111"; -- -0.12208510394930129
	pesos_i(5723) := b"1111111111111111_1111111111111111_1111001001011110_0001110011001011"; -- -0.05325145769742293
	pesos_i(5724) := b"0000000000000000_0000000000000000_0001110110001000_1111010100011001"; -- 0.11537105433244926
	pesos_i(5725) := b"0000000000000000_0000000000000000_0010000000000000_0010010001110001"; -- 0.1250021721497118
	pesos_i(5726) := b"1111111111111111_1111111111111111_1111101011010100_0010101110000101"; -- -0.020200042692990076
	pesos_i(5727) := b"0000000000000000_0000000000000000_0000101110110011_0110001011101011"; -- 0.045705969132037366
	pesos_i(5728) := b"1111111111111111_1111111111111111_1101111010100001_1001000000110101"; -- -0.13034723959247294
	pesos_i(5729) := b"1111111111111111_1111111111111111_1110111011001000_0010100111001000"; -- -0.06725825188735449
	pesos_i(5730) := b"1111111111111111_1111111111111111_1111000010110100_1001101010111000"; -- -0.05974419600427409
	pesos_i(5731) := b"1111111111111111_1111111111111111_1111001011100111_1101011101000100"; -- -0.051149888805451335
	pesos_i(5732) := b"0000000000000000_0000000000000000_0001011000001101_1111100000101011"; -- 0.08615065630439267
	pesos_i(5733) := b"1111111111111111_1111111111111111_1111111100101010_0001000110110101"; -- -0.003264325438064428
	pesos_i(5734) := b"1111111111111111_1111111111111111_1101110101010000_0000111101100000"; -- -0.13549713055884424
	pesos_i(5735) := b"1111111111111111_1111111111111111_1111010001001110_0011011001011000"; -- -0.04568157540880681
	pesos_i(5736) := b"0000000000000000_0000000000000000_0001101110101100_1101111110110111"; -- 0.10810659618598872
	pesos_i(5737) := b"0000000000000000_0000000000000000_0000010010100000_0000011000110000"; -- 0.01806677511271454
	pesos_i(5738) := b"1111111111111111_1111111111111111_1111000000100110_0011010010111100"; -- -0.06191702286293121
	pesos_i(5739) := b"1111111111111111_1111111111111111_1101000000011001_0101101111011011"; -- -0.18711305526131689
	pesos_i(5740) := b"0000000000000000_0000000000000000_0001110000111000_0101111101111000"; -- 0.11023518245218977
	pesos_i(5741) := b"0000000000000000_0000000000000000_0001001011111001_1101110110001010"; -- 0.07412514331857037
	pesos_i(5742) := b"1111111111111111_1111111111111111_1110111111000100_0000101010010110"; -- -0.06341489631599528
	pesos_i(5743) := b"0000000000000000_0000000000000000_0001000111011000_1100010101000101"; -- 0.06971390666724789
	pesos_i(5744) := b"0000000000000000_0000000000000000_0010011011100100_1100111011001110"; -- 0.15192883046497094
	pesos_i(5745) := b"0000000000000000_0000000000000000_0010011101100010_1110110101000101"; -- 0.1538532536740917
	pesos_i(5746) := b"1111111111111111_1111111111111111_1111010011011011_0101111010111011"; -- -0.04352767871389905
	pesos_i(5747) := b"0000000000000000_0000000000000000_0000011111100011_1001011101101011"; -- 0.03081652027601984
	pesos_i(5748) := b"1111111111111111_1111111111111111_1110111010011001_0011000001011000"; -- -0.06797502382306275
	pesos_i(5749) := b"0000000000000000_0000000000000000_0001011110101100_0001000001010000"; -- 0.09246923399819502
	pesos_i(5750) := b"1111111111111111_1111111111111111_1101000111111010_0100101111101110"; -- -0.17977452691368892
	pesos_i(5751) := b"1111111111111111_1111111111111111_1101100111010111_1111000110101110"; -- -0.14904870521289632
	pesos_i(5752) := b"0000000000000000_0000000000000000_0001010101000110_0010101111100100"; -- 0.08310198141860757
	pesos_i(5753) := b"0000000000000000_0000000000000000_0000111011000001_1010101100001101"; -- 0.05764264173664966
	pesos_i(5754) := b"1111111111111111_1111111111111111_1101001100010100_1110011111000010"; -- -0.1754622604247723
	pesos_i(5755) := b"0000000000000000_0000000000000000_0000111011110010_1001110000100000"; -- 0.05838943266758406
	pesos_i(5756) := b"1111111111111111_1111111111111111_1111011011101010_1001100100010111"; -- -0.03548281855641109
	pesos_i(5757) := b"0000000000000000_0000000000000000_0000010010001111_0100011100100100"; -- 0.017811247185143424
	pesos_i(5758) := b"0000000000000000_0000000000000000_0000110000101110_1110001100100000"; -- 0.04759044193260049
	pesos_i(5759) := b"1111111111111111_1111111111111111_1101101110000100_1100110011000110"; -- -0.14250488435703654
	pesos_i(5760) := b"0000000000000000_0000000000000000_0000011011110100_1100111010110001"; -- 0.02717296421834519
	pesos_i(5761) := b"0000000000000000_0000000000000000_0011000110101111_0111111110001010"; -- 0.1940841399010711
	pesos_i(5762) := b"0000000000000000_0000000000000000_0001011111000111_1100110111011000"; -- 0.09289251828437184
	pesos_i(5763) := b"1111111111111111_1111111111111111_1110000100100000_1101110111010110"; -- -0.12059224620902408
	pesos_i(5764) := b"1111111111111111_1111111111111111_1101000110010000_1011001101000100"; -- -0.18138579928587292
	pesos_i(5765) := b"0000000000000000_0000000000000000_0000000100111011_0100000100011110"; -- 0.004810399856233023
	pesos_i(5766) := b"0000000000000000_0000000000000000_0001101110101011_0011011011011110"; -- 0.1080812731771443
	pesos_i(5767) := b"0000000000000000_0000000000000000_0001100101001111_1110001000101000"; -- 0.09887517441233425
	pesos_i(5768) := b"0000000000000000_0000000000000000_0000111000101010_1100000101010000"; -- 0.05533989153622326
	pesos_i(5769) := b"1111111111111111_1111111111111111_1111010000010110_1111110101001010"; -- -0.04652420952353703
	pesos_i(5770) := b"1111111111111111_1111111111111111_1110011110001001_1101010111111011"; -- -0.09555304171671135
	pesos_i(5771) := b"1111111111111111_1111111111111111_1100110001001101_1001001000001001"; -- -0.20194136880956773
	pesos_i(5772) := b"0000000000000000_0000000000000000_0001000000101010_0111001100100010"; -- 0.0631477316075332
	pesos_i(5773) := b"1111111111111111_1111111111111111_1101011000010010_1000110111000101"; -- -0.1637793916802417
	pesos_i(5774) := b"1111111111111111_1111111111111111_1110101011010100_1011011010010010"; -- -0.0826917546877366
	pesos_i(5775) := b"0000000000000000_0000000000000000_0001110110010111_1110111011110110"; -- 0.11559957029925252
	pesos_i(5776) := b"0000000000000000_0000000000000000_0011001101011010_0110110011101100"; -- 0.20059853317829118
	pesos_i(5777) := b"0000000000000000_0000000000000000_0010011011111111_1010000001100011"; -- 0.15233805090819996
	pesos_i(5778) := b"1111111111111111_1111111111111111_1101111101101011_0011101011000010"; -- -0.12727005744467051
	pesos_i(5779) := b"1111111111111111_1111111111111111_1110001101101100_0010010001011101"; -- -0.11163113327157952
	pesos_i(5780) := b"0000000000000000_0000000000000000_0011001110011110_0001110111011001"; -- 0.2016314177776072
	pesos_i(5781) := b"0000000000000000_0000000000000000_0001001001111001_0011011011001100"; -- 0.07216207964608083
	pesos_i(5782) := b"1111111111111111_1111111111111111_1101001011100001_1110100101000000"; -- -0.17624036970672166
	pesos_i(5783) := b"1111111111111111_1111111111111111_1111110001100000_1100111101101101"; -- -0.014147792742664297
	pesos_i(5784) := b"1111111111111111_1111111111111111_1101011001001101_1011011001011011"; -- -0.16287670411718416
	pesos_i(5785) := b"1111111111111111_1111111111111111_1110011001010100_1011111111111100"; -- -0.10026931860929672
	pesos_i(5786) := b"0000000000000000_0000000000000000_0000100111100000_1111011110010001"; -- 0.0385889749507074
	pesos_i(5787) := b"1111111111111111_1111111111111111_1111110001010111_1001001000000000"; -- -0.01428878298538529
	pesos_i(5788) := b"0000000000000000_0000000000000000_0001010001111110_1101110111011011"; -- 0.08006083101031072
	pesos_i(5789) := b"1111111111111111_1111111111111111_1110001011000000_1101011001000111"; -- -0.11424504064171864
	pesos_i(5790) := b"1111111111111111_1111111111111111_1111100110101000_1000110100010111"; -- -0.02477186381739752
	pesos_i(5791) := b"1111111111111111_1111111111111111_1111011101111101_1111110001110101"; -- -0.03323385380457198
	pesos_i(5792) := b"0000000000000000_0000000000000000_0000001000100010_1100001001110110"; -- 0.00834288949861574
	pesos_i(5793) := b"1111111111111111_1111111111111111_1111101000101001_0001011001000000"; -- -0.022810563535113394
	pesos_i(5794) := b"1111111111111111_1111111111111111_1110000000110000_1100011110011111"; -- -0.12425567977770134
	pesos_i(5795) := b"0000000000000000_0000000000000000_0001011101100010_1010001110010001"; -- 0.09134886055660778
	pesos_i(5796) := b"1111111111111111_1111111111111111_1101000101110011_1111011011000100"; -- -0.18182428082798374
	pesos_i(5797) := b"0000000000000000_0000000000000000_0000011000001011_0010011001011101"; -- 0.023607633240445264
	pesos_i(5798) := b"1111111111111111_1111111111111111_1111011000000001_0010001101000100"; -- -0.039045139185671277
	pesos_i(5799) := b"1111111111111111_1111111111111111_1110110101011100_1011011110101110"; -- -0.07280399320250429
	pesos_i(5800) := b"1111111111111111_1111111111111111_1101001000111010_1110011001111110"; -- -0.1787887518659286
	pesos_i(5801) := b"0000000000000000_0000000000000000_0001110000000000_0101011011001100"; -- 0.10938017344851164
	pesos_i(5802) := b"0000000000000000_0000000000000000_0000000011011111_1110110110011000"; -- 0.0034168716217224566
	pesos_i(5803) := b"1111111111111111_1111111111111111_1111010011001000_1001010111100000"; -- -0.04381430897502863
	pesos_i(5804) := b"0000000000000000_0000000000000000_0000000001010110_1111101001111111"; -- 0.0013271866252436027
	pesos_i(5805) := b"1111111111111111_1111111111111111_1110111001011101_0011011011010010"; -- -0.06889016498267338
	pesos_i(5806) := b"1111111111111111_1111111111111111_1111000100001011_1101110110110010"; -- -0.058412689334014764
	pesos_i(5807) := b"0000000000000000_0000000000000000_0000101111101111_1101000110010001"; -- 0.046628091677431864
	pesos_i(5808) := b"0000000000000000_0000000000000000_0001111110110110_0001010101010001"; -- 0.12387212023153293
	pesos_i(5809) := b"1111111111111111_1111111111111111_1101110100010101_0110110110110001"; -- -0.136391777210815
	pesos_i(5810) := b"1111111111111111_1111111111111111_1101110001011011_0101101100001111"; -- -0.13923102274209317
	pesos_i(5811) := b"0000000000000000_0000000000000000_0000000000111000_1100010110111100"; -- 0.0008662781242243789
	pesos_i(5812) := b"1111111111111111_1111111111111111_1111101011010101_0011001101111110"; -- -0.02018430869339864
	pesos_i(5813) := b"1111111111111111_1111111111111111_1110000101000111_1010011101101010"; -- -0.12000039731750012
	pesos_i(5814) := b"0000000000000000_0000000000000000_0000000101100110_0010001010101111"; -- 0.005464713735707458
	pesos_i(5815) := b"0000000000000000_0000000000000000_0001111110000011_1010001111001010"; -- 0.12310241386831443
	pesos_i(5816) := b"1111111111111111_1111111111111111_1101011000101110_0001001010100100"; -- -0.16335948459248797
	pesos_i(5817) := b"0000000000000000_0000000000000000_0001000000100010_0101000000000101"; -- 0.06302356837630632
	pesos_i(5818) := b"1111111111111111_1111111111111111_1100110101110111_1100000101111010"; -- -0.19739142193752
	pesos_i(5819) := b"1111111111111111_1111111111111111_1110101001001110_0101010001111101"; -- -0.08474227858014735
	pesos_i(5820) := b"0000000000000000_0000000000000000_0000100001110011_0101111001001011"; -- 0.0330103810327315
	pesos_i(5821) := b"1111111111111111_1111111111111111_1110001100101111_0111001001000100"; -- -0.11255727621974664
	pesos_i(5822) := b"1111111111111111_1111111111111111_1111000111011000_0010001111010111"; -- -0.055295715429553915
	pesos_i(5823) := b"0000000000000000_0000000000000000_0010110000100100_1010010011101011"; -- 0.17243414617378597
	pesos_i(5824) := b"1111111111111111_1111111111111111_1101000011010110_1001001110011110"; -- -0.1842258205412826
	pesos_i(5825) := b"0000000000000000_0000000000000000_0010010101000110_1111101010000000"; -- 0.1456142963065737
	pesos_i(5826) := b"1111111111111111_1111111111111111_1110010000100111_1111100000010010"; -- -0.108765121045485
	pesos_i(5827) := b"0000000000000000_0000000000000000_0010001000110111_1001100011000110"; -- 0.1336608394660271
	pesos_i(5828) := b"1111111111111111_1111111111111111_1101111110100010_0100110010101011"; -- -0.12642975633873757
	pesos_i(5829) := b"0000000000000000_0000000000000000_0000110000010010_0011110010000111"; -- 0.04715326581987661
	pesos_i(5830) := b"1111111111111111_1111111111111111_1111000100011101_0000011101101011"; -- -0.0581508029850145
	pesos_i(5831) := b"1111111111111111_1111111111111111_1111011111110001_0100100101001010"; -- -0.031474513397282904
	pesos_i(5832) := b"0000000000000000_0000000000000000_0001111011101110_1110000010100001"; -- 0.12083248066671036
	pesos_i(5833) := b"0000000000000000_0000000000000000_0000100110110101_0101110011011001"; -- 0.037923624999069296
	pesos_i(5834) := b"1111111111111111_1111111111111111_1110101110111011_0100101000000001"; -- -0.0791734454173612
	pesos_i(5835) := b"1111111111111111_1111111111111111_1110101001011001_1111100111010100"; -- -0.08456457680034851
	pesos_i(5836) := b"0000000000000000_0000000000000000_0010111010101001_1000101010111100"; -- 0.1822745045840183
	pesos_i(5837) := b"0000000000000000_0000000000000000_0010001111001111_0000100100111001"; -- 0.13987786908201652
	pesos_i(5838) := b"0000000000000000_0000000000000000_0001010100111100_0010011111011110"; -- 0.08294915355587877
	pesos_i(5839) := b"1111111111111111_1111111111111111_1111100010010000_0100110001000110"; -- -0.02904818821219301
	pesos_i(5840) := b"1111111111111111_1111111111111111_1101111101100011_0001110111001001"; -- -0.12739385445790094
	pesos_i(5841) := b"1111111111111111_1111111111111111_1111010001110001_0110101010011111"; -- -0.04514440162309903
	pesos_i(5842) := b"1111111111111111_1111111111111111_1110000100110000_0011100011101110"; -- -0.12035793490190762
	pesos_i(5843) := b"0000000000000000_0000000000000000_0000110000001001_0110110110110000"; -- 0.04701886689122583
	pesos_i(5844) := b"0000000000000000_0000000000000000_0001000000010000_1001100001000000"; -- 0.06275321536463646
	pesos_i(5845) := b"0000000000000000_0000000000000000_0000000001111010_1011011100100011"; -- 0.0018724879877251252
	pesos_i(5846) := b"1111111111111111_1111111111111111_1111111100100100_0001000100010111"; -- -0.003355914934828489
	pesos_i(5847) := b"1111111111111111_1111111111111111_1111111111101111_0001101101101100"; -- -0.0002577649147595953
	pesos_i(5848) := b"0000000000000000_0000000000000000_0001111000100001_0010011110101010"; -- 0.11769340415790523
	pesos_i(5849) := b"1111111111111111_1111111111111111_1111110011010101_0001110100000101"; -- -0.01237314817260875
	pesos_i(5850) := b"1111111111111111_1111111111111111_1110100010000111_1011000101000101"; -- -0.09167949744541186
	pesos_i(5851) := b"1111111111111111_1111111111111111_1110010000110011_0001011001111001"; -- -0.10859546239097335
	pesos_i(5852) := b"0000000000000000_0000000000000000_0010101101111001_1111100101110101"; -- 0.1698299323555368
	pesos_i(5853) := b"0000000000000000_0000000000000000_0000011011001110_1100001010000100"; -- 0.026592404541997607
	pesos_i(5854) := b"0000000000000000_0000000000000000_0000010100101100_1010011001010011"; -- 0.020212550468775056
	pesos_i(5855) := b"1111111111111111_1111111111111111_1101000000100001_0000001001110110"; -- -0.18699631322016136
	pesos_i(5856) := b"1111111111111111_1111111111111111_1101010101011000_0001101000111011"; -- -0.1666244130644833
	pesos_i(5857) := b"0000000000000000_0000000000000000_0000111010000011_0010011000010010"; -- 0.05668867046469812
	pesos_i(5858) := b"0000000000000000_0000000000000000_0000100110010010_0101100001111000"; -- 0.037389306407636325
	pesos_i(5859) := b"0000000000000000_0000000000000000_0001011110101010_0111111000101100"; -- 0.092445264575159
	pesos_i(5860) := b"1111111111111111_1111111111111111_1111101111001001_1110111111111101"; -- -0.016449929086980456
	pesos_i(5861) := b"1111111111111111_1111111111111111_1101111100100100_0000101000110110"; -- -0.1283563249409474
	pesos_i(5862) := b"0000000000000000_0000000000000000_0010111000001100_1000100100011000"; -- 0.17987877698823077
	pesos_i(5863) := b"1111111111111111_1111111111111111_1110011111010110_1100100000001100"; -- -0.09437894542882379
	pesos_i(5864) := b"0000000000000000_0000000000000000_0000011101010110_1010001001000011"; -- 0.028665677353904902
	pesos_i(5865) := b"0000000000000000_0000000000000000_0001010110011110_0000001110011111"; -- 0.08444235452218893
	pesos_i(5866) := b"1111111111111111_1111111111111111_1110110110101101_0000000111111010"; -- -0.07157886158617448
	pesos_i(5867) := b"1111111111111111_1111111111111111_1110111111110100_1110101001101101"; -- -0.06266913257590274
	pesos_i(5868) := b"1111111111111111_1111111111111111_1101100011111010_1000101100010111"; -- -0.15242701232683464
	pesos_i(5869) := b"1111111111111111_1111111111111111_1101100001010010_0000001011000001"; -- -0.15499861514138885
	pesos_i(5870) := b"0000000000000000_0000000000000000_0000110101110100_1010101101110100"; -- 0.05256148897846598
	pesos_i(5871) := b"0000000000000000_0000000000000000_0000010110100110_1101100111011101"; -- 0.022077194640721824
	pesos_i(5872) := b"1111111111111111_1111111111111111_1110001110001111_1111001111110100"; -- -0.11108470241294223
	pesos_i(5873) := b"1111111111111111_1111111111111111_1101100011111011_0101000111001000"; -- -0.15241516942387923
	pesos_i(5874) := b"1111111111111111_1111111111111111_1110011110001000_1110101100101111"; -- -0.0955670365977179
	pesos_i(5875) := b"1111111111111111_1111111111111111_1110111101000010_1100000111110011"; -- -0.06538760972595513
	pesos_i(5876) := b"1111111111111111_1111111111111111_1111111100111000_0111101110000110"; -- -0.0030443952992292287
	pesos_i(5877) := b"1111111111111111_1111111111111111_1110000101010010_1100100000001000"; -- -0.11983060658150164
	pesos_i(5878) := b"0000000000000000_0000000000000000_0000100110010010_1110001011111111"; -- 0.0373975631492221
	pesos_i(5879) := b"1111111111111111_1111111111111111_1110011111111011_1001100101101100"; -- -0.09381714933544151
	pesos_i(5880) := b"1111111111111111_1111111111111111_1111001001001101_1110100011111110"; -- -0.053498685877163374
	pesos_i(5881) := b"0000000000000000_0000000000000000_0001101101000101_0110111111000000"; -- 0.10652826720991487
	pesos_i(5882) := b"0000000000000000_0000000000000000_0001110101010010_0101000111000111"; -- 0.11453734510104448
	pesos_i(5883) := b"1111111111111111_1111111111111111_1110110111011101_0100111011000010"; -- -0.07084186318740526
	pesos_i(5884) := b"1111111111111111_1111111111111111_1110100000010001_1100100111011011"; -- -0.09347856901429363
	pesos_i(5885) := b"1111111111111111_1111111111111111_1101001000000011_1110001010011011"; -- -0.1796282169337559
	pesos_i(5886) := b"0000000000000000_0000000000000000_0001110111100001_1111110010110000"; -- 0.11672953892374931
	pesos_i(5887) := b"1111111111111111_1111111111111111_1101011101111010_1010011100101000"; -- -0.15828471447121448
	pesos_i(5888) := b"0000000000000000_0000000000000000_0010100001110010_1101011111010111"; -- 0.15800236703830348
	pesos_i(5889) := b"1111111111111111_1111111111111111_1111000111010111_0100001110111101"; -- -0.055309072842475215
	pesos_i(5890) := b"1111111111111111_1111111111111111_1101011110010110_1001111011001000"; -- -0.15785796752309425
	pesos_i(5891) := b"0000000000000000_0000000000000000_0001010111010000_1100001100011000"; -- 0.08521670668897195
	pesos_i(5892) := b"0000000000000000_0000000000000000_0010010001100111_1110100100100101"; -- 0.1422105518805731
	pesos_i(5893) := b"0000000000000000_0000000000000000_0000101011110110_0110101011011011"; -- 0.0428225311951072
	pesos_i(5894) := b"1111111111111111_1111111111111111_1101000011100100_0010101010110010"; -- -0.18401845117276588
	pesos_i(5895) := b"1111111111111111_1111111111111111_1110011110011100_0101101100110011"; -- -0.0952704430158381
	pesos_i(5896) := b"1111111111111111_1111111111111111_1111100001111010_1000001011001101"; -- -0.029380631482015612
	pesos_i(5897) := b"0000000000000000_0000000000000000_0010110100110100_1101001110001111"; -- 0.17658731695169183
	pesos_i(5898) := b"1111111111111111_1111111111111111_1111011100000110_0111010111001000"; -- -0.0350576769803682
	pesos_i(5899) := b"0000000000000000_0000000000000000_0000101010111110_1111111100110000"; -- 0.04197688021231039
	pesos_i(5900) := b"0000000000000000_0000000000000000_0010010000101010_1001111110110101"; -- 0.14127538834439712
	pesos_i(5901) := b"1111111111111111_1111111111111111_1101100010011010_0110000101001000"; -- -0.15389434798683746
	pesos_i(5902) := b"1111111111111111_1111111111111111_1100101100100010_0110101011010111"; -- -0.2065060829743712
	pesos_i(5903) := b"0000000000000000_0000000000000000_0000100001110010_1100010010100101"; -- 0.03300122287697197
	pesos_i(5904) := b"0000000000000000_0000000000000000_0010010101111011_1011110000011100"; -- 0.14641929313609037
	pesos_i(5905) := b"0000000000000000_0000000000000000_0010100101010100_0111000001010111"; -- 0.16144468416545293
	pesos_i(5906) := b"1111111111111111_1111111111111111_1101111000001000_1011001111011000"; -- -0.13267971015409777
	pesos_i(5907) := b"0000000000000000_0000000000000000_0000110001110111_1101000001100110"; -- 0.048703217339561886
	pesos_i(5908) := b"0000000000000000_0000000000000000_0001000011010111_0011000001001111"; -- 0.06578351907922349
	pesos_i(5909) := b"0000000000000000_0000000000000000_0010100100001010_1101000100111010"; -- 0.16032130873691447
	pesos_i(5910) := b"0000000000000000_0000000000000000_0001111100000001_1110101110111010"; -- 0.12112305924722272
	pesos_i(5911) := b"1111111111111111_1111111111111111_1110110101001010_0000010111011000"; -- -0.0730892513288046
	pesos_i(5912) := b"1111111111111111_1111111111111111_1111000011001101_1101001100011111"; -- -0.05935936445689186
	pesos_i(5913) := b"1111111111111111_1111111111111111_1101110001100101_1001111011100010"; -- -0.13907439214345169
	pesos_i(5914) := b"1111111111111111_1111111111111111_1101011111001101_0110010011101001"; -- -0.15702218344326926
	pesos_i(5915) := b"1111111111111111_1111111111111111_1101000110011000_1011100000010010"; -- -0.18126344269471328
	pesos_i(5916) := b"0000000000000000_0000000000000000_0010111111011110_0010101110001111"; -- 0.1869837974873867
	pesos_i(5917) := b"1111111111111111_1111111111111111_1111110110001010_1111101010111000"; -- -0.00959809307458089
	pesos_i(5918) := b"1111111111111111_1111111111111111_1101110001011000_0101000010100101"; -- -0.13927741985728126
	pesos_i(5919) := b"1111111111111111_1111111111111111_1101001111100000_0101100101001011"; -- -0.17235795901326212
	pesos_i(5920) := b"1111111111111111_1111111111111111_1110001100000100_0001110001001011"; -- -0.1132185284563126
	pesos_i(5921) := b"0000000000000000_0000000000000000_0001010010011110_1001001001010101"; -- 0.08054461077306882
	pesos_i(5922) := b"1111111111111111_1111111111111111_1110000110101110_1011111110000100"; -- -0.1184273054138783
	pesos_i(5923) := b"0000000000000000_0000000000000000_0000110000001001_0010000110100010"; -- 0.047014333752406774
	pesos_i(5924) := b"1111111111111111_1111111111111111_1110110110100101_0001000011001100"; -- -0.07170004866654478
	pesos_i(5925) := b"0000000000000000_0000000000000000_0000110110000111_0001100100101100"; -- 0.052842686803380515
	pesos_i(5926) := b"0000000000000000_0000000000000000_0001010101111101_1001100101011000"; -- 0.08394773866509925
	pesos_i(5927) := b"1111111111111111_1111111111111111_1110100011001000_0110010010000001"; -- -0.09069225165864052
	pesos_i(5928) := b"0000000000000000_0000000000000000_0001100001001000_0010110001000001"; -- 0.09485127058771453
	pesos_i(5929) := b"0000000000000000_0000000000000000_0000111100100100_0011111101010011"; -- 0.059146840779681645
	pesos_i(5930) := b"0000000000000000_0000000000000000_0010001001111111_1010011110001001"; -- 0.13476035211262302
	pesos_i(5931) := b"0000000000000000_0000000000000000_0001100111001010_1111000111110110"; -- 0.10075294727309059
	pesos_i(5932) := b"1111111111111111_1111111111111111_1101100110001100_0010010101011110"; -- -0.15020529226449825
	pesos_i(5933) := b"1111111111111111_1111111111111111_1101101111000000_0000001111001100"; -- -0.14160133618041193
	pesos_i(5934) := b"0000000000000000_0000000000000000_0000110001010100_0010101001000101"; -- 0.04815925785154703
	pesos_i(5935) := b"1111111111111111_1111111111111111_1110010100101000_1001011111101110"; -- -0.10484934272237373
	pesos_i(5936) := b"0000000000000000_0000000000000000_0000100100000001_1011111011101100"; -- 0.03518288870746378
	pesos_i(5937) := b"1111111111111111_1111111111111111_1110110110010100_1111100111010011"; -- -0.07194555850274775
	pesos_i(5938) := b"1111111111111111_1111111111111111_1101111011100111_0111011010110100"; -- -0.1292806443998047
	pesos_i(5939) := b"0000000000000000_0000000000000000_0000000001000100_0011100001000101"; -- 0.0010409516062548007
	pesos_i(5940) := b"0000000000000000_0000000000000000_0011000011110111_0100011011010101"; -- 0.19127314286130198
	pesos_i(5941) := b"0000000000000000_0000000000000000_0010110001101100_0001111010000011"; -- 0.17352476783371729
	pesos_i(5942) := b"1111111111111111_1111111111111111_1111000001101100_1111101001110100"; -- -0.06083712253545995
	pesos_i(5943) := b"1111111111111111_1111111111111111_1111101001000000_0001001011110001"; -- -0.02245980857901499
	pesos_i(5944) := b"0000000000000000_0000000000000000_0000010110011100_1101110111010011"; -- 0.021924842866705208
	pesos_i(5945) := b"0000000000000000_0000000000000000_0001010101001011_0111100001000010"; -- 0.08318282714932684
	pesos_i(5946) := b"1111111111111111_1111111111111111_1110011101110100_1010111001110101"; -- -0.09587583211136232
	pesos_i(5947) := b"1111111111111111_1111111111111111_1101001000100011_1000110010001110"; -- -0.1791450645848313
	pesos_i(5948) := b"0000000000000000_0000000000000000_0010010010010110_0010100101011010"; -- 0.1429162831233695
	pesos_i(5949) := b"0000000000000000_0000000000000000_0000110100101010_1110011111011100"; -- 0.05143593910534945
	pesos_i(5950) := b"0000000000000000_0000000000000000_0000001001010000_0011100001000011"; -- 0.009036556619124916
	pesos_i(5951) := b"1111111111111111_1111111111111111_1101000101001000_1001110100100111"; -- -0.18248575011834473
	pesos_i(5952) := b"0000000000000000_0000000000000000_0010001100001111_1010011100111101"; -- 0.13695759993173848
	pesos_i(5953) := b"1111111111111111_1111111111111111_1101000111100101_1100101001000111"; -- -0.18008743075151018
	pesos_i(5954) := b"0000000000000000_0000000000000000_0001100110110111_0110101110110101"; -- 0.10045502820525169
	pesos_i(5955) := b"1111111111111111_1111111111111111_1100110011000101_0100101001001110"; -- -0.20011458974066715
	pesos_i(5956) := b"0000000000000000_0000000000000000_0000000011010001_1000111111010000"; -- 0.0031976589215393135
	pesos_i(5957) := b"1111111111111111_1111111111111111_1101101111110101_1000000110111101"; -- -0.14078511375897568
	pesos_i(5958) := b"0000000000000000_0000000000000000_0010110000101101_0101011010110100"; -- 0.17256681352199557
	pesos_i(5959) := b"1111111111111111_1111111111111111_1111101111101011_0001010101010001"; -- -0.015944163911648813
	pesos_i(5960) := b"1111111111111111_1111111111111111_1111011110011100_0100000111101010"; -- -0.03277195017136506
	pesos_i(5961) := b"0000000000000000_0000000000000000_0001110000011001_0110101110011001"; -- 0.1097628829709602
	pesos_i(5962) := b"1111111111111111_1111111111111111_1101100111000000_0001101010100000"; -- -0.14941247549051279
	pesos_i(5963) := b"0000000000000000_0000000000000000_0001100001100101_0110101011100111"; -- 0.09529750945606906
	pesos_i(5964) := b"0000000000000000_0000000000000000_0000000111100010_0111001101001001"; -- 0.007361607788515202
	pesos_i(5965) := b"1111111111111111_1111111111111111_1111011110110011_0011010010001000"; -- -0.03242179571256137
	pesos_i(5966) := b"0000000000000000_0000000000000000_0000000100001100_0000010101011000"; -- 0.004089673942622322
	pesos_i(5967) := b"1111111111111111_1111111111111111_1110111111011000_0000001000101010"; -- -0.06311022252896044
	pesos_i(5968) := b"0000000000000000_0000000000000000_0010000010001111_0110110011001001"; -- 0.1271884909518952
	pesos_i(5969) := b"1111111111111111_1111111111111111_1101110111011011_0010011110010001"; -- -0.13337471681113125
	pesos_i(5970) := b"1111111111111111_1111111111111111_1110100001001100_0100010111110011"; -- -0.09258616270423241
	pesos_i(5971) := b"0000000000000000_0000000000000000_0001010110101011_0010110110000011"; -- 0.08464321572244712
	pesos_i(5972) := b"0000000000000000_0000000000000000_0001010110100011_1000101111101000"; -- 0.08452677174439498
	pesos_i(5973) := b"0000000000000000_0000000000000000_0010000111001100_0000101010101011"; -- 0.13201967885706492
	pesos_i(5974) := b"1111111111111111_1111111111111111_1101010110000101_1011110101001111"; -- -0.1659280474146689
	pesos_i(5975) := b"0000000000000000_0000000000000000_0001110101011110_1101010100110110"; -- 0.11472828442012455
	pesos_i(5976) := b"0000000000000000_0000000000000000_0000000110110001_0010000011010001"; -- 0.006609011634988865
	pesos_i(5977) := b"0000000000000000_0000000000000000_0001001110101101_0001011100001111"; -- 0.0768598949551222
	pesos_i(5978) := b"1111111111111111_1111111111111111_1110110011111111_0110100110000001"; -- -0.0742277203278744
	pesos_i(5979) := b"0000000000000000_0000000000000000_0001010101111000_1111110110111110"; -- 0.08387742897553756
	pesos_i(5980) := b"1111111111111111_1111111111111111_1101011111100110_1100001010101110"; -- -0.15663512475144928
	pesos_i(5981) := b"0000000000000000_0000000000000000_0000000011011101_0111111111101101"; -- 0.0033798174543899612
	pesos_i(5982) := b"0000000000000000_0000000000000000_0001010110000000_0001110010001001"; -- 0.08398607585670989
	pesos_i(5983) := b"1111111111111111_1111111111111111_1101001110101110_0111011011101100"; -- -0.17311913230980897
	pesos_i(5984) := b"1111111111111111_1111111111111111_1110001001011110_0111101111101110"; -- -0.11574578713878705
	pesos_i(5985) := b"1111111111111111_1111111111111111_1111010000010010_0000011010011000"; -- -0.04659994884125855
	pesos_i(5986) := b"0000000000000000_0000000000000000_0000111000010110_0100000101100000"; -- 0.055027090030808766
	pesos_i(5987) := b"0000000000000000_0000000000000000_0000101100001001_0100110100110010"; -- 0.04311068032446958
	pesos_i(5988) := b"0000000000000000_0000000000000000_0001000111110011_1101111100000001"; -- 0.07012742773766269
	pesos_i(5989) := b"1111111111111111_1111111111111111_1111010101000000_0110010010001110"; -- -0.0419861938952106
	pesos_i(5990) := b"0000000000000000_0000000000000000_0000011001001000_0000001100111001"; -- 0.02453632493828234
	pesos_i(5991) := b"0000000000000000_0000000000000000_0001100111110010_1001111110101011"; -- 0.10135839394878322
	pesos_i(5992) := b"1111111111111111_1111111111111111_1101111111001011_1000110101001100"; -- -0.125800293823687
	pesos_i(5993) := b"1111111111111111_1111111111111111_1110100110001011_0101011011101110"; -- -0.0877175969158551
	pesos_i(5994) := b"0000000000000000_0000000000000000_0000010011000000_1001000011011101"; -- 0.018563322056565745
	pesos_i(5995) := b"0000000000000000_0000000000000000_0001101100010100_1101111011110011"; -- 0.10578721454425845
	pesos_i(5996) := b"0000000000000000_0000000000000000_0000010001000101_1001001110101011"; -- 0.016686658257503345
	pesos_i(5997) := b"1111111111111111_1111111111111111_1101110011111101_1010011000010111"; -- -0.13675462656817727
	pesos_i(5998) := b"0000000000000000_0000000000000000_0010000110000010_0100100011100110"; -- 0.13089423769474812
	pesos_i(5999) := b"1111111111111111_1111111111111111_1101100100111001_1111100001100001"; -- -0.15145919437181646
	pesos_i(6000) := b"0000000000000000_0000000000000000_0001111010001110_0001110000111011"; -- 0.11935593063955179
	pesos_i(6001) := b"1111111111111111_1111111111111111_1101100110111101_0000011010101101"; -- -0.1494594410340987
	pesos_i(6002) := b"0000000000000000_0000000000000000_0000110000101010_1111010110001101"; -- 0.04753050504739823
	pesos_i(6003) := b"1111111111111111_1111111111111111_1111101100101000_1110011000000000"; -- -0.018907189364282675
	pesos_i(6004) := b"0000000000000000_0000000000000000_0010001100100010_1010001010011111"; -- 0.1372472417858722
	pesos_i(6005) := b"0000000000000000_0000000000000000_0001001000011000_0100011000001101"; -- 0.07068288627039537
	pesos_i(6006) := b"1111111111111111_1111111111111111_1100110111110000_0001001000111000"; -- -0.19555555475134564
	pesos_i(6007) := b"1111111111111111_1111111111111111_1101101101000001_1011101111101010"; -- -0.1435282280978695
	pesos_i(6008) := b"1111111111111111_1111111111111111_1111110101101011_0101111011111100"; -- -0.010080398070332668
	pesos_i(6009) := b"1111111111111111_1111111111111111_1110011010101100_1111100000001110"; -- -0.09892320303673782
	pesos_i(6010) := b"1111111111111111_1111111111111111_1110100101000111_1011011100100000"; -- -0.08874946083773437
	pesos_i(6011) := b"1111111111111111_1111111111111111_1101101011111100_0100000110111110"; -- -0.14458836650723858
	pesos_i(6012) := b"1111111111111111_1111111111111111_1101001101010001_0000100101001001"; -- -0.17454473459751194
	pesos_i(6013) := b"1111111111111111_1111111111111111_1110100111010101_0111110100001100"; -- -0.08658617458421607
	pesos_i(6014) := b"1111111111111111_1111111111111111_1110110001111000_0101100000100001"; -- -0.07628869235027352
	pesos_i(6015) := b"1111111111111111_1111111111111111_1111011111000101_0001000100001100"; -- -0.03214925238959723
	pesos_i(6016) := b"1111111111111111_1111111111111111_1111111100000100_1010001101111100"; -- -0.003835470393709102
	pesos_i(6017) := b"0000000000000000_0000000000000000_0000110111001000_1000101011010100"; -- 0.053841282621416395
	pesos_i(6018) := b"0000000000000000_0000000000000000_0000010011010111_0001101001011011"; -- 0.018907210509538367
	pesos_i(6019) := b"1111111111111111_1111111111111111_1101110001001101_1111011101001000"; -- -0.13943533403763955
	pesos_i(6020) := b"1111111111111111_1111111111111111_1111011110100001_1010101010000101"; -- -0.03268942119694954
	pesos_i(6021) := b"1111111111111111_1111111111111111_1101000000111111_1010000011111001"; -- -0.18652910156963942
	pesos_i(6022) := b"0000000000000000_0000000000000000_0010011100001111_0000001011111000"; -- 0.1525728087467222
	pesos_i(6023) := b"1111111111111111_1111111111111111_1101111000100011_0001111110001100"; -- -0.1322765620635733
	pesos_i(6024) := b"0000000000000000_0000000000000000_0001011011101111_1111001100110000"; -- 0.08959884563797187
	pesos_i(6025) := b"1111111111111111_1111111111111111_1110101000100110_1001101000110011"; -- -0.08534847513713748
	pesos_i(6026) := b"0000000000000000_0000000000000000_0010101010100111_0010111110101001"; -- 0.16661355843960135
	pesos_i(6027) := b"1111111111111111_1111111111111111_1110110101000011_0110100011101100"; -- -0.07319015730320443
	pesos_i(6028) := b"1111111111111111_1111111111111111_1110010111100010_1111010010100100"; -- -0.10200568191391583
	pesos_i(6029) := b"1111111111111111_1111111111111111_1101110010110000_1110010001100001"; -- -0.13792584076595468
	pesos_i(6030) := b"1111111111111111_1111111111111111_1111010101111101_1010101011100111"; -- -0.04105121476014837
	pesos_i(6031) := b"1111111111111111_1111111111111111_1110000100111110_1100011101110000"; -- -0.12013581775847422
	pesos_i(6032) := b"0000000000000000_0000000000000000_0001110011111010_1111110011111111"; -- 0.11320477706794937
	pesos_i(6033) := b"1111111111111111_1111111111111111_1111001010110111_1101001000000111"; -- -0.0518826231099035
	pesos_i(6034) := b"0000000000000000_0000000000000000_0010001000100000_1100010010001001"; -- 0.1333124956153297
	pesos_i(6035) := b"1111111111111111_1111111111111111_1101111110111001_1110001100010110"; -- -0.12606983865523683
	pesos_i(6036) := b"0000000000000000_0000000000000000_0001100101000001_0111000000001111"; -- 0.09865475044186263
	pesos_i(6037) := b"0000000000000000_0000000000000000_0010000100101000_0101010011010111"; -- 0.1295216584693
	pesos_i(6038) := b"1111111111111111_1111111111111111_1111001001101110_1001100111001000"; -- -0.05299986703842231
	pesos_i(6039) := b"1111111111111111_1111111111111111_1110001111110011_1100110000111000"; -- -0.1095611918955443
	pesos_i(6040) := b"1111111111111111_1111111111111111_1111100011101001_1011111001000111"; -- -0.027683360802954218
	pesos_i(6041) := b"1111111111111111_1111111111111111_1111001000110000_1101010100011010"; -- -0.053942376291629776
	pesos_i(6042) := b"1111111111111111_1111111111111111_1110000111000000_0000111111011011"; -- -0.11816311754849239
	pesos_i(6043) := b"1111111111111111_1111111111111111_1111111010001100_0110110011001011"; -- -0.005669784912776739
	pesos_i(6044) := b"0000000000000000_0000000000000000_0000101111101011_0000010001111010"; -- 0.04655483231583382
	pesos_i(6045) := b"0000000000000000_0000000000000000_0010010010000100_0011111101110110"; -- 0.14264294264029004
	pesos_i(6046) := b"0000000000000000_0000000000000000_0010111000001000_0100111011010110"; -- 0.17981426925820362
	pesos_i(6047) := b"0000000000000000_0000000000000000_0010000100001101_0111000000011110"; -- 0.1291112968810971
	pesos_i(6048) := b"1111111111111111_1111111111111111_1110011111011011_1100101110110001"; -- -0.09430243423931405
	pesos_i(6049) := b"1111111111111111_1111111111111111_1110110101001110_0111111100000000"; -- -0.07302099455419309
	pesos_i(6050) := b"0000000000000000_0000000000000000_0001001010111010_1100000111010010"; -- 0.07316218731667397
	pesos_i(6051) := b"1111111111111111_1111111111111111_1111100000110011_1101101010011010"; -- -0.030458772193928927
	pesos_i(6052) := b"0000000000000000_0000000000000000_0000011110001011_0001000110110101"; -- 0.029465777159341525
	pesos_i(6053) := b"1111111111111111_1111111111111111_1110101011110011_1110101000111011"; -- -0.08221565308848665
	pesos_i(6054) := b"1111111111111111_1111111111111111_1101010001011001_1010010110000111"; -- -0.17050710156020657
	pesos_i(6055) := b"0000000000000000_0000000000000000_0010010011110100_1010100110001000"; -- 0.14435824926836233
	pesos_i(6056) := b"0000000000000000_0000000000000000_0000000010111100_0000001100001111"; -- 0.002868834753796127
	pesos_i(6057) := b"0000000000000000_0000000000000000_0010011100100001_0101101010101000"; -- 0.15285269357822379
	pesos_i(6058) := b"1111111111111111_1111111111111111_1110111101101001_0010100000010011"; -- -0.06480168864019803
	pesos_i(6059) := b"1111111111111111_1111111111111111_1101110110111110_0000001111001100"; -- -0.13381935381444995
	pesos_i(6060) := b"0000000000000000_0000000000000000_0001111101100000_0110111011000011"; -- 0.12256519556584776
	pesos_i(6061) := b"0000000000000000_0000000000000000_0001010000001001_0111111101011101"; -- 0.0782699206336588
	pesos_i(6062) := b"0000000000000000_0000000000000000_0000010010001010_1111010001000001"; -- 0.01774527164841124
	pesos_i(6063) := b"1111111111111111_1111111111111111_1111011101010111_0110100001001101"; -- -0.03382251862741207
	pesos_i(6064) := b"0000000000000000_0000000000000000_0001011001110010_0011010000110001"; -- 0.08768011289892304
	pesos_i(6065) := b"0000000000000000_0000000000000000_0001010110110101_1100001001001101"; -- 0.08480467208171602
	pesos_i(6066) := b"0000000000000000_0000000000000000_0010000100110001_0000110100000111"; -- 0.12965470703813595
	pesos_i(6067) := b"0000000000000000_0000000000000000_0010001011111010_0111001110000101"; -- 0.13663408268894484
	pesos_i(6068) := b"1111111111111111_1111111111111111_1111011100001000_1111101011110000"; -- -0.035019222596113835
	pesos_i(6069) := b"0000000000000000_0000000000000000_0000010011010101_0100111101111011"; -- 0.01887985941807346
	pesos_i(6070) := b"1111111111111111_1111111111111111_1110011110000111_0100100100010010"; -- -0.09559195810279869
	pesos_i(6071) := b"0000000000000000_0000000000000000_0001100100010111_0010001010110100"; -- 0.09800927053207072
	pesos_i(6072) := b"0000000000000000_0000000000000000_0001010011001111_0011000000110111"; -- 0.08128644326554979
	pesos_i(6073) := b"0000000000000000_0000000000000000_0000110001001111_1011111110101110"; -- 0.04809186933981024
	pesos_i(6074) := b"1111111111111111_1111111111111111_1111000100110111_0010010001000000"; -- -0.0577523558199781
	pesos_i(6075) := b"1111111111111111_1111111111111111_1111011001000110_1011111011000111"; -- -0.03798301345742545
	pesos_i(6076) := b"0000000000000000_0000000000000000_0000111100010000_0111101100000011"; -- 0.058845222764863106
	pesos_i(6077) := b"1111111111111111_1111111111111111_1101111110011111_1101110100010001"; -- -0.1264669259647906
	pesos_i(6078) := b"0000000000000000_0000000000000000_0010001011101001_1100000100100111"; -- 0.13637931058014569
	pesos_i(6079) := b"0000000000000000_0000000000000000_0010001110101101_0111110100001000"; -- 0.13936597304255216
	pesos_i(6080) := b"1111111111111111_1111111111111111_1111101110011001_1010111111111000"; -- -0.01718616677703694
	pesos_i(6081) := b"1111111111111111_1111111111111111_1110101010110010_1011111000000011"; -- -0.08321011000902645
	pesos_i(6082) := b"1111111111111111_1111111111111111_1110101110111100_1111000001011111"; -- -0.0791482703989584
	pesos_i(6083) := b"1111111111111111_1111111111111111_1110001100010000_1010011100100011"; -- -0.11302714735538047
	pesos_i(6084) := b"0000000000000000_0000000000000000_0001010111001001_0101111001101011"; -- 0.08510389431105092
	pesos_i(6085) := b"1111111111111111_1111111111111111_1111001110001110_0011111111101110"; -- -0.04861069136541067
	pesos_i(6086) := b"0000000000000000_0000000000000000_0001111011100101_1000100100010100"; -- 0.1206899331087987
	pesos_i(6087) := b"0000000000000000_0000000000000000_0000111010101110_1010100001100110"; -- 0.05735256656974273
	pesos_i(6088) := b"0000000000000000_0000000000000000_0001100100111000_0110101010101000"; -- 0.09851709928173265
	pesos_i(6089) := b"0000000000000000_0000000000000000_0001010110111101_1110010100011011"; -- 0.08492881679504301
	pesos_i(6090) := b"0000000000000000_0000000000000000_0001100011001111_1010110010010011"; -- 0.09691885567672999
	pesos_i(6091) := b"0000000000000000_0000000000000000_0001101110111111_0001010110101001"; -- 0.10838446976421427
	pesos_i(6092) := b"0000000000000000_0000000000000000_0000110100100010_0011111100110111"; -- 0.05130381672104875
	pesos_i(6093) := b"1111111111111111_1111111111111111_1111010011011001_0100110000101011"; -- -0.04355930280855448
	pesos_i(6094) := b"1111111111111111_1111111111111111_1101110100001100_1101010101101011"; -- -0.13652292394323595
	pesos_i(6095) := b"0000000000000000_0000000000000000_0000001000001000_1000101011101101"; -- 0.00794285101644971
	pesos_i(6096) := b"0000000000000000_0000000000000000_0001000011101001_1101001100101100"; -- 0.06606788474930408
	pesos_i(6097) := b"1111111111111111_1111111111111111_1111110000110000_0011011101101010"; -- -0.014889275201551894
	pesos_i(6098) := b"0000000000000000_0000000000000000_0001110111001111_1011011100001010"; -- 0.11645072934346153
	pesos_i(6099) := b"1111111111111111_1111111111111111_1111001011111010_1010000101110111"; -- -0.05086317863270405
	pesos_i(6100) := b"0000000000000000_0000000000000000_0000110011011001_1100011010001110"; -- 0.050197992062349366
	pesos_i(6101) := b"0000000000000000_0000000000000000_0000001001100010_0010001001000000"; -- 0.009309902842780013
	pesos_i(6102) := b"0000000000000000_0000000000000000_0001100101010011_1101001001111011"; -- 0.0989352751152939
	pesos_i(6103) := b"0000000000000000_0000000000000000_0000101001001001_1101011111101011"; -- 0.04018926122795535
	pesos_i(6104) := b"1111111111111111_1111111111111111_1110111100111111_0001000100001110"; -- -0.06544392975460238
	pesos_i(6105) := b"0000000000000000_0000000000000000_0001110000110010_1100010000101100"; -- 0.11014963225910925
	pesos_i(6106) := b"0000000000000000_0000000000000000_0010001101011010_1111000100000001"; -- 0.13810640597013113
	pesos_i(6107) := b"1111111111111111_1111111111111111_1111000101110011_1101101000001111"; -- -0.056825992014925955
	pesos_i(6108) := b"0000000000000000_0000000000000000_0000011111110000_1011111110110000"; -- 0.031017284785887615
	pesos_i(6109) := b"1111111111111111_1111111111111111_1111001010010011_0001010100100000"; -- -0.052443198830294226
	pesos_i(6110) := b"0000000000000000_0000000000000000_0001110100111110_0011101100010001"; -- 0.1142308155113688
	pesos_i(6111) := b"0000000000000000_0000000000000000_0000000100100010_1100000010000000"; -- 0.004436522802719195
	pesos_i(6112) := b"1111111111111111_1111111111111111_1110100001111011_0010110110111011"; -- -0.09187044321141323
	pesos_i(6113) := b"0000000000000000_0000000000000000_0000110110111010_1001010010001100"; -- 0.05362823874944213
	pesos_i(6114) := b"0000000000000000_0000000000000000_0010001010111100_0000001011010110"; -- 0.135681321431866
	pesos_i(6115) := b"1111111111111111_1111111111111111_1110010100010010_1100001100110000"; -- -0.10518245777059625
	pesos_i(6116) := b"1111111111111111_1111111111111111_1110011010100011_0010100011101100"; -- -0.09907287826903796
	pesos_i(6117) := b"0000000000000000_0000000000000000_0010101101010010_0100110101100110"; -- 0.16922458392709436
	pesos_i(6118) := b"0000000000000000_0000000000000000_0000001011010000_1101110000010110"; -- 0.010999446268412387
	pesos_i(6119) := b"0000000000000000_0000000000000000_0010000101111100_0011001010010000"; -- 0.13080135349178842
	pesos_i(6120) := b"0000000000000000_0000000000000000_0001011101001101_0101000000011100"; -- 0.09102345163969985
	pesos_i(6121) := b"1111111111111111_1111111111111111_1110100100000101_0001011011011011"; -- -0.08976609377493125
	pesos_i(6122) := b"1111111111111111_1111111111111111_1101111010101110_0011011001001001"; -- -0.1301542350710084
	pesos_i(6123) := b"1111111111111111_1111111111111111_1101110000100111_0010101100110110"; -- -0.14002733164761166
	pesos_i(6124) := b"1111111111111111_1111111111111111_1100110010100011_0010001011000001"; -- -0.20063574597140887
	pesos_i(6125) := b"0000000000000000_0000000000000000_0000011010011110_0100111101101110"; -- 0.025853123016336483
	pesos_i(6126) := b"0000000000000000_0000000000000000_0010111100000100_0001001011111000"; -- 0.18365591579295004
	pesos_i(6127) := b"1111111111111111_1111111111111111_1111101001010100_0000110011101001"; -- -0.022154992273550073
	pesos_i(6128) := b"1111111111111111_1111111111111111_1111011011001110_0111110101111110"; -- -0.03591170956599632
	pesos_i(6129) := b"1111111111111111_1111111111111111_1101010101010011_0001111001000111"; -- -0.16670046574765054
	pesos_i(6130) := b"0000000000000000_0000000000000000_0001101111101100_0000110011110101"; -- 0.1090705966075419
	pesos_i(6131) := b"1111111111111111_1111111111111111_1101111001100110_1001010001101001"; -- -0.13124725759706166
	pesos_i(6132) := b"0000000000000000_0000000000000000_0000000111101111_0001100100100001"; -- 0.007554598413586303
	pesos_i(6133) := b"1111111111111111_1111111111111111_1111011111001011_1100100001101111"; -- -0.03204676906153066
	pesos_i(6134) := b"1111111111111111_1111111111111111_1111110100011001_0010110111110010"; -- -0.01133454180875938
	pesos_i(6135) := b"0000000000000000_0000000000000000_0000110111110001_1001001011111001"; -- 0.054467378394161665
	pesos_i(6136) := b"1111111111111111_1111111111111111_1111101100001000_1111010110101010"; -- -0.019394537031896912
	pesos_i(6137) := b"1111111111111111_1111111111111111_1101100100111001_0000110001011011"; -- -0.15147326250167847
	pesos_i(6138) := b"0000000000000000_0000000000000000_0000111011110001_0010111111010101"; -- 0.05836771917376922
	pesos_i(6139) := b"0000000000000000_0000000000000000_0000011110000111_1011101000110100"; -- 0.02941478504257788
	pesos_i(6140) := b"0000000000000000_0000000000000000_0001010111101101_1111001111000011"; -- 0.08566211243038682
	pesos_i(6141) := b"0000000000000000_0000000000000000_0010011101100000_1010010011101010"; -- 0.15381842339120996
	pesos_i(6142) := b"0000000000000000_0000000000000000_0001101001110101_1110110010111011"; -- 0.10336188845688071
	pesos_i(6143) := b"1111111111111111_1111111111111111_1110011111000000_1010100001101000"; -- -0.09471652468094181
	pesos_i(6144) := b"1111111111111111_1111111111111111_1111000110000001_1101010100101001"; -- -0.056612660922838086
	pesos_i(6145) := b"1111111111111111_1111111111111111_1110011101001101_0001011100011010"; -- -0.0964799461926964
	pesos_i(6146) := b"1111111111111111_1111111111111111_1110110010111011_0100101100110011"; -- -0.07526712411184736
	pesos_i(6147) := b"1111111111111111_1111111111111111_1101111000001110_1101010001001001"; -- -0.13258622373093304
	pesos_i(6148) := b"0000000000000000_0000000000000000_0001011000000000_0100010110011011"; -- 0.08594164870932729
	pesos_i(6149) := b"0000000000000000_0000000000000000_0000010100011111_0000111100000011"; -- 0.020005167247888794
	pesos_i(6150) := b"0000000000000000_0000000000000000_0000101001101111_1011110110111101"; -- 0.040767534824148306
	pesos_i(6151) := b"1111111111111111_1111111111111111_1110001010000111_1110000110010000"; -- -0.11511411897574726
	pesos_i(6152) := b"1111111111111111_1111111111111111_1110111100010011_0011100111100111"; -- -0.06611288182292163
	pesos_i(6153) := b"1111111111111111_1111111111111111_1111111001111111_1111100011100001"; -- -0.005859799391755067
	pesos_i(6154) := b"0000000000000000_0000000000000000_0010011111001011_0001011110110111"; -- 0.15544269761274168
	pesos_i(6155) := b"0000000000000000_0000000000000000_0000100000011110_1101111000000111"; -- 0.03172099764795988
	pesos_i(6156) := b"1111111111111111_1111111111111111_1101010110100010_1010100100101100"; -- -0.16548674269647454
	pesos_i(6157) := b"1111111111111111_1111111111111111_1101010100010100_0101100101001110"; -- -0.16765825125110823
	pesos_i(6158) := b"0000000000000000_0000000000000000_0000100101011110_0001011110111110"; -- 0.036591991357821256
	pesos_i(6159) := b"0000000000000000_0000000000000000_0001010100011110_0001110111111100"; -- 0.0824908008787678
	pesos_i(6160) := b"0000000000000000_0000000000000000_0000011000000010_1100101010001001"; -- 0.02348008962208411
	pesos_i(6161) := b"1111111111111111_1111111111111111_1110001011101010_1100010011011110"; -- -0.11360520925044845
	pesos_i(6162) := b"0000000000000000_0000000000000000_0001011111100010_1000110010010001"; -- 0.09330061473275601
	pesos_i(6163) := b"0000000000000000_0000000000000000_0010000111101110_1000010001100000"; -- 0.1325457319336304
	pesos_i(6164) := b"1111111111111111_1111111111111111_1101110110000110_1100010101000000"; -- -0.13466231535646697
	pesos_i(6165) := b"1111111111111111_1111111111111111_1101100100001110_1010111001011000"; -- -0.15211973535773293
	pesos_i(6166) := b"1111111111111111_1111111111111111_1111001011101110_0111101001111111"; -- -0.05104860692703011
	pesos_i(6167) := b"1111111111111111_1111111111111111_1110001001111000_1111010110101000"; -- -0.11534180296110827
	pesos_i(6168) := b"1111111111111111_1111111111111111_1110100011110011_0011010000000101"; -- -0.09003901365787445
	pesos_i(6169) := b"1111111111111111_1111111111111111_1110101111111011_0000011101010011"; -- -0.07820085749080626
	pesos_i(6170) := b"0000000000000000_0000000000000000_0010000000011011_0001001011111101"; -- 0.12541311899519003
	pesos_i(6171) := b"1111111111111111_1111111111111111_1100010010001011_1000101111001010"; -- -0.23224569627543812
	pesos_i(6172) := b"0000000000000000_0000000000000000_0000010101101111_1110001000110110"; -- 0.021238458894299213
	pesos_i(6173) := b"0000000000000000_0000000000000000_0001000101100001_0000000000010111"; -- 0.06788635789166184
	pesos_i(6174) := b"1111111111111111_1111111111111111_1101101110011010_1001010000111011"; -- -0.14217256120986543
	pesos_i(6175) := b"0000000000000000_0000000000000000_0001101110001111_1001000000000000"; -- 0.1076593399832033
	pesos_i(6176) := b"0000000000000000_0000000000000000_0000010010001110_0111100100101111"; -- 0.017798971091208905
	pesos_i(6177) := b"0000000000000000_0000000000000000_0001001011000011_1111101001110001"; -- 0.0733028914451578
	pesos_i(6178) := b"1111111111111111_1111111111111111_1110110100010101_1010101100100010"; -- -0.07388811521786304
	pesos_i(6179) := b"1111111111111111_1111111111111111_1111001111111110_0111001101000110"; -- -0.046898646837285916
	pesos_i(6180) := b"0000000000000000_0000000000000000_0000000001000100_0010111100101100"; -- 0.001040409279412299
	pesos_i(6181) := b"1111111111111111_1111111111111111_1110011001000110_0010001111011010"; -- -0.10049224792258042
	pesos_i(6182) := b"1111111111111111_1111111111111111_1101111101100001_0100010011010100"; -- -0.1274220449418031
	pesos_i(6183) := b"0000000000000000_0000000000000000_0010010001010110_1010110101111100"; -- 0.14194759644659094
	pesos_i(6184) := b"1111111111111111_1111111111111111_1101101001110011_1011100100110101"; -- -0.14667170009211236
	pesos_i(6185) := b"1111111111111111_1111111111111111_1100111001011001_1111100011000111"; -- -0.19393963950461823
	pesos_i(6186) := b"1111111111111111_1111111111111111_1111110011101001_1100000101100011"; -- -0.012058175303732547
	pesos_i(6187) := b"1111111111111111_1111111111111111_1101100110001100_1001100100111000"; -- -0.15019838690175957
	pesos_i(6188) := b"1111111111111111_1111111111111111_1111010101011111_1010011010000111"; -- -0.04150923932974582
	pesos_i(6189) := b"1111111111111111_1111111111111111_1100101101110101_1011010111101011"; -- -0.20523512844706118
	pesos_i(6190) := b"0000000000000000_0000000000000000_0001010111101010_0111010010001010"; -- 0.08560875292338022
	pesos_i(6191) := b"0000000000000000_0000000000000000_0000100000010001_0000010011100111"; -- 0.03150969158528573
	pesos_i(6192) := b"1111111111111111_1111111111111111_1100111011111111_1011011010001111"; -- -0.1914106275082013
	pesos_i(6193) := b"1111111111111111_1111111111111111_1111110101100000_1011011000111011"; -- -0.010243044576825618
	pesos_i(6194) := b"0000000000000000_0000000000000000_0001100100100000_0111110110111111"; -- 0.09815202621903624
	pesos_i(6195) := b"0000000000000000_0000000000000000_0000010111000111_0011101000011011"; -- 0.022571212395211548
	pesos_i(6196) := b"1111111111111111_1111111111111111_1110111101110110_1001110100001010"; -- -0.06459635269841077
	pesos_i(6197) := b"0000000000000000_0000000000000000_0001101101111100_0110110101100000"; -- 0.10736735907880923
	pesos_i(6198) := b"0000000000000000_0000000000000000_0001001000101111_0100110111001010"; -- 0.07103429965506147
	pesos_i(6199) := b"0000000000000000_0000000000000000_0000001010100100_0000000010101001"; -- 0.010314980815881678
	pesos_i(6200) := b"0000000000000000_0000000000000000_0001110010001010_0010110000011001"; -- 0.11148334141595309
	pesos_i(6201) := b"1111111111111111_1111111111111111_1110011101111101_0011101110111010"; -- -0.09574534137793818
	pesos_i(6202) := b"0000000000000000_0000000000000000_0001110001010110_1110011101010111"; -- 0.11070104487208599
	pesos_i(6203) := b"0000000000000000_0000000000000000_0000011011011001_0111001110101101"; -- 0.026755552098435803
	pesos_i(6204) := b"0000000000000000_0000000000000000_0010110110111010_0010010101001010"; -- 0.17862160734680282
	pesos_i(6205) := b"0000000000000000_0000000000000000_0001110010000111_0010111101010010"; -- 0.11143775714064158
	pesos_i(6206) := b"0000000000000000_0000000000000000_0010000001111001_0101111101010001"; -- 0.12685199470651312
	pesos_i(6207) := b"1111111111111111_1111111111111111_1101100000100101_0000001011110110"; -- -0.15568524822551635
	pesos_i(6208) := b"1111111111111111_1111111111111111_1111110100010101_1111011010100001"; -- -0.011383615253905351
	pesos_i(6209) := b"0000000000000000_0000000000000000_0001100110011000_1110101011101001"; -- 0.09998958776533044
	pesos_i(6210) := b"0000000000000000_0000000000000000_0001010101010110_1100111001001010"; -- 0.0833558015432626
	pesos_i(6211) := b"0000000000000000_0000000000000000_0000101101010011_1111101111101110"; -- 0.044250245743136574
	pesos_i(6212) := b"1111111111111111_1111111111111111_1111001000000110_1101001011110011"; -- -0.0545833736637806
	pesos_i(6213) := b"1111111111111111_1111111111111111_1101100101010101_0110101101100011"; -- -0.15104035223371945
	pesos_i(6214) := b"1111111111111111_1111111111111111_1110001001110001_0110001100011110"; -- -0.11545734910443871
	pesos_i(6215) := b"0000000000000000_0000000000000000_0000101010100001_1111110111100101"; -- 0.0415342982211663
	pesos_i(6216) := b"1111111111111111_1111111111111111_1110110011110000_1000010000110010"; -- -0.07445501126802952
	pesos_i(6217) := b"1111111111111111_1111111111111111_1111111100001101_0000011011101000"; -- -0.003707474013172309
	pesos_i(6218) := b"1111111111111111_1111111111111111_1111000000010100_1110110100100011"; -- -0.062180689805309844
	pesos_i(6219) := b"0000000000000000_0000000000000000_0001100001011011_0110100010100110"; -- 0.09514478726939404
	pesos_i(6220) := b"1111111111111111_1111111111111111_1111011001110010_1011110000100011"; -- -0.037311784335118496
	pesos_i(6221) := b"0000000000000000_0000000000000000_0000010111110011_0010001000001110"; -- 0.023241165607464587
	pesos_i(6222) := b"1111111111111111_1111111111111111_1111001100000000_1011110111111000"; -- -0.05076992704247171
	pesos_i(6223) := b"1111111111111111_1111111111111111_1111111011000110_0100101010110111"; -- -0.0047868063026824115
	pesos_i(6224) := b"1111111111111111_1111111111111111_1100110100001111_1010001111100101"; -- -0.19898009926927757
	pesos_i(6225) := b"0000000000000000_0000000000000000_0001111100111011_0100100010111100"; -- 0.12199835390681955
	pesos_i(6226) := b"1111111111111111_1111111111111111_1110010110111010_1101001101000101"; -- -0.10261802264196988
	pesos_i(6227) := b"0000000000000000_0000000000000000_0010011100100010_0000111001010000"; -- 0.15286340195776507
	pesos_i(6228) := b"1111111111111111_1111111111111111_1111110111011001_1011101110110011"; -- -0.008396405015886352
	pesos_i(6229) := b"0000000000000000_0000000000000000_0010101001110001_1011001001010101"; -- 0.1657973725925928
	pesos_i(6230) := b"0000000000000000_0000000000000000_0000111000000001_1000111000100011"; -- 0.05471123083347136
	pesos_i(6231) := b"0000000000000000_0000000000000000_0001110011011110_0100110000000010"; -- 0.11276698154573966
	pesos_i(6232) := b"0000000000000000_0000000000000000_0010100110101110_1101001111111110"; -- 0.1628239149223504
	pesos_i(6233) := b"0000000000000000_0000000000000000_0000110111101000_1111000001100101"; -- 0.054335617701100604
	pesos_i(6234) := b"0000000000000000_0000000000000000_0000011000110011_0111011111000000"; -- 0.024222835840787046
	pesos_i(6235) := b"1111111111111111_1111111111111111_1111111111100010_1101011010110101"; -- -0.0004449660676218211
	pesos_i(6236) := b"1111111111111111_1111111111111111_1111100110100010_0001011010000100"; -- -0.024870484095323424
	pesos_i(6237) := b"0000000000000000_0000000000000000_0001101110001101_1000111000000111"; -- 0.10762870472712999
	pesos_i(6238) := b"1111111111111111_1111111111111111_1100111010101101_0101101000011111"; -- -0.1926673578747404
	pesos_i(6239) := b"1111111111111111_1111111111111111_1110011001010111_1001111111000110"; -- -0.1002254621250184
	pesos_i(6240) := b"0000000000000000_0000000000000000_0000000100010110_0011101010010011"; -- 0.004245434742758347
	pesos_i(6241) := b"0000000000000000_0000000000000000_0001111111001011_1001101111010010"; -- 0.12420057177799529
	pesos_i(6242) := b"0000000000000000_0000000000000000_0010101111110000_0101000100001100"; -- 0.17163569010620888
	pesos_i(6243) := b"0000000000000000_0000000000000000_0000110110000110_0000101100110111"; -- 0.05282659628713648
	pesos_i(6244) := b"1111111111111111_1111111111111111_1110111000110000_0101111111001101"; -- -0.0695743680554763
	pesos_i(6245) := b"1111111111111111_1111111111111111_1111100010100010_0000100011011101"; -- -0.02877754795744996
	pesos_i(6246) := b"1111111111111111_1111111111111111_1111010101111100_0100101100101110"; -- -0.04107217906511698
	pesos_i(6247) := b"1111111111111111_1111111111111111_1111011111010101_1000011011000100"; -- -0.031898095369672225
	pesos_i(6248) := b"1111111111111111_1111111111111111_1111101111000110_1000110100011100"; -- -0.016501598917345327
	pesos_i(6249) := b"1111111111111111_1111111111111111_1111010101111110_1101011000101100"; -- -0.04103337695446838
	pesos_i(6250) := b"0000000000000000_0000000000000000_0001001100110110_0101111100010000"; -- 0.07504839066304152
	pesos_i(6251) := b"1111111111111111_1111111111111111_1110000100100110_0111001011101011"; -- -0.12050706637685223
	pesos_i(6252) := b"1111111111111111_1111111111111111_1111010011010110_1101111101010111"; -- -0.04359630703447679
	pesos_i(6253) := b"1111111111111111_1111111111111111_1100111101000011_0111110111011000"; -- -0.19037641015595647
	pesos_i(6254) := b"0000000000000000_0000000000000000_0001111110001001_1011001000100111"; -- 0.12319482280545813
	pesos_i(6255) := b"0000000000000000_0000000000000000_0001100111101010_0011110011000011"; -- 0.10123042826333338
	pesos_i(6256) := b"1111111111111111_1111111111111111_1110100100111011_1010011101101100"; -- -0.0889335024153706
	pesos_i(6257) := b"1111111111111111_1111111111111111_1101101000001100_1100100000111101"; -- -0.14824245948048384
	pesos_i(6258) := b"0000000000000000_0000000000000000_0010011000001111_1000111001000111"; -- 0.1486748623298391
	pesos_i(6259) := b"1111111111111111_1111111111111111_1111110011111101_1110010101011100"; -- -0.011750855577525164
	pesos_i(6260) := b"0000000000000000_0000000000000000_0010100010101000_0111011010000001"; -- 0.15882053984516242
	pesos_i(6261) := b"0000000000000000_0000000000000000_0011000101111101_1000011000000101"; -- 0.19332158684618925
	pesos_i(6262) := b"1111111111111111_1111111111111111_1110110001001000_1101110110110100"; -- -0.07701315261381012
	pesos_i(6263) := b"1111111111111111_1111111111111111_1100100010001101_1100000100000111"; -- -0.21658700535039102
	pesos_i(6264) := b"1111111111111111_1111111111111111_1110111010010101_1000010001101100"; -- -0.06803104742197871
	pesos_i(6265) := b"1111111111111111_1111111111111111_1111110011110001_0001110101001100"; -- -0.011945885558309893
	pesos_i(6266) := b"1111111111111111_1111111111111111_1101111010001100_0001101110011001"; -- -0.1306746246933479
	pesos_i(6267) := b"0000000000000000_0000000000000000_0000000111111111_1011010110101111"; -- 0.007808070293005603
	pesos_i(6268) := b"1111111111111111_1111111111111111_1111101010100100_1010011010100100"; -- -0.02092512604269446
	pesos_i(6269) := b"1111111111111111_1111111111111111_1110010000010011_0110100011111010"; -- -0.1090788260053473
	pesos_i(6270) := b"1111111111111111_1111111111111111_1110000010110010_0110100111010110"; -- -0.12227762730270587
	pesos_i(6271) := b"1111111111111111_1111111111111111_1101010011100010_0110100110101000"; -- -0.16842021608796262
	pesos_i(6272) := b"1111111111111111_1111111111111111_1100111111111101_0101111000001001"; -- -0.18754017149724725
	pesos_i(6273) := b"1111111111111111_1111111111111111_1110100001000011_0111110100011110"; -- -0.0927202036238701
	pesos_i(6274) := b"0000000000000000_0000000000000000_0001100100111110_1000101110000101"; -- 0.09861061096613044
	pesos_i(6275) := b"1111111111111111_1111111111111111_1111110000011011_1010010101000000"; -- -0.015203163121751358
	pesos_i(6276) := b"1111111111111111_1111111111111111_1101100111011010_1001010010100101"; -- -0.14900847415952354
	pesos_i(6277) := b"1111111111111111_1111111111111111_1111100110000100_1011100110010110"; -- -0.025318527964650842
	pesos_i(6278) := b"0000000000000000_0000000000000000_0010100100111110_1010110011110011"; -- 0.16111260355122242
	pesos_i(6279) := b"0000000000000000_0000000000000000_0001000110111100_1001001010000011"; -- 0.06928363516646585
	pesos_i(6280) := b"1111111111111111_1111111111111111_1111000000110111_0100100111110110"; -- -0.06165635808888906
	pesos_i(6281) := b"0000000000000000_0000000000000000_0011100110100110_0010101110011110"; -- 0.22519180884719958
	pesos_i(6282) := b"0000000000000000_0000000000000000_0000100000010111_0111001110110110"; -- 0.03160784911734549
	pesos_i(6283) := b"0000000000000000_0000000000000000_0000110010011101_1110100010101100"; -- 0.049284498122049734
	pesos_i(6284) := b"0000000000000000_0000000000000000_0010100100011101_1010101000011101"; -- 0.16060889442365042
	pesos_i(6285) := b"0000000000000000_0000000000000000_0000000111010111_1001110110111000"; -- 0.007196290494960913
	pesos_i(6286) := b"0000000000000000_0000000000000000_0000101111100110_1011010110000100"; -- 0.04648909071325007
	pesos_i(6287) := b"1111111111111111_1111111111111111_1101111001010001_1101001101010100"; -- -0.13156394187169915
	pesos_i(6288) := b"1111111111111111_1111111111111111_1101100110001001_1101001001111000"; -- -0.1502407509398315
	pesos_i(6289) := b"1111111111111111_1111111111111111_1100101101100110_1010111011001100"; -- -0.20546443473259854
	pesos_i(6290) := b"0000000000000000_0000000000000000_0001010010000010_1000001110111001"; -- 0.08011649375580726
	pesos_i(6291) := b"0000000000000000_0000000000000000_0000000000011011_1001110111010010"; -- 0.00042139405274426036
	pesos_i(6292) := b"1111111111111111_1111111111111111_1111010011111001_0111111011001011"; -- -0.04306800401737721
	pesos_i(6293) := b"1111111111111111_1111111111111111_1111000101101101_1111100111100000"; -- -0.056915648254474545
	pesos_i(6294) := b"1111111111111111_1111111111111111_1111011011000110_1010110111001111"; -- -0.036030899958380325
	pesos_i(6295) := b"1111111111111111_1111111111111111_1101110101011000_0100100010010010"; -- -0.13537165095217293
	pesos_i(6296) := b"1111111111111111_1111111111111111_1111011010110111_0100010001010110"; -- -0.03626606850376199
	pesos_i(6297) := b"1111111111111111_1111111111111111_1110000011100001_1000100100101001"; -- -0.12155859705185904
	pesos_i(6298) := b"1111111111111111_1111111111111111_1111100101110010_0001010100011100"; -- -0.02560298976300232
	pesos_i(6299) := b"1111111111111111_1111111111111111_1111100100010110_0011001110010101"; -- -0.027004982167627697
	pesos_i(6300) := b"0000000000000000_0000000000000000_0000101111000100_1101101011010111"; -- 0.045972516524071555
	pesos_i(6301) := b"1111111111111111_1111111111111111_1101110000011001_0000011111011111"; -- -0.1402430610979489
	pesos_i(6302) := b"1111111111111111_1111111111111111_1110110000010101_0101000001111001"; -- -0.07779976883790553
	pesos_i(6303) := b"0000000000000000_0000000000000000_0001011100100111_1100011100001010"; -- 0.09045070644211518
	pesos_i(6304) := b"1111111111111111_1111111111111111_1110110010110111_0111011101100011"; -- -0.0753255256380205
	pesos_i(6305) := b"1111111111111111_1111111111111111_1111110000000101_0111101000010101"; -- -0.01554142930321498
	pesos_i(6306) := b"1111111111111111_1111111111111111_1111011000110011_0110100001001001"; -- -0.03827808592614704
	pesos_i(6307) := b"1111111111111111_1111111111111111_1110001111100110_0000011101000001"; -- -0.10977129618401724
	pesos_i(6308) := b"1111111111111111_1111111111111111_1110100110100101_1100100100000000"; -- -0.08731406934567387
	pesos_i(6309) := b"1111111111111111_1111111111111111_1101100111010100_1111100010011110"; -- -0.14909406788053123
	pesos_i(6310) := b"0000000000000000_0000000000000000_0010010000110000_1110111110001110"; -- 0.14137170041558172
	pesos_i(6311) := b"1111111111111111_1111111111111111_1110011110011110_0011101100100101"; -- -0.09524183596639925
	pesos_i(6312) := b"1111111111111111_1111111111111111_1110011100110011_0110111001100111"; -- -0.09687147131215715
	pesos_i(6313) := b"1111111111111111_1111111111111111_1111001010100111_0110010110101100"; -- -0.05213322218579538
	pesos_i(6314) := b"1111111111111111_1111111111111111_1110101111010011_1101000101110001"; -- -0.0787991618304081
	pesos_i(6315) := b"1111111111111111_1111111111111111_1101010100100000_0011011110011011"; -- -0.1674771545116907
	pesos_i(6316) := b"0000000000000000_0000000000000000_0000111001001111_0010100100011010"; -- 0.055895394117171426
	pesos_i(6317) := b"0000000000000000_0000000000000000_0000100110011010_1000000110011101"; -- 0.037513829182585556
	pesos_i(6318) := b"0000000000000000_0000000000000000_0000100000010111_0111010100001101"; -- 0.03160792895318227
	pesos_i(6319) := b"0000000000000000_0000000000000000_0010101000001000_1001001100111110"; -- 0.16419334667636099
	pesos_i(6320) := b"1111111111111111_1111111111111111_1111101100110001_1101111010101011"; -- -0.018770297287879358
	pesos_i(6321) := b"0000000000000000_0000000000000000_0010000001100010_1001100110011001"; -- 0.12650451648241684
	pesos_i(6322) := b"1111111111111111_1111111111111111_1110110111100010_1111111111001110"; -- -0.07075501663409596
	pesos_i(6323) := b"1111111111111111_1111111111111111_1111010011100111_0001000011111111"; -- -0.04334920664755801
	pesos_i(6324) := b"1111111111111111_1111111111111111_1111110010101010_1011110100110011"; -- -0.013019728770355427
	pesos_i(6325) := b"0000000000000000_0000000000000000_0000000010110101_1110010001000111"; -- 0.0027754470986908566
	pesos_i(6326) := b"1111111111111111_1111111111111111_1100000010010100_1111010011100000"; -- -0.24772710357003952
	pesos_i(6327) := b"0000000000000000_0000000000000000_0001001011000101_1101101110101010"; -- 0.07333157454527814
	pesos_i(6328) := b"0000000000000000_0000000000000000_0000100001110001_0100010011111001"; -- 0.03297835431420885
	pesos_i(6329) := b"1111111111111111_1111111111111111_1111101111110011_0101101001100101"; -- -0.015817976288290958
	pesos_i(6330) := b"1111111111111111_1111111111111111_1011110010110100_1101001000010001"; -- -0.26286589706801894
	pesos_i(6331) := b"0000000000000000_0000000000000000_0001110000100110_0000100001110100"; -- 0.10995533794268628
	pesos_i(6332) := b"0000000000000000_0000000000000000_0001000101010110_0100011100100100"; -- 0.06772274608435888
	pesos_i(6333) := b"0000000000000000_0000000000000000_0001011010100111_1111111010110100"; -- 0.08850089931978883
	pesos_i(6334) := b"1111111111111111_1111111111111111_1111100010100110_1010100101110011"; -- -0.028706940987607305
	pesos_i(6335) := b"1111111111111111_1111111111111111_1010110110000011_1101010110111010"; -- -0.3222071095395587
	pesos_i(6336) := b"1111111111111111_1111111111111111_1100110010101011_0010110100111111"; -- -0.20051305019117446
	pesos_i(6337) := b"0000000000000000_0000000000000000_0001101010100000_0011011010110101"; -- 0.10400716703611823
	pesos_i(6338) := b"0000000000000000_0000000000000000_0000100101011001_0011101010100010"; -- 0.036517777070242244
	pesos_i(6339) := b"1111111111111111_1111111111111111_1111001100001010_1000111110111110"; -- -0.050620094470977484
	pesos_i(6340) := b"1111111111111111_1111111111111111_1110111011010010_0000000001111000"; -- -0.06710812633462035
	pesos_i(6341) := b"1111111111111111_1111111111111111_1011001011110011_1101100100111011"; -- -0.30096666624970103
	pesos_i(6342) := b"0000000000000000_0000000000000000_0001001111001011_0101001100010000"; -- 0.07732123506565913
	pesos_i(6343) := b"0000000000000000_0000000000000000_0010000001011010_1110010001110001"; -- 0.12638690727424287
	pesos_i(6344) := b"1111111111111111_1111111111111111_1100001101001010_0110111100110001"; -- -0.2371454720005807
	pesos_i(6345) := b"1111111111111111_1111111111111111_1110101011100100_0010111010101010"; -- -0.08245571480562196
	pesos_i(6346) := b"1111111111111111_1111111111111111_1110101101000110_0100110011101000"; -- -0.08095855087383623
	pesos_i(6347) := b"1111111111111111_1111111111111111_1110000100011111_1001101001001011"; -- -0.12061153103686263
	pesos_i(6348) := b"0000000000000000_0000000000000000_0010110010011011_1010010001101100"; -- 0.1742499125100464
	pesos_i(6349) := b"1111111111111111_1111111111111111_1110111001111001_1011110111010101"; -- -0.0684548717012998
	pesos_i(6350) := b"1111111111111111_1111111111111111_1011111010000100_1011000011100111"; -- -0.2557877956334145
	pesos_i(6351) := b"1111111111111111_1111111111111111_1110101000010101_0101111100000101"; -- -0.0856114017941303
	pesos_i(6352) := b"0000000000000000_0000000000000000_0011011101111101_0001110011111011"; -- 0.2167528259776927
	pesos_i(6353) := b"1111111111111111_1111111111111111_1101000001001001_0001100101000011"; -- -0.18638460256972536
	pesos_i(6354) := b"0000000000000000_0000000000000000_0010000001110000_1011110011001100"; -- 0.12672023759311216
	pesos_i(6355) := b"1111111111111111_1111111111111111_1110111010110110_1001100011010111"; -- -0.06752629053465879
	pesos_i(6356) := b"1111111111111111_1111111111111111_1101011110011010_0110111000100010"; -- -0.1577998319949377
	pesos_i(6357) := b"1111111111111111_1111111111111111_1111000100110001_1101101011010001"; -- -0.057833026884951476
	pesos_i(6358) := b"1111111111111111_1111111111111111_1110010011001101_1110100010010111"; -- -0.10623308478586754
	pesos_i(6359) := b"0000000000000000_0000000000000000_0001100101101100_1011101110100010"; -- 0.0993153830194614
	pesos_i(6360) := b"0000000000000000_0000000000000000_0010101001110000_1110000000010011"; -- 0.16578484016917772
	pesos_i(6361) := b"0000000000000000_0000000000000000_0001101100100110_0010010001101101"; -- 0.10605075511578471
	pesos_i(6362) := b"0000000000000000_0000000000000000_0100010011000111_0110001101011110"; -- 0.2686674216791829
	pesos_i(6363) := b"0000000000000000_0000000000000000_0000101101011101_1001111110010010"; -- 0.0443973284259619
	pesos_i(6364) := b"1111111111111111_1111111111111111_1110100001110100_1110111000000010"; -- -0.0919657940312183
	pesos_i(6365) := b"0000000000000000_0000000000000000_0000111001010010_0000110010010100"; -- 0.05593947044568677
	pesos_i(6366) := b"0000000000000000_0000000000000000_0010011111100000_1111010100011100"; -- 0.15577632829735674
	pesos_i(6367) := b"0000000000000000_0000000000000000_0001111111100001_0110000101110111"; -- 0.12453278695612449
	pesos_i(6368) := b"1111111111111111_1111111111111111_1110111000010001_0011000111111001"; -- -0.07005012195792001
	pesos_i(6369) := b"0000000000000000_0000000000000000_0001100111100110_1101111101110110"; -- 0.10117909084107857
	pesos_i(6370) := b"0000000000000000_0000000000000000_0010100001101101_1010110110100000"; -- 0.1579235569508627
	pesos_i(6371) := b"1111111111111111_1111111111111111_1100101101101101_1011001101010000"; -- -0.20535735423850118
	pesos_i(6372) := b"1111111111111111_1111111111111111_1101001011011110_1100111110011110"; -- -0.17628767395117562
	pesos_i(6373) := b"1111111111111111_1111111111111111_1101101010001001_1010101011110001"; -- -0.1463368569947415
	pesos_i(6374) := b"1111111111111111_1111111111111111_1111001010010101_0110110001110110"; -- -0.05240747576587271
	pesos_i(6375) := b"0000000000000000_0000000000000000_0000101001100101_0100101111001110"; -- 0.040608155944924854
	pesos_i(6376) := b"0000000000000000_0000000000000000_0001100111000011_0110001000000000"; -- 0.10063755518188788
	pesos_i(6377) := b"1111111111111111_1111111111111111_1110100100100111_1110001000100110"; -- -0.08923517769849362
	pesos_i(6378) := b"0000000000000000_0000000000000000_0000000101010101_1110000100110110"; -- 0.005216670600302805
	pesos_i(6379) := b"1111111111111111_1111111111111111_1110111101010000_0101100101101010"; -- -0.06518021732414642
	pesos_i(6380) := b"1111111111111111_1111111111111111_1110001000111101_1000111110111100"; -- -0.11624814665142219
	pesos_i(6381) := b"1111111111111111_1111111111111111_1110001100111000_1101100010111000"; -- -0.11241384044392344
	pesos_i(6382) := b"1111111111111111_1111111111111111_1101011110011101_1110001010000110"; -- -0.15774711830838217
	pesos_i(6383) := b"1111111111111111_1111111111111111_1100110110111111_1010001011001100"; -- -0.1962946178188272
	pesos_i(6384) := b"1111111111111111_1111111111111111_1100111111111110_1100001001110111"; -- -0.1875189265835304
	pesos_i(6385) := b"0000000000000000_0000000000000000_0010101000011010_0010011010000000"; -- 0.16446152336097883
	pesos_i(6386) := b"0000000000000000_0000000000000000_0100011000011010_1110101000110011"; -- 0.27384818780997483
	pesos_i(6387) := b"1111111111111111_1111111111111111_1111010011011110_0011001010010110"; -- -0.04348453360709083
	pesos_i(6388) := b"1111111111111111_1111111111111111_1101101110001100_1110000101001011"; -- -0.1423815910434416
	pesos_i(6389) := b"1111111111111111_1111111111111111_1111111101010011_0000000000100011"; -- -0.00263976232905632
	pesos_i(6390) := b"1111111111111111_1111111111111111_1111111010101001_1110111001100100"; -- -0.005219555407267744
	pesos_i(6391) := b"0000000000000000_0000000000000000_0010001110000101_0110001010010000"; -- 0.1387540436926264
	pesos_i(6392) := b"1111111111111111_1111111111111111_1110001000000111_0101110011110101"; -- -0.11707514784731887
	pesos_i(6393) := b"0000000000000000_0000000000000000_0010011000100101_1000011101011111"; -- 0.14901014400245377
	pesos_i(6394) := b"1111111111111111_1111111111111111_1110000100000010_0001011110101001"; -- -0.12106182227254711
	pesos_i(6395) := b"1111111111111111_1111111111111111_1111110100101110_1000101111101101"; -- -0.011008505375597583
	pesos_i(6396) := b"1111111111111111_1111111111111111_1101000111010111_1111101010101010"; -- -0.18029816967410267
	pesos_i(6397) := b"1111111111111111_1111111111111111_1111011010101011_0011100101110111"; -- -0.03644982191649318
	pesos_i(6398) := b"0000000000000000_0000000000000000_0001111011111101_0001111101011100"; -- 0.12104984278057175
	pesos_i(6399) := b"0000000000000000_0000000000000000_0001001111001010_0110010000110010"; -- 0.07730699752153043
	pesos_i(6400) := b"1111111111111111_1111111111111111_1111110001101101_0010100011001100"; -- -0.013959360194386051
	pesos_i(6401) := b"0000000000000000_0000000000000000_0001100110101101_1110100100110100"; -- 0.10030992045738668
	pesos_i(6402) := b"0000000000000000_0000000000000000_0010101100010101_0110010010111000"; -- 0.1682951878265823
	pesos_i(6403) := b"0000000000000000_0000000000000000_0000000111111110_1000011010110101"; -- 0.007790011625566622
	pesos_i(6404) := b"0000000000000000_0000000000000000_0010011010000000_1011010010101001"; -- 0.15040139310435455
	pesos_i(6405) := b"0000000000000000_0000000000000000_0000010100111001_0001101101001011"; -- 0.02040262777346459
	pesos_i(6406) := b"0000000000000000_0000000000000000_0000101111111100_0001111110011110"; -- 0.046815849395001996
	pesos_i(6407) := b"0000000000000000_0000000000000000_0000011000101101_1010100010011001"; -- 0.024134194721988283
	pesos_i(6408) := b"1111111111111111_1111111111111111_1111001011100100_1100000111111001"; -- -0.05119693433892191
	pesos_i(6409) := b"1111111111111111_1111111111111111_1110010101000001_1010001000100110"; -- -0.10446726379716988
	pesos_i(6410) := b"1111111111111111_1111111111111111_1111111101110011_1001000111000101"; -- -0.0021428007315503314
	pesos_i(6411) := b"1111111111111111_1111111111111111_1100110000000100_0101111000011011"; -- -0.20305835571838565
	pesos_i(6412) := b"1111111111111111_1111111111111111_1100111010111110_0001100110001101"; -- -0.19241180711233521
	pesos_i(6413) := b"1111111111111111_1111111111111111_1110100001000001_0111011110010100"; -- -0.09275105124934166
	pesos_i(6414) := b"0000000000000000_0000000000000000_0011100000010000_1011100101010000"; -- 0.21900518602624766
	pesos_i(6415) := b"0000000000000000_0000000000000000_0010010111011100_1011100100001011"; -- 0.14789921302590125
	pesos_i(6416) := b"0000000000000000_0000000000000000_0001000111011100_1001100010110101"; -- 0.06977228566841477
	pesos_i(6417) := b"0000000000000000_0000000000000000_0000001001110101_0001111100111001"; -- 0.009599639232765182
	pesos_i(6418) := b"1111111111111111_1111111111111111_1101110111100001_1010101011001100"; -- -0.1332753420928115
	pesos_i(6419) := b"0000000000000000_0000000000000000_0000110010010110_1111110111000001"; -- 0.04917894321879154
	pesos_i(6420) := b"1111111111111111_1111111111111111_1111100111111001_1101010101110101"; -- -0.023531588605626146
	pesos_i(6421) := b"1111111111111111_1111111111111111_1110100010111110_0000001111110111"; -- -0.0908505937500187
	pesos_i(6422) := b"0000000000000000_0000000000000000_0000111101110000_0110111000000110"; -- 0.06030929220059093
	pesos_i(6423) := b"1111111111111111_1111111111111111_1110101001100100_0011000101010000"; -- -0.08440868174979992
	pesos_i(6424) := b"0000000000000000_0000000000000000_0001100110001000_0010001110100101"; -- 0.0997335699435704
	pesos_i(6425) := b"0000000000000000_0000000000000000_0000111001010100_1101110101011011"; -- 0.05598243212481388
	pesos_i(6426) := b"0000000000000000_0000000000000000_0000000011011101_1011101101111100"; -- 0.003383367268689608
	pesos_i(6427) := b"0000000000000000_0000000000000000_0000110010100010_1111100110000111"; -- 0.04936179691324762
	pesos_i(6428) := b"1111111111111111_1111111111111111_1111001000000001_1100100000000101"; -- -0.054660319152173925
	pesos_i(6429) := b"1111111111111111_1111111111111111_1100100111110001_1110111100000111"; -- -0.21115213468446958
	pesos_i(6430) := b"1111111111111111_1111111111111111_1100111100101111_0011001001010000"; -- -0.19068608793973998
	pesos_i(6431) := b"0000000000000000_0000000000000000_0000111111110001_1011011001000010"; -- 0.062281981646941036
	pesos_i(6432) := b"0000000000000000_0000000000000000_0010100111010010_0010100100000111"; -- 0.16336304112522881
	pesos_i(6433) := b"1111111111111111_1111111111111111_1110001001001100_1110111001100011"; -- -0.11601362303068893
	pesos_i(6434) := b"1111111111111111_1111111111111111_1100011000101101_0111001110110000"; -- -0.22586895909595403
	pesos_i(6435) := b"1111111111111111_1111111111111111_1101110100001101_0111010110110001"; -- -0.1365133706771632
	pesos_i(6436) := b"1111111111111111_1111111111111111_1110001011110101_1011100101111101"; -- -0.11343804081813788
	pesos_i(6437) := b"0000000000000000_0000000000000000_0010011101111111_0001011111010100"; -- 0.15428303637842453
	pesos_i(6438) := b"0000000000000000_0000000000000000_0000100011111100_1110001011010011"; -- 0.03510873465914121
	pesos_i(6439) := b"1111111111111111_1111111111111111_1100111000001011_1100001100101101"; -- -0.1951330200230963
	pesos_i(6440) := b"1111111111111111_1111111111111111_1100011001101011_0110111000011011"; -- -0.224923246759961
	pesos_i(6441) := b"1111111111111111_1111111111111111_1110000010101010_0111110010011101"; -- -0.1223985784039257
	pesos_i(6442) := b"0000000000000000_0000000000000000_0011000111000001_0011101100110011"; -- 0.19435472491623237
	pesos_i(6443) := b"1111111111111111_1111111111111111_1101010010011101_0000100101001001"; -- -0.16947881662969486
	pesos_i(6444) := b"0000000000000000_0000000000000000_0011001100110110_0010111000101010"; -- 0.2000454762242926
	pesos_i(6445) := b"1111111111111111_1111111111111111_1111110101011111_0110000000111000"; -- -0.010263430017316538
	pesos_i(6446) := b"1111111111111111_1111111111111111_1110101010100000_0111001011111010"; -- -0.08348924054063826
	pesos_i(6447) := b"1111111111111111_1111111111111111_1111111100100000_1001111001101000"; -- -0.0034085269736168814
	pesos_i(6448) := b"0000000000000000_0000000000000000_0001101001000001_1001100011111101"; -- 0.10256344003611677
	pesos_i(6449) := b"0000000000000000_0000000000000000_0011010000101111_1010001100101001"; -- 0.2038518880905515
	pesos_i(6450) := b"1111111111111111_1111111111111111_1101000100111010_0111001011101011"; -- -0.18270189067687698
	pesos_i(6451) := b"0000000000000000_0000000000000000_0010100100110010_0100101101111000"; -- 0.16092368779682717
	pesos_i(6452) := b"0000000000000000_0000000000000000_0001111010001101_0011000110100001"; -- 0.11934194732599679
	pesos_i(6453) := b"1111111111111111_1111111111111111_1101001111010011_1001101011000110"; -- -0.17255242025694126
	pesos_i(6454) := b"1111111111111111_1111111111111111_1111110101011010_0000010111000100"; -- -0.010345115291664068
	pesos_i(6455) := b"0000000000000000_0000000000000000_0000001001011000_1011101101111000"; -- 0.009166447404277366
	pesos_i(6456) := b"1111111111111111_1111111111111111_1111000110110101_1001000010011101"; -- -0.055823289475760776
	pesos_i(6457) := b"0000000000000000_0000000000000000_0001010111111101_0010111011011001"; -- 0.0858945160252628
	pesos_i(6458) := b"0000000000000000_0000000000000000_0010101111100010_0111110100111010"; -- 0.1714247004116212
	pesos_i(6459) := b"0000000000000000_0000000000000000_0010100011001100_1001010111111110"; -- 0.15937173308742164
	pesos_i(6460) := b"1111111111111111_1111111111111111_1111110010011101_1010101011010111"; -- -0.01321918738138479
	pesos_i(6461) := b"0000000000000000_0000000000000000_0011001100111011_0001101000101110"; -- 0.20012057905364122
	pesos_i(6462) := b"1111111111111111_1111111111111111_1110100100111010_0001101101100100"; -- -0.08895710768344901
	pesos_i(6463) := b"1111111111111111_1111111111111111_1110101101101100_1010010001100001"; -- -0.08037350300404247
	pesos_i(6464) := b"0000000000000000_0000000000000000_0010000000001011_1101111111011011"; -- 0.12518118961342553
	pesos_i(6465) := b"0000000000000000_0000000000000000_0000010111000011_0101000100011010"; -- 0.022511547860662003
	pesos_i(6466) := b"1111111111111111_1111111111111111_1101101101101110_0011110010110101"; -- -0.14284916475375303
	pesos_i(6467) := b"1111111111111111_1111111111111111_1111011100101001_0111100101110001"; -- -0.034523401139532825
	pesos_i(6468) := b"1111111111111111_1111111111111111_1110011000011100_1001000001010110"; -- -0.10112665086315466
	pesos_i(6469) := b"0000000000000000_0000000000000000_0001110001000011_1011010001111101"; -- 0.11040809676613625
	pesos_i(6470) := b"0000000000000000_0000000000000000_0010101001001000_1010000110100010"; -- 0.16517076677089956
	pesos_i(6471) := b"1111111111111111_1111111111111111_1110100011000000_1101100100011000"; -- -0.09080737277808441
	pesos_i(6472) := b"1111111111111111_1111111111111111_1110011010101110_1111101000100110"; -- -0.09889256060317983
	pesos_i(6473) := b"0000000000000000_0000000000000000_0011000000001111_0101111001100010"; -- 0.18773450758277146
	pesos_i(6474) := b"1111111111111111_1111111111111111_1111011000001101_1111111110100100"; -- -0.038848898282862386
	pesos_i(6475) := b"1111111111111111_1111111111111111_1111110111100011_1110111001011110"; -- -0.008240797081101833
	pesos_i(6476) := b"0000000000000000_0000000000000000_0001000011111111_1001011111000000"; -- 0.06640003614481037
	pesos_i(6477) := b"1111111111111111_1111111111111111_1111101001110001_0111001100001111"; -- -0.021706398885245868
	pesos_i(6478) := b"0000000000000000_0000000000000000_0000010110100010_1000101011000100"; -- 0.022011444985100072
	pesos_i(6479) := b"0000000000000000_0000000000000000_0011010011101001_1010001010001011"; -- 0.206689986199717
	pesos_i(6480) := b"0000000000000000_0000000000000000_0000111100001000_1001000010101101"; -- 0.05872444355467454
	pesos_i(6481) := b"0000000000000000_0000000000000000_0010001101011101_0101111100111000"; -- 0.1381434928779346
	pesos_i(6482) := b"0000000000000000_0000000000000000_0000110000101010_0000100001111101"; -- 0.047516374966623004
	pesos_i(6483) := b"0000000000000000_0000000000000000_0001100001010101_0011001100011101"; -- 0.09505004377087789
	pesos_i(6484) := b"1111111111111111_1111111111111111_1111111100111001_0100111110100111"; -- -0.0030317512868238417
	pesos_i(6485) := b"1111111111111111_1111111111111111_1111010010100100_0000100100011110"; -- -0.04437201518989884
	pesos_i(6486) := b"1111111111111111_1111111111111111_1110111100000000_1110011110010001"; -- -0.06639244764956588
	pesos_i(6487) := b"1111111111111111_1111111111111111_1111100001101100_0011101100111011"; -- -0.029598520458632982
	pesos_i(6488) := b"1111111111111111_1111111111111111_1101010111111000_1100001000101100"; -- -0.16417299683786046
	pesos_i(6489) := b"1111111111111111_1111111111111111_1011101001111100_0111110011111110"; -- -0.271537960149915
	pesos_i(6490) := b"0000000000000000_0000000000000000_0010110010010100_0001001100011110"; -- 0.17413444035017414
	pesos_i(6491) := b"1111111111111111_1111111111111111_1101011111011110_0110010000110100"; -- -0.1567628262544229
	pesos_i(6492) := b"1111111111111111_1111111111111111_1111011000110101_1100011000011011"; -- -0.03824197608631085
	pesos_i(6493) := b"1111111111111111_1111111111111111_1100111100101011_1010100111010101"; -- -0.1907399993978621
	pesos_i(6494) := b"0000000000000000_0000000000000000_0000001011010100_0111100101011110"; -- 0.011054597392508024
	pesos_i(6495) := b"0000000000000000_0000000000000000_0000000101010101_0100001100111001"; -- 0.005207253827754103
	pesos_i(6496) := b"1111111111111111_1111111111111111_1111101000011100_0000011100011110"; -- -0.023009829581376897
	pesos_i(6497) := b"0000000000000000_0000000000000000_0010101010001001_0000000001001101"; -- 0.16615297199726733
	pesos_i(6498) := b"1111111111111111_1111111111111111_1111110001111110_0011010101110001"; -- -0.013699207181276237
	pesos_i(6499) := b"1111111111111111_1111111111111111_1101110000110001_0111111000010100"; -- -0.13986980451111827
	pesos_i(6500) := b"1111111111111111_1111111111111111_1111011011001001_1100111101110010"; -- -0.03598311874564295
	pesos_i(6501) := b"0000000000000000_0000000000000000_0000110001001001_0101000001100110"; -- 0.047993683682596974
	pesos_i(6502) := b"1111111111111111_1111111111111111_1110001001011111_0011110100100111"; -- -0.11573426999662471
	pesos_i(6503) := b"0000000000000000_0000000000000000_0010000100010011_1100101101110000"; -- 0.12920829275493068
	pesos_i(6504) := b"1111111111111111_1111111111111111_1110101010010110_0110101110110111"; -- -0.08364226136231305
	pesos_i(6505) := b"0000000000000000_0000000000000000_0010100101110011_1011101110000011"; -- 0.16192218725785584
	pesos_i(6506) := b"0000000000000000_0000000000000000_0001100110111000_1011010101101010"; -- 0.10047468025843738
	pesos_i(6507) := b"1111111111111111_1111111111111111_1110101101011110_0100001011000000"; -- -0.08059294521927578
	pesos_i(6508) := b"1111111111111111_1111111111111111_1111010111000101_1101110100100100"; -- -0.03994958761715776
	pesos_i(6509) := b"0000000000000000_0000000000000000_0010100010101111_0100011010011011"; -- 0.1589244965665701
	pesos_i(6510) := b"1111111111111111_1111111111111111_1110000101101110_0111001101110101"; -- -0.11940840136969251
	pesos_i(6511) := b"1111111111111111_1111111111111111_1111000110101111_1000011011010100"; -- -0.05591542553552575
	pesos_i(6512) := b"1111111111111111_1111111111111111_1111110010000000_0000100111110111"; -- -0.01367128106659285
	pesos_i(6513) := b"0000000000000000_0000000000000000_0001001110110100_1001011010110010"; -- 0.0769743141588154
	pesos_i(6514) := b"1111111111111111_1111111111111111_1101101111000100_0100001101001000"; -- -0.14153651713247997
	pesos_i(6515) := b"1111111111111111_1111111111111111_1111100100111001_0111111000001101"; -- -0.026466485893604508
	pesos_i(6516) := b"0000000000000000_0000000000000000_0001100100101001_0111111111000001"; -- 0.09828947510147745
	pesos_i(6517) := b"1111111111111111_1111111111111111_1111011010011000_1011101001010001"; -- -0.03673205863171958
	pesos_i(6518) := b"0000000000000000_0000000000000000_0010100100110001_0011100001000010"; -- 0.16090728378051217
	pesos_i(6519) := b"0000000000000000_0000000000000000_0010101110000101_1010110110110011"; -- 0.17000852233854036
	pesos_i(6520) := b"1111111111111111_1111111111111111_1110000101001111_1001110011010001"; -- -0.11987895865072073
	pesos_i(6521) := b"0000000000000000_0000000000000000_0001111110101111_1101110110101100"; -- 0.1237772508664533
	pesos_i(6522) := b"1111111111111111_1111111111111111_1110000110111010_0001111101001100"; -- -0.11825374990960962
	pesos_i(6523) := b"0000000000000000_0000000000000000_0010000111101001_1111011100101110"; -- 0.13247628101159495
	pesos_i(6524) := b"0000000000000000_0000000000000000_0011001101100010_0110010011100111"; -- 0.2007201255414816
	pesos_i(6525) := b"1111111111111111_1111111111111111_1100110001000110_0001010110100001"; -- -0.20205559569784162
	pesos_i(6526) := b"1111111111111111_1111111111111111_1100101000111100_1011011110101111"; -- -0.2100110242487218
	pesos_i(6527) := b"1111111111111111_1111111111111111_1101000100001100_0110000101000101"; -- -0.1834048467723789
	pesos_i(6528) := b"1111111111111111_1111111111111111_1110111000000100_1111001101101111"; -- -0.07023695505165096
	pesos_i(6529) := b"0000000000000000_0000000000000000_0010000001111010_1011000001001000"; -- 0.1268720794230611
	pesos_i(6530) := b"0000000000000000_0000000000000000_0000110101111101_1011111001101110"; -- 0.052699949030338214
	pesos_i(6531) := b"1111111111111111_1111111111111111_1111100111101111_0101101110100001"; -- -0.02369143790966639
	pesos_i(6532) := b"1111111111111111_1111111111111111_1111101010001100_1011001101110011"; -- -0.021290573586036227
	pesos_i(6533) := b"0000000000000000_0000000000000000_0001010000101111_0000101000010100"; -- 0.07884276373076551
	pesos_i(6534) := b"0000000000000000_0000000000000000_0001100010011110_1011011111101001"; -- 0.09617185066472955
	pesos_i(6535) := b"0000000000000000_0000000000000000_0001011111111110_1000011011011001"; -- 0.09372752007857973
	pesos_i(6536) := b"1111111111111111_1111111111111111_1111101111001000_1100111001010001"; -- -0.016467194779672328
	pesos_i(6537) := b"0000000000000000_0000000000000000_0010111100111111_1001000111111010"; -- 0.1845637545814215
	pesos_i(6538) := b"0000000000000000_0000000000000000_0001110011110101_0110000001001011"; -- 0.11311914273010308
	pesos_i(6539) := b"0000000000000000_0000000000000000_0001110111111111_1001000001110100"; -- 0.11718085135473272
	pesos_i(6540) := b"1111111111111111_1111111111111111_1110000100101001_1100011010000110"; -- -0.12045630673349074
	pesos_i(6541) := b"1111111111111111_1111111111111111_1111000011100011_1010110111101111"; -- -0.05902588764905444
	pesos_i(6542) := b"1111111111111111_1111111111111111_1111010011001100_1101111100100110"; -- -0.04374890626987542
	pesos_i(6543) := b"1111111111111111_1111111111111111_1101001111111110_0111110100100110"; -- -0.1718980582250091
	pesos_i(6544) := b"0000000000000000_0000000000000000_0000111101100110_1011111110011010"; -- 0.06016156681716945
	pesos_i(6545) := b"1111111111111111_1111111111111111_1101001001100101_0001011101110010"; -- -0.178144964793913
	pesos_i(6546) := b"1111111111111111_1111111111111111_1110100110110100_1110110001011110"; -- -0.08708307937445983
	pesos_i(6547) := b"0000000000000000_0000000000000000_0001011111001001_1110010000000001"; -- 0.09292435674772885
	pesos_i(6548) := b"1111111111111111_1111111111111111_1101111001110101_1010001110010100"; -- -0.13101747164375646
	pesos_i(6549) := b"0000000000000000_0000000000000000_0001011011110111_0100111101111111"; -- 0.0897111592736109
	pesos_i(6550) := b"0000000000000000_0000000000000000_0001100100110111_0100100110011000"; -- 0.09849986985767267
	pesos_i(6551) := b"1111111111111111_1111111111111111_1101101001000100_1000100101001100"; -- -0.1473917187512726
	pesos_i(6552) := b"1111111111111111_1111111111111111_1111110110110010_0110000011100100"; -- -0.008996910332016175
	pesos_i(6553) := b"0000000000000000_0000000000000000_0001111100110100_1101001000011111"; -- 0.12189973117750653
	pesos_i(6554) := b"0000000000000000_0000000000000000_0010010001011110_0010100110001100"; -- 0.14206180263827012
	pesos_i(6555) := b"0000000000000000_0000000000000000_0000111010010000_1000010011100000"; -- 0.056892685557224106
	pesos_i(6556) := b"0000000000000000_0000000000000000_0000011011111101_0001001101111010"; -- 0.027299134621117754
	pesos_i(6557) := b"1111111111111111_1111111111111111_1111101011011110_1010100001010010"; -- -0.020040016247673254
	pesos_i(6558) := b"1111111111111111_1111111111111111_1110000010001010_0100000110101011"; -- -0.1228903729852024
	pesos_i(6559) := b"0000000000000000_0000000000000000_0001100000011100_1101001001111000"; -- 0.09418979095631408
	pesos_i(6560) := b"0000000000000000_0000000000000000_0000010010011100_1011101000010000"; -- 0.018016461368059275
	pesos_i(6561) := b"0000000000000000_0000000000000000_0001001001100001_1111100010011110"; -- 0.07180742125799132
	pesos_i(6562) := b"0000000000000000_0000000000000000_0001001100010010_0110100101101001"; -- 0.07449969120825972
	pesos_i(6563) := b"1111111111111111_1111111111111111_1100100111100101_0000101100000010"; -- -0.2113488312256736
	pesos_i(6564) := b"1111111111111111_1111111111111111_1110010110111111_0100100011110110"; -- -0.10254997250695172
	pesos_i(6565) := b"0000000000000000_0000000000000000_0000010100001001_0111100100001110"; -- 0.01967579450775766
	pesos_i(6566) := b"0000000000000000_0000000000000000_0001110110011001_0010010000110101"; -- 0.11561800276485766
	pesos_i(6567) := b"0000000000000000_0000000000000000_0011000001101010_1001001011010011"; -- 0.18912618306430698
	pesos_i(6568) := b"0000000000000000_0000000000000000_0010011100110000_0101100011101111"; -- 0.15308147273470946
	pesos_i(6569) := b"0000000000000000_0000000000000000_0001100011011110_0101000110011010"; -- 0.09714231501635491
	pesos_i(6570) := b"1111111111111111_1111111111111111_1110011000010010_0001100000010001"; -- -0.10128640734085927
	pesos_i(6571) := b"0000000000000000_0000000000000000_0001111100111111_0101101110000110"; -- 0.12206050891534605
	pesos_i(6572) := b"0000000000000000_0000000000000000_0010000011011111_1001010101111111"; -- 0.1284116205150092
	pesos_i(6573) := b"0000000000000000_0000000000000000_0010000011000010_1000110001110101"; -- 0.1279685769488265
	pesos_i(6574) := b"1111111111111111_1111111111111111_1111111011111011_0010010111111111"; -- -0.0039802792871462675
	pesos_i(6575) := b"0000000000000000_0000000000000000_0001010001111010_1001100011001001"; -- 0.07999567887010386
	pesos_i(6576) := b"1111111111111111_1111111111111111_1101101101011011_0111110011110010"; -- -0.14313525297895352
	pesos_i(6577) := b"1111111111111111_1111111111111111_1110111010111000_0111101101101100"; -- -0.0674975263902665
	pesos_i(6578) := b"0000000000000000_0000000000000000_0011010001110000_1010011110001110"; -- 0.20484397136662758
	pesos_i(6579) := b"0000000000000000_0000000000000000_0011011100010011_0010011111001011"; -- 0.21513603888777755
	pesos_i(6580) := b"0000000000000000_0000000000000000_0000110100010111_1001011101001101"; -- 0.05114122042538978
	pesos_i(6581) := b"0000000000000000_0000000000000000_0001010001010000_1000101100000111"; -- 0.07935398977662193
	pesos_i(6582) := b"0000000000000000_0000000000000000_0001101000111111_1100110100101100"; -- 0.10253603299502197
	pesos_i(6583) := b"0000000000000000_0000000000000000_0011010101000010_0001000010111011"; -- 0.2080393272111597
	pesos_i(6584) := b"0000000000000000_0000000000000000_0011000101000000_0000010110100011"; -- 0.1923831485895847
	pesos_i(6585) := b"1111111111111111_1111111111111111_1111000110100010_1100011100101000"; -- -0.056109955418416964
	pesos_i(6586) := b"0000000000000000_0000000000000000_0001011110100011_1111101111100100"; -- 0.09234594638876781
	pesos_i(6587) := b"1111111111111111_1111111111111111_1111100001111100_0110010011110110"; -- -0.029351892335806044
	pesos_i(6588) := b"1111111111111111_1111111111111111_1110011000011010_1010111100010101"; -- -0.10115533576536896
	pesos_i(6589) := b"1111111111111111_1111111111111111_1111100000010001_1100011001111100"; -- -0.03097877009336805
	pesos_i(6590) := b"1111111111111111_1111111111111111_1110110010000000_0010100011001101"; -- -0.07616944303627352
	pesos_i(6591) := b"1111111111111111_1111111111111111_1110110010111111_1110110010110001"; -- -0.07519646327677239
	pesos_i(6592) := b"0000000000000000_0000000000000000_0010110001010110_1000111000000010"; -- 0.17319572009267223
	pesos_i(6593) := b"1111111111111111_1111111111111111_1101001110000010_1001010001111000"; -- -0.1737887579291752
	pesos_i(6594) := b"1111111111111111_1111111111111111_1101011101001111_0010011101010010"; -- -0.15894846198921644
	pesos_i(6595) := b"0000000000000000_0000000000000000_0001001001111111_1110100010111100"; -- 0.0722642383289405
	pesos_i(6596) := b"0000000000000000_0000000000000000_0001110000100100_0010111011111010"; -- 0.10992711642040093
	pesos_i(6597) := b"0000000000000000_0000000000000000_0000011010010111_1111011001100111"; -- 0.025756263824410663
	pesos_i(6598) := b"0000000000000000_0000000000000000_0001101011011110_1110111011011011"; -- 0.1049641880338476
	pesos_i(6599) := b"1111111111111111_1111111111111111_1111001100101000_0100111100101010"; -- -0.050166179913438136
	pesos_i(6600) := b"1111111111111111_1111111111111111_1110001100100101_1001000000010100"; -- -0.1127080871695684
	pesos_i(6601) := b"1111111111111111_1111111111111111_1110101001100101_1101110110110100"; -- -0.08438314778093538
	pesos_i(6602) := b"0000000000000000_0000000000000000_0000100101101110_1000011100110111"; -- 0.036842776152998795
	pesos_i(6603) := b"1111111111111111_1111111111111111_1101001110110101_1011101011110010"; -- -0.17300826630760435
	pesos_i(6604) := b"1111111111111111_1111111111111111_1111101110000100_1001010101110001"; -- -0.017508182515066226
	pesos_i(6605) := b"1111111111111111_1111111111111111_1110011100100110_0101010111110101"; -- -0.09707129264533863
	pesos_i(6606) := b"1111111111111111_1111111111111111_1111101001111101_0110111001101001"; -- -0.0215235705234785
	pesos_i(6607) := b"0000000000000000_0000000000000000_0010111101110101_1010110111111110"; -- 0.18538939901258455
	pesos_i(6608) := b"1111111111111111_1111111111111111_1111110001100111_1100101000111000"; -- -0.014041291547749649
	pesos_i(6609) := b"0000000000000000_0000000000000000_0011000100101111_0111011111101011"; -- 0.19213056069148068
	pesos_i(6610) := b"0000000000000000_0000000000000000_0011010100111011_1011111011101100"; -- 0.20794289841125363
	pesos_i(6611) := b"0000000000000000_0000000000000000_0000000111111100_1111101010011111"; -- 0.007766403087451259
	pesos_i(6612) := b"1111111111111111_1111111111111111_1101010111100100_0011100010111010"; -- -0.16448636489285728
	pesos_i(6613) := b"0000000000000000_0000000000000000_0011000001001011_1100111000001101"; -- 0.18865669079281663
	pesos_i(6614) := b"1111111111111111_1111111111111111_1101000010001001_0101000010001101"; -- -0.1854047446336157
	pesos_i(6615) := b"0000000000000000_0000000000000000_0011010010010010_1011001001110001"; -- 0.20536341922501428
	pesos_i(6616) := b"0000000000000000_0000000000000000_0011000011001111_1011100010110011"; -- 0.19066957828052203
	pesos_i(6617) := b"0000000000000000_0000000000000000_0001101000101101_1100110001010111"; -- 0.10226132506488866
	pesos_i(6618) := b"1111111111111111_1111111111111111_1101101111011100_0011111110100001"; -- -0.14117052377574923
	pesos_i(6619) := b"1111111111111111_1111111111111111_1111110010000001_0100010010111000"; -- -0.013652520196340069
	pesos_i(6620) := b"0000000000000000_0000000000000000_0001101001011001_1001101011000000"; -- 0.10292975595248816
	pesos_i(6621) := b"1111111111111111_1111111111111111_1101010001001100_1010000110111100"; -- -0.17070569181261253
	pesos_i(6622) := b"1111111111111111_1111111111111111_1110100011011010_0001110010010100"; -- -0.09042188055567751
	pesos_i(6623) := b"1111111111111111_1111111111111111_1111001010110010_1101110110001100"; -- -0.051958230440319914
	pesos_i(6624) := b"1111111111111111_1111111111111111_1111000100111000_1101101010101111"; -- -0.05772622334647656
	pesos_i(6625) := b"0000000000000000_0000000000000000_0010111011100010_1001110110000000"; -- 0.18314537395865987
	pesos_i(6626) := b"1111111111111111_1111111111111111_1100110001001101_0110001010001011"; -- -0.20194419970882313
	pesos_i(6627) := b"1111111111111111_1111111111111111_1101100010100110_1000011100000110"; -- -0.1537089930873481
	pesos_i(6628) := b"1111111111111111_1111111111111111_1101101110100100_1101010100110111"; -- -0.14201610004932913
	pesos_i(6629) := b"1111111111111111_1111111111111111_1100111111110100_0001010111101100"; -- -0.18768179887701944
	pesos_i(6630) := b"1111111111111111_1111111111111111_1111011000100101_1111111001010110"; -- -0.03848276512232177
	pesos_i(6631) := b"1111111111111111_1111111111111111_1111110010001000_0101101001110001"; -- -0.013544413985240821
	pesos_i(6632) := b"1111111111111111_1111111111111111_1111011101011000_1101001011001010"; -- -0.03380091245033492
	pesos_i(6633) := b"1111111111111111_1111111111111111_1101100110001111_1010000010110010"; -- -0.1501521649353812
	pesos_i(6634) := b"0000000000000000_0000000000000000_0001000100110110_1100101101110011"; -- 0.06724235105699113
	pesos_i(6635) := b"0000000000000000_0000000000000000_0010000110100011_1001011101010001"; -- 0.13140245179038412
	pesos_i(6636) := b"1111111111111111_1111111111111111_1101011001000010_1001000010001101"; -- -0.16304680403379795
	pesos_i(6637) := b"1111111111111111_1111111111111111_1111001111110011_1110100100110001"; -- -0.04705946492406842
	pesos_i(6638) := b"0000000000000000_0000000000000000_0000101101110101_0101111000100001"; -- 0.04475963882766624
	pesos_i(6639) := b"1111111111111111_1111111111111111_1110110001111101_0001011110011111"; -- -0.07621624350984436
	pesos_i(6640) := b"1111111111111111_1111111111111111_1100100101111100_1110101010000111"; -- -0.21293768114729367
	pesos_i(6641) := b"1111111111111111_1111111111111111_1100101010100001_1001011000001001"; -- -0.20847189217003995
	pesos_i(6642) := b"0000000000000000_0000000000000000_0000100011111100_1010101011011111"; -- 0.035105399561360356
	pesos_i(6643) := b"0000000000000000_0000000000000000_0010101010101110_1100000001101101"; -- 0.16672899887615186
	pesos_i(6644) := b"1111111111111111_1111111111111111_1101001010101100_1000000000110100"; -- -0.1770553467147262
	pesos_i(6645) := b"1111111111111111_1111111111111111_1111111000111101_0010010010110100"; -- -0.006879526251458313
	pesos_i(6646) := b"0000000000000000_0000000000000000_0000001101001011_1100011110011110"; -- 0.012875057367329315
	pesos_i(6647) := b"1111111111111111_1111111111111111_1111000111000000_0011111101000100"; -- -0.05566029163887053
	pesos_i(6648) := b"0000000000000000_0000000000000000_0000000011100000_1011001010100010"; -- 0.0034286160404762627
	pesos_i(6649) := b"1111111111111111_1111111111111111_1110011110000010_0101110110000010"; -- -0.09566703400378744
	pesos_i(6650) := b"1111111111111111_1111111111111111_1101111100101100_0010000100101100"; -- -0.12823288619806789
	pesos_i(6651) := b"0000000000000000_0000000000000000_0000010001101010_1000100011001001"; -- 0.01725058473503988
	pesos_i(6652) := b"0000000000000000_0000000000000000_0001111100001101_0110111100001001"; -- 0.12129873244515861
	pesos_i(6653) := b"1111111111111111_1111111111111111_1111111101100100_0100011011101011"; -- -0.0023761440100550507
	pesos_i(6654) := b"1111111111111111_1111111111111111_1110000001011111_1000110000111100"; -- -0.12354205644527971
	pesos_i(6655) := b"0000000000000000_0000000000000000_0011110110101111_0111011111100001"; -- 0.24095868336021573
	pesos_i(6656) := b"1111111111111111_1111111111111111_1111000100010101_0101110111000111"; -- -0.05826772597167126
	pesos_i(6657) := b"0000000000000000_0000000000000000_0000100101111101_0010110110101010"; -- 0.037066320351779716
	pesos_i(6658) := b"0000000000000000_0000000000000000_0010100110011110_1011101000001110"; -- 0.16257822838918862
	pesos_i(6659) := b"1111111111111111_1111111111111111_1101001011100100_0000101011010100"; -- -0.1762078507843518
	pesos_i(6660) := b"0000000000000000_0000000000000000_0000010100110100_1110011100010001"; -- 0.02033847956417917
	pesos_i(6661) := b"1111111111111111_1111111111111111_1101101000101111_1111011001001101"; -- -0.14770565616228035
	pesos_i(6662) := b"1111111111111111_1111111111111111_1100110001111101_0000101110010001"; -- -0.20121696201138295
	pesos_i(6663) := b"0000000000000000_0000000000000000_0010100000010111_1101101010101011"; -- 0.1566139857515831
	pesos_i(6664) := b"0000000000000000_0000000000000000_0010011110100011_1010001111010000"; -- 0.15484069659961716
	pesos_i(6665) := b"1111111111111111_1111111111111111_1110011010011010_0101110010100101"; -- -0.09920712449654892
	pesos_i(6666) := b"1111111111111111_1111111111111111_1111100000000011_0011101011110010"; -- -0.031200710220910054
	pesos_i(6667) := b"1111111111111111_1111111111111111_1101100110100111_0011111010111101"; -- -0.14979179265588502
	pesos_i(6668) := b"0000000000000000_0000000000000000_0000001011111001_1101110111100111"; -- 0.011625164874275482
	pesos_i(6669) := b"0000000000000000_0000000000000000_0000010111100000_1111011101110001"; -- 0.022963967319771315
	pesos_i(6670) := b"1111111111111111_1111111111111111_1101011010010000_1011110001011010"; -- -0.1618540076741481
	pesos_i(6671) := b"0000000000000000_0000000000000000_0001000011010110_1011001010110101"; -- 0.06577603253138832
	pesos_i(6672) := b"0000000000000000_0000000000000000_0011011110100110_1011110001010101"; -- 0.21738793447939375
	pesos_i(6673) := b"1111111111111111_1111111111111111_1110010110111111_1111101110001111"; -- -0.10253932726314126
	pesos_i(6674) := b"0000000000000000_0000000000000000_0001100000010011_0000111100011101"; -- 0.0940408178717443
	pesos_i(6675) := b"0000000000000000_0000000000000000_0000111000011111_0010110101011100"; -- 0.0551632260711078
	pesos_i(6676) := b"0000000000000000_0000000000000000_0000111111100000_0110011010011000"; -- 0.06201783372328884
	pesos_i(6677) := b"1111111111111111_1111111111111111_1101010110100110_0101101000111111"; -- -0.16543041185254892
	pesos_i(6678) := b"0000000000000000_0000000000000000_0000010001000010_0011011100110000"; -- 0.016635369418056125
	pesos_i(6679) := b"0000000000000000_0000000000000000_0001101111100110_1100011000111101"; -- 0.1089900873316548
	pesos_i(6680) := b"0000000000000000_0000000000000000_0010000000010000_1111101100101111"; -- 0.1252591122778164
	pesos_i(6681) := b"1111111111111111_1111111111111111_1110100001001101_1011111111000010"; -- -0.09256364365661111
	pesos_i(6682) := b"0000000000000000_0000000000000000_0001101001000100_0100111000100110"; -- 0.102604755748417
	pesos_i(6683) := b"0000000000000000_0000000000000000_0001000101000000_0011111110001011"; -- 0.06738660003031602
	pesos_i(6684) := b"1111111111111111_1111111111111111_1111001110110110_1101000100001000"; -- -0.04799169106023596
	pesos_i(6685) := b"0000000000000000_0000000000000000_0010001011100111_1010110011001101"; -- 0.1363475799140367
	pesos_i(6686) := b"0000000000000000_0000000000000000_0001000101101111_1010110000101001"; -- 0.06811023720411807
	pesos_i(6687) := b"0000000000000000_0000000000000000_0001110101101111_1011000111101000"; -- 0.11498557961496018
	pesos_i(6688) := b"1111111111111111_1111111111111111_1101001111101000_0001110001101101"; -- -0.17223951670919366
	pesos_i(6689) := b"1111111111111111_1111111111111111_1111100100011011_0101011110110001"; -- -0.026926535829863887
	pesos_i(6690) := b"0000000000000000_0000000000000000_0001110010000100_0001110000000110"; -- 0.11139083050552832
	pesos_i(6691) := b"0000000000000000_0000000000000000_0011001100010011_0010110011100110"; -- 0.19951134319241703
	pesos_i(6692) := b"0000000000000000_0000000000000000_0000010101111111_1111001000011011"; -- 0.021483546855598425
	pesos_i(6693) := b"1111111111111111_1111111111111111_1110011111100111_1101011110011000"; -- -0.09411861936686304
	pesos_i(6694) := b"1111111111111111_1111111111111111_1110111010011011_0101110011000011"; -- -0.06794185860285783
	pesos_i(6695) := b"1111111111111111_1111111111111111_1110111010000101_1101100100100011"; -- -0.06827013880421386
	pesos_i(6696) := b"1111111111111111_1111111111111111_1110100001010111_0011010011010011"; -- -0.09241933678541737
	pesos_i(6697) := b"1111111111111111_1111111111111111_1111111011001100_0101110100111000"; -- -0.004694150796491075
	pesos_i(6698) := b"1111111111111111_1111111111111111_1111111100010111_1100101001100010"; -- -0.0035432348771272672
	pesos_i(6699) := b"1111111111111111_1111111111111111_1110011011001000_0110011111000001"; -- -0.09850455799025758
	pesos_i(6700) := b"0000000000000000_0000000000000000_0001110111011111_0000101101110011"; -- 0.11668464249944932
	pesos_i(6701) := b"0000000000000000_0000000000000000_0000110110010111_0011001000010010"; -- 0.05308831165745617
	pesos_i(6702) := b"1111111111111111_1111111111111111_1100011011100101_1110100001011101"; -- -0.2230543874019338
	pesos_i(6703) := b"0000000000000000_0000000000000000_0011101110100000_0011110101111001"; -- 0.23291382040812997
	pesos_i(6704) := b"0000000000000000_0000000000000000_0001101010000010_1000101101010110"; -- 0.10355444776181019
	pesos_i(6705) := b"0000000000000000_0000000000000000_0001111110011001_0000111010011011"; -- 0.12342921519636281
	pesos_i(6706) := b"0000000000000000_0000000000000000_0000100010100000_1001010011110010"; -- 0.03370028397330647
	pesos_i(6707) := b"0000000000000000_0000000000000000_0010011000110010_1000000101001111"; -- 0.14920814691270423
	pesos_i(6708) := b"0000000000000000_0000000000000000_0010010110111100_1001100101010110"; -- 0.14740904184118342
	pesos_i(6709) := b"1111111111111111_1111111111111111_1100101010010101_0011011011111101"; -- -0.20866066278363787
	pesos_i(6710) := b"0000000000000000_0000000000000000_0010011111110100_0100101100101100"; -- 0.1560713751642982
	pesos_i(6711) := b"1111111111111111_1111111111111111_1101110011001011_1111001011011010"; -- -0.13751299070044437
	pesos_i(6712) := b"0000000000000000_0000000000000000_0001100111111110_0001000101010011"; -- 0.1015330149252121
	pesos_i(6713) := b"1111111111111111_1111111111111111_1111110101010010_0111001000000011"; -- -0.010460733667899832
	pesos_i(6714) := b"0000000000000000_0000000000000000_0011100001110001_1010000001100010"; -- 0.2204838026446964
	pesos_i(6715) := b"0000000000000000_0000000000000000_0000000001100111_1100001011010100"; -- 0.0015832678516329482
	pesos_i(6716) := b"0000000000000000_0000000000000000_0000001000110111_1111100111011001"; -- 0.008666625522851567
	pesos_i(6717) := b"1111111111111111_1111111111111111_1111011000011111_0000100011010011"; -- -0.03858895146007166
	pesos_i(6718) := b"0000000000000000_0000000000000000_0010100110111100_1010000001001100"; -- 0.1630344567457525
	pesos_i(6719) := b"1111111111111111_1111111111111111_1101011100101011_1000101101001000"; -- -0.15949182037334242
	pesos_i(6720) := b"1111111111111111_1111111111111111_1110000011110001_0011111011101010"; -- -0.12131888174936521
	pesos_i(6721) := b"0000000000000000_0000000000000000_0010011001110000_1100000010110110"; -- 0.1501579709101427
	pesos_i(6722) := b"1111111111111111_1111111111111111_1101101000010111_0100110111001111"; -- -0.14808191008242777
	pesos_i(6723) := b"1111111111111111_1111111111111111_1110000101000110_0101111101010101"; -- -0.12001995261240576
	pesos_i(6724) := b"0000000000000000_0000000000000000_0001010010101110_1010110111100011"; -- 0.08079039377973873
	pesos_i(6725) := b"1111111111111111_1111111111111111_1110001101000001_0111110111111010"; -- -0.11228191983716809
	pesos_i(6726) := b"0000000000000000_0000000000000000_0010001011010101_1111100100010101"; -- 0.1360774684546965
	pesos_i(6727) := b"1111111111111111_1111111111111111_1111110000111100_0001010001111001"; -- -0.01470825235783803
	pesos_i(6728) := b"0000000000000000_0000000000000000_0010100011110110_0100110110111000"; -- 0.16000829454345658
	pesos_i(6729) := b"1111111111111111_1111111111111111_1101000001001010_0001101100111011"; -- -0.18636922653541316
	pesos_i(6730) := b"1111111111111111_1111111111111111_1101101010110100_1011010011101011"; -- -0.14568013433963842
	pesos_i(6731) := b"0000000000000000_0000000000000000_0000010010111111_0101100010000000"; -- 0.018544703740923783
	pesos_i(6732) := b"1111111111111111_1111111111111111_1110000110011010_0101110010000010"; -- -0.11873838264769172
	pesos_i(6733) := b"1111111111111111_1111111111111111_1111101010101100_0101110000000001"; -- -0.02080750437251364
	pesos_i(6734) := b"1111111111111111_1111111111111111_1111110000110101_0110100110000110"; -- -0.014809994541793626
	pesos_i(6735) := b"1111111111111111_1111111111111111_1111001101100010_0010011000000101"; -- -0.04928362246647809
	pesos_i(6736) := b"1111111111111111_1111111111111111_1111110000010010_0100111101001000"; -- -0.015345616245408129
	pesos_i(6737) := b"1111111111111111_1111111111111111_1100011001100101_0110000001111010"; -- -0.22501561177903334
	pesos_i(6738) := b"1111111111111111_1111111111111111_1111111001110000_1111011111001101"; -- -0.0060887454349091135
	pesos_i(6739) := b"1111111111111111_1111111111111111_1101101001110000_1110110101111011"; -- -0.14671436075127384
	pesos_i(6740) := b"1111111111111111_1111111111111111_1110011000100100_1000010001110100"; -- -0.10100528875214658
	pesos_i(6741) := b"0000000000000000_0000000000000000_0000001101010010_1111101101011000"; -- 0.01298495189292392
	pesos_i(6742) := b"1111111111111111_1111111111111111_1111110100001010_1111000110000110"; -- -0.01155176622933971
	pesos_i(6743) := b"1111111111111111_1111111111111111_1101110100010110_0011111010001111"; -- -0.1363793278338109
	pesos_i(6744) := b"0000000000000000_0000000000000000_0001001001100110_1111001001110011"; -- 0.07188334766287229
	pesos_i(6745) := b"0000000000000000_0000000000000000_0001011011000001_1101000011101000"; -- 0.08889489812099904
	pesos_i(6746) := b"1111111111111111_1111111111111111_1110011111110011_0011101100110101"; -- -0.09394483521653062
	pesos_i(6747) := b"0000000000000000_0000000000000000_0011001000011111_1001110100100010"; -- 0.19579488834418138
	pesos_i(6748) := b"0000000000000000_0000000000000000_0000000010101000_0101100001101100"; -- 0.0025687470030953314
	pesos_i(6749) := b"1111111111111111_1111111111111111_1110000011100011_0110110000111001"; -- -0.12152980419517269
	pesos_i(6750) := b"0000000000000000_0000000000000000_0001110010011000_1010000000101001"; -- 0.11170388219179743
	pesos_i(6751) := b"1111111111111111_1111111111111111_1101100000101110_0110001010001001"; -- -0.1555422225738988
	pesos_i(6752) := b"1111111111111111_1111111111111111_1101001011001011_1100011101101011"; -- -0.17657807952347646
	pesos_i(6753) := b"0000000000000000_0000000000000000_0010000100101110_0000010011000110"; -- 0.12960843883631062
	pesos_i(6754) := b"0000000000000000_0000000000000000_0000100101011000_1011010010101000"; -- 0.03650979137571513
	pesos_i(6755) := b"0000000000000000_0000000000000000_0011011011011111_1110011111100010"; -- 0.2143540312831122
	pesos_i(6756) := b"1111111111111111_1111111111111111_1110001101100101_1100001010000110"; -- -0.11172851777175724
	pesos_i(6757) := b"0000000000000000_0000000000000000_0000100000010000_1011001101101010"; -- 0.03150483447437796
	pesos_i(6758) := b"1111111111111111_1111111111111111_1110010100101000_0010111100110010"; -- -0.1048555854030095
	pesos_i(6759) := b"0000000000000000_0000000000000000_0001111010000010_1010111100001111"; -- 0.1191815768150464
	pesos_i(6760) := b"1111111111111111_1111111111111111_1111101111000000_0000100110011010"; -- -0.016600990238814874
	pesos_i(6761) := b"1111111111111111_1111111111111111_1101011111000111_1110000101100000"; -- -0.15710631748983192
	pesos_i(6762) := b"0000000000000000_0000000000000000_0001010100010111_1100100011110111"; -- 0.08239418058047548
	pesos_i(6763) := b"0000000000000000_0000000000000000_0000100111011100_1110101101010001"; -- 0.038527209530362004
	pesos_i(6764) := b"1111111111111111_1111111111111111_1110001111111011_1111111110001101"; -- -0.10943606186833263
	pesos_i(6765) := b"1111111111111111_1111111111111111_1110110101100100_1001000110101101"; -- -0.07268418815514796
	pesos_i(6766) := b"1111111111111111_1111111111111111_1111110011001101_1010011100011111"; -- -0.012486986966325468
	pesos_i(6767) := b"0000000000000000_0000000000000000_0000001100011101_0110000110111010"; -- 0.012167079782097074
	pesos_i(6768) := b"1111111111111111_1111111111111111_1111001100001001_0000011010010100"; -- -0.05064352892396101
	pesos_i(6769) := b"1111111111111111_1111111111111111_1111011111111000_0000100100001000"; -- -0.0313715319686529
	pesos_i(6770) := b"1111111111111111_1111111111111111_1101111010011110_1110110111010000"; -- -0.13038743656216584
	pesos_i(6771) := b"1111111111111111_1111111111111111_1110001111100011_0111001000100101"; -- -0.1098107012803107
	pesos_i(6772) := b"1111111111111111_1111111111111111_1110100101000011_0111001010010100"; -- -0.08881458176372296
	pesos_i(6773) := b"1111111111111111_1111111111111111_1110001010111001_0101001010110110"; -- -0.11435969406586918
	pesos_i(6774) := b"1111111111111111_1111111111111111_1110100011101100_0111001010000101"; -- -0.09014209991015008
	pesos_i(6775) := b"1111111111111111_1111111111111111_1101001001010110_0000010000010000"; -- -0.17837500209654217
	pesos_i(6776) := b"1111111111111111_1111111111111111_1110110101011110_1101101011001100"; -- -0.07277138257054964
	pesos_i(6777) := b"1111111111111111_1111111111111111_1110101010101101_1011110100101000"; -- -0.08328645495351693
	pesos_i(6778) := b"0000000000000000_0000000000000000_0010000011011000_0100101110101001"; -- 0.12830040809828575
	pesos_i(6779) := b"1111111111111111_1111111111111111_1101100111000101_0101110100101100"; -- -0.14933221507803338
	pesos_i(6780) := b"0000000000000000_0000000000000000_0010100110100111_0010110011111001"; -- 0.16270714836865738
	pesos_i(6781) := b"1111111111111111_1111111111111111_1110101101111111_1100110111010011"; -- -0.08008111564529481
	pesos_i(6782) := b"0000000000000000_0000000000000000_0010001111110100_1010101000000100"; -- 0.14045202832795278
	pesos_i(6783) := b"0000000000000000_0000000000000000_0001101110000011_0111110011100111"; -- 0.10747509617566135
	pesos_i(6784) := b"0000000000000000_0000000000000000_0001101010001000_1101011011001100"; -- 0.10365049822992149
	pesos_i(6785) := b"0000000000000000_0000000000000000_0000110000101110_1010011010011010"; -- 0.04758683443674266
	pesos_i(6786) := b"0000000000000000_0000000000000000_0010001101101010_1011011111010001"; -- 0.13834713794090783
	pesos_i(6787) := b"1111111111111111_1111111111111111_1110011111110110_0100011100010111"; -- -0.09389835063735492
	pesos_i(6788) := b"0000000000000000_0000000000000000_0000001010110101_1111000101101010"; -- 0.01058873031000266
	pesos_i(6789) := b"0000000000000000_0000000000000000_0001101111001111_0100100100011001"; -- 0.10863167641046713
	pesos_i(6790) := b"1111111111111111_1111111111111111_1111011000000000_1110001111010110"; -- -0.03904891981840864
	pesos_i(6791) := b"0000000000000000_0000000000000000_0010011010111110_0000010110001100"; -- 0.1513370004490123
	pesos_i(6792) := b"1111111111111111_1111111111111111_1110111011000000_1000100000101110"; -- -0.0673746954478755
	pesos_i(6793) := b"1111111111111111_1111111111111111_1101011001011000_0101001010001111"; -- -0.1627148056012988
	pesos_i(6794) := b"0000000000000000_0000000000000000_0010101011001111_1110100101111000"; -- 0.16723498504501239
	pesos_i(6795) := b"1111111111111111_1111111111111111_1101001110111110_1000100000111111"; -- -0.17287395909170836
	pesos_i(6796) := b"0000000000000000_0000000000000000_0001010001010100_0011110001011010"; -- 0.07941033555444145
	pesos_i(6797) := b"0000000000000000_0000000000000000_0010001001010101_1110111000010101"; -- 0.13412368780727643
	pesos_i(6798) := b"1111111111111111_1111111111111111_1101000010001101_0111001110000110"; -- -0.1853416250659978
	pesos_i(6799) := b"1111111111111111_1111111111111111_1101100111101110_0110010110001010"; -- -0.14870610594447103
	pesos_i(6800) := b"0000000000000000_0000000000000000_0001010111000010_1111101000001110"; -- 0.08500635945916668
	pesos_i(6801) := b"0000000000000000_0000000000000000_0000111000010011_1001001110100000"; -- 0.05498621622845252
	pesos_i(6802) := b"0000000000000000_0000000000000000_0001110110101000_1010101100011111"; -- 0.11585492613284919
	pesos_i(6803) := b"0000000000000000_0000000000000000_0000000001111101_0001011010101101"; -- 0.0019087002433662722
	pesos_i(6804) := b"0000000000000000_0000000000000000_0000001110100101_0011101011110111"; -- 0.014239964732938653
	pesos_i(6805) := b"1111111111111111_1111111111111111_1110101001011001_0001000000101100"; -- -0.08457850395266396
	pesos_i(6806) := b"0000000000000000_0000000000000000_0001000101110101_1001001111010100"; -- 0.06820033957205124
	pesos_i(6807) := b"1111111111111111_1111111111111111_1111000100010111_0001100111110000"; -- -0.05824125180862417
	pesos_i(6808) := b"1111111111111111_1111111111111111_1101111100011111_1110101000001101"; -- -0.1284192769906065
	pesos_i(6809) := b"0000000000000000_0000000000000000_0010001110101010_0100100111100010"; -- 0.13931714788647412
	pesos_i(6810) := b"1111111111111111_1111111111111111_1110111010000000_1101100111010101"; -- -0.06834639113467939
	pesos_i(6811) := b"0000000000000000_0000000000000000_0010101101111100_1111101111101000"; -- 0.16987585464632168
	pesos_i(6812) := b"0000000000000000_0000000000000000_0010000010001001_0111100001001101"; -- 0.12709762467434307
	pesos_i(6813) := b"0000000000000000_0000000000000000_0000110101000010_0110101110101111"; -- 0.05179474848394687
	pesos_i(6814) := b"1111111111111111_1111111111111111_1101110110101011_1000110110101110"; -- -0.1341010521900134
	pesos_i(6815) := b"0000000000000000_0000000000000000_0001001001010110_0001111100111100"; -- 0.07162661754732462
	pesos_i(6816) := b"1111111111111111_1111111111111111_1111000100110100_0000110100110001"; -- -0.057799506592920796
	pesos_i(6817) := b"1111111111111111_1111111111111111_1111010010111100_1001001010011110"; -- -0.04399760863257368
	pesos_i(6818) := b"1111111111111111_1111111111111111_1101010001111010_1011101100001011"; -- -0.17000227899730336
	pesos_i(6819) := b"1111111111111111_1111111111111111_1100111010100100_1010111010000010"; -- -0.19279965717290923
	pesos_i(6820) := b"1111111111111111_1111111111111111_1110101010010110_0110010010110100"; -- -0.08364267919038959
	pesos_i(6821) := b"0000000000000000_0000000000000000_0010010010010111_1101100110010100"; -- 0.1429420457442484
	pesos_i(6822) := b"1111111111111111_1111111111111111_1110101000001111_1001000111001010"; -- -0.08569992854510111
	pesos_i(6823) := b"0000000000000000_0000000000000000_0001100111101110_0101111011001110"; -- 0.10129349256779474
	pesos_i(6824) := b"1111111111111111_1111111111111111_1100111100110011_0011100100101111"; -- -0.19062464342313318
	pesos_i(6825) := b"0000000000000000_0000000000000000_0001011011101000_0100001001100001"; -- 0.08948149560007695
	pesos_i(6826) := b"0000000000000000_0000000000000000_0011101100001011_1011011000101001"; -- 0.23064745438555712
	pesos_i(6827) := b"1111111111111111_1111111111111111_1101101011110001_1010100011010100"; -- -0.14475006892963424
	pesos_i(6828) := b"1111111111111111_1111111111111111_1111111101111111_1000110111011001"; -- -0.0019599290669641833
	pesos_i(6829) := b"0000000000000000_0000000000000000_0001100011110011_0001111111110010"; -- 0.09745978979133935
	pesos_i(6830) := b"1111111111111111_1111111111111111_1110100110010001_0111111110010110"; -- -0.08762362077277916
	pesos_i(6831) := b"0000000000000000_0000000000000000_0001011001010110_1010010011110110"; -- 0.08725958826028378
	pesos_i(6832) := b"0000000000000000_0000000000000000_0000100100010000_0011111011001111"; -- 0.03540413436046622
	pesos_i(6833) := b"1111111111111111_1111111111111111_1111111100101101_1101100000110011"; -- -0.003206717946932315
	pesos_i(6834) := b"1111111111111111_1111111111111111_1101001100010000_1000010100111011"; -- -0.17552916816017214
	pesos_i(6835) := b"0000000000000000_0000000000000000_0000011011101100_0010100100001110"; -- 0.027041021258827607
	pesos_i(6836) := b"0000000000000000_0000000000000000_0010011000000110_1110100010110101"; -- 0.1485429231785247
	pesos_i(6837) := b"1111111111111111_1111111111111111_1110010010100000_1101010110101010"; -- -0.10692085849516374
	pesos_i(6838) := b"0000000000000000_0000000000000000_0000110110010010_0011111010111010"; -- 0.05301277192949417
	pesos_i(6839) := b"1111111111111111_1111111111111111_1110101110101010_0111100001101101"; -- -0.07943007802104388
	pesos_i(6840) := b"0000000000000000_0000000000000000_0010000111100100_0101001011011011"; -- 0.13239019242396455
	pesos_i(6841) := b"0000000000000000_0000000000000000_0000001111110011_1111100001111001"; -- 0.015441445948456986
	pesos_i(6842) := b"0000000000000000_0000000000000000_0000110001101000_1110101101000101"; -- 0.048475937141869485
	pesos_i(6843) := b"1111111111111111_1111111111111111_1111101011011001_1010000011001011"; -- -0.020116758719188787
	pesos_i(6844) := b"1111111111111111_1111111111111111_1111111110110100_1001000001001101"; -- -0.0011510670145234683
	pesos_i(6845) := b"1111111111111111_1111111111111111_1111110100101111_0101010100111111"; -- -0.010996505826662503
	pesos_i(6846) := b"1111111111111111_1111111111111111_1101100001100010_0010110100110100"; -- -0.15475194424394176
	pesos_i(6847) := b"0000000000000000_0000000000000000_0010000000111011_1011110111000110"; -- 0.12591157984297183
	pesos_i(6848) := b"1111111111111111_1111111111111111_1101110101111101_1001000110111100"; -- -0.1348027148836201
	pesos_i(6849) := b"1111111111111111_1111111111111111_1101010010100111_1100000111110110"; -- -0.16931522117018077
	pesos_i(6850) := b"0000000000000000_0000000000000000_0000111110001111_0111010111011101"; -- 0.06078278206071949
	pesos_i(6851) := b"1111111111111111_1111111111111111_1110101001111011_1101001100011101"; -- -0.0840480856622028
	pesos_i(6852) := b"0000000000000000_0000000000000000_0001001111010011_1000101110011110"; -- 0.07744667626488805
	pesos_i(6853) := b"0000000000000000_0000000000000000_0001100110110111_0010011100111001"; -- 0.10045094629521253
	pesos_i(6854) := b"0000000000000000_0000000000000000_0001111000111010_0011010101001010"; -- 0.11807568605332136
	pesos_i(6855) := b"1111111111111111_1111111111111111_1111100111010010_0010001111100101"; -- -0.024137264837234343
	pesos_i(6856) := b"1111111111111111_1111111111111111_1111101011011000_1000010000100000"; -- -0.02013372626077511
	pesos_i(6857) := b"0000000000000000_0000000000000000_0000011111011110_0001110101101010"; -- 0.0307329544730855
	pesos_i(6858) := b"1111111111111111_1111111111111111_1111110101001011_1000100001011001"; -- -0.010566213915972218
	pesos_i(6859) := b"1111111111111111_1111111111111111_1101110101001111_0111111000000110"; -- -0.1355057940496184
	pesos_i(6860) := b"1111111111111111_1111111111111111_1101000110010100_1011010110011110"; -- -0.18132462405327074
	pesos_i(6861) := b"0000000000000000_0000000000000000_0000111101110100_1010100010110111"; -- 0.06037382562265111
	pesos_i(6862) := b"1111111111111111_1111111111111111_1110110110000101_1111101110011100"; -- -0.07217433386011067
	pesos_i(6863) := b"1111111111111111_1111111111111111_1110110011100011_0001111001010101"; -- -0.07465944702325461
	pesos_i(6864) := b"1111111111111111_1111111111111111_1101010010110001_0011110100100011"; -- -0.16917055027360417
	pesos_i(6865) := b"0000000000000000_0000000000000000_0001001001001100_1010101011011011"; -- 0.07148235184330469
	pesos_i(6866) := b"1111111111111111_1111111111111111_1110110000010110_0101111110010001"; -- -0.07778361032876006
	pesos_i(6867) := b"1111111111111111_1111111111111111_1110001101000010_0110001011110100"; -- -0.11226827194899308
	pesos_i(6868) := b"0000000000000000_0000000000000000_0001011100001000_0110111101010011"; -- 0.0899724556935785
	pesos_i(6869) := b"1111111111111111_1111111111111111_1100110101111101_0110011011100000"; -- -0.1973052695470454
	pesos_i(6870) := b"0000000000000000_0000000000000000_0001011001110101_1110011001010000"; -- 0.08773650598030816
	pesos_i(6871) := b"0000000000000000_0000000000000000_0001000010100000_0100100010000100"; -- 0.06494572842401253
	pesos_i(6872) := b"0000000000000000_0000000000000000_0001000101111100_0010101101100100"; -- 0.06830092615975816
	pesos_i(6873) := b"0000000000000000_0000000000000000_0011110110001100_0100110010010101"; -- 0.24042204501365505
	pesos_i(6874) := b"0000000000000000_0000000000000000_0001111111101010_0111101001111110"; -- 0.12467160776812576
	pesos_i(6875) := b"1111111111111111_1111111111111111_1101011101000110_0010010000001011"; -- -0.1590859863672124
	pesos_i(6876) := b"0000000000000000_0000000000000000_0010101101110001_1111100101011101"; -- 0.1697078564710339
	pesos_i(6877) := b"0000000000000000_0000000000000000_0001111100101011_1000011101110010"; -- 0.12175795117701767
	pesos_i(6878) := b"1111111111111111_1111111111111111_1101100110001100_1101101110110011"; -- -0.15019442446656053
	pesos_i(6879) := b"1111111111111111_1111111111111111_1110000101010100_0001001101110110"; -- -0.11981085170950896
	pesos_i(6880) := b"1111111111111111_1111111111111111_1111100110100110_0110011101110001"; -- -0.02480462546736663
	pesos_i(6881) := b"1111111111111111_1111111111111111_1101110110111011_1101001101100011"; -- -0.13385275676909567
	pesos_i(6882) := b"1111111111111111_1111111111111111_1100110101111011_1010111000111011"; -- -0.1973315340835273
	pesos_i(6883) := b"1111111111111111_1111111111111111_1101001011000111_0011100101000101"; -- -0.1766475875063511
	pesos_i(6884) := b"1111111111111111_1111111111111111_1111111101111000_0110101001010101"; -- -0.002068857446838491
	pesos_i(6885) := b"1111111111111111_1111111111111111_1110111110100110_1000011011111010"; -- -0.063865245721319
	pesos_i(6886) := b"1111111111111111_1111111111111111_1101000101001101_0000111111111101"; -- -0.18241787037384216
	pesos_i(6887) := b"0000000000000000_0000000000000000_0010100110111110_1111001000010110"; -- 0.1630698493704435
	pesos_i(6888) := b"0000000000000000_0000000000000000_0010000100111111_0111000001001100"; -- 0.12987424714467086
	pesos_i(6889) := b"1111111111111111_1111111111111111_1111110111001101_0011100001101000"; -- -0.008587336229884536
	pesos_i(6890) := b"0000000000000000_0000000000000000_0001111011000101_1100100101010010"; -- 0.120205481113268
	pesos_i(6891) := b"1111111111111111_1111111111111111_1101111110111111_1110100110111000"; -- -0.1259778905605856
	pesos_i(6892) := b"1111111111111111_1111111111111111_1100110010110101_0000010011110110"; -- -0.20036286339875317
	pesos_i(6893) := b"0000000000000000_0000000000000000_0000100000101000_0001001000101111"; -- 0.03186143535474882
	pesos_i(6894) := b"0000000000000000_0000000000000000_0000101001000110_0111111111100101"; -- 0.04013823840963088
	pesos_i(6895) := b"0000000000000000_0000000000000000_0000011000011011_1100101001000111"; -- 0.023861543888369245
	pesos_i(6896) := b"0000000000000000_0000000000000000_0010000001110101_1111011101111110"; -- 0.1268000300310192
	pesos_i(6897) := b"0000000000000000_0000000000000000_0000100001000111_1001000101101100"; -- 0.032342041883464234
	pesos_i(6898) := b"1111111111111111_1111111111111111_1110010000100111_0010101110001110"; -- -0.10877731114119082
	pesos_i(6899) := b"0000000000000000_0000000000000000_0000010000101111_1010010001101100"; -- 0.01635196340895388
	pesos_i(6900) := b"0000000000000000_0000000000000000_0000000011001110_0011110001100110"; -- 0.003146910565561937
	pesos_i(6901) := b"1111111111111111_1111111111111111_1101100010100010_1000111100100111"; -- -0.15376954369348486
	pesos_i(6902) := b"0000000000000000_0000000000000000_0010010110000001_1010011001010101"; -- 0.1465095479321988
	pesos_i(6903) := b"1111111111111111_1111111111111111_1110110010111010_1101101111011010"; -- -0.07527376096915439
	pesos_i(6904) := b"0000000000000000_0000000000000000_0000111001010110_0101010011001011"; -- 0.05600480984867777
	pesos_i(6905) := b"0000000000000000_0000000000000000_0000000011101110_0001001000011100"; -- 0.003632671119341026
	pesos_i(6906) := b"0000000000000000_0000000000000000_0001000100010000_1100100110001000"; -- 0.06666240280908824
	pesos_i(6907) := b"1111111111111111_1111111111111111_1111110100110111_1101000110110100"; -- -0.010867017206604079
	pesos_i(6908) := b"1111111111111111_1111111111111111_1110000011101110_0110000101011011"; -- -0.1213626052527345
	pesos_i(6909) := b"0000000000000000_0000000000000000_0001101110110001_1100001001101100"; -- 0.108181144167811
	pesos_i(6910) := b"0000000000000000_0000000000000000_0010101010010101_1111010010100000"; -- 0.16635064026568333
	pesos_i(6911) := b"1111111111111111_1111111111111111_1111100010001101_0010001000111100"; -- -0.029096470190864556
	pesos_i(6912) := b"0000000000000000_0000000000000000_0011001110000110_0100101011010110"; -- 0.2012678881960376
	pesos_i(6913) := b"0000000000000000_0000000000000000_0000000001110111_0110100011001111"; -- 0.0018220430667774275
	pesos_i(6914) := b"1111111111111111_1111111111111111_1110011101000101_1111110111110011"; -- -0.09658825704211432
	pesos_i(6915) := b"0000000000000000_0000000000000000_0000010100100100_1001001100000111"; -- 0.020089329861795267
	pesos_i(6916) := b"1111111111111111_1111111111111111_1101110101100011_0110110000001001"; -- -0.13520169045025393
	pesos_i(6917) := b"0000000000000000_0000000000000000_0000110101101000_1001111010100110"; -- 0.05237762023360067
	pesos_i(6918) := b"0000000000000000_0000000000000000_0000011011000001_1000101011111010"; -- 0.02639072999209676
	pesos_i(6919) := b"1111111111111111_1111111111111111_1101111101001110_0101010100111001"; -- -0.12771098489273905
	pesos_i(6920) := b"0000000000000000_0000000000000000_0010100110101011_1111010000100000"; -- 0.16278005385282363
	pesos_i(6921) := b"0000000000000000_0000000000000000_0010111111110101_1110100110011100"; -- 0.1873460774388052
	pesos_i(6922) := b"0000000000000000_0000000000000000_0000101110111100_1110001000100111"; -- 0.04585088207351271
	pesos_i(6923) := b"1111111111111111_1111111111111111_1111101011010001_0100101101011101"; -- -0.020243921054490577
	pesos_i(6924) := b"0000000000000000_0000000000000000_0001001010010011_1100111111000110"; -- 0.07256792624535804
	pesos_i(6925) := b"0000000000000000_0000000000000000_0001111101110111_0100100100000011"; -- 0.12291389784160682
	pesos_i(6926) := b"0000000000000000_0000000000000000_0001100000100101_1100101100111001"; -- 0.09432668816082285
	pesos_i(6927) := b"1111111111111111_1111111111111111_1100101001001001_1000001100001111"; -- -0.20981579673224002
	pesos_i(6928) := b"1111111111111111_1111111111111111_1111000111011100_0001010000001011"; -- -0.055235621756679676
	pesos_i(6929) := b"0000000000000000_0000000000000000_0010001111010100_0101010111000010"; -- 0.1399587247523398
	pesos_i(6930) := b"0000000000000000_0000000000000000_0000111110010110_1111110100010001"; -- 0.060897652208460086
	pesos_i(6931) := b"1111111111111111_1111111111111111_1100100010011011_0010011111000011"; -- -0.2163825176473621
	pesos_i(6932) := b"0000000000000000_0000000000000000_0011001100000100_1000110001110110"; -- 0.19928815720868773
	pesos_i(6933) := b"1111111111111111_1111111111111111_1111000001010110_0111110010001011"; -- -0.061180320713425135
	pesos_i(6934) := b"0000000000000000_0000000000000000_0001010111001111_0001101001110110"; -- 0.08519139663865263
	pesos_i(6935) := b"1111111111111111_1111111111111111_1111100011001000_0110000011010001"; -- -0.028192471449456274
	pesos_i(6936) := b"0000000000000000_0000000000000000_0000111110110011_1010001110001111"; -- 0.06133482197843369
	pesos_i(6937) := b"0000000000000000_0000000000000000_0000011110010011_1001111111110001"; -- 0.02959632514534774
	pesos_i(6938) := b"0000000000000000_0000000000000000_0001010110010111_0111110100100111"; -- 0.08434278691315047
	pesos_i(6939) := b"1111111111111111_1111111111111111_1111111100100101_1010010100101101"; -- -0.0033318295449163058
	pesos_i(6940) := b"1111111111111111_1111111111111111_1110010101010111_1110110111111001"; -- -0.10412705115318123
	pesos_i(6941) := b"1111111111111111_1111111111111111_1111011100101000_1100101110100000"; -- -0.03453376144187453
	pesos_i(6942) := b"0000000000000000_0000000000000000_0001001100000011_1110100110010101"; -- 0.07427844882504096
	pesos_i(6943) := b"0000000000000000_0000000000000000_0010101001010011_1100110110001000"; -- 0.16534123002671544
	pesos_i(6944) := b"1111111111111111_1111111111111111_1111010100001101_1001011010100001"; -- -0.04276140750042341
	pesos_i(6945) := b"0000000000000000_0000000000000000_0000010111011100_1101010000001001"; -- 0.022900821928874417
	pesos_i(6946) := b"1111111111111111_1111111111111111_1110110100111110_1000010111001010"; -- -0.07326473071453714
	pesos_i(6947) := b"1111111111111111_1111111111111111_1110101011000111_0001111111101101"; -- -0.08289909801362694
	pesos_i(6948) := b"0000000000000000_0000000000000000_0000011001011111_0100111101001000"; -- 0.02489181053651111
	pesos_i(6949) := b"0000000000000000_0000000000000000_0001011000111110_0000011010000100"; -- 0.08688393325361489
	pesos_i(6950) := b"0000000000000000_0000000000000000_0011010001001101_0010010000011010"; -- 0.20430207865849376
	pesos_i(6951) := b"1111111111111111_1111111111111111_1100110111110101_0000000011110001"; -- -0.1954802904703073
	pesos_i(6952) := b"1111111111111111_1111111111111111_1110000010111101_0011011100011100"; -- -0.12211280410506405
	pesos_i(6953) := b"1111111111111111_1111111111111111_1111110100110001_1100100110000011"; -- -0.01095905839924841
	pesos_i(6954) := b"1111111111111111_1111111111111111_1111011101001101_0011110111110100"; -- -0.03397763043672321
	pesos_i(6955) := b"0000000000000000_0000000000000000_0000101000010111_1110011000111011"; -- 0.039427174881137284
	pesos_i(6956) := b"0000000000000000_0000000000000000_0010110001101100_0110011111110101"; -- 0.1735291456542883
	pesos_i(6957) := b"0000000000000000_0000000000000000_0000011011110000_0101101110110000"; -- 0.02710507426754106
	pesos_i(6958) := b"0000000000000000_0000000000000000_0001010010110001_0000010001010001"; -- 0.08082606303912533
	pesos_i(6959) := b"0000000000000000_0000000000000000_0001001000100100_1001010101001011"; -- 0.07087071504742068
	pesos_i(6960) := b"1111111111111111_1111111111111111_1111110111101000_1100000000000011"; -- -0.008167266105997465
	pesos_i(6961) := b"1111111111111111_1111111111111111_1111111101111100_1101101100101000"; -- -0.002001097515052968
	pesos_i(6962) := b"0000000000000000_0000000000000000_0000111010000101_0111100011111001"; -- 0.056724129529863825
	pesos_i(6963) := b"0000000000000000_0000000000000000_0000011001100011_1000111010101011"; -- 0.024956623754047426
	pesos_i(6964) := b"1111111111111111_1111111111111111_1110011111110010_0111110101100111"; -- -0.09395614841945876
	pesos_i(6965) := b"0000000000000000_0000000000000000_0011010111111100_1100110010001001"; -- 0.21088865601396217
	pesos_i(6966) := b"1111111111111111_1111111111111111_1101010001010001_1110010010111100"; -- -0.1706254044867064
	pesos_i(6967) := b"1111111111111111_1111111111111111_1111100001000011_1110001111101001"; -- -0.03021407660513456
	pesos_i(6968) := b"0000000000000000_0000000000000000_0011001110110110_1111101001100000"; -- 0.20201077318441163
	pesos_i(6969) := b"1111111111111111_1111111111111111_1111111010011010_1101100100010001"; -- -0.005449708408194579
	pesos_i(6970) := b"0000000000000000_0000000000000000_0000010001100110_0001111100011100"; -- 0.017183250658717272
	pesos_i(6971) := b"1111111111111111_1111111111111111_1100010111111101_1000110000011100"; -- -0.2265999252024778
	pesos_i(6972) := b"1111111111111111_1111111111111111_1110111101000010_1100101111011110"; -- -0.06538701849971112
	pesos_i(6973) := b"0000000000000000_0000000000000000_0011010100100000_0110101101110110"; -- 0.2075259365008984
	pesos_i(6974) := b"1111111111111111_1111111111111111_1111101111101101_1110111000111110"; -- -0.015900716619926054
	pesos_i(6975) := b"1111111111111111_1111111111111111_1110001100011000_1100110000101110"; -- -0.11290286899460522
	pesos_i(6976) := b"1111111111111111_1111111111111111_1110111110100010_0010101001000001"; -- -0.06393180768003656
	pesos_i(6977) := b"0000000000000000_0000000000000000_0000010000100111_1010111011110011"; -- 0.016230520502899127
	pesos_i(6978) := b"1111111111111111_1111111111111111_1111001001110010_0100100101001011"; -- -0.05294362948002185
	pesos_i(6979) := b"0000000000000000_0000000000000000_0001110110110010_0001111101100001"; -- 0.11599918472801635
	pesos_i(6980) := b"0000000000000000_0000000000000000_0001011101000101_0110110100111011"; -- 0.09090311700736561
	pesos_i(6981) := b"1111111111111111_1111111111111111_1110101000111011_0001010100110001"; -- -0.08503596843981796
	pesos_i(6982) := b"1111111111111111_1111111111111111_1111000110000101_1010011100100000"; -- -0.05655436965179272
	pesos_i(6983) := b"1111111111111111_1111111111111111_1111010110011110_1010010010010010"; -- -0.04054805206916356
	pesos_i(6984) := b"0000000000000000_0000000000000000_0010111101100010_0000011010110101"; -- 0.1850895110813437
	pesos_i(6985) := b"1111111111111111_1111111111111111_1111010010000101_0001000111011010"; -- -0.04484451705250323
	pesos_i(6986) := b"1111111111111111_1111111111111111_1110101100100000_0001101001100000"; -- -0.08154139657119189
	pesos_i(6987) := b"1111111111111111_1111111111111111_1100011101111101_0010010010001011"; -- -0.22074672326631128
	pesos_i(6988) := b"0000000000000000_0000000000000000_0001111100110010_0111101011100000"; -- 0.1218640133192932
	pesos_i(6989) := b"0000000000000000_0000000000000000_0001011100110000_0110100111101011"; -- 0.09058248516205489
	pesos_i(6990) := b"0000000000000000_0000000000000000_0010010000000001_0111101111001010"; -- 0.14064763726775503
	pesos_i(6991) := b"1111111111111111_1111111111111111_1101010110000011_1101010101101011"; -- -0.16595712803981316
	pesos_i(6992) := b"0000000000000000_0000000000000000_0001111101100100_1110001011111010"; -- 0.12263315773587104
	pesos_i(6993) := b"1111111111111111_1111111111111111_1111101101011111_1010010100111100"; -- -0.01807181641895993
	pesos_i(6994) := b"1111111111111111_1111111111111111_1111011110110100_0000101100100001"; -- -0.03240900454560657
	pesos_i(6995) := b"1111111111111111_1111111111111111_1111110001000001_1010010010001110"; -- -0.014623370602710649
	pesos_i(6996) := b"0000000000000000_0000000000000000_0010110111101010_0001111100111011"; -- 0.17935366820596868
	pesos_i(6997) := b"0000000000000000_0000000000000000_0000101011110010_0000111010000011"; -- 0.04275599184505091
	pesos_i(6998) := b"0000000000000000_0000000000000000_0000000110111101_1011000111111111"; -- 0.006800770574303231
	pesos_i(6999) := b"0000000000000000_0000000000000000_0001010001001011_0010010011101010"; -- 0.07927160937953322
	pesos_i(7000) := b"0000000000000000_0000000000000000_0001111010010110_1111101101101011"; -- 0.11949130405459979
	pesos_i(7001) := b"0000000000000000_0000000000000000_0001100011001100_0000111011100000"; -- 0.09686367949403686
	pesos_i(7002) := b"1111111111111111_1111111111111111_1111010100100111_0110001111100110"; -- -0.0423677029290991
	pesos_i(7003) := b"0000000000000000_0000000000000000_0001001000000001_0110001111101011"; -- 0.07033371445019079
	pesos_i(7004) := b"1111111111111111_1111111111111111_1011100101001011_0000001001011001"; -- -0.2761992008771634
	pesos_i(7005) := b"0000000000000000_0000000000000000_0000011100101000_0001101101000111"; -- 0.02795572748910733
	pesos_i(7006) := b"0000000000000000_0000000000000000_0001000110111111_1000010110001100"; -- 0.06932863881401863
	pesos_i(7007) := b"0000000000000000_0000000000000000_0000011100011101_1011011110000101"; -- 0.02779719357375449
	pesos_i(7008) := b"1111111111111111_1111111111111111_1110100111111100_1001100000101101"; -- -0.08598946465865773
	pesos_i(7009) := b"0000000000000000_0000000000000000_0010110010000011_0100100001011111"; -- 0.17387821501125963
	pesos_i(7010) := b"0000000000000000_0000000000000000_0001101100101110_0000110100110011"; -- 0.10617144097456314
	pesos_i(7011) := b"1111111111111111_1111111111111111_1110011100010001_1001111110010011"; -- -0.09738733933707669
	pesos_i(7012) := b"1111111111111111_1111111111111111_1101001101010011_1011111110011001"; -- -0.1745033504805972
	pesos_i(7013) := b"0000000000000000_0000000000000000_0001111011011101_1110101101100001"; -- 0.12057372213040787
	pesos_i(7014) := b"0000000000000000_0000000000000000_0001110100011000_1001101010001010"; -- 0.11365667209131533
	pesos_i(7015) := b"1111111111111111_1111111111111111_1101111110000101_1111110101010101"; -- -0.1268617312467164
	pesos_i(7016) := b"0000000000000000_0000000000000000_0000010000001010_1010100101110001"; -- 0.015787687387991432
	pesos_i(7017) := b"1111111111111111_1111111111111111_1110111110000111_1001011111101001"; -- -0.06433725890028184
	pesos_i(7018) := b"1111111111111111_1111111111111111_1110000011110011_1110101100111101"; -- -0.12127809288182416
	pesos_i(7019) := b"0000000000000000_0000000000000000_0011011000010101_0011100110100011"; -- 0.21126136998374095
	pesos_i(7020) := b"0000000000000000_0000000000000000_0010011110111111_1011111001100010"; -- 0.1552695264053099
	pesos_i(7021) := b"0000000000000000_0000000000000000_0010010100101110_0110011010000101"; -- 0.14523926489510555
	pesos_i(7022) := b"0000000000000000_0000000000000000_0010100110001111_1110000100111111"; -- 0.16235168245475837
	pesos_i(7023) := b"1111111111111111_1111111111111111_1100111001101101_1000100010101010"; -- -0.19364114611637956
	pesos_i(7024) := b"1111111111111111_1111111111111111_1101000101011101_1101110111000100"; -- -0.18216146434402425
	pesos_i(7025) := b"0000000000000000_0000000000000000_0000000010101011_1001001001010000"; -- 0.0026179737985228763
	pesos_i(7026) := b"0000000000000000_0000000000000000_0010111001010001_1111111110110101"; -- 0.18093870317181518
	pesos_i(7027) := b"1111111111111111_1111111111111111_1110101010000001_1010110111010000"; -- -0.08395875616999633
	pesos_i(7028) := b"1111111111111111_1111111111111111_1111010011001110_0001011011110010"; -- -0.0437303218746033
	pesos_i(7029) := b"0000000000000000_0000000000000000_0010110000110000_0101000110001010"; -- 0.17261228201372245
	pesos_i(7030) := b"0000000000000000_0000000000000000_0011001010101011_0010011100100001"; -- 0.1979240852741212
	pesos_i(7031) := b"0000000000000000_0000000000000000_0001101110110101_0001111000010000"; -- 0.10823238272290116
	pesos_i(7032) := b"0000000000000000_0000000000000000_0000011011101100_1111001110111101"; -- 0.02705310211661216
	pesos_i(7033) := b"0000000000000000_0000000000000000_0010110011011001_0011000001001001"; -- 0.17518903530006963
	pesos_i(7034) := b"0000000000000000_0000000000000000_0010100110111011_1100001100010011"; -- 0.16302127095129107
	pesos_i(7035) := b"0000000000000000_0000000000000000_0000011101101000_1010000000000101"; -- 0.02894020188882232
	pesos_i(7036) := b"0000000000000000_0000000000000000_0000110010000010_1110101000010010"; -- 0.048872594273319796
	pesos_i(7037) := b"1111111111111111_1111111111111111_1110101101010011_1011000101011000"; -- -0.0807542000132663
	pesos_i(7038) := b"0000000000000000_0000000000000000_0011001000111010_1100000000100111"; -- 0.19620896295279758
	pesos_i(7039) := b"1111111111111111_1111111111111111_1110010111100011_1100011000100000"; -- -0.10199319573763384
	pesos_i(7040) := b"1111111111111111_1111111111111111_1101010000110010_0111001111000001"; -- -0.1711051611860155
	pesos_i(7041) := b"1111111111111111_1111111111111111_1110001111100001_1000011011000011"; -- -0.10983999007766915
	pesos_i(7042) := b"1111111111111111_1111111111111111_1111100010101110_1100000010001000"; -- -0.028583494884060087
	pesos_i(7043) := b"0000000000000000_0000000000000000_0010100100010001_1011110001001101"; -- 0.16042687292867583
	pesos_i(7044) := b"0000000000000000_0000000000000000_0000001010110010_0000110001010100"; -- 0.010529299279139655
	pesos_i(7045) := b"1111111111111111_1111111111111111_1110110110011010_0011111101011110"; -- -0.07186511945879358
	pesos_i(7046) := b"0000000000000000_0000000000000000_0011100101110111_0111011000101010"; -- 0.2244790889220787
	pesos_i(7047) := b"1111111111111111_1111111111111111_1110110110111010_1000000011100110"; -- -0.0713729323258747
	pesos_i(7048) := b"0000000000000000_0000000000000000_0001001110101011_1101111110001100"; -- 0.0768413272769029
	pesos_i(7049) := b"1111111111111111_1111111111111111_1110010101011011_0111000011101010"; -- -0.10407346988250299
	pesos_i(7050) := b"0000000000000000_0000000000000000_0000100010110011_1001110100101010"; -- 0.03399069089125758
	pesos_i(7051) := b"1111111111111111_1111111111111111_1101100010111000_1001110100110101"; -- -0.1534330125141998
	pesos_i(7052) := b"0000000000000000_0000000000000000_0010010110001000_1000110111101010"; -- 0.14661490411658581
	pesos_i(7053) := b"0000000000000000_0000000000000000_0010011000001000_0110100101101110"; -- 0.14856585433352917
	pesos_i(7054) := b"0000000000000000_0000000000000000_0010101001100101_1100100011110011"; -- 0.16561561525136642
	pesos_i(7055) := b"1111111111111111_1111111111111111_1111000111000000_0100101010000010"; -- -0.05565962155778023
	pesos_i(7056) := b"1111111111111111_1111111111111111_1110010100100111_1111001111011000"; -- -0.10485912300880385
	pesos_i(7057) := b"1111111111111111_1111111111111111_1110101100011101_0110111101011110"; -- -0.08158210700987358
	pesos_i(7058) := b"1111111111111111_1111111111111111_1101001101110110_1101010101100010"; -- -0.17396799420765055
	pesos_i(7059) := b"0000000000000000_0000000000000000_0010111011001011_1110100100000011"; -- 0.18279892269528317
	pesos_i(7060) := b"1111111111111111_1111111111111111_1111100110010000_0001000000100010"; -- -0.0251455228639518
	pesos_i(7061) := b"0000000000000000_0000000000000000_0001000101010001_0010000100101110"; -- 0.06764418949325841
	pesos_i(7062) := b"1111111111111111_1111111111111111_1110001100000100_1000001000100111"; -- -0.1132124572567223
	pesos_i(7063) := b"1111111111111111_1111111111111111_1100100111111110_0100001010111101"; -- -0.21096403957367105
	pesos_i(7064) := b"1111111111111111_1111111111111111_1101011111010001_0101100111011111"; -- -0.15696180644664048
	pesos_i(7065) := b"1111111111111111_1111111111111111_1111001101101011_0011111101111110"; -- -0.049144775104316855
	pesos_i(7066) := b"1111111111111111_1111111111111111_1110001010101100_0010010000010010"; -- -0.1145608382086639
	pesos_i(7067) := b"1111111111111111_1111111111111111_1101000000110101_0101010010110001"; -- -0.18668623607086224
	pesos_i(7068) := b"0000000000000000_0000000000000000_0010100111101001_1010101100100011"; -- 0.16372174833535505
	pesos_i(7069) := b"1111111111111111_1111111111111111_1110001100111011_1101100010011110"; -- -0.11236807002973777
	pesos_i(7070) := b"1111111111111111_1111111111111111_1110011001110101_1101001000100100"; -- -0.0997646962647188
	pesos_i(7071) := b"1111111111111111_1111111111111111_1110011111011100_1001111010111110"; -- -0.09428985463348212
	pesos_i(7072) := b"0000000000000000_0000000000000000_0010001100001111_0100000001000011"; -- 0.13695146203717834
	pesos_i(7073) := b"1111111111111111_1111111111111111_1111010101111101_0001001101010001"; -- -0.041060249999045645
	pesos_i(7074) := b"0000000000000000_0000000000000000_0010000010001000_0111101100001110"; -- 0.12708252994417962
	pesos_i(7075) := b"1111111111111111_1111111111111111_1111110001101001_1111000001001000"; -- -0.01400850527788334
	pesos_i(7076) := b"0000000000000000_0000000000000000_0000100101101010_0110001111010100"; -- 0.03677963181013168
	pesos_i(7077) := b"1111111111111111_1111111111111111_1101011101101000_1100011001010001"; -- -0.15855751533916757
	pesos_i(7078) := b"1111111111111111_1111111111111111_1100101101001001_1100101000011110"; -- -0.20590531128499975
	pesos_i(7079) := b"0000000000000000_0000000000000000_0010110011111111_0001100111010000"; -- 0.17576752967211215
	pesos_i(7080) := b"0000000000000000_0000000000000000_0000101010001111_0101100001101111"; -- 0.04124977788881418
	pesos_i(7081) := b"1111111111111111_1111111111111111_1101100100110110_1000000001010000"; -- -0.151512127256034
	pesos_i(7082) := b"1111111111111111_1111111111111111_1101100001100010_0010100010101000"; -- -0.1547522153226598
	pesos_i(7083) := b"0000000000000000_0000000000000000_0000000101110110_0010101000001101"; -- 0.00570929348813781
	pesos_i(7084) := b"1111111111111111_1111111111111111_1110000100101010_1111110000110100"; -- -0.12043784842186646
	pesos_i(7085) := b"1111111111111111_1111111111111111_1111001000011110_1111101110000100"; -- -0.05421474481717628
	pesos_i(7086) := b"0000000000000000_0000000000000000_0010010101111111_1010011101101100"; -- 0.1464790952802639
	pesos_i(7087) := b"1111111111111111_1111111111111111_1111011001000010_1000101010000110"; -- -0.038047163328650706
	pesos_i(7088) := b"1111111111111111_1111111111111111_1110100000110101_0111010111101111"; -- -0.0929342548087629
	pesos_i(7089) := b"0000000000000000_0000000000000000_0001010001001100_1111100101111111"; -- 0.07929953906630643
	pesos_i(7090) := b"1111111111111111_1111111111111111_1110001000101111_1001110011101010"; -- -0.11646098415761608
	pesos_i(7091) := b"0000000000000000_0000000000000000_0000111111010101_1000010001101001"; -- 0.06185176435021854
	pesos_i(7092) := b"0000000000000000_0000000000000000_0000111011000100_1000011100101011"; -- 0.05768627933266816
	pesos_i(7093) := b"0000000000000000_0000000000000000_0001110101101011_1100111110000100"; -- 0.11492630922604125
	pesos_i(7094) := b"0000000000000000_0000000000000000_0000001100011101_1110100011101011"; -- 0.01217513781767428
	pesos_i(7095) := b"0000000000000000_0000000000000000_0001011010100010_0111101100100001"; -- 0.08841676295071005
	pesos_i(7096) := b"0000000000000000_0000000000000000_0001000100011111_0010101101011101"; -- 0.06688185723002295
	pesos_i(7097) := b"1111111111111111_1111111111111111_1111001010010110_1110000001111111"; -- -0.05238530071796857
	pesos_i(7098) := b"1111111111111111_1111111111111111_1111000001000110_0110010001011010"; -- -0.06142590337625509
	pesos_i(7099) := b"1111111111111111_1111111111111111_1100001101001010_0010100010111100"; -- -0.23714967159446412
	pesos_i(7100) := b"0000000000000000_0000000000000000_0000110010111111_1100100100101100"; -- 0.04980141939999484
	pesos_i(7101) := b"1111111111111111_1111111111111111_1110101010100101_0001001010000011"; -- -0.08341869631205456
	pesos_i(7102) := b"0000000000000000_0000000000000000_0000001011100011_1110011000001110"; -- 0.011289957518784956
	pesos_i(7103) := b"1111111111111111_1111111111111111_1111011111101100_0111100001001010"; -- -0.03154800591384274
	pesos_i(7104) := b"0000000000000000_0000000000000000_0011101001110001_1101110111001101"; -- 0.22829996350489715
	pesos_i(7105) := b"1111111111111111_1111111111111111_1110100001010001_0001100010011000"; -- -0.09251257211003149
	pesos_i(7106) := b"1111111111111111_1111111111111111_1111010100011001_0111100010010100"; -- -0.04258009329500206
	pesos_i(7107) := b"0000000000000000_0000000000000000_0011010000110101_0010000111001001"; -- 0.20393572951080924
	pesos_i(7108) := b"0000000000000000_0000000000000000_0011101111001001_0110001101010001"; -- 0.23354168631213765
	pesos_i(7109) := b"1111111111111111_1111111111111111_1101000001010001_0111000000111000"; -- -0.186257349424472
	pesos_i(7110) := b"0000000000000000_0000000000000000_0000101111100110_0010101000000011"; -- 0.04648077554190224
	pesos_i(7111) := b"0000000000000000_0000000000000000_0011011001010010_0111110111100100"; -- 0.21219622439180572
	pesos_i(7112) := b"0000000000000000_0000000000000000_0010110010101001_1000100101100110"; -- 0.17446192490723705
	pesos_i(7113) := b"0000000000000000_0000000000000000_0011010011010010_1100101001001010"; -- 0.2063414030826
	pesos_i(7114) := b"0000000000000000_0000000000000000_0011000000111101_1000010101111011"; -- 0.1884387421362958
	pesos_i(7115) := b"1111111111111111_1111111111111111_1110100101011111_0111010011100100"; -- -0.08838719774885179
	pesos_i(7116) := b"1111111111111111_1111111111111111_1111001011000010_1011110110010000"; -- -0.05171599617388511
	pesos_i(7117) := b"0000000000000000_0000000000000000_0001101110010011_1100000010011100"; -- 0.10772327239705895
	pesos_i(7118) := b"1111111111111111_1111111111111111_1101000001001001_1000010111001000"; -- -0.18637813448067006
	pesos_i(7119) := b"0000000000000000_0000000000000000_0010000101100011_1100100000000000"; -- 0.1304287911484685
	pesos_i(7120) := b"1111111111111111_1111111111111111_1111010110111111_0111101110100010"; -- -0.04004695222610448
	pesos_i(7121) := b"1111111111111111_1111111111111111_1110111111010100_0110111111000010"; -- -0.06316472534896753
	pesos_i(7122) := b"0000000000000000_0000000000000000_0001001100100001_1000000011000000"; -- 0.07472996416512263
	pesos_i(7123) := b"0000000000000000_0000000000000000_0010011110000101_0110111100101100"; -- 0.15437979534158686
	pesos_i(7124) := b"1111111111111111_1111111111111111_1110000001100110_1111101100111010"; -- -0.12342862929822657
	pesos_i(7125) := b"1111111111111111_1111111111111111_1110100101000001_0010001010111000"; -- -0.08884985941153571
	pesos_i(7126) := b"0000000000000000_0000000000000000_0010110000111000_1000001011010100"; -- 0.1727372901608185
	pesos_i(7127) := b"1111111111111111_1111111111111111_1100111100110000_0100001100100110"; -- -0.19066982583722974
	pesos_i(7128) := b"0000000000000000_0000000000000000_0001100110101000_1010001101101011"; -- 0.10022946711999275
	pesos_i(7129) := b"1111111111111111_1111111111111111_1110101011001101_0001010110001111"; -- -0.08280816316551493
	pesos_i(7130) := b"0000000000000000_0000000000000000_0010011011101110_0000000010100000"; -- 0.15206912898665603
	pesos_i(7131) := b"0000000000000000_0000000000000000_0000110000010100_0010110011010110"; -- 0.04718284824313328
	pesos_i(7132) := b"0000000000000000_0000000000000000_0000100000110110_0101111100010101"; -- 0.03207964183843566
	pesos_i(7133) := b"1111111111111111_1111111111111111_1101110000010010_0010000010001010"; -- -0.14034840224928802
	pesos_i(7134) := b"1111111111111111_1111111111111111_1101011111000110_0000011100111101"; -- -0.1571345783703801
	pesos_i(7135) := b"1111111111111111_1111111111111111_1110101101011000_1000001011001101"; -- -0.08068068016940193
	pesos_i(7136) := b"1111111111111111_1111111111111111_1110101001010111_1000011001001101"; -- -0.08460198032614281
	pesos_i(7137) := b"0000000000000000_0000000000000000_0000110010111111_1010111011010100"; -- 0.04979984918560872
	pesos_i(7138) := b"1111111111111111_1111111111111111_1100110010111111_0010000111001010"; -- -0.20020855724000536
	pesos_i(7139) := b"1111111111111111_1111111111111111_1110110010000000_1011111111100010"; -- -0.07616043794689684
	pesos_i(7140) := b"0000000000000000_0000000000000000_0011010110000110_1000010001100000"; -- 0.20908381799110487
	pesos_i(7141) := b"0000000000000000_0000000000000000_0011001001011110_1110111110000101"; -- 0.196761102683165
	pesos_i(7142) := b"0000000000000000_0000000000000000_0000111111001111_0011100111011110"; -- 0.06175576842699456
	pesos_i(7143) := b"1111111111111111_1111111111111111_1111111010001010_0111010110110000"; -- -0.0056997722851547744
	pesos_i(7144) := b"1111111111111111_1111111111111111_1101010110001100_1001101000000111"; -- -0.16582333869404337
	pesos_i(7145) := b"1111111111111111_1111111111111111_1100101101100000_0101100101111011"; -- -0.20556107287444195
	pesos_i(7146) := b"1111111111111111_1111111111111111_1111001100010011_1001010110010000"; -- -0.05048241831536377
	pesos_i(7147) := b"1111111111111111_1111111111111111_1100100010001000_1100101011010101"; -- -0.21666271490125544
	pesos_i(7148) := b"1111111111111111_1111111111111111_1100111110000011_0011101101001010"; -- -0.1894038146193725
	pesos_i(7149) := b"0000000000000000_0000000000000000_0010011110110100_1010101010000101"; -- 0.15510049581530094
	pesos_i(7150) := b"0000000000000000_0000000000000000_0000101010100000_1101010010101000"; -- 0.04151658155692205
	pesos_i(7151) := b"1111111111111111_1111111111111111_1101011100010010_1100011111100000"; -- -0.15986967833617477
	pesos_i(7152) := b"0000000000000000_0000000000000000_0000101110000110_0101111101110101"; -- 0.04501911746249425
	pesos_i(7153) := b"0000000000000000_0000000000000000_0010101000011101_0010011001011000"; -- 0.1645072903716477
	pesos_i(7154) := b"1111111111111111_1111111111111111_1110011000111001_0001000100000001"; -- -0.10069173550911055
	pesos_i(7155) := b"1111111111111111_1111111111111111_1101010101101010_0111010011110000"; -- -0.16634434828514325
	pesos_i(7156) := b"0000000000000000_0000000000000000_0001111100111111_1110100110110110"; -- 0.12206898385200389
	pesos_i(7157) := b"0000000000000000_0000000000000000_0010010001010000_0001001111000110"; -- 0.1418468817564868
	pesos_i(7158) := b"1111111111111111_1111111111111111_1110100010000100_0010000010100010"; -- -0.09173389487199099
	pesos_i(7159) := b"1111111111111111_1111111111111111_1101110011110101_1101011001101101"; -- -0.13687381594789622
	pesos_i(7160) := b"0000000000000000_0000000000000000_0010010111101010_1111001010110101"; -- 0.14811627312888942
	pesos_i(7161) := b"1111111111111111_1111111111111111_1110111101010100_1011000100001110"; -- -0.0651139584151772
	pesos_i(7162) := b"1111111111111111_1111111111111111_1101011010010001_1000000000111100"; -- -0.16184233233529183
	pesos_i(7163) := b"0000000000000000_0000000000000000_0001000100001001_0010110100011001"; -- 0.06654626707106136
	pesos_i(7164) := b"0000000000000000_0000000000000000_0001100100111100_1000110110100001"; -- 0.09858021905925614
	pesos_i(7165) := b"1111111111111111_1111111111111111_1111000000001000_1101001011001000"; -- -0.06236536624225016
	pesos_i(7166) := b"0000000000000000_0000000000000000_0010010000010000_1101110110100110"; -- 0.14088235194829027
	pesos_i(7167) := b"0000000000000000_0000000000000000_0010011111000010_0010000011000101"; -- 0.15530590839349598
	pesos_i(7168) := b"1111111111111111_1111111111111111_1101111010010000_0100000011000001"; -- -0.13061137470508485
	pesos_i(7169) := b"0000000000000000_0000000000000000_0001111111001110_0100011001100010"; -- 0.12424125571344591
	pesos_i(7170) := b"1111111111111111_1111111111111111_1110110010101111_1000110110010010"; -- -0.07544627370858681
	pesos_i(7171) := b"0000000000000000_0000000000000000_0010001110101001_1011010000000111"; -- 0.1393082157138554
	pesos_i(7172) := b"0000000000000000_0000000000000000_0010110100001011_1011011111100011"; -- 0.1759600572088742
	pesos_i(7173) := b"0000000000000000_0000000000000000_0010000110101100_0111010010000111"; -- 0.13153770731777914
	pesos_i(7174) := b"0000000000000000_0000000000000000_0000010110000111_1110101101011110"; -- 0.021605215425472803
	pesos_i(7175) := b"0000000000000000_0000000000000000_0000100101011011_1010000010101011"; -- 0.036554376296924644
	pesos_i(7176) := b"1111111111111111_1111111111111111_1110111101000101_0111100010110000"; -- -0.06534619993377824
	pesos_i(7177) := b"1111111111111111_1111111111111111_1110011111101010_0010100010011000"; -- -0.09408327383351778
	pesos_i(7178) := b"0000000000000000_0000000000000000_0000101100001001_1110100001110101"; -- 0.04311993454360052
	pesos_i(7179) := b"1111111111111111_1111111111111111_1111001001000101_1111001011000011"; -- -0.05362017388619245
	pesos_i(7180) := b"1111111111111111_1111111111111111_1100111101011011_0111001000100111"; -- -0.19001089618032177
	pesos_i(7181) := b"0000000000000000_0000000000000000_0000000010010100_0001010011000011"; -- 0.002259538168348109
	pesos_i(7182) := b"0000000000000000_0000000000000000_0001010101000001_1111011011100111"; -- 0.08303778782646543
	pesos_i(7183) := b"0000000000000000_0000000000000000_0010011001010110_1000110011111001"; -- 0.1497581584953665
	pesos_i(7184) := b"0000000000000000_0000000000000000_0011000111000011_1100110001000010"; -- 0.19439388863953902
	pesos_i(7185) := b"1111111111111111_1111111111111111_1110111101000011_0110100111100011"; -- -0.0653775998365171
	pesos_i(7186) := b"1111111111111111_1111111111111111_1100010001110011_1011100010101000"; -- -0.23260923281614118
	pesos_i(7187) := b"1111111111111111_1111111111111111_1111101110011000_1110111011101110"; -- -0.017197672693949402
	pesos_i(7188) := b"1111111111111111_1111111111111111_1101010111011111_1010000001001011"; -- -0.16455648590228766
	pesos_i(7189) := b"1111111111111111_1111111111111111_1101000110110010_1111001010000101"; -- -0.18086323027610585
	pesos_i(7190) := b"0000000000000000_0000000000000000_0010111110110010_1101100100000111"; -- 0.18632275024952724
	pesos_i(7191) := b"1111111111111111_1111111111111111_1111001010011100_0111011110011010"; -- -0.052300000022786085
	pesos_i(7192) := b"1111111111111111_1111111111111111_1100010110011011_1001101110100000"; -- -0.22809436168296884
	pesos_i(7193) := b"0000000000000000_0000000000000000_0001101011010110_1011111110001110"; -- 0.10483929841648466
	pesos_i(7194) := b"0000000000000000_0000000000000000_0010011010101000_0000111101010000"; -- 0.15100188927202635
	pesos_i(7195) := b"0000000000000000_0000000000000000_0000011001111110_0011100010000001"; -- 0.025363475298328584
	pesos_i(7196) := b"0000000000000000_0000000000000000_0000001111011110_0010001001111100"; -- 0.015108256486804085
	pesos_i(7197) := b"1111111111111111_1111111111111111_1110110100101010_0001110001110000"; -- -0.0735761858632134
	pesos_i(7198) := b"0000000000000000_0000000000000000_0001001111100011_0001001101111011"; -- 0.07768365618995092
	pesos_i(7199) := b"0000000000000000_0000000000000000_0001010111101110_1101011001000111"; -- 0.08567561368862102
	pesos_i(7200) := b"0000000000000000_0000000000000000_0000101001000110_1101111000011101"; -- 0.040143854323746946
	pesos_i(7201) := b"0000000000000000_0000000000000000_0010011111101100_0000110000111010"; -- 0.15594555301563975
	pesos_i(7202) := b"1111111111111111_1111111111111111_1101011100100010_0111101011010100"; -- -0.15963012999534884
	pesos_i(7203) := b"0000000000000000_0000000000000000_0000101000001000_1010011111101100"; -- 0.039194579247695066
	pesos_i(7204) := b"1111111111111111_1111111111111111_1111001100101000_0011100111011001"; -- -0.05016745036469399
	pesos_i(7205) := b"0000000000000000_0000000000000000_0011100000110111_1000110110011001"; -- 0.21959767338152075
	pesos_i(7206) := b"1111111111111111_1111111111111111_1111110101001101_0001011010011110"; -- -0.010542475039410217
	pesos_i(7207) := b"1111111111111111_1111111111111111_1110111010010110_0101010100101000"; -- -0.06801860594611701
	pesos_i(7208) := b"0000000000000000_0000000000000000_0011001101011011_1100101101000101"; -- 0.20061941554728563
	pesos_i(7209) := b"0000000000000000_0000000000000000_0010100000011111_0010100011111010"; -- 0.15672546475764362
	pesos_i(7210) := b"1111111111111111_1111111111111111_1110001100001011_1001110010100100"; -- -0.11310406687356192
	pesos_i(7211) := b"1111111111111111_1111111111111111_1110101011110000_1101101010010001"; -- -0.08226236311944556
	pesos_i(7212) := b"1111111111111111_1111111111111111_1101010000001011_0101000100000100"; -- -0.17170232449271086
	pesos_i(7213) := b"1111111111111111_1111111111111111_1110110000010100_1111010110001110"; -- -0.07780518809087092
	pesos_i(7214) := b"1111111111111111_1111111111111111_1110011010111100_1101010100101000"; -- -0.09868114260713667
	pesos_i(7215) := b"0000000000000000_0000000000000000_0001001100011000_1110011000101100"; -- 0.07459868018222883
	pesos_i(7216) := b"1111111111111111_1111111111111111_1110110100001110_0001011001010101"; -- -0.07400379591169363
	pesos_i(7217) := b"0000000000000000_0000000000000000_0010001100010011_0001011111000101"; -- 0.13701008375023122
	pesos_i(7218) := b"1111111111111111_1111111111111111_1110010001010010_0101010000010001"; -- -0.10811876858399387
	pesos_i(7219) := b"1111111111111111_1111111111111111_1111110110001110_0011100000100010"; -- -0.009548656091760473
	pesos_i(7220) := b"1111111111111111_1111111111111111_1100011101010101_1000100010011110"; -- -0.22135110993937845
	pesos_i(7221) := b"0000000000000000_0000000000000000_0001001001000011_1010000001010000"; -- 0.0713443941482587
	pesos_i(7222) := b"0000000000000000_0000000000000000_0010000110010000_0111001100100011"; -- 0.13111037821588525
	pesos_i(7223) := b"0000000000000000_0000000000000000_0001101011010000_1110001111101000"; -- 0.10474991230435411
	pesos_i(7224) := b"1111111111111111_1111111111111111_1110001011100110_0000111110111001"; -- -0.11367704140224853
	pesos_i(7225) := b"1111111111111111_1111111111111111_1111111000010000_1111110111001001"; -- -0.0075532327094186774
	pesos_i(7226) := b"1111111111111111_1111111111111111_1110111110000000_1100001001000101"; -- -0.06444154570083675
	pesos_i(7227) := b"1111111111111111_1111111111111111_1110001011110010_0110101101101100"; -- -0.11348847016090415
	pesos_i(7228) := b"1111111111111111_1111111111111111_1100011001000000_1111110111111100"; -- -0.2255707987949689
	pesos_i(7229) := b"0000000000000000_0000000000000000_0000111001101110_0101010000111110"; -- 0.056370987957446654
	pesos_i(7230) := b"0000000000000000_0000000000000000_0001110000000101_1100110001111000"; -- 0.10946348113963894
	pesos_i(7231) := b"1111111111111111_1111111111111111_1100000010100011_1010110011101001"; -- -0.24750251116172345
	pesos_i(7232) := b"0000000000000000_0000000000000000_0010100000001000_1111100101001110"; -- 0.15638692994619693
	pesos_i(7233) := b"1111111111111111_1111111111111111_1110001011000100_0111001100000001"; -- -0.11418992262673373
	pesos_i(7234) := b"1111111111111111_1111111111111111_1110011011011110_0011110111100010"; -- -0.09817136025999043
	pesos_i(7235) := b"0000000000000000_0000000000000000_0010110010000011_0101100100111000"; -- 0.1738792191605053
	pesos_i(7236) := b"1111111111111111_1111111111111111_1110010010001110_1011010100011110"; -- -0.10719745645441842
	pesos_i(7237) := b"0000000000000000_0000000000000000_0011000011011011_1101101111011010"; -- 0.19085477898149023
	pesos_i(7238) := b"1111111111111111_1111111111111111_1111000001001011_1000010100110101"; -- -0.061347651060746036
	pesos_i(7239) := b"0000000000000000_0000000000000000_0001001101101011_1001010000010101"; -- 0.07586026682085
	pesos_i(7240) := b"1111111111111111_1111111111111111_1101101100011101_1101011100111010"; -- -0.1440759165815678
	pesos_i(7241) := b"0000000000000000_0000000000000000_0010000100010101_1010010011100111"; -- 0.12923651344342243
	pesos_i(7242) := b"1111111111111111_1111111111111111_1101000110000100_0011101101001110"; -- -0.1815760550078036
	pesos_i(7243) := b"0000000000000000_0000000000000000_0010010010010011_1110100011100101"; -- 0.14288192357500298
	pesos_i(7244) := b"1111111111111111_1111111111111111_1101100011110000_0110000010111001"; -- -0.15258212543689811
	pesos_i(7245) := b"1111111111111111_1111111111111111_1101011101001011_0110101111010101"; -- -0.15900541354866862
	pesos_i(7246) := b"1111111111111111_1111111111111111_1110001111000010_0101110110111101"; -- -0.11031545759487624
	pesos_i(7247) := b"0000000000000000_0000000000000000_0000110010101110_0001110000110011"; -- 0.04953171005611236
	pesos_i(7248) := b"0000000000000000_0000000000000000_0011001011101101_1101101000110001"; -- 0.19894183830147294
	pesos_i(7249) := b"1111111111111111_1111111111111111_1111001011011000_0110010000011100"; -- -0.05138563461908506
	pesos_i(7250) := b"1111111111111111_1111111111111111_1101011110101101_0100010100000100"; -- -0.15751236579883068
	pesos_i(7251) := b"0000000000000000_0000000000000000_0000010101110111_1110011011010110"; -- 0.02136080475581674
	pesos_i(7252) := b"0000000000000000_0000000000000000_0010001100010110_1010101001100101"; -- 0.1370645996571331
	pesos_i(7253) := b"1111111111111111_1111111111111111_1101100010101100_1000110101101001"; -- -0.15361705963985556
	pesos_i(7254) := b"0000000000000000_0000000000000000_0001100110111110_0101000001100001"; -- 0.10056021097638124
	pesos_i(7255) := b"1111111111111111_1111111111111111_1101110100010011_1111100010010101"; -- -0.13641401641913123
	pesos_i(7256) := b"1111111111111111_1111111111111111_1111000000110001_1011101111011110"; -- -0.06174112158984556
	pesos_i(7257) := b"0000000000000000_0000000000000000_0000110110001111_1101001100001110"; -- 0.05297583659839004
	pesos_i(7258) := b"1111111111111111_1111111111111111_1110110000010111_1010000101111000"; -- -0.07776442356559571
	pesos_i(7259) := b"0000000000000000_0000000000000000_0001001100111110_0010011010111000"; -- 0.07516710264342762
	pesos_i(7260) := b"1111111111111111_1111111111111111_1110011010001000_0110010101010010"; -- -0.09948126544365327
	pesos_i(7261) := b"1111111111111111_1111111111111111_1111111110110110_0101110101001000"; -- -0.001123590378983138
	pesos_i(7262) := b"1111111111111111_1111111111111111_1101010010010000_1000100100000111"; -- -0.16966956695159527
	pesos_i(7263) := b"1111111111111111_1111111111111111_1110100011010100_1000011011101011"; -- -0.09050709496425867
	pesos_i(7264) := b"1111111111111111_1111111111111111_1111011010011101_1100001100001011"; -- -0.036655244683760746
	pesos_i(7265) := b"1111111111111111_1111111111111111_1110110011000010_0001000011010101"; -- -0.0751637915449106
	pesos_i(7266) := b"1111111111111111_1111111111111111_1110011100101100_1110110101110101"; -- -0.09697070970070576
	pesos_i(7267) := b"0000000000000000_0000000000000000_0001101111010111_0010101010001001"; -- 0.10875192490380325
	pesos_i(7268) := b"0000000000000000_0000000000000000_0010101111100010_1001111110010011"; -- 0.17142674780110614
	pesos_i(7269) := b"0000000000000000_0000000000000000_0000100011110010_0100100100000010"; -- 0.034946978509842845
	pesos_i(7270) := b"1111111111111111_1111111111111111_1101111111000011_0000110111100110"; -- -0.12592995782196956
	pesos_i(7271) := b"0000000000000000_0000000000000000_0010000100111010_0011101000110000"; -- 0.12979472804239295
	pesos_i(7272) := b"1111111111111111_1111111111111111_1111110111111100_1011000100101010"; -- -0.007862975268479113
	pesos_i(7273) := b"1111111111111111_1111111111111111_1100100111001100_1100010000100001"; -- -0.21171926688251116
	pesos_i(7274) := b"1111111111111111_1111111111111111_1110001000111010_1001110010000110"; -- -0.11629316065628752
	pesos_i(7275) := b"0000000000000000_0000000000000000_0001001111010011_1011001011101101"; -- 0.07744901935021475
	pesos_i(7276) := b"1111111111111111_1111111111111111_1110001100010100_1110100111101111"; -- -0.11296213068193028
	pesos_i(7277) := b"1111111111111111_1111111111111111_1111011010001000_1000010011100111"; -- -0.03697938302795668
	pesos_i(7278) := b"1111111111111111_1111111111111111_1101110101001010_1110101100110001"; -- -0.13557558121223492
	pesos_i(7279) := b"0000000000000000_0000000000000000_0001101110100011_1111100111001101"; -- 0.10797082178772882
	pesos_i(7280) := b"1111111111111111_1111111111111111_1101110100101011_0010010010100101"; -- -0.13606043797406356
	pesos_i(7281) := b"0000000000000000_0000000000000000_0000011110010111_0101100000000101"; -- 0.02965307343280551
	pesos_i(7282) := b"1111111111111111_1111111111111111_1111000001011001_0000111110001110"; -- -0.06114104053034035
	pesos_i(7283) := b"0000000000000000_0000000000000000_0001001111010101_0101110100011101"; -- 0.07747442216384916
	pesos_i(7284) := b"0000000000000000_0000000000000000_0001101010111101_1010001000011111"; -- 0.10445607421047769
	pesos_i(7285) := b"1111111111111111_1111111111111111_1111011101110010_1110011100101010"; -- -0.03340296970049836
	pesos_i(7286) := b"0000000000000000_0000000000000000_0010011111110101_0010110110011010"; -- 0.15608487133986107
	pesos_i(7287) := b"1111111111111111_1111111111111111_1111101000110101_1010101110001101"; -- -0.02261855907253606
	pesos_i(7288) := b"0000000000000000_0000000000000000_0010101011101010_0011011010001101"; -- 0.16763630819936384
	pesos_i(7289) := b"0000000000000000_0000000000000000_0000011100101001_0111000101111000"; -- 0.027976123512254803
	pesos_i(7290) := b"1111111111111111_1111111111111111_1111000110001011_0110010110110111"; -- -0.05646671556632376
	pesos_i(7291) := b"0000000000000000_0000000000000000_0010000010010011_1010101111011011"; -- 0.12725328547278203
	pesos_i(7292) := b"0000000000000000_0000000000000000_0010100101110110_1000100111011001"; -- 0.1619650033872
	pesos_i(7293) := b"1111111111111111_1111111111111111_1100110111111110_1111100011001000"; -- -0.19532818894766069
	pesos_i(7294) := b"1111111111111111_1111111111111111_1110101000111001_1011110011011000"; -- -0.08505649297653262
	pesos_i(7295) := b"1111111111111111_1111111111111111_1101110111001010_1010001110000000"; -- -0.13362672919294766
	pesos_i(7296) := b"0000000000000000_0000000000000000_0001111000011110_1111001000110011"; -- 0.11765969988398686
	pesos_i(7297) := b"0000000000000000_0000000000000000_0010100110001100_1101011101100111"; -- 0.16230531938047307
	pesos_i(7298) := b"0000000000000000_0000000000000000_0000111011011111_0110111011100010"; -- 0.05809681913578474
	pesos_i(7299) := b"1111111111111111_1111111111111111_1101011001011110_1001000011001010"; -- -0.16261954377847312
	pesos_i(7300) := b"0000000000000000_0000000000000000_0011001100011110_1111000111110111"; -- 0.1996909359864964
	pesos_i(7301) := b"1111111111111111_1111111111111111_1100111111111101_0100001100101010"; -- -0.18754177311852988
	pesos_i(7302) := b"1111111111111111_1111111111111111_1111111111100111_1010001011011111"; -- -0.00037176173721546117
	pesos_i(7303) := b"1111111111111111_1111111111111111_1101011001010111_0100110101110101"; -- -0.16273036853793307
	pesos_i(7304) := b"1111111111111111_1111111111111111_1111001000110011_0101111100000010"; -- -0.05390363878212719
	pesos_i(7305) := b"1111111111111111_1111111111111111_1111100000000100_1000110011100000"; -- -0.031180568074189275
	pesos_i(7306) := b"0000000000000000_0000000000000000_0001001110110110_0011110000010100"; -- 0.07699943050296781
	pesos_i(7307) := b"1111111111111111_1111111111111111_1111010101110011_1111100101010010"; -- -0.041199128718016544
	pesos_i(7308) := b"1111111111111111_1111111111111111_1101001111110111_0101000001111010"; -- -0.17200753235338076
	pesos_i(7309) := b"0000000000000000_0000000000000000_0010111110101111_0001001100100000"; -- 0.18626517792677955
	pesos_i(7310) := b"0000000000000000_0000000000000000_0001001111011110_1010011010110101"; -- 0.07761613772619651
	pesos_i(7311) := b"0000000000000000_0000000000000000_0001110010000011_0001000001101000"; -- 0.11137487920853724
	pesos_i(7312) := b"0000000000000000_0000000000000000_0011010001101001_0111110110100000"; -- 0.20473466069144786
	pesos_i(7313) := b"1111111111111111_1111111111111111_1110000010011001_0011010010111011"; -- -0.12266226228933672
	pesos_i(7314) := b"1111111111111111_1111111111111111_1110110100110010_1110110100100100"; -- -0.07344167574906328
	pesos_i(7315) := b"0000000000000000_0000000000000000_0010011011111100_0100001110111001"; -- 0.15228675139287948
	pesos_i(7316) := b"1111111111111111_1111111111111111_1101001011011111_0000101000110111"; -- -0.1762841811882434
	pesos_i(7317) := b"0000000000000000_0000000000000000_0010010101000110_1000000110110001"; -- 0.14560709537587213
	pesos_i(7318) := b"1111111111111111_1111111111111111_1111101101000011_1100000001110101"; -- -0.018497439900418813
	pesos_i(7319) := b"0000000000000000_0000000000000000_0011010110100101_0011100011110100"; -- 0.20955234480766105
	pesos_i(7320) := b"1111111111111111_1111111111111111_1110001110100101_0000011111101011"; -- -0.11076307784286797
	pesos_i(7321) := b"1111111111111111_1111111111111111_1111110100010011_1000101111010000"; -- -0.01142049941995036
	pesos_i(7322) := b"0000000000000000_0000000000000000_0001000011010100_0101011110100010"; -- 0.06574008649335512
	pesos_i(7323) := b"0000000000000000_0000000000000000_0010011011110101_1111111100011100"; -- 0.15219110898586447
	pesos_i(7324) := b"0000000000000000_0000000000000000_0000011111101000_0101110101011001"; -- 0.030889352917917893
	pesos_i(7325) := b"0000000000000000_0000000000000000_0001110111111000_1110010101110110"; -- 0.11707910661588863
	pesos_i(7326) := b"1111111111111111_1111111111111111_1110000010101000_0010110001000001"; -- -0.12243388564853336
	pesos_i(7327) := b"0000000000000000_0000000000000000_0001110111010010_1011111101001001"; -- 0.11649699715066615
	pesos_i(7328) := b"1111111111111111_1111111111111111_1110110110001010_0110010111111010"; -- -0.07210695886101966
	pesos_i(7329) := b"0000000000000000_0000000000000000_0000100101010111_1101100001101110"; -- 0.03649666480523817
	pesos_i(7330) := b"1111111111111111_1111111111111111_1110110000011010_1100010110111001"; -- -0.07771648641102046
	pesos_i(7331) := b"0000000000000000_0000000000000000_0010010011010010_1001011000110000"; -- 0.1438382975066413
	pesos_i(7332) := b"0000000000000000_0000000000000000_0001110101110001_1110100011110011"; -- 0.11501937802200558
	pesos_i(7333) := b"0000000000000000_0000000000000000_0010010111100010_1101100111011110"; -- 0.14799272217995094
	pesos_i(7334) := b"0000000000000000_0000000000000000_0000001001011111_0111111011101011"; -- 0.009269649914964302
	pesos_i(7335) := b"0000000000000000_0000000000000000_0000111011100010_1110010010101011"; -- 0.05814961598662412
	pesos_i(7336) := b"1111111111111111_1111111111111111_1110010011000100_1001111101101100"; -- -0.10637477498308742
	pesos_i(7337) := b"1111111111111111_1111111111111111_1111110001111111_0100101000111110"; -- -0.013682708714600525
	pesos_i(7338) := b"0000000000000000_0000000000000000_0010111011100011_1011010101110000"; -- 0.18316205964947121
	pesos_i(7339) := b"0000000000000000_0000000000000000_0000110111100111_0001100110000110"; -- 0.0543075516588828
	pesos_i(7340) := b"1111111111111111_1111111111111111_1110100000100010_1101110011010100"; -- -0.09321803884408247
	pesos_i(7341) := b"0000000000000000_0000000000000000_0010101111101010_1100011100010111"; -- 0.17155117325974634
	pesos_i(7342) := b"0000000000000000_0000000000000000_0010110000101110_1100110100000101"; -- 0.1725891244065847
	pesos_i(7343) := b"1111111111111111_1111111111111111_1100110000000001_0111010011010100"; -- -0.2031027777268107
	pesos_i(7344) := b"1111111111111111_1111111111111111_1110111100100111_0101010011010111"; -- -0.06580610033280174
	pesos_i(7345) := b"1111111111111111_1111111111111111_1101011001100011_1001101000000111"; -- -0.16254269903233892
	pesos_i(7346) := b"1111111111111111_1111111111111111_1110111011001110_1100101011000110"; -- -0.06715710318869333
	pesos_i(7347) := b"1111111111111111_1111111111111111_1100010100111111_1100110000100101"; -- -0.2294952782992493
	pesos_i(7348) := b"0000000000000000_0000000000000000_0010101011111001_0110111110110110"; -- 0.16786859686491817
	pesos_i(7349) := b"1111111111111111_1111111111111111_1110001100110000_0101111110010101"; -- -0.11254313107375372
	pesos_i(7350) := b"0000000000000000_0000000000000000_0000111101000010_0010000000001101"; -- 0.059602740472757605
	pesos_i(7351) := b"0000000000000000_0000000000000000_0000111110111000_1001010010010010"; -- 0.06141022264563922
	pesos_i(7352) := b"0000000000000000_0000000000000000_0000011000100001_1011110010010011"; -- 0.023952279849378942
	pesos_i(7353) := b"1111111111111111_1111111111111111_1100111001011110_0000111001111111"; -- -0.19387730978061568
	pesos_i(7354) := b"0000000000000000_0000000000000000_0001001001010111_0111111100010010"; -- 0.07164758871351969
	pesos_i(7355) := b"1111111111111111_1111111111111111_1110100001001001_1001001101011100"; -- -0.09262732519824143
	pesos_i(7356) := b"1111111111111111_1111111111111111_1111010101010000_0100100100101000"; -- -0.04174368650993516
	pesos_i(7357) := b"1111111111111111_1111111111111111_1110101100100010_0101110010101101"; -- -0.08150692727539964
	pesos_i(7358) := b"1111111111111111_1111111111111111_1101011101100100_0010010010101111"; -- -0.15862818461177133
	pesos_i(7359) := b"1111111111111111_1111111111111111_1101110010100110_1011110001010000"; -- -0.13808081663650462
	pesos_i(7360) := b"0000000000000000_0000000000000000_0000001100101011_1001111000101100"; -- 0.012384305819575392
	pesos_i(7361) := b"0000000000000000_0000000000000000_0001100101110001_1010100111010010"; -- 0.0993906153068142
	pesos_i(7362) := b"1111111111111111_1111111111111111_1100111100000010_1001001010001110"; -- -0.191366997071364
	pesos_i(7363) := b"0000000000000000_0000000000000000_0010110101101100_0010011010110110"; -- 0.17743150657932838
	pesos_i(7364) := b"0000000000000000_0000000000000000_0000100111000010_0011001010110001"; -- 0.03811947651074793
	pesos_i(7365) := b"0000000000000000_0000000000000000_0001011111101011_1110000110011111"; -- 0.09344301342813155
	pesos_i(7366) := b"0000000000000000_0000000000000000_0010111001011010_0000110011101110"; -- 0.18106156167586784
	pesos_i(7367) := b"1111111111111111_1111111111111111_1111011100001011_1111001101101100"; -- -0.03497389418405486
	pesos_i(7368) := b"1111111111111111_1111111111111111_1111100111101100_0111010011001000"; -- -0.02373571499780111
	pesos_i(7369) := b"1111111111111111_1111111111111111_1111001110010100_1100110101010110"; -- -0.04851071034785917
	pesos_i(7370) := b"1111111111111111_1111111111111111_1110001010001000_1010110110000001"; -- -0.11510196299740637
	pesos_i(7371) := b"0000000000000000_0000000000000000_0000110111000101_0000111011011101"; -- 0.05378811747589968
	pesos_i(7372) := b"0000000000000000_0000000000000000_0000101111101101_1111100011011110"; -- 0.04659991675397429
	pesos_i(7373) := b"0000000000000000_0000000000000000_0000011001001011_0011011110000111"; -- 0.024585218912573037
	pesos_i(7374) := b"1111111111111111_1111111111111111_1101011110111110_1010101100010000"; -- -0.15724688400525252
	pesos_i(7375) := b"1111111111111111_1111111111111111_1100111010010010_1101001010101100"; -- -0.1930721597291568
	pesos_i(7376) := b"0000000000000000_0000000000000000_0011010000001000_1101001101000010"; -- 0.20325966230893228
	pesos_i(7377) := b"1111111111111111_1111111111111111_1110001100010111_1100111001110111"; -- -0.11291799162250024
	pesos_i(7378) := b"1111111111111111_1111111111111111_1101000010001101_1111011101101000"; -- -0.1853337642880925
	pesos_i(7379) := b"1111111111111111_1111111111111111_1100011001010001_1111110000100000"; -- -0.22531151025829096
	pesos_i(7380) := b"0000000000000000_0000000000000000_0001011100000000_1010001111110110"; -- 0.08985352289604662
	pesos_i(7381) := b"0000000000000000_0000000000000000_0010010001010101_0111101110100101"; -- 0.14192936677516577
	pesos_i(7382) := b"0000000000000000_0000000000000000_0010100010101001_1111000111101100"; -- 0.15884315499416157
	pesos_i(7383) := b"1111111111111111_1111111111111111_1100100101111001_1010011000100011"; -- -0.21298753401128276
	pesos_i(7384) := b"1111111111111111_1111111111111111_1110101000111111_0000100111000000"; -- -0.0849756151866622
	pesos_i(7385) := b"0000000000000000_0000000000000000_0001111101111011_0101111000111100"; -- 0.12297619778375259
	pesos_i(7386) := b"1111111111111111_1111111111111111_1110101100001110_1111101110011010"; -- -0.08180263032736458
	pesos_i(7387) := b"0000000000000000_0000000000000000_0001100111001111_1100111011100110"; -- 0.10082715152157139
	pesos_i(7388) := b"0000000000000000_0000000000000000_0000010001111101_1110001101111100"; -- 0.017545907724518164
	pesos_i(7389) := b"1111111111111111_1111111111111111_1101010010111001_1001011100000001"; -- -0.1690431235028953
	pesos_i(7390) := b"0000000000000000_0000000000000000_0010111000011111_0101011001010100"; -- 0.18016566806444032
	pesos_i(7391) := b"0000000000000000_0000000000000000_0010001000100011_1001110101010100"; -- 0.1333559351464479
	pesos_i(7392) := b"0000000000000000_0000000000000000_0000010100111111_1011111100101000"; -- 0.020503947462236913
	pesos_i(7393) := b"1111111111111111_1111111111111111_1100101100011101_1010101100010010"; -- -0.20657854855057156
	pesos_i(7394) := b"0000000000000000_0000000000000000_0010001011010001_1011110100000100"; -- 0.13601285304476274
	pesos_i(7395) := b"1111111111111111_1111111111111111_1110110010011111_1010010011011101"; -- -0.07568902584664321
	pesos_i(7396) := b"0000000000000000_0000000000000000_0001100111000001_0110100000110111"; -- 0.1006074080728255
	pesos_i(7397) := b"0000000000000000_0000000000000000_0000111011001011_1000100011100010"; -- 0.05779319294559522
	pesos_i(7398) := b"1111111111111111_1111111111111111_1100111011011110_1011100000110111"; -- -0.19191406883139578
	pesos_i(7399) := b"1111111111111111_1111111111111111_1110110011101100_0000010101101100"; -- -0.07452360255001539
    return pesos_i;
    end function;
end package body mnist_weights;
    